* NGSPICE file created from mux4onehot_parax.ext - technology: sky130A

.subckt mux4onehot_parax select0 select1 A1 Z4 Z3 Z2 A2 Z1 A4 A3 VGND VPWR
X0 VGND.t97 passgatesCtrl_0.net2.t2 a_n597_n2040# VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND.t140 VPWR.t176 VGND.t139 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2 VPWR.t66 VGND.t177 VPWR.t65 VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3 VGND.t142 VPWR.t177 VGND.t141 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4 VPWR.t64 VGND.t178 VPWR.t63 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5 VGND.t41 a_n1361_n1429# passgatex4_0.GN3 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6 a_n1361_n1429# passgatesCtrl_0.net5 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7 VGND.t99 select1.t0 a_n2480_n4368# VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VGND.t157 VPWR.t178 VGND.t156 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X9 VGND.t53 a_n2189_n1429# passgatex4_0.GP3 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10 a_n2189_n1429# passgatesCtrl_0.net9 VPWR.t134 VPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11 passgatesCtrl_0.net6 a_n2975_n2192# VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12 a_n1084_n4216# a_n988_n4394# VGND.t112 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X13 VGND.t160 VPWR.t179 VGND.t159 VGND.t158 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X14 VPWR.t117 passgatesCtrl_0.net2.t3 a_n2161_n4368# VPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 VPWR.t138 a_n715_n3850# passgatesCtrl_0._04_ VPWR.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR.t62 VGND.t179 VPWR.t61 VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X17 a_n1913_n1429# passgatesCtrl_0.net10.t3 VGND.t68 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X18 a_n1173_n2218# a_n1003_n2040# a_n1045_n1942# VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 passgatex4_0.GN2 a_n951_n2736# VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X20 a_n801_n4216# passgatesCtrl_0.net1.t2 VGND.t168 VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X21 VPWR.t98 a_n1085_n1429# passgatex4_0.GP2 VPWR.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X22 Z3.t1 passgatex4_0.GN3 A3.t1 VGND.t154 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X23 VPWR.t60 VGND.t180 VPWR.t59 VPWR.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X24 Z3.t0 passgatex4_0.GN3 A3.t0 VGND.t154 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X25 VPWR.t175 a_n1459_n3306# a_n1635_n3306# VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X26 passgatesCtrl_0.net10.t2 passgatesCtrl_0.net1.t3 a_n2429_n1328# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VGND.t7 passgatesCtrl_0._01_ a_n1503_n2192# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X28 VGND.t137 passgatesCtrl_0.net3 a_n1227_n2736# VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X29 VPWR.t4 a_n995_n3605# passgatesCtrl_0.net4 VPWR.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X30 passgatex4_0.GP1 a_n491_n3280# VGND.t145 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X31 VGND.t105 passgatesCtrl_0.net7 a_n491_n3280# VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X32 VPWR.t74 passgatesCtrl_0._00_ a_n2883_n1648# VPWR.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X33 VGND.t173 VPWR.t180 VGND.t172 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X34 a_n715_n3850# passgatesCtrl_0.net1.t4 VPWR.t8 VPWR.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X35 VPWR.t125 a_n1637_n1429# passgatex4_0.GN4 VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X36 passgatex4_0.GN1 a_n1227_n2736# VPWR.t159 VPWR.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X37 passgatesCtrl_0.net7 a_n675_n1648# VPWR.t121 VPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X38 VGND.t155 passgatesCtrl_0._02_ a_n675_n1648# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X39 A3.t2 passgatex4_0.GP3 Z3.t3 VPWR.t172 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X40 VPWR.t58 VGND.t181 VPWR.t57 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X41 a_n482_n4216# select0.t0 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X42 VGND.t175 VPWR.t181 VGND.t174 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X43 a_n2185_n2218# a_n2015_n2040# a_n2057_n1942# VPWR.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 VPWR.t56 VGND.t182 VPWR.t55 VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X45 VGND.t107 a_n1635_n3306# passgatesCtrl_0._03_ VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X46 VPWR.t54 VGND.t183 VPWR.t53 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X47 VPWR.t52 VGND.t184 VPWR.t51 VPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X48 VPWR.t140 passgatesCtrl_0._05_ a_n2975_n2192# VPWR.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X49 VGND.t119 VPWR.t182 VGND.t118 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X50 VPWR.t128 a_n1635_n3306# passgatesCtrl_0._03_ VPWR.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X51 A2.t1 passgatex4_0.GP2 Z2.t0 VPWR.t85 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X52 VGND.t122 VPWR.t183 VGND.t121 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X53 VGND.t55 a_n1984_n4368# a_n1878_n4368# VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X54 VPWR.t49 VGND.t185 VPWR.t48 VPWR.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X55 a_n2189_n1429# passgatesCtrl_0.net9 VGND.t113 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X56 VPWR.t146 a_n1173_n2218# passgatesCtrl_0._01_ VPWR.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X57 VGND.t76 VPWR.t184 VGND.t75 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X58 VGND.t52 a_n1003_n2040# a_n1173_n2218# VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X59 a_n2429_n1328# passgatesCtrl_0.net2.t4 VGND.t95 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 VGND.t131 a_n1173_n2218# passgatesCtrl_0._01_ VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1755 ps=1.84 w=0.65 l=0.15
X61 VGND.t5 a_n995_n3605# passgatesCtrl_0.net4 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X62 VGND.t79 VPWR.t185 VGND.t78 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X63 a_n1003_n2040# passgatesCtrl_0.net1.t5 VGND.t135 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1575 ps=1.17 w=0.42 l=0.15
X64 VGND.t65 a_n1085_n1429# passgatex4_0.GP2 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X65 passgatesCtrl_0.net2.t1 a_n2480_n4368# VGND.t134 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X66 a_n1459_n3306# passgatesCtrl_0.net1.t6 VPWR.t155 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X67 VPWR.t47 VGND.t186 VPWR.t46 VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X68 a_n1085_n1429# passgatesCtrl_0.net8 VPWR.t84 VPWR.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X69 a_n715_n3850# a_n539_n3518# a_n587_n3458# VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X70 a_n587_n3458# passgatesCtrl_0.net1.t7 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X71 VGND.t21 VPWR.t186 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X72 passgatesCtrl_0.net2.t0 a_n2480_n4368# VPWR.t150 VPWR.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X73 passgatesCtrl_0.net8 a_n1503_n2192# VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X74 passgatex4_0.GN1 a_n1227_n2736# VGND.t153 VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X75 A4.t3 passgatex4_0.GP4 Z4.t2 VPWR.t163 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X76 Z4.t0 passgatex4_0.GN4 A4.t1 VGND.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X77 Z2.t2 passgatex4_0.GN2 A2.t3 VGND.t108 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X78 VPWR.t2 passgatesCtrl_0._03_ a_n1963_n3280# VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X79 VGND.t38 a_n801_n4216# a_n988_n4394# VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X80 passgatesCtrl_0.net9 a_n2883_n1648# VPWR.t144 VPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X81 VGND.t24 VPWR.t187 VGND.t23 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X82 VPWR.t153 a_n539_n3518# a_n715_n3850# VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X83 VGND.t36 passgatesCtrl_0._00_ a_n2883_n1648# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X84 a_n1637_n1429# passgatesCtrl_0.net6 VPWR.t148 VPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X85 VPWR.t76 a_n801_n4216# a_n988_n4394# VPWR.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X86 VGND.t103 a_n1637_n1429# passgatex4_0.GN4 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X87 VPWR.t45 VGND.t187 VPWR.t44 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X88 VPWR.t119 a_n2185_n2218# passgatesCtrl_0._00_ VPWR.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X89 Z2.t3 passgatex4_0.GN2 A2.t2 VGND.t108 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X90 VGND.t149 a_n1084_n4216# a_n1135_n4368# VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X91 passgatesCtrl_0.net7 a_n675_n1648# VGND.t102 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X92 VPWR.t123 passgatesCtrl_0.net1.t8 passgatesCtrl_0.net10.t1 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X93 VPWR.t157 a_n1084_n4216# a_n1135_n4368# VPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X94 VGND.t101 a_n2185_n2218# passgatesCtrl_0._00_ VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1755 ps=1.84 w=0.65 l=0.15
X95 VGND.t93 passgatesCtrl_0.net2.t5 a_n539_n3518# VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X96 a_n1173_n2218# passgatesCtrl_0.net2.t6 VGND.t91 VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X97 VGND.t89 passgatesCtrl_0.net2.t7 a_n2161_n4368# VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X98 VGND.t14 VPWR.t188 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X99 passgatesCtrl_0.net6 a_n2975_n2192# VPWR.t78 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X100 VPWR.t43 VGND.t188 VPWR.t42 VPWR.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X101 VGND.t17 VPWR.t189 VGND.t16 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X102 VPWR.t82 a_n2639_n2040# passgatesCtrl_0._05_ VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X103 VGND.t61 VPWR.t190 VGND.t60 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X104 VGND.t64 VPWR.t191 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X105 a_n2465_n2164# passgatesCtrl_0.net2.t8 VGND.t87 VGND.t86 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X106 VGND.t49 a_n2639_n2040# passgatesCtrl_0._05_ VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X107 VPWR.t158 passgatesCtrl_0.net4 a_n951_n2736# VPWR.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X108 a_n2015_n2040# passgatesCtrl_0.net2.t9 VGND.t85 VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1575 ps=1.17 w=0.42 l=0.15
X109 VPWR.t40 VGND.t189 VPWR.t39 VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X110 VPWR.t68 a_n1913_n1429# passgatex4_0.GP4 VPWR.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X111 VPWR.t6 passgatesCtrl_0._01_ a_n1503_n2192# VPWR.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X112 VPWR.t38 VGND.t190 VPWR.t37 VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X113 VGND.t83 passgatesCtrl_0.net2.t10 passgatesCtrl_0.net3 VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X114 A1.t3 passgatex4_0.GP1 Z1.t2 VPWR.t171 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X115 VGND.t128 a_n482_n4216# passgatesCtrl_0.net1.t0 VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X116 VPWR.t136 select1.t1 a_n2480_n4368# VPWR.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X117 a_n2185_n2218# passgatesCtrl_0.net1.t9 VGND.t126 VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X118 a_n1701_n4368# a_n1878_n4368# VGND.t162 VGND.t161 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X119 VPWR.t142 a_n482_n4216# passgatesCtrl_0.net1.t1 VPWR.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X120 a_n1085_n1429# passgatesCtrl_0.net8 VGND.t50 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X121 VPWR.t35 VGND.t191 VPWR.t34 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X122 VGND.t44 VPWR.t192 VGND.t43 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X123 Z4.t1 passgatex4_0.GN4 A4.t0 VGND.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X124 a_n1701_n4368# a_n1878_n4368# VPWR.t169 VPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X125 passgatesCtrl_0.net10.t0 passgatesCtrl_0.net2.t11 VPWR.t115 VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X126 a_n2639_n2040# passgatesCtrl_0.net2.t12 VPWR.t113 VPWR.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X127 VPWR.t102 passgatesCtrl_0.net1.t10 a_n1003_n2040# VPWR.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1176 ps=1.4 w=0.42 l=0.15
X128 VGND.t3 passgatesCtrl_0._03_ a_n1963_n3280# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X129 passgatesCtrl_0.net5 a_n1963_n3280# VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X130 a_n1084_n4216# a_n988_n4394# VPWR.t132 VPWR.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X131 a_n539_n3518# passgatesCtrl_0.net2.t13 VPWR.t111 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X132 passgatesCtrl_0.net9 a_n2883_n1648# VGND.t129 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X133 a_n1637_n1429# passgatesCtrl_0.net6 VGND.t132 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X134 a_n801_n4216# passgatesCtrl_0.net1.t11 VPWR.t174 VPWR.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X135 a_n2639_n2040# passgatesCtrl_0.net1.t12 a_n2465_n2164# VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X136 A3.t3 passgatex4_0.GP3 Z3.t2 VPWR.t172 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X137 VPWR.t12 a_n597_n2040# passgatesCtrl_0._02_ VPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X138 VPWR.t33 VGND.t192 VPWR.t32 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X139 VGND.t47 VPWR.t193 VGND.t46 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X140 a_n995_n3605# passgatesCtrl_0._04_ VPWR.t96 VPWR.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X141 a_n1507_n3280# passgatesCtrl_0.net2.t14 VGND.t81 VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X142 a_n1635_n3306# a_n1459_n3306# a_n1507_n3280# VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X143 VGND.t11 a_n597_n2040# passgatesCtrl_0._02_ VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X144 VGND.t32 VPWR.t194 VGND.t31 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X145 A2.t0 passgatex4_0.GP2 Z2.t1 VPWR.t85 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X146 VPWR.t30 VGND.t193 VPWR.t29 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X147 VGND.t151 passgatesCtrl_0.net4 a_n951_n2736# VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X148 VGND.t117 a_n715_n3850# passgatesCtrl_0._04_ VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X149 VPWR.t80 a_n1361_n1429# passgatex4_0.GN3 VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X150 a_n1361_n1429# passgatesCtrl_0.net5 VPWR.t10 VPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X151 VGND.t164 a_n2015_n2040# a_n2185_n2218# VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X152 VGND.t35 VPWR.t195 VGND.t34 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X153 VPWR.t27 VGND.t194 VPWR.t26 VPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X154 VGND.t71 VPWR.t196 VGND.t70 VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X155 VPWR.t90 passgatesCtrl_0.net1.t13 a_n2639_n2040# VPWR.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X156 a_n1045_n1942# passgatesCtrl_0.net2.t15 VPWR.t109 VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14825 ps=1.34 w=0.42 l=0.15
X157 VPWR.t92 a_n2189_n1429# passgatex4_0.GP3 VPWR.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X158 VGND.t124 passgatesCtrl_0._05_ a_n2975_n2192# VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X159 a_n482_n4216# select0.t1 VPWR.t162 VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X160 passgatesCtrl_0.net3 passgatesCtrl_0.net1.t14 VGND.t59 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X161 A1.t2 passgatex4_0.GP1 Z1.t3 VPWR.t171 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X162 VPWR.t24 VGND.t195 VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X163 VGND.t74 VPWR.t197 VGND.t73 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X164 VGND.t147 passgatesCtrl_0.net1.t15 a_n1459_n3306# VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X165 a_n1984_n4368# a_n2161_n4368# VGND.t110 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X166 VGND.t18 a_n1913_n1429# passgatex4_0.GP4 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X167 a_n1913_n1429# passgatesCtrl_0.net10.t4 VPWR.t72 VPWR.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X168 a_n1984_n4368# a_n2161_n4368# VPWR.t130 VPWR.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X169 passgatesCtrl_0.net8 a_n1503_n2192# VPWR.t70 VPWR.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X170 a_n597_n2040# passgatesCtrl_0.net2.t16 a_n434_n1942# VPWR.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X171 VPWR.t106 passgatesCtrl_0.net2.t17 a_n2015_n2040# VPWR.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1176 ps=1.4 w=0.42 l=0.15
X172 VPWR.t94 a_n1984_n4368# a_n1878_n4368# VPWR.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X173 a_n1635_n3306# passgatesCtrl_0.net2.t18 VPWR.t105 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X174 passgatex4_0.GN2 a_n951_n2736# VPWR.t100 VPWR.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X175 VPWR.t21 VGND.t196 VPWR.t20 VPWR.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X176 passgatesCtrl_0.net5 a_n1963_n3280# VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X177 a_n434_n1942# passgatesCtrl_0.net1.t16 VPWR.t167 VPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X178 passgatex4_0.GP1 a_n491_n3280# VPWR.t154 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X179 A4.t2 passgatex4_0.GP4 Z4.t3 VPWR.t163 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X180 VPWR.t126 passgatesCtrl_0.net7 a_n491_n3280# VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X181 a_n2057_n1942# passgatesCtrl_0.net1.t17 VPWR.t88 VPWR.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14825 ps=1.34 w=0.42 l=0.15
X182 Z1.t0 passgatex4_0.GN1 A1.t1 VGND.t166 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X183 a_n995_n3605# passgatesCtrl_0._04_ VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X184 VPWR.t18 VGND.t197 VPWR.t17 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X185 a_n597_n2040# passgatesCtrl_0.net1.t18 VGND.t170 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X186 passgatesCtrl_0.net3 passgatesCtrl_0.net2.t19 a_n485_n2736# VPWR.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X187 VPWR.t151 passgatesCtrl_0.net3 a_n1227_n2736# VPWR.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X188 Z1.t1 passgatex4_0.GN1 A1.t0 VGND.t165 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X189 VPWR.t165 passgatesCtrl_0._02_ a_n675_n1648# VPWR.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X190 VPWR.t15 VGND.t198 VPWR.t14 VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X191 a_n485_n2736# passgatesCtrl_0.net1.t19 VPWR.t160 VPWR.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
R0 passgatesCtrl_0.net2.n5 passgatesCtrl_0.net2.t15 562.236
R1 passgatesCtrl_0.net2.t15 passgatesCtrl_0.net2.t6 392.027
R2 passgatesCtrl_0.net2.n21 passgatesCtrl_0.net2.t13 327.99
R3 passgatesCtrl_0.net2.n2 passgatesCtrl_0.net2.t3 323.55
R4 passgatesCtrl_0.net2.n1 passgatesCtrl_0.net2.t0 319.171
R5 passgatesCtrl_0.net2.n18 passgatesCtrl_0.net2.t14 293.969
R6 passgatesCtrl_0.net2.n13 passgatesCtrl_0.net2.t12 261.887
R7 passgatesCtrl_0.net2.n6 passgatesCtrl_0.net2.t19 230.363
R8 passgatesCtrl_0.net2.n15 passgatesCtrl_0.net2.t11 229.369
R9 passgatesCtrl_0.net2 passgatesCtrl_0.net2.t1 209.923
R10 passgatesCtrl_0.net2.n21 passgatesCtrl_0.net2.t5 199.457
R11 passgatesCtrl_0.net2.n2 passgatesCtrl_0.net2.t7 195.017
R12 passgatesCtrl_0.net2.n8 passgatesCtrl_0.net2.t2 192.639
R13 passgatesCtrl_0.net2.n11 passgatesCtrl_0.net2.t9 185.376
R14 passgatesCtrl_0.net2.n6 passgatesCtrl_0.net2.t10 158.064
R15 passgatesCtrl_0.net2.n15 passgatesCtrl_0.net2.t4 157.07
R16 passgatesCtrl_0.net2.n13 passgatesCtrl_0.net2.t8 155.847
R17 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n8 154.286
R18 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n18 154.065
R19 passgatesCtrl_0.net2.n16 passgatesCtrl_0.net2.n15 153.66
R20 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n2 153.409
R21 passgatesCtrl_0.net2.n7 passgatesCtrl_0.net2.n6 153.097
R22 passgatesCtrl_0.net2.n22 passgatesCtrl_0.net2.n21 152
R23 passgatesCtrl_0.net2.n14 passgatesCtrl_0.net2.n13 152
R24 passgatesCtrl_0.net2.n12 passgatesCtrl_0.net2.n11 152
R25 passgatesCtrl_0.net2.n18 passgatesCtrl_0.net2.t18 138.338
R26 passgatesCtrl_0.net2.n11 passgatesCtrl_0.net2.t17 137.177
R27 passgatesCtrl_0.net2.n8 passgatesCtrl_0.net2.t16 134.799
R28 passgatesCtrl_0.net2.n10 passgatesCtrl_0.net2.n5 26.6879
R29 passgatesCtrl_0.net2.n23 passgatesCtrl_0.net2 24.7034
R30 passgatesCtrl_0.net2.n17 passgatesCtrl_0.net2.n16 21.1865
R31 passgatesCtrl_0.net2.n9 passgatesCtrl_0.net2.n7 21.1676
R32 passgatesCtrl_0.net2.n24 passgatesCtrl_0.net2.n23 17.5163
R33 passgatesCtrl_0.net2.n4 passgatesCtrl_0.net2 16.0005
R34 passgatesCtrl_0.net2.n19 passgatesCtrl_0.net2 15.4844
R35 passgatesCtrl_0.net2.n9 passgatesCtrl_0.net2 11.2434
R36 passgatesCtrl_0.net2.n0 passgatesCtrl_0.net2.n12 10.8365
R37 passgatesCtrl_0.net2.n17 passgatesCtrl_0.net2.n14 10.1066
R38 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n19 10.0713
R39 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n22 9.6005
R40 passgatesCtrl_0.net2.n0 passgatesCtrl_0.net2.n10 9.15538
R41 passgatesCtrl_0.net2.n5 passgatesCtrl_0.net2 8.92171
R42 passgatesCtrl_0.net2.n24 passgatesCtrl_0.net2.n4 8.88939
R43 passgatesCtrl_0.net2.n20 passgatesCtrl_0.net2.n0 8.61863
R44 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n24 7.82272
R45 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n1 7.73474
R46 passgatesCtrl_0.net2.n10 passgatesCtrl_0.net2.n9 7.03724
R47 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n3 6.34564
R48 passgatesCtrl_0.net2.n4 passgatesCtrl_0.net2 6.0165
R49 passgatesCtrl_0.net2.n4 passgatesCtrl_0.net2 5.7605
R50 passgatesCtrl_0.net2.n20 passgatesCtrl_0.net2 5.25599
R51 passgatesCtrl_0.net2.n22 passgatesCtrl_0.net2 4.90717
R52 passgatesCtrl_0.net2.n16 passgatesCtrl_0.net2 4.26717
R53 passgatesCtrl_0.net2.n14 passgatesCtrl_0.net2 3.8405
R54 passgatesCtrl_0.net2.n19 passgatesCtrl_0.net2 3.51018
R55 passgatesCtrl_0.net2.n7 passgatesCtrl_0.net2 3.10907
R56 passgatesCtrl_0.net2.n12 passgatesCtrl_0.net2 3.0725
R57 passgatesCtrl_0.net2.n0 passgatesCtrl_0.net2.n17 2.62704
R58 passgatesCtrl_0.net2.n1 passgatesCtrl_0.net2 2.48634
R59 passgatesCtrl_0.net2.n23 passgatesCtrl_0.net2.n20 2.2972
R60 passgatesCtrl_0.net2.n3 passgatesCtrl_0.net2 2.19479
R61 passgatesCtrl_0.net2.n3 passgatesCtrl_0.net2 1.80756
R62 VGND.t165 VGND.n7 13018.9
R63 VGND.n115 VGND.n114 12462.1
R64 VGND.n108 VGND.n92 12047.7
R65 VGND.n135 VGND.n94 11744.7
R66 VGND.n135 VGND.n95 11744.7
R67 VGND.n94 VGND.n93 11744.7
R68 VGND.n95 VGND.n93 11744.7
R69 VGND.n121 VGND.n100 11744.7
R70 VGND.n121 VGND.n101 11744.7
R71 VGND.n120 VGND.n100 11744.7
R72 VGND.n120 VGND.n101 11744.7
R73 VGND.n113 VGND.n102 11744.7
R74 VGND.n109 VGND.n102 11744.7
R75 VGND.n113 VGND.n103 11744.7
R76 VGND.n109 VGND.n103 11744.7
R77 VGND.n562 VGND.n4 11744.7
R78 VGND.n562 VGND.n5 11744.7
R79 VGND.n560 VGND.n5 11744.7
R80 VGND.n560 VGND.n4 11744.7
R81 VGND.n387 VGND 10843
R82 VGND.n387 VGND.n386 10123.6
R83 VGND.n386 VGND.n385 10123.6
R84 VGND.n137 VGND.n136 3869.02
R85 VGND.n136 VGND.n91 3771.63
R86 VGND.n116 VGND.n91 3735.78
R87 VGND.n561 VGND.n6 3570.22
R88 VGND.n558 VGND.t165 2593.05
R89 VGND.t165 VGND 2390.62
R90 VGND.n561 VGND.n558 2369.23
R91 VGND.t69 VGND.t138 2326.44
R92 VGND.n388 VGND.t19 1938.7
R93 VGND VGND.t12 1694.25
R94 VGND VGND.t15 1601.53
R95 VGND.n386 VGND 1601.53
R96 VGND VGND.n387 1601.53
R97 VGND.t176 VGND.t146 1584.67
R98 VGND.t0 VGND.t77 1567.82
R99 VGND.t163 VGND.t84 1517.24
R100 VGND VGND.t30 1407.66
R101 VGND.t166 VGND.n6 1392.06
R102 VGND VGND.t100 1340.23
R103 VGND VGND.t4 1230.65
R104 VGND.t120 VGND.t158 1219.28
R105 VGND.n384 VGND.n383 1194.5
R106 VGND.n254 VGND.t48 1194.5
R107 VGND.n557 VGND.n556 1194.5
R108 VGND.n389 VGND.n388 1194.5
R109 VGND VGND.t62 1019.92
R110 VGND.t19 VGND 1019.92
R111 VGND VGND.t10 977.779
R112 VGND.t48 VGND 918.774
R113 VGND.t30 VGND 918.774
R114 VGND.n388 VGND 918.774
R115 VGND.t138 VGND 918.774
R116 VGND.t48 VGND.t86 910.346
R117 VGND.t22 VGND 893.633
R118 VGND VGND.n6 851.341
R119 VGND.n558 VGND 851.341
R120 VGND.t127 VGND.t167 848.193
R121 VGND.t88 VGND.t133 848.193
R122 VGND.t100 VGND.t125 826.054
R123 VGND.t116 VGND.t114 826.054
R124 VGND.t106 VGND.t80 826.054
R125 VGND.t42 VGND.t116 792.337
R126 VGND.n112 VGND.n111 767.294
R127 VGND.n559 VGND.n3 767.294
R128 VGND.n131 VGND.n130 763.106
R129 VGND.n119 VGND.n99 763.106
R130 VGND.t33 VGND 742.169
R131 VGND.t150 VGND.t66 741.763
R132 VGND.t6 VGND.t25 741.763
R133 VGND.t39 VGND.t123 741.763
R134 VGND.t104 VGND.t92 741.763
R135 VGND.t4 VGND.t56 741.763
R136 VGND.t2 VGND.t0 741.763
R137 VGND.n130 VGND.n96 732.236
R138 VGND.n123 VGND.n99 732.236
R139 VGND.n112 VGND.n104 732.236
R140 VGND.n559 VGND.n1 732.236
R141 VGND.t130 VGND.t152 724.904
R142 VGND.t37 VGND.t111 711.876
R143 VGND.t54 VGND.t109 711.876
R144 VGND.t90 VGND.t51 708.047
R145 VGND.t125 VGND.t163 708.047
R146 VGND.t80 VGND.t176 657.471
R147 VGND.t15 VGND 632.184
R148 VGND.t12 VGND 632.184
R149 VGND.t148 VGND 594.492
R150 VGND.t144 VGND 564.751
R151 VGND VGND.t6 547.894
R152 VGND.t123 VGND 547.894
R153 VGND VGND.t2 547.894
R154 VGND.t58 VGND.t169 531.034
R155 VGND VGND.t150 531.034
R156 VGND VGND.t136 531.034
R157 VGND VGND.t104 531.034
R158 VGND VGND.t42 531.034
R159 VGND VGND.t161 507.401
R160 VGND.t96 VGND 505.748
R161 VGND.t86 VGND 497.318
R162 VGND VGND.t143 480.461
R163 VGND.n385 VGND.t166 479.757
R164 VGND VGND.t22 458.176
R165 VGND.t158 VGND 458.176
R166 VGND.n557 VGND 412.738
R167 VGND VGND.t120 412.738
R168 VGND.t98 VGND 397.591
R169 VGND.t72 VGND.t69 387.74
R170 VGND.t28 VGND.t127 359.726
R171 VGND.t167 VGND.t37 359.726
R172 VGND.t111 VGND.t148 359.726
R173 VGND.t161 VGND.t54 359.726
R174 VGND.t109 VGND.t88 359.726
R175 VGND.t133 VGND.t98 359.726
R176 VGND.n111 VGND.n110 325.502
R177 VGND.n563 VGND.n3 325.502
R178 VGND.t143 VGND 311.877
R179 VGND.n132 VGND.n131 304.204
R180 VGND.n119 VGND.n118 304.204
R181 VGND.t10 VGND.t58 286.591
R182 VGND VGND.t33 283.993
R183 VGND VGND.t96 278.161
R184 VGND.n226 VGND.t173 273.171
R185 VGND.n431 VGND.t79 273.171
R186 VGND VGND.t28 268.848
R187 VGND VGND.n557 265.06
R188 VGND.n158 VGND.t191 262.719
R189 VGND.n70 VGND.t195 262.719
R190 VGND.t25 VGND 261.303
R191 VGND.t92 VGND 261.303
R192 VGND.t56 VGND 261.303
R193 VGND.t146 VGND 261.303
R194 VGND.n393 VGND.t186 259.082
R195 VGND.n49 VGND.t179 259.082
R196 VGND.n48 VGND.t177 259.082
R197 VGND.n395 VGND.t189 259.082
R198 VGND.n394 VGND.t188 259.082
R199 VGND.n372 VGND.t197 259.082
R200 VGND.n304 VGND.t187 259.082
R201 VGND.n175 VGND.t193 259.082
R202 VGND.n174 VGND.t192 259.082
R203 VGND.n243 VGND.t183 259.082
R204 VGND.n242 VGND.t181 259.082
R205 VGND.n468 VGND.t190 259.082
R206 VGND.n544 VGND.t180 259.082
R207 VGND.t82 VGND 252.875
R208 VGND.t66 VGND 252.875
R209 VGND.n158 VGND.t172 251.564
R210 VGND.n70 VGND.t78 251.564
R211 VGND.t51 VGND 244.445
R212 VGND VGND.t72 244.445
R213 VGND.n133 VGND.n132 242.448
R214 VGND.n118 VGND.n98 242.448
R215 VGND.n110 VGND.n107 242.448
R216 VGND.n564 VGND.n563 242.448
R217 VGND.n179 VGND.t97 241.971
R218 VGND.n411 VGND.t21 240.72
R219 VGND.n439 VGND.t147 237.327
R220 VGND.n53 VGND.t93 237.327
R221 VGND.t171 VGND 236.016
R222 VGND.n64 VGND.t44 233.073
R223 VGND.n241 VGND.t64 225.427
R224 VGND.n504 VGND.t24 225.427
R225 VGND.n551 VGND.t160 225.427
R226 VGND.n411 VGND.t76 225.427
R227 VGND.n391 VGND.t74 225.427
R228 VGND.n89 VGND.t20 225.261
R229 VGND.n401 VGND.t71 221.793
R230 VGND.n51 VGND.t14 221.793
R231 VGND.n51 VGND.t61 221.793
R232 VGND.n396 VGND.t139 221.793
R233 VGND.n396 VGND.t156 221.793
R234 VGND.n373 VGND.t174 221.793
R235 VGND.n305 VGND.t47 221.793
R236 VGND.n177 VGND.t17 221.793
R237 VGND.n177 VGND.t119 221.793
R238 VGND.n244 VGND.t141 221.793
R239 VGND.n244 VGND.t31 221.793
R240 VGND.n469 VGND.t35 221.793
R241 VGND.n545 VGND.t121 221.793
R242 VGND.n42 VGND.t43 221.603
R243 VGND.n240 VGND.t178 218.308
R244 VGND.n24 VGND.t184 218.308
R245 VGND.n542 VGND.t196 218.308
R246 VGND.n90 VGND.t194 218.308
R247 VGND.n390 VGND.t185 218.308
R248 VGND.n240 VGND.t63 217.78
R249 VGND.n24 VGND.t23 217.78
R250 VGND.n542 VGND.t159 217.78
R251 VGND.n90 VGND.t75 217.78
R252 VGND.n390 VGND.t73 217.78
R253 VGND.n393 VGND.t70 215.905
R254 VGND.n49 VGND.t13 215.905
R255 VGND.n48 VGND.t60 215.905
R256 VGND.n395 VGND.t140 215.905
R257 VGND.n394 VGND.t157 215.905
R258 VGND.n372 VGND.t175 215.905
R259 VGND.n304 VGND.t46 215.905
R260 VGND.n175 VGND.t16 215.905
R261 VGND.n174 VGND.t118 215.905
R262 VGND.n243 VGND.t142 215.905
R263 VGND.n242 VGND.t32 215.905
R264 VGND.n468 VGND.t34 215.905
R265 VGND.n544 VGND.t122 215.905
R266 VGND VGND.t144 210.728
R267 VGND.n185 VGND.n184 205.541
R268 VGND.n236 VGND.n235 200.105
R269 VGND.n433 VGND.n69 197.476
R270 VGND.n44 VGND.n43 197.476
R271 VGND.n426 VGND.n73 196.442
R272 VGND.n445 VGND.n41 196.442
R273 VGND.n46 VGND.n45 196.442
R274 VGND.n379 VGND.n370 196.442
R275 VGND.n142 VGND.n141 196.442
R276 VGND.n281 VGND.n280 196.442
R277 VGND.n341 VGND.n283 196.442
R278 VGND.n336 VGND.n286 196.442
R279 VGND.n331 VGND.n289 196.442
R280 VGND.n301 VGND.n300 196.442
R281 VGND.n249 VGND.n239 196.442
R282 VGND.n161 VGND.n160 196.442
R283 VGND.n163 VGND.n162 196.442
R284 VGND.n192 VGND.n191 196.442
R285 VGND.n210 VGND.n209 195.612
R286 VGND.n232 VGND.n155 195.612
R287 VGND.n111 VGND.n103 195
R288 VGND.n103 VGND.t154 195
R289 VGND.n106 VGND.n102 195
R290 VGND.n102 VGND.t154 195
R291 VGND.n120 VGND.n119 195
R292 VGND.t27 VGND.n120 195
R293 VGND.n122 VGND.n121 195
R294 VGND.n121 VGND.t27 195
R295 VGND.n131 VGND.n93 195
R296 VGND.t108 VGND.n93 195
R297 VGND.n135 VGND.n134 195
R298 VGND.t108 VGND.n135 195
R299 VGND.n4 VGND.n2 195
R300 VGND.n137 VGND.n4 195
R301 VGND.n5 VGND.n3 195
R302 VGND.t165 VGND.n5 195
R303 VGND.n475 VGND.n466 194.809
R304 VGND.n481 VGND.n463 194.809
R305 VGND.n497 VGND.n27 194.809
R306 VGND.n512 VGND.n511 194.809
R307 VGND.n519 VGND.n518 194.809
R308 VGND.n537 VGND.n11 194.809
R309 VGND.t169 VGND.t82 177.012
R310 VGND.t114 VGND 177.012
R311 VGND.n117 VGND.n100 172.754
R312 VGND.n114 VGND.t154 161.819
R313 VGND.t108 VGND.n92 161.685
R314 VGND.n172 VGND.t83 152.381
R315 VGND.n171 VGND.t59 150.101
R316 VGND.n365 VGND.t95 147.411
R317 VGND VGND.n137 133.785
R318 VGND.n385 VGND.n384 131.803
R319 VGND.n42 VGND.t182 116.734
R320 VGND.n116 VGND.n115 103.636
R321 VGND.t152 VGND.t90 101.15
R322 VGND.n89 VGND.t198 99.7822
R323 VGND.n108 VGND.n91 97.2732
R324 VGND.n136 VGND.n7 97.1929
R325 VGND.n165 VGND.t135 89.3384
R326 VGND.n156 VGND.t85 89.3384
R327 VGND.n165 VGND.t52 88.7758
R328 VGND.n156 VGND.t164 88.7758
R329 VGND.t8 VGND 81.2618
R330 VGND.n235 VGND.t87 72.8576
R331 VGND.n166 VGND.n165 70.4565
R332 VGND.n157 VGND.n156 70.4565
R333 VGND.t154 VGND.n91 64.546
R334 VGND.n136 VGND.t108 64.4927
R335 VGND.n69 VGND.t81 58.5719
R336 VGND.n43 VGND.t115 58.5719
R337 VGND.n117 VGND.n116 58.1458
R338 VGND.n184 VGND.t170 55.7148
R339 VGND.n209 VGND.t91 52.8576
R340 VGND.n155 VGND.t126 52.8576
R341 VGND.n466 VGND.t29 45.7148
R342 VGND.n463 VGND.t168 45.7148
R343 VGND.n27 VGND.t112 45.7148
R344 VGND.n511 VGND.t55 45.7148
R345 VGND.n518 VGND.t89 45.7148
R346 VGND.n11 VGND.t99 45.7148
R347 VGND.n305 VGND.n303 34.6358
R348 VGND.n309 VGND.n303 34.6358
R349 VGND.n310 VGND.n309 34.6358
R350 VGND.n311 VGND.n310 34.6358
R351 VGND.n311 VGND.n301 34.6358
R352 VGND.n315 VGND.n301 34.6358
R353 VGND.n316 VGND.n315 34.6358
R354 VGND.n316 VGND.n290 34.6358
R355 VGND.n330 VGND.n290 34.6358
R356 VGND.n331 VGND.n330 34.6358
R357 VGND.n331 VGND.n287 34.6358
R358 VGND.n335 VGND.n287 34.6358
R359 VGND.n336 VGND.n335 34.6358
R360 VGND.n337 VGND.n336 34.6358
R361 VGND.n337 VGND.n284 34.6358
R362 VGND.n341 VGND.n284 34.6358
R363 VGND.n342 VGND.n341 34.6358
R364 VGND.n343 VGND.n342 34.6358
R365 VGND.n343 VGND.n281 34.6358
R366 VGND.n347 VGND.n281 34.6358
R367 VGND.n348 VGND.n347 34.6358
R368 VGND.n348 VGND.n142 34.6358
R369 VGND.n363 VGND.n142 34.6358
R370 VGND.n364 VGND.n363 34.6358
R371 VGND.n366 VGND.n364 34.6358
R372 VGND.n383 VGND.n138 34.6358
R373 VGND.n383 VGND.n139 34.6358
R374 VGND.n379 VGND.n139 34.6358
R375 VGND.n379 VGND.n378 34.6358
R376 VGND.n378 VGND.n377 34.6358
R377 VGND.n377 VGND.n371 34.6358
R378 VGND.n373 VGND.n371 34.6358
R379 VGND.n178 VGND.n177 34.6358
R380 VGND.n180 VGND.n178 34.6358
R381 VGND.n186 VGND.n183 34.6358
R382 VGND.n190 VGND.n171 34.6358
R383 VGND.n193 VGND.n190 34.6358
R384 VGND.n193 VGND.n192 34.6358
R385 VGND.n211 VGND.n208 34.6358
R386 VGND.n215 VGND.n163 34.6358
R387 VGND.n216 VGND.n215 34.6358
R388 VGND.n216 VGND.n161 34.6358
R389 VGND.n220 VGND.n161 34.6358
R390 VGND.n221 VGND.n220 34.6358
R391 VGND.n221 VGND.n159 34.6358
R392 VGND.n225 VGND.n159 34.6358
R393 VGND.n231 VGND.n230 34.6358
R394 VGND.n269 VGND.n268 34.6358
R395 VGND.n268 VGND.n233 34.6358
R396 VGND.n258 VGND.n233 34.6358
R397 VGND.n258 VGND.n257 34.6358
R398 VGND.n254 VGND.n253 34.6358
R399 VGND.n253 VGND.n237 34.6358
R400 VGND.n249 VGND.n248 34.6358
R401 VGND.n248 VGND.n247 34.6358
R402 VGND.n247 VGND.n244 34.6358
R403 VGND.n469 VGND.n467 34.6358
R404 VGND.n473 VGND.n467 34.6358
R405 VGND.n474 VGND.n473 34.6358
R406 VGND.n476 VGND.n464 34.6358
R407 VGND.n480 VGND.n464 34.6358
R408 VGND.n482 VGND.n28 34.6358
R409 VGND.n496 VGND.n28 34.6358
R410 VGND.n498 VGND.n25 34.6358
R411 VGND.n502 VGND.n25 34.6358
R412 VGND.n503 VGND.n502 34.6358
R413 VGND.n505 VGND.n22 34.6358
R414 VGND.n509 VGND.n22 34.6358
R415 VGND.n510 VGND.n509 34.6358
R416 VGND.n513 VGND.n510 34.6358
R417 VGND.n517 VGND.n20 34.6358
R418 VGND.n520 VGND.n517 34.6358
R419 VGND.n535 VGND.n12 34.6358
R420 VGND.n536 VGND.n535 34.6358
R421 VGND.n538 VGND.n8 34.6358
R422 VGND.n556 VGND.n8 34.6358
R423 VGND.n556 VGND.n9 34.6358
R424 VGND.n552 VGND.n9 34.6358
R425 VGND.n550 VGND.n549 34.6358
R426 VGND.n549 VGND.n543 34.6358
R427 VGND.n545 VGND.n543 34.6358
R428 VGND.n52 VGND.n51 34.6358
R429 VGND.n54 VGND.n52 34.6358
R430 VGND.n58 VGND.n46 34.6358
R431 VGND.n59 VGND.n58 34.6358
R432 VGND.n63 VGND.n62 34.6358
R433 VGND.n445 VGND.n65 34.6358
R434 VGND.n445 VGND.n444 34.6358
R435 VGND.n444 VGND.n66 34.6358
R436 VGND.n440 VGND.n66 34.6358
R437 VGND.n438 VGND.n67 34.6358
R438 VGND.n434 VGND.n67 34.6358
R439 VGND.n430 VGND.n71 34.6358
R440 VGND.n426 VGND.n71 34.6358
R441 VGND.n426 VGND.n425 34.6358
R442 VGND.n425 VGND.n424 34.6358
R443 VGND.n424 VGND.n74 34.6358
R444 VGND.n88 VGND.n74 34.6358
R445 VGND.n412 VGND.n88 34.6358
R446 VGND.n410 VGND.n409 34.6358
R447 VGND.n409 VGND.n389 34.6358
R448 VGND.n405 VGND.n389 34.6358
R449 VGND.n405 VGND.n404 34.6358
R450 VGND.n401 VGND.n400 34.6358
R451 VGND.n400 VGND.n399 34.6358
R452 VGND.n399 VGND.n396 34.6358
R453 VGND.n466 VGND.t128 34.506
R454 VGND.n463 VGND.t38 34.506
R455 VGND.n27 VGND.t149 34.506
R456 VGND.n511 VGND.t162 34.506
R457 VGND.n518 VGND.t110 34.506
R458 VGND.n11 VGND.t134 34.506
R459 VGND.n366 VGND.n365 33.8829
R460 VGND.n497 VGND.n496 33.5064
R461 VGND.n73 VGND.t1 33.462
R462 VGND.n73 VGND.t3 33.462
R463 VGND.n41 VGND.t57 33.462
R464 VGND.n41 VGND.t5 33.462
R465 VGND.n45 VGND.t145 33.462
R466 VGND.n45 VGND.t105 33.462
R467 VGND.n370 VGND.t129 33.462
R468 VGND.n370 VGND.t36 33.462
R469 VGND.n141 VGND.t113 33.462
R470 VGND.n141 VGND.t53 33.462
R471 VGND.n280 VGND.t68 33.462
R472 VGND.n280 VGND.t18 33.462
R473 VGND.n283 VGND.t132 33.462
R474 VGND.n283 VGND.t103 33.462
R475 VGND.n286 VGND.t9 33.462
R476 VGND.n286 VGND.t41 33.462
R477 VGND.n289 VGND.t50 33.462
R478 VGND.n289 VGND.t65 33.462
R479 VGND.n300 VGND.t102 33.462
R480 VGND.n300 VGND.t155 33.462
R481 VGND.n239 VGND.t40 33.462
R482 VGND.n239 VGND.t124 33.462
R483 VGND.n160 VGND.t26 33.462
R484 VGND.n160 VGND.t7 33.462
R485 VGND.n162 VGND.t153 33.462
R486 VGND.n162 VGND.t137 33.462
R487 VGND.n191 VGND.t67 33.462
R488 VGND.n191 VGND.t151 33.462
R489 VGND.n512 VGND.n20 33.1299
R490 VGND.n59 VGND.n44 33.1299
R491 VGND.n434 VGND.n433 33.1299
R492 VGND.n53 VGND.n46 32.377
R493 VGND.n439 VGND.n438 32.377
R494 VGND.n211 VGND.n210 31.2476
R495 VGND.n232 VGND.n231 31.2476
R496 VGND.n134 VGND.n96 30.8711
R497 VGND.n123 VGND.n122 30.8711
R498 VGND.n106 VGND.n104 30.8711
R499 VGND.n481 VGND.n480 30.8711
R500 VGND.n2 VGND.n1 30.8711
R501 VGND.n519 VGND.n12 30.4946
R502 VGND.n209 VGND.t131 28.3166
R503 VGND.n155 VGND.t101 28.3166
R504 VGND.n184 VGND.t11 26.8576
R505 VGND.n69 VGND.t107 25.4291
R506 VGND.n43 VGND.t117 25.4291
R507 VGND.n185 VGND.n171 24.0946
R508 VGND.n179 VGND.n172 23.7181
R509 VGND.n235 VGND.t49 22.3257
R510 VGND.n226 VGND.n158 21.6078
R511 VGND.n431 VGND.n70 21.6078
R512 VGND.n192 VGND.n166 20.3299
R513 VGND.n227 VGND.n157 20.3299
R514 VGND.n537 VGND.n536 20.3299
R515 VGND.n476 VGND.n475 19.9534
R516 VGND.n254 VGND.n236 18.824
R517 VGND.n226 VGND.n225 17.3181
R518 VGND.n227 VGND.n226 17.3181
R519 VGND.n241 VGND.n237 17.3181
R520 VGND.n249 VGND.n241 17.3181
R521 VGND.n504 VGND.n503 17.3181
R522 VGND.n505 VGND.n504 17.3181
R523 VGND.n552 VGND.n551 17.3181
R524 VGND.n551 VGND.n550 17.3181
R525 VGND.n64 VGND.n63 17.3181
R526 VGND.n65 VGND.n64 17.3181
R527 VGND.n432 VGND.n431 17.3181
R528 VGND.n431 VGND.n430 17.3181
R529 VGND.n412 VGND.n411 17.3181
R530 VGND.n411 VGND.n410 17.3181
R531 VGND.n404 VGND.n391 17.3181
R532 VGND.n401 VGND.n391 17.3181
R533 VGND.t136 VGND.t130 16.8587
R534 VGND.t84 VGND.t171 16.8587
R535 VGND.t62 VGND.t39 16.8587
R536 VGND.t77 VGND.t106 16.8587
R537 VGND.n384 VGND.t94 15.8564
R538 VGND.n257 VGND.n236 15.8123
R539 VGND.n411 VGND.n89 15.4602
R540 VGND.n475 VGND.n474 14.6829
R541 VGND.n208 VGND.n166 14.3064
R542 VGND.n230 VGND.n157 14.3064
R543 VGND.n538 VGND.n537 14.3064
R544 VGND.n81 VGND 13.1605
R545 VGND.n64 VGND.n42 11.4706
R546 VGND.n110 VGND.n109 11.0382
R547 VGND.n109 VGND.n108 11.0382
R548 VGND.n113 VGND.n112 11.0382
R549 VGND.n114 VGND.n113 11.0382
R550 VGND.n118 VGND.n101 11.0382
R551 VGND.n115 VGND.n101 11.0382
R552 VGND.n100 VGND.n99 11.0382
R553 VGND.n132 VGND.n95 11.0382
R554 VGND.n95 VGND.n7 11.0382
R555 VGND.n130 VGND.n94 11.0382
R556 VGND.n94 VGND.n92 11.0382
R557 VGND.n560 VGND.n559 11.0382
R558 VGND.n561 VGND.n560 11.0382
R559 VGND.n563 VGND.n562 11.0382
R560 VGND.n562 VGND.n561 11.0382
R561 VGND.n134 VGND.n133 10.9181
R562 VGND.n122 VGND.n98 10.9181
R563 VGND.n107 VGND.n106 10.9181
R564 VGND.n564 VGND.n2 10.9181
R565 VGND.n180 VGND.n179 10.5417
R566 VGND.n186 VGND.n185 10.5417
R567 VGND.n129 VGND.n96 10.4476
R568 VGND.n124 VGND.n123 10.4476
R569 VGND.n105 VGND.n104 10.4476
R570 VGND.n565 VGND.n1 10.4476
R571 VGND.t94 VGND.t45 9.91041
R572 VGND.n307 VGND.n303 9.3005
R573 VGND.n309 VGND.n308 9.3005
R574 VGND.n310 VGND.n302 9.3005
R575 VGND.n312 VGND.n311 9.3005
R576 VGND.n313 VGND.n301 9.3005
R577 VGND.n315 VGND.n314 9.3005
R578 VGND.n317 VGND.n316 9.3005
R579 VGND.n291 VGND.n290 9.3005
R580 VGND.n330 VGND.n329 9.3005
R581 VGND.n332 VGND.n331 9.3005
R582 VGND.n333 VGND.n287 9.3005
R583 VGND.n335 VGND.n334 9.3005
R584 VGND.n336 VGND.n285 9.3005
R585 VGND.n338 VGND.n337 9.3005
R586 VGND.n339 VGND.n284 9.3005
R587 VGND.n341 VGND.n340 9.3005
R588 VGND.n342 VGND.n282 9.3005
R589 VGND.n344 VGND.n343 9.3005
R590 VGND.n345 VGND.n281 9.3005
R591 VGND.n347 VGND.n346 9.3005
R592 VGND.n349 VGND.n348 9.3005
R593 VGND.n353 VGND.n142 9.3005
R594 VGND.n363 VGND.n362 9.3005
R595 VGND.n364 VGND.n140 9.3005
R596 VGND.n367 VGND.n366 9.3005
R597 VGND.n368 VGND.n138 9.3005
R598 VGND.n383 VGND.n382 9.3005
R599 VGND.n381 VGND.n139 9.3005
R600 VGND.n380 VGND.n379 9.3005
R601 VGND.n378 VGND.n369 9.3005
R602 VGND.n377 VGND.n376 9.3005
R603 VGND.n375 VGND.n371 9.3005
R604 VGND.n247 VGND.n246 9.3005
R605 VGND.n178 VGND.n173 9.3005
R606 VGND.n181 VGND.n180 9.3005
R607 VGND.n183 VGND.n182 9.3005
R608 VGND.n187 VGND.n186 9.3005
R609 VGND.n188 VGND.n171 9.3005
R610 VGND.n190 VGND.n189 9.3005
R611 VGND.n194 VGND.n193 9.3005
R612 VGND.n192 VGND.n167 9.3005
R613 VGND.n208 VGND.n207 9.3005
R614 VGND.n212 VGND.n211 9.3005
R615 VGND.n213 VGND.n163 9.3005
R616 VGND.n215 VGND.n214 9.3005
R617 VGND.n217 VGND.n216 9.3005
R618 VGND.n218 VGND.n161 9.3005
R619 VGND.n220 VGND.n219 9.3005
R620 VGND.n222 VGND.n221 9.3005
R621 VGND.n223 VGND.n159 9.3005
R622 VGND.n225 VGND.n224 9.3005
R623 VGND.n228 VGND.n227 9.3005
R624 VGND.n230 VGND.n229 9.3005
R625 VGND.n231 VGND.n153 9.3005
R626 VGND.n270 VGND.n269 9.3005
R627 VGND.n268 VGND.n267 9.3005
R628 VGND.n260 VGND.n233 9.3005
R629 VGND.n259 VGND.n258 9.3005
R630 VGND.n257 VGND.n256 9.3005
R631 VGND.n255 VGND.n254 9.3005
R632 VGND.n253 VGND.n252 9.3005
R633 VGND.n251 VGND.n237 9.3005
R634 VGND.n250 VGND.n249 9.3005
R635 VGND.n248 VGND.n238 9.3005
R636 VGND.n547 VGND.n543 9.3005
R637 VGND.n471 VGND.n467 9.3005
R638 VGND.n473 VGND.n472 9.3005
R639 VGND.n474 VGND.n465 9.3005
R640 VGND.n477 VGND.n476 9.3005
R641 VGND.n478 VGND.n464 9.3005
R642 VGND.n480 VGND.n479 9.3005
R643 VGND.n483 VGND.n482 9.3005
R644 VGND.n29 VGND.n28 9.3005
R645 VGND.n496 VGND.n495 9.3005
R646 VGND.n499 VGND.n498 9.3005
R647 VGND.n500 VGND.n25 9.3005
R648 VGND.n502 VGND.n501 9.3005
R649 VGND.n503 VGND.n23 9.3005
R650 VGND.n506 VGND.n505 9.3005
R651 VGND.n507 VGND.n22 9.3005
R652 VGND.n509 VGND.n508 9.3005
R653 VGND.n510 VGND.n21 9.3005
R654 VGND.n514 VGND.n513 9.3005
R655 VGND.n515 VGND.n20 9.3005
R656 VGND.n517 VGND.n516 9.3005
R657 VGND.n521 VGND.n520 9.3005
R658 VGND.n525 VGND.n12 9.3005
R659 VGND.n535 VGND.n534 9.3005
R660 VGND.n536 VGND.n10 9.3005
R661 VGND.n539 VGND.n538 9.3005
R662 VGND.n540 VGND.n8 9.3005
R663 VGND.n556 VGND.n555 9.3005
R664 VGND.n554 VGND.n9 9.3005
R665 VGND.n553 VGND.n552 9.3005
R666 VGND.n550 VGND.n541 9.3005
R667 VGND.n549 VGND.n548 9.3005
R668 VGND.n399 VGND.n398 9.3005
R669 VGND.n52 VGND.n47 9.3005
R670 VGND.n55 VGND.n54 9.3005
R671 VGND.n56 VGND.n46 9.3005
R672 VGND.n58 VGND.n57 9.3005
R673 VGND.n60 VGND.n59 9.3005
R674 VGND.n62 VGND.n61 9.3005
R675 VGND.n63 VGND.n37 9.3005
R676 VGND.n65 VGND.n38 9.3005
R677 VGND.n446 VGND.n445 9.3005
R678 VGND.n444 VGND.n443 9.3005
R679 VGND.n442 VGND.n66 9.3005
R680 VGND.n441 VGND.n440 9.3005
R681 VGND.n438 VGND.n437 9.3005
R682 VGND.n436 VGND.n67 9.3005
R683 VGND.n435 VGND.n434 9.3005
R684 VGND.n432 VGND.n68 9.3005
R685 VGND.n430 VGND.n429 9.3005
R686 VGND.n428 VGND.n71 9.3005
R687 VGND.n427 VGND.n426 9.3005
R688 VGND.n425 VGND.n72 9.3005
R689 VGND.n424 VGND.n423 9.3005
R690 VGND.n76 VGND.n74 9.3005
R691 VGND.n88 VGND.n87 9.3005
R692 VGND.n413 VGND.n412 9.3005
R693 VGND.n410 VGND.n84 9.3005
R694 VGND.n409 VGND.n408 9.3005
R695 VGND.n407 VGND.n389 9.3005
R696 VGND.n406 VGND.n405 9.3005
R697 VGND.n404 VGND.n403 9.3005
R698 VGND.n402 VGND.n401 9.3005
R699 VGND.n400 VGND.n392 9.3005
R700 VGND.n126 VGND.n125 8.45078
R701 VGND.n566 VGND.n0 8.30267
R702 VGND.n128 VGND.n127 7.97888
R703 VGND.n126 VGND.n97 7.97601
R704 VGND.n306 VGND.n305 7.66295
R705 VGND.n177 VGND.n176 7.66295
R706 VGND.n470 VGND.n469 7.66295
R707 VGND.n51 VGND.n50 7.66295
R708 VGND.n374 VGND.n373 7.65909
R709 VGND.n245 VGND.n244 7.65909
R710 VGND.n546 VGND.n545 7.65909
R711 VGND.n397 VGND.n396 7.65909
R712 VGND.n241 VGND.n240 7.64725
R713 VGND.n504 VGND.n24 7.64725
R714 VGND.n551 VGND.n542 7.64725
R715 VGND.n411 VGND.n90 7.64725
R716 VGND.n391 VGND.n390 7.64725
R717 VGND.n129 VGND.n128 7.16724
R718 VGND.n125 VGND.n124 7.16724
R719 VGND.n105 VGND.n97 7.16724
R720 VGND.n566 VGND.n565 7.16724
R721 VGND.n401 VGND.n393 5.8885
R722 VGND.n51 VGND.n48 5.8885
R723 VGND.n51 VGND.n49 5.8885
R724 VGND.n396 VGND.n394 5.8885
R725 VGND.n396 VGND.n395 5.8885
R726 VGND.n373 VGND.n372 5.8885
R727 VGND.n305 VGND.n304 5.8885
R728 VGND.n177 VGND.n174 5.8885
R729 VGND.n177 VGND.n175 5.8885
R730 VGND.n244 VGND.n242 5.8885
R731 VGND.n244 VGND.n243 5.8885
R732 VGND.n469 VGND.n468 5.8885
R733 VGND.n545 VGND.n544 5.8885
R734 VGND.n133 VGND.n129 4.73093
R735 VGND.n124 VGND.n98 4.73093
R736 VGND.n107 VGND.n105 4.73093
R737 VGND.n565 VGND.n564 4.73093
R738 VGND.n356 VGND.n278 4.51401
R739 VGND.n361 VGND.n360 4.51401
R740 VGND.n322 VGND.n298 4.51401
R741 VGND.n326 VGND.n288 4.51401
R742 VGND.n273 VGND.n151 4.51401
R743 VGND.n266 VGND.n265 4.51401
R744 VGND.n199 VGND.n170 4.51401
R745 VGND.n204 VGND.n164 4.51401
R746 VGND.n455 VGND.n35 4.51401
R747 VGND.n40 VGND.n39 4.51401
R748 VGND.n528 VGND.n18 4.51401
R749 VGND.n533 VGND.n532 4.51401
R750 VGND.n488 VGND.n461 4.51401
R751 VGND.n492 VGND.n26 4.51401
R752 VGND.n77 VGND.n75 4.51401
R753 VGND.n415 VGND.n414 4.51401
R754 VGND.n144 VGND.n143 4.5005
R755 VGND.n355 VGND.n354 4.5005
R756 VGND.n352 VGND.n351 4.5005
R757 VGND.n321 VGND.n320 4.5005
R758 VGND.n319 VGND.n318 4.5005
R759 VGND.n328 VGND.n327 4.5005
R760 VGND.n264 VGND.n234 4.5005
R761 VGND.n272 VGND.n271 4.5005
R762 VGND.n261 VGND.n154 4.5005
R763 VGND.n198 VGND.n197 4.5005
R764 VGND.n196 VGND.n195 4.5005
R765 VGND.n206 VGND.n205 4.5005
R766 VGND.n14 VGND.n13 4.5005
R767 VGND.n527 VGND.n526 4.5005
R768 VGND.n524 VGND.n523 4.5005
R769 VGND.n487 VGND.n486 4.5005
R770 VGND.n485 VGND.n484 4.5005
R771 VGND.n494 VGND.n493 4.5005
R772 VGND.n86 VGND.n83 4.5005
R773 VGND.n454 VGND.n453 4.5005
R774 VGND.n452 VGND.n451 4.5005
R775 VGND.n448 VGND.n447 4.5005
R776 VGND.n422 VGND.n421 4.5005
R777 VGND.n85 VGND.n78 4.5005
R778 VGND.n520 VGND.n519 4.14168
R779 VGND.n146 VGND 4.01425
R780 VGND.n482 VGND.n481 3.76521
R781 VGND.n360 VGND.n359 3.43925
R782 VGND.n357 VGND.n356 3.43925
R783 VGND.n326 VGND.n325 3.43925
R784 VGND.n323 VGND.n322 3.43925
R785 VGND.n265 VGND.n149 3.43925
R786 VGND.n274 VGND.n273 3.43925
R787 VGND.n204 VGND.n203 3.43925
R788 VGND.n200 VGND.n199 3.43925
R789 VGND.n39 VGND.n33 3.43925
R790 VGND.n456 VGND.n455 3.43925
R791 VGND.n532 VGND.n531 3.43925
R792 VGND.n529 VGND.n528 3.43925
R793 VGND.n492 VGND.n491 3.43925
R794 VGND.n489 VGND.n488 3.43925
R795 VGND.n279 VGND.n277 3.4105
R796 VGND.n350 VGND.n145 3.4105
R797 VGND.n299 VGND.n297 3.4105
R798 VGND.n293 VGND.n292 3.4105
R799 VGND.n152 VGND.n150 3.4105
R800 VGND.n263 VGND.n262 3.4105
R801 VGND.n201 VGND.n169 3.4105
R802 VGND.n202 VGND.n168 3.4105
R803 VGND.n36 VGND.n34 3.4105
R804 VGND.n450 VGND.n449 3.4105
R805 VGND.n19 VGND.n17 3.4105
R806 VGND.n522 VGND.n15 3.4105
R807 VGND.n462 VGND.n460 3.4105
R808 VGND.n31 VGND.n30 3.4105
R809 VGND.n417 VGND.n416 3.4105
R810 VGND.n417 VGND.n79 3.4105
R811 VGND.n416 VGND.n415 3.4105
R812 VGND.n79 VGND.n77 3.4105
R813 VGND.n420 VGND.n419 3.4105
R814 VGND.n82 VGND.n80 3.4105
R815 VGND.n210 VGND.n163 3.38874
R816 VGND.n269 VGND.n232 3.38874
R817 VGND.t45 VGND.t8 2.97347
R818 VGND.n54 VGND.n53 2.25932
R819 VGND.n440 VGND.n439 2.25932
R820 VGND.n491 VGND.n490 1.69188
R821 VGND.n490 VGND.n489 1.69188
R822 VGND.n457 VGND.n33 1.69188
R823 VGND.n457 VGND.n456 1.69188
R824 VGND.n203 VGND.n32 1.69188
R825 VGND.n200 VGND.n32 1.69188
R826 VGND.n325 VGND.n324 1.69188
R827 VGND.n324 VGND.n323 1.69188
R828 VGND.n531 VGND.n530 1.69188
R829 VGND.n530 VGND.n529 1.69188
R830 VGND.n275 VGND.n149 1.69188
R831 VGND.n275 VGND.n274 1.69188
R832 VGND.n359 VGND.n358 1.69188
R833 VGND.n358 VGND.n357 1.69188
R834 VGND.n418 VGND.n417 1.69188
R835 VGND.n513 VGND.n512 1.50638
R836 VGND.n62 VGND.n44 1.50638
R837 VGND.n433 VGND.n432 1.50638
R838 VGND.n498 VGND.n497 1.12991
R839 VGND.n358 VGND.n148 0.867399
R840 VGND.n365 VGND.n138 0.753441
R841 VGND.n324 VGND.n148 0.659756
R842 VGND.n147 VGND.n146 0.595833
R843 VGND.n459 VGND.n458 0.500125
R844 VGND.n295 VGND.n294 0.500125
R845 VGND.n296 VGND 0.478236
R846 VGND.n127 VGND.n126 0.467019
R847 VGND.n294 VGND.n276 0.3805
R848 VGND.n458 VGND.n16 0.3805
R849 VGND.n183 VGND.n172 0.376971
R850 VGND.n146 VGND.n0 0.195328
R851 VGND.n530 VGND.n16 0.162755
R852 VGND.n457 VGND.n32 0.1603
R853 VGND.n490 VGND.n459 0.159712
R854 VGND.n375 VGND.n374 0.141672
R855 VGND.n246 VGND.n245 0.141672
R856 VGND.n547 VGND.n546 0.141672
R857 VGND.n398 VGND.n397 0.141672
R858 VGND.n307 VGND.n306 0.137814
R859 VGND.n176 VGND.n173 0.137814
R860 VGND.n471 VGND.n470 0.137814
R861 VGND.n50 VGND.n47 0.137814
R862 VGND.n148 VGND.n147 0.13699
R863 VGND.n358 VGND.n276 0.129226
R864 VGND.n374 VGND 0.121778
R865 VGND.n245 VGND 0.121778
R866 VGND.n546 VGND 0.121778
R867 VGND.n397 VGND 0.121778
R868 VGND.n296 VGND.n295 0.121084
R869 VGND.n308 VGND.n307 0.120292
R870 VGND.n312 VGND.n302 0.120292
R871 VGND.n313 VGND.n312 0.120292
R872 VGND.n314 VGND.n313 0.120292
R873 VGND.n333 VGND.n332 0.120292
R874 VGND.n334 VGND.n333 0.120292
R875 VGND.n338 VGND.n285 0.120292
R876 VGND.n339 VGND.n338 0.120292
R877 VGND.n340 VGND.n282 0.120292
R878 VGND.n344 VGND.n282 0.120292
R879 VGND.n346 VGND.n345 0.120292
R880 VGND.n367 VGND.n140 0.120292
R881 VGND.n368 VGND.n367 0.120292
R882 VGND.n381 VGND.n380 0.120292
R883 VGND.n380 VGND.n369 0.120292
R884 VGND.n181 VGND.n173 0.120292
R885 VGND.n188 VGND.n187 0.120292
R886 VGND.n189 VGND.n188 0.120292
R887 VGND.n213 VGND.n212 0.120292
R888 VGND.n214 VGND.n213 0.120292
R889 VGND.n219 VGND.n218 0.120292
R890 VGND.n224 VGND.n223 0.120292
R891 VGND.n229 VGND.n228 0.120292
R892 VGND.n256 VGND.n255 0.120292
R893 VGND.n251 VGND.n250 0.120292
R894 VGND.n250 VGND.n238 0.120292
R895 VGND.n472 VGND.n471 0.120292
R896 VGND.n477 VGND.n465 0.120292
R897 VGND.n478 VGND.n477 0.120292
R898 VGND.n479 VGND.n478 0.120292
R899 VGND.n500 VGND.n499 0.120292
R900 VGND.n501 VGND.n500 0.120292
R901 VGND.n506 VGND.n23 0.120292
R902 VGND.n507 VGND.n506 0.120292
R903 VGND.n508 VGND.n507 0.120292
R904 VGND.n514 VGND.n21 0.120292
R905 VGND.n515 VGND.n514 0.120292
R906 VGND.n516 VGND.n515 0.120292
R907 VGND.n539 VGND.n10 0.120292
R908 VGND.n540 VGND.n539 0.120292
R909 VGND.n553 VGND.n541 0.120292
R910 VGND.n548 VGND.n541 0.120292
R911 VGND.n548 VGND.n547 0.120292
R912 VGND.n55 VGND.n47 0.120292
R913 VGND.n57 VGND.n56 0.120292
R914 VGND.n443 VGND.n442 0.120292
R915 VGND.n437 VGND.n436 0.120292
R916 VGND.n436 VGND.n435 0.120292
R917 VGND.n435 VGND.n68 0.120292
R918 VGND.n429 VGND.n68 0.120292
R919 VGND.n429 VGND.n428 0.120292
R920 VGND.n428 VGND.n427 0.120292
R921 VGND.n427 VGND.n72 0.120292
R922 VGND.n413 VGND.n84 0.120292
R923 VGND.n408 VGND.n84 0.120292
R924 VGND.n408 VGND.n407 0.120292
R925 VGND.n402 VGND.n392 0.120292
R926 VGND.n398 VGND.n392 0.120292
R927 VGND.n458 VGND 0.107437
R928 VGND.n294 VGND 0.107437
R929 VGND VGND.n375 0.104667
R930 VGND VGND.n465 0.104667
R931 VGND.n217 VGND 0.10076
R932 VGND.n60 VGND 0.10076
R933 VGND.n376 VGND 0.0981562
R934 VGND.n182 VGND 0.0981562
R935 VGND.n218 VGND 0.0981562
R936 VGND.n222 VGND 0.0981562
R937 VGND VGND.n259 0.0981562
R938 VGND VGND.n251 0.0981562
R939 VGND.n246 VGND 0.0981562
R940 VGND VGND.n23 0.0981562
R941 VGND VGND.n553 0.0981562
R942 VGND.n56 VGND 0.0981562
R943 VGND.n61 VGND 0.0981562
R944 VGND VGND.n441 0.0981562
R945 VGND.n437 VGND 0.0981562
R946 VGND.n403 VGND 0.0981562
R947 VGND VGND.n402 0.0981562
R948 VGND.n346 VGND.n278 0.0968542
R949 VGND.n382 VGND 0.0968542
R950 VGND.n187 VGND 0.0968542
R951 VGND.n228 VGND 0.0968542
R952 VGND.n229 VGND.n151 0.0968542
R953 VGND.n516 VGND.n18 0.0968542
R954 VGND VGND.n285 0.0955521
R955 VGND.n340 VGND 0.0955521
R956 VGND.n345 VGND 0.0955521
R957 VGND.n356 VGND.n355 0.0950946
R958 VGND.n360 VGND.n144 0.0950946
R959 VGND.n322 VGND.n321 0.0950946
R960 VGND.n327 VGND.n326 0.0950946
R961 VGND.n273 VGND.n272 0.0950946
R962 VGND.n265 VGND.n264 0.0950946
R963 VGND.n199 VGND.n198 0.0950946
R964 VGND.n205 VGND.n204 0.0950946
R965 VGND.n455 VGND.n454 0.0950946
R966 VGND.n448 VGND.n39 0.0950946
R967 VGND.n528 VGND.n527 0.0950946
R968 VGND.n532 VGND.n14 0.0950946
R969 VGND.n488 VGND.n487 0.0950946
R970 VGND.n493 VGND.n492 0.0950946
R971 VGND.n421 VGND.n77 0.0950946
R972 VGND.n415 VGND.n83 0.0950946
R973 VGND.n332 VGND.n288 0.0916458
R974 VGND.n212 VGND.n164 0.0916458
R975 VGND.n499 VGND.n26 0.0916458
R976 VGND.n555 VGND 0.0916458
R977 VGND.n443 VGND.n40 0.0916458
R978 VGND VGND.n381 0.0864375
R979 VGND.n252 VGND 0.0864375
R980 VGND VGND.n554 0.0864375
R981 VGND VGND.n406 0.0864375
R982 VGND VGND.n302 0.0851354
R983 VGND.n223 VGND 0.0851354
R984 VGND.n256 VGND 0.0851354
R985 VGND.n352 VGND.n143 0.0838333
R986 VGND.n234 VGND.n154 0.0838333
R987 VGND.n486 VGND.n485 0.0838333
R988 VGND.n524 VGND.n13 0.0838333
R989 VGND.n453 VGND.n452 0.0838333
R990 VGND.n86 VGND.n85 0.0838333
R991 VGND.n275 VGND.n81 0.0819267
R992 VGND.n417 VGND.n81 0.0819267
R993 VGND.n306 VGND 0.0814556
R994 VGND.n176 VGND 0.0814556
R995 VGND.n470 VGND 0.0814556
R996 VGND.n50 VGND 0.0814556
R997 VGND VGND.n196 0.078625
R998 VGND.n127 VGND.n0 0.0766574
R999 VGND.n75 VGND 0.0747188
R1000 VGND.n362 VGND.n361 0.0708125
R1001 VGND.n267 VGND.n266 0.0708125
R1002 VGND.n534 VGND.n533 0.0708125
R1003 VGND.n351 VGND.n279 0.0680676
R1004 VGND.n351 VGND.n350 0.0680676
R1005 VGND.n318 VGND.n299 0.0680676
R1006 VGND.n318 VGND.n292 0.0680676
R1007 VGND.n261 VGND.n152 0.0680676
R1008 VGND.n263 VGND.n261 0.0680676
R1009 VGND.n195 VGND.n169 0.0680676
R1010 VGND.n195 VGND.n168 0.0680676
R1011 VGND.n451 VGND.n36 0.0680676
R1012 VGND.n451 VGND.n450 0.0680676
R1013 VGND.n523 VGND.n19 0.0680676
R1014 VGND.n523 VGND.n522 0.0680676
R1015 VGND.n484 VGND.n462 0.0680676
R1016 VGND.n484 VGND.n30 0.0680676
R1017 VGND.n420 VGND.n78 0.0680676
R1018 VGND.n82 VGND.n78 0.0680676
R1019 VGND VGND.n319 0.0669062
R1020 VGND.n317 VGND.n298 0.0656042
R1021 VGND.n328 VGND.n291 0.0656042
R1022 VGND.n194 VGND.n170 0.0656042
R1023 VGND.n206 VGND.n167 0.0656042
R1024 VGND.n483 VGND.n461 0.0656042
R1025 VGND.n494 VGND.n29 0.0656042
R1026 VGND.n37 VGND.n35 0.0656042
R1027 VGND.n128 VGND 0.064875
R1028 VGND.n97 VGND 0.064875
R1029 VGND VGND.n566 0.064875
R1030 VGND.n125 VGND 0.063625
R1031 VGND.n354 VGND.n353 0.0603958
R1032 VGND.n271 VGND.n153 0.0603958
R1033 VGND.n271 VGND.n270 0.0603958
R1034 VGND VGND.n21 0.0603958
R1035 VGND.n526 VGND.n521 0.0603958
R1036 VGND.n526 VGND.n525 0.0603958
R1037 VGND.n422 VGND.n76 0.0603958
R1038 VGND.n277 VGND.n145 0.0574697
R1039 VGND.n297 VGND.n293 0.0574697
R1040 VGND.n262 VGND.n150 0.0574697
R1041 VGND.n202 VGND.n201 0.0574697
R1042 VGND.n449 VGND.n34 0.0574697
R1043 VGND.n17 VGND.n15 0.0574697
R1044 VGND.n460 VGND.n31 0.0574697
R1045 VGND.n419 VGND.n79 0.0574697
R1046 VGND.n416 VGND.n80 0.0574697
R1047 VGND.n329 VGND.n328 0.0551875
R1048 VGND.n207 VGND.n206 0.0551875
R1049 VGND.n479 VGND.n461 0.0551875
R1050 VGND.n495 VGND.n494 0.0551875
R1051 VGND.n61 VGND.n35 0.0551875
R1052 VGND.n447 VGND.n446 0.0551875
R1053 VGND.n361 VGND.n140 0.0499792
R1054 VGND.n266 VGND.n260 0.0499792
R1055 VGND.n533 VGND.n10 0.0499792
R1056 VGND.n414 VGND.n413 0.0499792
R1057 VGND.n414 VGND 0.0486771
R1058 VGND.n447 VGND 0.0434688
R1059 VGND.n355 VGND.n279 0.0410405
R1060 VGND.n350 VGND.n144 0.0410405
R1061 VGND.n321 VGND.n299 0.0410405
R1062 VGND.n327 VGND.n292 0.0410405
R1063 VGND.n272 VGND.n152 0.0410405
R1064 VGND.n264 VGND.n263 0.0410405
R1065 VGND.n198 VGND.n169 0.0410405
R1066 VGND.n205 VGND.n168 0.0410405
R1067 VGND.n454 VGND.n36 0.0410405
R1068 VGND.n450 VGND.n448 0.0410405
R1069 VGND.n527 VGND.n19 0.0410405
R1070 VGND.n522 VGND.n14 0.0410405
R1071 VGND.n487 VGND.n462 0.0410405
R1072 VGND.n493 VGND.n30 0.0410405
R1073 VGND.n421 VGND.n420 0.0410405
R1074 VGND.n83 VGND.n82 0.0410405
R1075 VGND VGND.n170 0.0395625
R1076 VGND VGND.n422 0.0382604
R1077 VGND.n308 VGND 0.0356562
R1078 VGND.n354 VGND 0.0356562
R1079 VGND VGND.n222 0.0356562
R1080 VGND.n259 VGND 0.0356562
R1081 VGND.n276 VGND.n275 0.0346274
R1082 VGND.n382 VGND 0.0343542
R1083 VGND.n255 VGND 0.0343542
R1084 VGND.n555 VGND 0.0343542
R1085 VGND.n407 VGND 0.0343542
R1086 VGND.n295 VGND.n32 0.0339875
R1087 VGND VGND.n298 0.0330521
R1088 VGND.n489 VGND.n460 0.0292489
R1089 VGND.n491 VGND.n31 0.0292489
R1090 VGND.n456 VGND.n34 0.0292489
R1091 VGND.n449 VGND.n33 0.0292489
R1092 VGND.n201 VGND.n200 0.0292489
R1093 VGND.n203 VGND.n202 0.0292489
R1094 VGND.n323 VGND.n297 0.0292489
R1095 VGND.n325 VGND.n293 0.0292489
R1096 VGND.n529 VGND.n17 0.0292489
R1097 VGND.n531 VGND.n15 0.0292489
R1098 VGND.n274 VGND.n150 0.0292489
R1099 VGND.n262 VGND.n149 0.0292489
R1100 VGND.n357 VGND.n277 0.0292489
R1101 VGND.n359 VGND.n145 0.0292489
R1102 VGND.n418 VGND.n80 0.0292489
R1103 VGND.n419 VGND.n418 0.0292489
R1104 VGND.n495 VGND.n26 0.0291458
R1105 VGND VGND.n540 0.0291458
R1106 VGND.n446 VGND.n40 0.0291458
R1107 VGND.t27 VGND.n117 0.0282554
R1108 VGND.n329 VGND 0.0252396
R1109 VGND.n334 VGND 0.0252396
R1110 VGND VGND.n339 0.0252396
R1111 VGND VGND.n344 0.0252396
R1112 VGND VGND.n349 0.0252396
R1113 VGND.n349 VGND.n278 0.0239375
R1114 VGND.n353 VGND.n352 0.0239375
R1115 VGND VGND.n368 0.0239375
R1116 VGND.n182 VGND 0.0239375
R1117 VGND.n224 VGND 0.0239375
R1118 VGND.n153 VGND.n151 0.0239375
R1119 VGND.n270 VGND.n154 0.0239375
R1120 VGND.n521 VGND.n18 0.0239375
R1121 VGND.n525 VGND.n524 0.0239375
R1122 VGND.n423 VGND.n75 0.0239375
R1123 VGND.n85 VGND.n76 0.0239375
R1124 VGND.n314 VGND 0.0226354
R1125 VGND VGND.n369 0.0226354
R1126 VGND VGND.n217 0.0226354
R1127 VGND.n219 VGND 0.0226354
R1128 VGND.n260 VGND 0.0226354
R1129 VGND.n252 VGND 0.0226354
R1130 VGND VGND.n238 0.0226354
R1131 VGND.n501 VGND 0.0226354
R1132 VGND.n554 VGND 0.0226354
R1133 VGND VGND.n55 0.0226354
R1134 VGND VGND.n60 0.0226354
R1135 VGND VGND.n38 0.0226354
R1136 VGND.n441 VGND 0.0226354
R1137 VGND VGND.n72 0.0226354
R1138 VGND.n423 VGND 0.0226354
R1139 VGND.n87 VGND 0.0226354
R1140 VGND.n406 VGND 0.0226354
R1141 VGND.n403 VGND 0.0226354
R1142 VGND.n147 VGND 0.0223384
R1143 VGND.n207 VGND 0.0200312
R1144 VGND.n214 VGND 0.0200312
R1145 VGND.n57 VGND 0.0200312
R1146 VGND.n320 VGND.n317 0.0187292
R1147 VGND.n319 VGND.n291 0.0187292
R1148 VGND.n197 VGND.n194 0.0187292
R1149 VGND.n196 VGND.n167 0.0187292
R1150 VGND.n486 VGND.n483 0.0187292
R1151 VGND.n485 VGND.n29 0.0187292
R1152 VGND.n453 VGND.n37 0.0187292
R1153 VGND.n452 VGND.n38 0.0187292
R1154 VGND.n320 VGND 0.0174271
R1155 VGND.n376 VGND 0.016125
R1156 VGND VGND.n181 0.016125
R1157 VGND.n189 VGND 0.016125
R1158 VGND.n472 VGND 0.016125
R1159 VGND.n508 VGND 0.016125
R1160 VGND.n442 VGND 0.016125
R1161 VGND.n362 VGND.n143 0.0135208
R1162 VGND.n267 VGND.n234 0.0135208
R1163 VGND.n534 VGND.n13 0.0135208
R1164 VGND.n87 VGND.n86 0.0135208
R1165 VGND VGND.n164 0.00961458
R1166 VGND.n530 VGND 0.00768471
R1167 VGND.n490 VGND 0.00755
R1168 VGND.n324 VGND.n296 0.00619255
R1169 VGND.n197 VGND 0.00570833
R1170 VGND VGND.n288 0.00440625
R1171 VGND.n417 VGND.n16 0.00109873
R1172 VGND.n459 VGND.n457 0.0010875
R1173 VPWR.n488 VPWR.n487 8629.41
R1174 VPWR.n490 VPWR.n484 8629.41
R1175 VPWR.n506 VPWR.n500 8629.41
R1176 VPWR.n509 VPWR.n499 8629.41
R1177 VPWR.n523 VPWR.n517 8629.41
R1178 VPWR.n526 VPWR.n516 8629.41
R1179 VPWR.n537 VPWR.n535 8629.41
R1180 VPWR.n540 VPWR.n534 8629.41
R1181 VPWR.n491 VPWR.n483 920.471
R1182 VPWR.n505 VPWR.n501 920.471
R1183 VPWR.n522 VPWR.n518 920.471
R1184 VPWR.n536 VPWR.n533 920.471
R1185 VPWR.n492 VPWR.n491 914.447
R1186 VPWR.n501 VPWR.n497 914.447
R1187 VPWR.n518 VPWR.n514 914.447
R1188 VPWR.n542 VPWR.n533 914.447
R1189 VPWR.n53 VPWR.t45 804.731
R1190 VPWR.n57 VPWR.t30 804.731
R1191 VPWR.n120 VPWR.t18 804.731
R1192 VPWR.n123 VPWR.t54 804.731
R1193 VPWR.n280 VPWR.t47 804.731
R1194 VPWR.n276 VPWR.t15 804.731
R1195 VPWR.n14 VPWR.t35 804.731
R1196 VPWR.n243 VPWR.t34 804.731
R1197 VPWR.n204 VPWR.t33 804.731
R1198 VPWR.n209 VPWR.t62 804.731
R1199 VPWR.n287 VPWR.t58 804.731
R1200 VPWR.n290 VPWR.t40 804.731
R1201 VPWR.n431 VPWR.t24 804.731
R1202 VPWR.n395 VPWR.t23 804.731
R1203 VPWR.n345 VPWR.t66 804.731
R1204 VPWR.n348 VPWR.t38 804.731
R1205 VPWR.n320 VPWR.t49 804.731
R1206 VPWR.n456 VPWR.t21 804.731
R1207 VPWR.n459 VPWR.t43 804.731
R1208 VPWR.n462 VPWR.t60 804.731
R1209 VPWR.t15 VPWR.n275 751.692
R1210 VPWR.t49 VPWR.n319 751.692
R1211 VPWR.t21 VPWR.n455 751.692
R1212 VPWR.t45 VPWR.n52 725.173
R1213 VPWR.t30 VPWR.n56 725.173
R1214 VPWR.t18 VPWR.n119 725.173
R1215 VPWR.t54 VPWR.n122 725.173
R1216 VPWR.t47 VPWR.n279 725.173
R1217 VPWR.t33 VPWR.n203 725.173
R1218 VPWR.t62 VPWR.n208 725.173
R1219 VPWR.t58 VPWR.n286 725.173
R1220 VPWR.t40 VPWR.n289 725.173
R1221 VPWR.t66 VPWR.n344 725.173
R1222 VPWR.t38 VPWR.n347 725.173
R1223 VPWR.t43 VPWR.n458 725.173
R1224 VPWR.t60 VPWR.n461 725.173
R1225 VPWR.n63 VPWR.t102 701.529
R1226 VPWR VPWR.t106 697.264
R1227 VPWR.n96 VPWR.t90 671.408
R1228 VPWR.n370 VPWR.n342 599.159
R1229 VPWR.n341 VPWR.n340 594.144
R1230 VPWR.n430 VPWR.n327 594.144
R1231 VPWR.n423 VPWR.n330 594.144
R1232 VPWR.n437 VPWR.n324 594.144
R1233 VPWR.n33 VPWR.n32 590.973
R1234 VPWR.n247 VPWR.n246 585
R1235 VPWR.n249 VPWR.n248 585
R1236 VPWR.n379 VPWR.n378 585
R1237 VPWR.n377 VPWR.n376 585
R1238 VPWR.n381 VPWR.n380 585
R1239 VPWR.n389 VPWR.n388 585
R1240 VPWR.t19 VPWR.t41 540.46
R1241 VPWR.n485 VPWR.n483 480.764
R1242 VPWR.n505 VPWR.n504 480.764
R1243 VPWR.n522 VPWR.n521 480.764
R1244 VPWR.n536 VPWR.n531 480.764
R1245 VPWR VPWR.t50 394.435
R1246 VPWR.n10 VPWR.t63 393.002
R1247 VPWR.n284 VPWR.t64 388.656
R1248 VPWR.n325 VPWR.t26 388.656
R1249 VPWR.n440 VPWR.t27 388.656
R1250 VPWR.n225 VPWR.t55 388.656
R1251 VPWR.n232 VPWR.t56 388.656
R1252 VPWR.n268 VPWR.t14 388.656
R1253 VPWR.n396 VPWR.t51 388.656
R1254 VPWR.n407 VPWR.t52 388.656
R1255 VPWR.n318 VPWR.t48 387.682
R1256 VPWR.n454 VPWR.t20 387.682
R1257 VPWR.n51 VPWR.t44 380.193
R1258 VPWR.n55 VPWR.t29 380.193
R1259 VPWR.n118 VPWR.t17 380.193
R1260 VPWR.n121 VPWR.t53 380.193
R1261 VPWR.n278 VPWR.t46 380.193
R1262 VPWR.n202 VPWR.t32 380.193
R1263 VPWR.n207 VPWR.t61 380.193
R1264 VPWR.n285 VPWR.t57 380.193
R1265 VPWR.n288 VPWR.t39 380.193
R1266 VPWR.n343 VPWR.t65 380.193
R1267 VPWR.n346 VPWR.t37 380.193
R1268 VPWR.n457 VPWR.t42 380.193
R1269 VPWR.n460 VPWR.t59 380.193
R1270 VPWR.n485 VPWR.n482 379.2
R1271 VPWR.n504 VPWR.n503 379.2
R1272 VPWR.n521 VPWR.n520 379.2
R1273 VPWR.n544 VPWR.n531 379.2
R1274 VPWR VPWR.t28 335.69
R1275 VPWR VPWR.t36 328.976
R1276 VPWR.n137 VPWR.n98 322.329
R1277 VPWR.n165 VPWR.n68 317.104
R1278 VPWR.n146 VPWR.n95 316.515
R1279 VPWR.t129 VPWR.t93 315.548
R1280 VPWR.n78 VPWR.n77 312.053
R1281 VPWR.n117 VPWR.n116 312.053
R1282 VPWR.n41 VPWR.n40 312.053
R1283 VPWR.n166 VPWR.n65 312.051
R1284 VPWR.n70 VPWR.n69 312.051
R1285 VPWR.n89 VPWR.n80 312.051
R1286 VPWR.n151 VPWR.n90 312.051
R1287 VPWR.n146 VPWR.n94 312.051
R1288 VPWR.n107 VPWR.n106 312.051
R1289 VPWR.n237 VPWR.n36 312.051
R1290 VPWR.n390 VPWR.n387 312.051
R1291 VPWR.n174 VPWR.n61 312.005
R1292 VPWR.n16 VPWR.t180 310.853
R1293 VPWR.n263 VPWR.n18 308.755
R1294 VPWR.n173 VPWR.n62 308.755
R1295 VPWR.n231 VPWR.n38 308.755
R1296 VPWR.n424 VPWR.t185 306.735
R1297 VPWR.n9 VPWR.t103 293.159
R1298 VPWR.t173 VPWR.t7 281.979
R1299 VPWR VPWR.t16 280.3
R1300 VPWR.n9 VPWR.n8 269.485
R1301 VPWR VPWR.t124 263.517
R1302 VPWR VPWR.t91 263.517
R1303 VPWR VPWR.t101 256.803
R1304 VPWR.n52 VPWR.t193 245.667
R1305 VPWR.n56 VPWR.t189 245.667
R1306 VPWR.n119 VPWR.t181 245.667
R1307 VPWR.n122 VPWR.t177 245.667
R1308 VPWR.n279 VPWR.t196 245.667
R1309 VPWR.n203 VPWR.t182 245.667
R1310 VPWR.n208 VPWR.t188 245.667
R1311 VPWR.n286 VPWR.t194 245.667
R1312 VPWR.n289 VPWR.t176 245.667
R1313 VPWR.n344 VPWR.t190 245.667
R1314 VPWR.n347 VPWR.t195 245.667
R1315 VPWR.n458 VPWR.t178 245.667
R1316 VPWR.n461 VPWR.t183 245.667
R1317 VPWR.n144 VPWR.t123 245.178
R1318 VPWR.n138 VPWR.t115 243.508
R1319 VPWR.n224 VPWR.t160 240.939
R1320 VPWR VPWR.t116 240.018
R1321 VPWR.t81 VPWR.t143 234.982
R1322 VPWR.n319 VPWR.t197 213.148
R1323 VPWR.n455 VPWR.t179 213.148
R1324 VPWR.n281 VPWR.t191 210.964
R1325 VPWR.n406 VPWR.t187 210.964
R1326 VPWR.n439 VPWR.t184 210.964
R1327 VPWR.n136 VPWR.t81 209.368
R1328 VPWR.t50 VPWR 203.093
R1329 VPWR VPWR.t19 203.093
R1330 VPWR.t16 VPWR 182.952
R1331 VPWR.n316 VPWR 182.952
R1332 VPWR.t41 VPWR 182.952
R1333 VPWR VPWR.t135 176.238
R1334 VPWR.t170 VPWR.t67 174.559
R1335 VPWR.n248 VPWR.n247 159.476
R1336 VPWR.n378 VPWR.n377 159.476
R1337 VPWR.t93 VPWR.t168 159.452
R1338 VPWR.t116 VPWR.t129 159.452
R1339 VPWR.t168 VPWR.t22 157.774
R1340 VPWR.t156 VPWR.t3 154.417
R1341 VPWR.t145 VPWR.t97 151.06
R1342 VPWR.t79 VPWR.t9 147.703
R1343 VPWR.t5 VPWR.t69 147.703
R1344 VPWR.t67 VPWR.t71 147.703
R1345 VPWR.t143 VPWR.t73 147.703
R1346 VPWR.t118 VPWR.t133 144.346
R1347 VPWR.t75 VPWR.t137 142.668
R1348 VPWR.t131 VPWR.t95 142.668
R1349 VPWR.t149 VPWR 135.954
R1350 VPWR.n34 VPWR.n33 132.268
R1351 VPWR.n233 VPWR.t192 129.344
R1352 VPWR.t28 VPWR 125.883
R1353 VPWR.t36 VPWR 125.883
R1354 VPWR.t81 VPWR 124.206
R1355 VPWR.t107 VPWR 120.849
R1356 VPWR.t166 VPWR.t107 120.849
R1357 VPWR.t108 VPWR.t86 120.849
R1358 VPWR VPWR.t75 120.849
R1359 VPWR.t120 VPWR.t166 119.171
R1360 VPWR.n275 VPWR.t186 118.853
R1361 VPWR.n316 VPWR 117.492
R1362 VPWR.n98 VPWR.t113 116.341
R1363 VPWR VPWR.t145 112.457
R1364 VPWR VPWR.t164 109.1
R1365 VPWR VPWR.t5 109.1
R1366 VPWR VPWR.t156 109.1
R1367 VPWR.n317 VPWR.n316 106.561
R1368 VPWR.t152 VPWR.t161 105.743
R1369 VPWR.t164 VPWR.t11 104.064
R1370 VPWR.t77 VPWR 102.385
R1371 VPWR VPWR.t147 100.707
R1372 VPWR.n68 VPWR.t109 98.5005
R1373 VPWR.n95 VPWR.t88 98.5005
R1374 VPWR.n61 VPWR.t167 96.1553
R1375 VPWR.n32 VPWR.t175 96.1553
R1376 VPWR.n342 VPWR.t153 96.1553
R1377 VPWR.t7 VPWR.t141 93.9934
R1378 VPWR.t135 VPWR.t25 92.315
R1379 VPWR VPWR.t170 88.9581
R1380 VPWR.t139 VPWR 88.9581
R1381 VPWR.n248 VPWR.t105 86.7743
R1382 VPWR.n377 VPWR.t8 86.7743
R1383 VPWR.t114 VPWR.t89 80.5659
R1384 VPWR.n388 VPWR.t132 77.3934
R1385 VPWR.n380 VPWR.t174 77.3934
R1386 VPWR.n340 VPWR.t162 77.3934
R1387 VPWR.n327 VPWR.t117 77.3934
R1388 VPWR.n330 VPWR.t94 77.3934
R1389 VPWR.n324 VPWR.t136 77.3934
R1390 VPWR.n10 VPWR.n9 72.8099
R1391 VPWR.t22 VPWR 68.8168
R1392 VPWR.t25 VPWR.t149 67.1383
R1393 VPWR.n247 VPWR.t128 66.8398
R1394 VPWR.n378 VPWR.t138 66.8398
R1395 VPWR.n493 VPWR.n492 66.6358
R1396 VPWR.n498 VPWR.n497 66.6358
R1397 VPWR.n515 VPWR.n514 66.6358
R1398 VPWR.n543 VPWR.n542 66.6358
R1399 VPWR.n32 VPWR.t155 63.3219
R1400 VPWR.n342 VPWR.t111 63.3219
R1401 VPWR.n488 VPWR.n483 61.6672
R1402 VPWR.n484 VPWR.n480 61.6672
R1403 VPWR.n506 VPWR.n505 61.6672
R1404 VPWR.n510 VPWR.n509 61.6672
R1405 VPWR.n523 VPWR.n522 61.6672
R1406 VPWR.n527 VPWR.n526 61.6672
R1407 VPWR.n537 VPWR.n536 61.6672
R1408 VPWR.n541 VPWR.n540 61.6672
R1409 VPWR.n489 VPWR.n488 60.9564
R1410 VPWR.n486 VPWR.n484 60.9564
R1411 VPWR.n507 VPWR.n506 60.9564
R1412 VPWR.n509 VPWR.n508 60.9564
R1413 VPWR.n524 VPWR.n523 60.9564
R1414 VPWR.n526 VPWR.n525 60.9564
R1415 VPWR.n538 VPWR.n537 60.9564
R1416 VPWR.n540 VPWR.n539 60.9564
R1417 VPWR.n510 VPWR.n498 60.6123
R1418 VPWR.n527 VPWR.n515 60.6123
R1419 VPWR.t89 VPWR.t122 60.4245
R1420 VPWR.t112 VPWR.t114 60.4245
R1421 VPWR.n494 VPWR.n493 59.4829
R1422 VPWR.t161 VPWR.t110 58.7461
R1423 VPWR.n543 VPWR.n532 58.7299
R1424 VPWR VPWR.t112 57.0676
R1425 VPWR.t141 VPWR.t152 53.7107
R1426 VPWR.t83 VPWR 52.0323
R1427 VPWR.t9 VPWR 52.0323
R1428 VPWR.t147 VPWR 52.0323
R1429 VPWR.t122 VPWR 52.0323
R1430 VPWR.t110 VPWR 52.0323
R1431 VPWR.t95 VPWR 52.0323
R1432 VPWR.t101 VPWR 50.3539
R1433 VPWR.t71 VPWR 50.3539
R1434 VPWR.t124 VPWR 46.997
R1435 VPWR VPWR.t139 45.3185
R1436 VPWR.t11 VPWR.t120 43.6401
R1437 VPWR.n388 VPWR.t157 41.0422
R1438 VPWR.n380 VPWR.t76 41.0422
R1439 VPWR.n340 VPWR.t142 41.0422
R1440 VPWR.n327 VPWR.t130 41.0422
R1441 VPWR.n330 VPWR.t169 41.0422
R1442 VPWR.n324 VPWR.t150 41.0422
R1443 VPWR.n490 VPWR.n489 38.5759
R1444 VPWR.n487 VPWR.n486 38.5759
R1445 VPWR.n507 VPWR.n499 38.5759
R1446 VPWR.n508 VPWR.n500 38.5759
R1447 VPWR.n524 VPWR.n516 38.5759
R1448 VPWR.n525 VPWR.n517 38.5759
R1449 VPWR.n538 VPWR.n534 38.5759
R1450 VPWR.n539 VPWR.n535 38.5759
R1451 VPWR.n62 VPWR.t121 36.1587
R1452 VPWR.n62 VPWR.t165 36.1587
R1453 VPWR.n65 VPWR.t84 36.1587
R1454 VPWR.n65 VPWR.t98 36.1587
R1455 VPWR.n69 VPWR.t10 36.1587
R1456 VPWR.n69 VPWR.t80 36.1587
R1457 VPWR.n77 VPWR.t70 36.1587
R1458 VPWR.n77 VPWR.t6 36.1587
R1459 VPWR.n80 VPWR.t148 36.1587
R1460 VPWR.n80 VPWR.t125 36.1587
R1461 VPWR.n90 VPWR.t72 36.1587
R1462 VPWR.n90 VPWR.t68 36.1587
R1463 VPWR.n94 VPWR.t134 36.1587
R1464 VPWR.n94 VPWR.t92 36.1587
R1465 VPWR.n106 VPWR.t144 36.1587
R1466 VPWR.n106 VPWR.t74 36.1587
R1467 VPWR.n116 VPWR.t78 36.1587
R1468 VPWR.n116 VPWR.t140 36.1587
R1469 VPWR.n18 VPWR.t1 36.1587
R1470 VPWR.n18 VPWR.t2 36.1587
R1471 VPWR.n38 VPWR.t100 36.1587
R1472 VPWR.n38 VPWR.t158 36.1587
R1473 VPWR.n40 VPWR.t154 36.1587
R1474 VPWR.n40 VPWR.t126 36.1587
R1475 VPWR.n36 VPWR.t159 36.1587
R1476 VPWR.n36 VPWR.t151 36.1587
R1477 VPWR.n387 VPWR.t96 36.1587
R1478 VPWR.n387 VPWR.t4 36.1587
R1479 VPWR.n173 VPWR.n172 34.6358
R1480 VPWR.n185 VPWR.n58 34.6358
R1481 VPWR.n175 VPWR.n58 34.6358
R1482 VPWR.n168 VPWR.n167 34.6358
R1483 VPWR.n150 VPWR.n92 34.6358
R1484 VPWR.n140 VPWR.n139 34.6358
R1485 VPWR.n136 VPWR.n99 34.6358
R1486 VPWR.n370 VPWR.n369 33.8829
R1487 VPWR.n145 VPWR.n144 33.5064
R1488 VPWR.t87 VPWR 31.891
R1489 VPWR.n8 VPWR 31.4055
R1490 VPWR.n98 VPWR.t82 28.4453
R1491 VPWR.n375 VPWR.n374 27.724
R1492 VPWR.n386 VPWR.n338 27.1064
R1493 VPWR.n168 VPWR.n63 25.977
R1494 VPWR.n61 VPWR.t12 25.6105
R1495 VPWR.n68 VPWR.t146 25.6105
R1496 VPWR.n95 VPWR.t119 25.6105
R1497 VPWR.n165 VPWR.n164 25.224
R1498 VPWR.n172 VPWR.n63 24.0946
R1499 VPWR.n153 VPWR.n152 24.0946
R1500 VPWR.n186 VPWR.n185 23.7181
R1501 VPWR.n126 VPWR.n125 23.7181
R1502 VPWR.n211 VPWR.n210 23.7181
R1503 VPWR.n369 VPWR.n349 23.7181
R1504 VPWR.n174 VPWR.n173 22.5887
R1505 VPWR.n167 VPWR.n166 22.2123
R1506 VPWR.n164 VPWR.n70 22.2123
R1507 VPWR.n79 VPWR.n78 22.2123
R1508 VPWR.n89 VPWR.n79 22.2123
R1509 VPWR.n153 VPWR.n89 22.2123
R1510 VPWR.n151 VPWR.n150 22.2123
R1511 VPWR.n146 VPWR.n92 22.2123
R1512 VPWR.n146 VPWR.n145 22.2123
R1513 VPWR.n107 VPWR.n99 22.2123
R1514 VPWR.n126 VPWR.n117 22.2123
R1515 VPWR.n210 VPWR.n41 22.2123
R1516 VPWR.n223 VPWR.n41 22.2123
R1517 VPWR.n238 VPWR.n237 22.2123
R1518 VPWR.n390 VPWR.n386 22.2123
R1519 VPWR.n238 VPWR.n34 21.4593
R1520 VPWR.n224 VPWR.n223 21.2076
R1521 VPWR VPWR.t104 20.1894
R1522 VPWR.t133 VPWR.t87 20.1418
R1523 VPWR.n140 VPWR.n96 19.9534
R1524 VPWR.n374 VPWR.n341 19.9534
R1525 VPWR.n138 VPWR.n137 18.4476
R1526 VPWR.n433 VPWR.n432 17.612
R1527 VPWR.n394 VPWR.n337 17.3741
R1528 VPWR.t137 VPWR.t173 16.785
R1529 VPWR.n137 VPWR.n136 15.8123
R1530 VPWR.n382 VPWR.n381 14.8543
R1531 VPWR.n143 VPWR.n96 14.6829
R1532 VPWR.n371 VPWR.n341 14.6829
R1533 VPWR.n292 VPWR.n291 14.2735
R1534 VPWR.n441 VPWR.n317 14.2735
R1535 VPWR.n152 VPWR.n151 13.5534
R1536 VPWR.t86 VPWR.t83 13.4281
R1537 VPWR.t97 VPWR.t108 13.4281
R1538 VPWR.n464 VPWR.n317 12.8005
R1539 VPWR.n464 VPWR.n463 12.8005
R1540 VPWR.n237 VPWR.n35 12.7676
R1541 VPWR.n175 VPWR.n174 12.0476
R1542 VPWR.n482 VPWR.n481 11.3235
R1543 VPWR.n503 VPWR.n502 11.3235
R1544 VPWR.n520 VPWR.n519 11.3235
R1545 VPWR.n545 VPWR.n544 11.3235
R1546 VPWR.n390 VPWR.n389 10.5955
R1547 VPWR.n166 VPWR.n165 10.5417
R1548 VPWR.t104 VPWR.t0 10.3754
R1549 VPWR.n78 VPWR.n70 9.78874
R1550 VPWR.n117 VPWR.n107 9.78874
R1551 VPWR.n262 VPWR.n19 9.73273
R1552 VPWR.n263 VPWR.n262 9.73273
R1553 VPWR.n264 VPWR.n263 9.73273
R1554 VPWR.n421 VPWR.n331 9.73273
R1555 VPWR.n422 VPWR.n421 9.73273
R1556 VPWR.n425 VPWR.n328 9.73273
R1557 VPWR.n429 VPWR.n328 9.73273
R1558 VPWR.n242 VPWR.n33 9.6005
R1559 VPWR.n186 VPWR 9.32264
R1560 VPWR.n211 VPWR 9.32264
R1561 VPWR VPWR.n349 9.32264
R1562 VPWR.n187 VPWR.n186 9.3005
R1563 VPWR.n186 VPWR.n54 9.3005
R1564 VPWR.n185 VPWR.n184 9.3005
R1565 VPWR.n177 VPWR.n58 9.3005
R1566 VPWR.n176 VPWR.n175 9.3005
R1567 VPWR.n173 VPWR.n60 9.3005
R1568 VPWR.n172 VPWR.n171 9.3005
R1569 VPWR.n170 VPWR.n63 9.3005
R1570 VPWR.n169 VPWR.n168 9.3005
R1571 VPWR.n167 VPWR.n64 9.3005
R1572 VPWR.n166 VPWR.n66 9.3005
R1573 VPWR.n165 VPWR.n67 9.3005
R1574 VPWR.n164 VPWR.n163 9.3005
R1575 VPWR.n162 VPWR.n70 9.3005
R1576 VPWR.n78 VPWR.n71 9.3005
R1577 VPWR.n82 VPWR.n79 9.3005
R1578 VPWR.n89 VPWR.n88 9.3005
R1579 VPWR.n154 VPWR.n153 9.3005
R1580 VPWR.n152 VPWR.n76 9.3005
R1581 VPWR.n151 VPWR.n91 9.3005
R1582 VPWR.n150 VPWR.n149 9.3005
R1583 VPWR.n148 VPWR.n92 9.3005
R1584 VPWR.n147 VPWR.n146 9.3005
R1585 VPWR.n145 VPWR.n93 9.3005
R1586 VPWR.n143 VPWR.n142 9.3005
R1587 VPWR.n141 VPWR.n140 9.3005
R1588 VPWR.n139 VPWR.n97 9.3005
R1589 VPWR.n136 VPWR.n135 9.3005
R1590 VPWR.n100 VPWR.n99 9.3005
R1591 VPWR.n109 VPWR.n107 9.3005
R1592 VPWR.n117 VPWR.n115 9.3005
R1593 VPWR.n127 VPWR.n126 9.3005
R1594 VPWR.n212 VPWR.n211 9.3005
R1595 VPWR.n211 VPWR.n206 9.3005
R1596 VPWR.n210 VPWR.n42 9.3005
R1597 VPWR.n221 VPWR.n41 9.3005
R1598 VPWR.n223 VPWR.n222 9.3005
R1599 VPWR.n227 VPWR.n226 9.3005
R1600 VPWR.n228 VPWR.n39 9.3005
R1601 VPWR.n230 VPWR.n229 9.3005
R1602 VPWR.n231 VPWR.n37 9.3005
R1603 VPWR.n234 VPWR.n233 9.3005
R1604 VPWR.n235 VPWR.n35 9.3005
R1605 VPWR.n237 VPWR.n236 9.3005
R1606 VPWR.n239 VPWR.n238 9.3005
R1607 VPWR.n241 VPWR.n240 9.3005
R1608 VPWR.n244 VPWR.n27 9.3005
R1609 VPWR.n251 VPWR.n250 9.3005
R1610 VPWR.n245 VPWR.n20 9.3005
R1611 VPWR.n260 VPWR.n19 9.3005
R1612 VPWR.n262 VPWR.n261 9.3005
R1613 VPWR.n263 VPWR.n17 9.3005
R1614 VPWR.n265 VPWR.n264 9.3005
R1615 VPWR.n267 VPWR.n266 9.3005
R1616 VPWR.n269 VPWR.n15 9.3005
R1617 VPWR.n271 VPWR.n270 9.3005
R1618 VPWR.n273 VPWR.n272 9.3005
R1619 VPWR.n277 VPWR.n13 9.3005
R1620 VPWR.n277 VPWR.n11 9.3005
R1621 VPWR.n304 VPWR.n303 9.3005
R1622 VPWR.n302 VPWR.n301 9.3005
R1623 VPWR.n293 VPWR.n292 9.3005
R1624 VPWR.n359 VPWR.n349 9.3005
R1625 VPWR.n360 VPWR.n349 9.3005
R1626 VPWR.n369 VPWR.n368 9.3005
R1627 VPWR.n372 VPWR.n371 9.3005
R1628 VPWR.n374 VPWR.n373 9.3005
R1629 VPWR.n375 VPWR.n339 9.3005
R1630 VPWR.n383 VPWR.n382 9.3005
R1631 VPWR.n384 VPWR.n338 9.3005
R1632 VPWR.n386 VPWR.n385 9.3005
R1633 VPWR.n391 VPWR.n390 9.3005
R1634 VPWR.n392 VPWR.n337 9.3005
R1635 VPWR.n394 VPWR.n393 9.3005
R1636 VPWR.n398 VPWR.n397 9.3005
R1637 VPWR.n399 VPWR.n336 9.3005
R1638 VPWR.n405 VPWR.n404 9.3005
R1639 VPWR.n409 VPWR.n408 9.3005
R1640 VPWR.n410 VPWR.n331 9.3005
R1641 VPWR.n421 VPWR.n420 9.3005
R1642 VPWR.n422 VPWR.n329 9.3005
R1643 VPWR.n426 VPWR.n425 9.3005
R1644 VPWR.n427 VPWR.n328 9.3005
R1645 VPWR.n429 VPWR.n428 9.3005
R1646 VPWR.n432 VPWR.n326 9.3005
R1647 VPWR.n434 VPWR.n433 9.3005
R1648 VPWR.n436 VPWR.n435 9.3005
R1649 VPWR.n438 VPWR.n323 9.3005
R1650 VPWR.n442 VPWR.n441 9.3005
R1651 VPWR.n443 VPWR.n317 9.3005
R1652 VPWR.n464 VPWR.n453 9.3005
R1653 VPWR.n464 VPWR.n322 9.3005
R1654 VPWR.n464 VPWR.n321 9.3005
R1655 VPWR.n465 VPWR.n464 9.3005
R1656 VPWR.n244 VPWR.n243 9.09802
R1657 VPWR.n245 VPWR.n19 8.80773
R1658 VPWR.n250 VPWR.n244 8.57648
R1659 VPWR.n532 VPWR.n530 8.23557
R1660 VPWR.n431 VPWR.n430 7.93438
R1661 VPWR.n408 VPWR.n331 7.75995
R1662 VPWR.n397 VPWR.n395 7.12524
R1663 VPWR.n379 VPWR.n376 6.8005
R1664 VPWR.t69 VPWR.t79 6.71428
R1665 VPWR.t73 VPWR.t77 6.71428
R1666 VPWR.n492 VPWR.n480 6.02403
R1667 VPWR.n542 VPWR.n541 6.02403
R1668 VPWR.n8 VPWR.t99 5.88893
R1669 VPWR.n425 VPWR.n424 5.18397
R1670 VPWR.t3 VPWR.t131 5.03584
R1671 VPWR.n511 VPWR.n510 4.89462
R1672 VPWR.n528 VPWR.n514 4.89462
R1673 VPWR.n230 VPWR.n39 4.67352
R1674 VPWR.n231 VPWR.n230 4.67352
R1675 VPWR.n233 VPWR.n231 4.67352
R1676 VPWR.n303 VPWR.n302 4.67352
R1677 VPWR.n277 VPWR.n12 4.62124
R1678 VPWR.n161 VPWR.n160 4.51401
R1679 VPWR.n156 VPWR.n155 4.51401
R1680 VPWR.n134 VPWR.n133 4.51401
R1681 VPWR.n129 VPWR.n128 4.51401
R1682 VPWR.n190 VPWR.n48 4.51401
R1683 VPWR.n183 VPWR.n182 4.51401
R1684 VPWR.n254 VPWR.n25 4.51401
R1685 VPWR.n259 VPWR.n258 4.51401
R1686 VPWR.n307 VPWR.n6 4.51401
R1687 VPWR.n298 VPWR.n294 4.51401
R1688 VPWR.n215 VPWR.n197 4.51401
R1689 VPWR.n220 VPWR.n219 4.51401
R1690 VPWR.n356 VPWR.n354 4.51401
R1691 VPWR.n367 VPWR.n366 4.51401
R1692 VPWR.n445 VPWR.n444 4.51401
R1693 VPWR.n467 VPWR.n466 4.51401
R1694 VPWR.n403 VPWR.n402 4.51401
R1695 VPWR.n81 VPWR.n72 4.5005
R1696 VPWR.n86 VPWR.n85 4.5005
R1697 VPWR.n87 VPWR.n75 4.5005
R1698 VPWR.n108 VPWR.n101 4.5005
R1699 VPWR.n113 VPWR.n112 4.5005
R1700 VPWR.n114 VPWR.n105 4.5005
R1701 VPWR.n189 VPWR.n188 4.5005
R1702 VPWR.n178 VPWR.n50 4.5005
R1703 VPWR.n181 VPWR.n59 4.5005
R1704 VPWR.n253 VPWR.n252 4.5005
R1705 VPWR.n31 VPWR.n30 4.5005
R1706 VPWR.n28 VPWR.n21 4.5005
R1707 VPWR.n306 VPWR.n305 4.5005
R1708 VPWR.n295 VPWR.n282 4.5005
R1709 VPWR.n300 VPWR.n299 4.5005
R1710 VPWR.n214 VPWR.n213 4.5005
R1711 VPWR.n201 VPWR.n200 4.5005
R1712 VPWR.n205 VPWR.n43 4.5005
R1713 VPWR.n358 VPWR.n357 4.5005
R1714 VPWR.n362 VPWR.n361 4.5005
R1715 VPWR.n351 VPWR.n350 4.5005
R1716 VPWR.n452 VPWR.n451 4.5005
R1717 VPWR.n448 VPWR.n447 4.5005
R1718 VPWR.n314 VPWR.n313 4.5005
R1719 VPWR.n400 VPWR.n335 4.5005
R1720 VPWR.n413 VPWR.n412 4.5005
R1721 VPWR.n411 VPWR.n332 4.5005
R1722 VPWR.n419 VPWR.n418 4.5005
R1723 VPWR.n264 VPWR.n16 4.47065
R1724 VPWR.n225 VPWR.n39 4.36875
R1725 VPWR.n233 VPWR.n232 4.36875
R1726 VPWR.n436 VPWR.n325 4.36875
R1727 VPWR.n152 VPWR 4.26717
R1728 VPWR.n424 VPWR.n423 4.12612
R1729 VPWR.n249 VPWR.n246 4.04887
R1730 VPWR.n186 VPWR.n53 4.02033
R1731 VPWR.n186 VPWR.n57 4.02033
R1732 VPWR.n125 VPWR.n120 4.02033
R1733 VPWR.n125 VPWR.n123 4.02033
R1734 VPWR.n211 VPWR.n204 4.02033
R1735 VPWR.n211 VPWR.n209 4.02033
R1736 VPWR.n291 VPWR.n287 4.02033
R1737 VPWR.n291 VPWR.n290 4.02033
R1738 VPWR.n349 VPWR.n345 4.02033
R1739 VPWR.n349 VPWR.n348 4.02033
R1740 VPWR.n463 VPWR.n459 4.02033
R1741 VPWR.n463 VPWR.n462 4.02033
R1742 VPWR.t31 VPWR.t103 3.64572
R1743 VPWR.t13 VPWR.t127 3.64572
R1744 VPWR.n270 VPWR.n269 3.47425
R1745 VPWR.n405 VPWR.n336 3.47425
R1746 VPWR.n157 VPWR.n156 3.43925
R1747 VPWR.n160 VPWR.n159 3.43925
R1748 VPWR.n130 VPWR.n129 3.43925
R1749 VPWR.n133 VPWR.n132 3.43925
R1750 VPWR.n182 VPWR.n46 3.43925
R1751 VPWR.n191 VPWR.n190 3.43925
R1752 VPWR.n258 VPWR.n257 3.43925
R1753 VPWR.n255 VPWR.n254 3.43925
R1754 VPWR.n298 VPWR.n4 3.43925
R1755 VPWR.n308 VPWR.n307 3.43925
R1756 VPWR.n219 VPWR.n218 3.43925
R1757 VPWR.n216 VPWR.n215 3.43925
R1758 VPWR.n366 VPWR.n365 3.43925
R1759 VPWR.n356 VPWR.n355 3.43925
R1760 VPWR.n417 VPWR.n416 3.43925
R1761 VPWR.n402 VPWR.n401 3.43925
R1762 VPWR.n83 VPWR.n73 3.4105
R1763 VPWR.n84 VPWR.n74 3.4105
R1764 VPWR.n110 VPWR.n102 3.4105
R1765 VPWR.n111 VPWR.n104 3.4105
R1766 VPWR.n49 VPWR.n47 3.4105
R1767 VPWR.n180 VPWR.n179 3.4105
R1768 VPWR.n26 VPWR.n24 3.4105
R1769 VPWR.n29 VPWR.n22 3.4105
R1770 VPWR.n7 VPWR.n5 3.4105
R1771 VPWR.n297 VPWR.n296 3.4105
R1772 VPWR.n198 VPWR.n196 3.4105
R1773 VPWR.n199 VPWR.n44 3.4105
R1774 VPWR.n353 VPWR.n352 3.4105
R1775 VPWR.n364 VPWR.n363 3.4105
R1776 VPWR.n469 VPWR.n468 3.4105
R1777 VPWR.n469 VPWR.n311 3.4105
R1778 VPWR.n468 VPWR.n467 3.4105
R1779 VPWR.n445 VPWR.n311 3.4105
R1780 VPWR.n450 VPWR.n449 3.4105
R1781 VPWR.n446 VPWR.n312 3.4105
R1782 VPWR.n334 VPWR.n333 3.4105
R1783 VPWR.n415 VPWR.n414 3.4105
R1784 VPWR.t91 VPWR.t118 3.35739
R1785 VPWR.n269 VPWR.n268 3.2477
R1786 VPWR.n270 VPWR.n14 3.2477
R1787 VPWR.n396 VPWR.n336 3.2477
R1788 VPWR.n512 VPWR.n511 3.23917
R1789 VPWR.n529 VPWR.n528 3.23136
R1790 VPWR.n495 VPWR.n494 3.22655
R1791 VPWR.n267 VPWR.n16 3.219
R1792 VPWR.n303 VPWR.n277 3.2005
R1793 VPWR.n302 VPWR.n280 3.12116
R1794 VPWR.n241 VPWR.n34 3.06827
R1795 VPWR.n125 VPWR.n124 3.04861
R1796 VPWR.n291 VPWR.n283 3.04861
R1797 VPWR.n463 VPWR.n315 3.04861
R1798 VPWR.n464 VPWR.n320 2.91308
R1799 VPWR.n464 VPWR.n456 2.91308
R1800 VPWR.n277 VPWR.n276 2.87861
R1801 VPWR.n491 VPWR.n490 2.84665
R1802 VPWR.n487 VPWR.n485 2.84665
R1803 VPWR.n501 VPWR.n499 2.84665
R1804 VPWR.n504 VPWR.n500 2.84665
R1805 VPWR.n518 VPWR.n516 2.84665
R1806 VPWR.n521 VPWR.n517 2.84665
R1807 VPWR.n534 VPWR.n533 2.84665
R1808 VPWR.n535 VPWR.n531 2.84665
R1809 VPWR.n437 VPWR.n436 2.74336
R1810 VPWR.n53 VPWR.n51 2.63539
R1811 VPWR.n57 VPWR.n55 2.63539
R1812 VPWR.n120 VPWR.n118 2.63539
R1813 VPWR.n123 VPWR.n121 2.63539
R1814 VPWR.n280 VPWR.n278 2.63539
R1815 VPWR.n204 VPWR.n202 2.63539
R1816 VPWR.n209 VPWR.n207 2.63539
R1817 VPWR.n287 VPWR.n285 2.63539
R1818 VPWR.n290 VPWR.n288 2.63539
R1819 VPWR.n345 VPWR.n343 2.63539
R1820 VPWR.n348 VPWR.n346 2.63539
R1821 VPWR.n459 VPWR.n457 2.63539
R1822 VPWR.n462 VPWR.n460 2.63539
R1823 VPWR.n274 VPWR.n273 2.63233
R1824 VPWR.n275 VPWR.n274 2.61352
R1825 VPWR.n56 VPWR.n55 2.37495
R1826 VPWR.n52 VPWR.n51 2.37495
R1827 VPWR.n122 VPWR.n121 2.37495
R1828 VPWR.n119 VPWR.n118 2.37495
R1829 VPWR.n279 VPWR.n278 2.37495
R1830 VPWR.n208 VPWR.n207 2.37495
R1831 VPWR.n203 VPWR.n202 2.37495
R1832 VPWR.n289 VPWR.n288 2.37495
R1833 VPWR.n286 VPWR.n285 2.37495
R1834 VPWR.n347 VPWR.n346 2.37495
R1835 VPWR.n344 VPWR.n343 2.37495
R1836 VPWR.n461 VPWR.n460 2.37495
R1837 VPWR.n458 VPWR.n457 2.37495
R1838 VPWR.n302 VPWR.n281 2.33701
R1839 VPWR.n439 VPWR.n438 2.33701
R1840 VPWR.n493 VPWR.n482 2.28169
R1841 VPWR.n503 VPWR.n498 2.28169
R1842 VPWR.n520 VPWR.n515 2.28169
R1843 VPWR.n544 VPWR.n543 2.28169
R1844 VPWR.t99 VPWR.t31 2.24371
R1845 VPWR.t0 VPWR.t13 2.24371
R1846 VPWR.n284 VPWR.n281 2.03225
R1847 VPWR.n440 VPWR.n439 2.03225
R1848 VPWR.n320 VPWR.n318 2.01703
R1849 VPWR.n456 VPWR.n454 2.01703
R1850 VPWR.n438 VPWR.n437 1.93066
R1851 VPWR.n455 VPWR.n454 1.88416
R1852 VPWR.n319 VPWR.n318 1.88416
R1853 VPWR.n541 VPWR.n532 1.88285
R1854 VPWR.n406 VPWR.n405 1.73737
R1855 VPWR.n365 VPWR.n0 1.69188
R1856 VPWR.n355 VPWR.n0 1.69188
R1857 VPWR.n218 VPWR.n217 1.69188
R1858 VPWR.n217 VPWR.n216 1.69188
R1859 VPWR.n192 VPWR.n46 1.69188
R1860 VPWR.n192 VPWR.n191 1.69188
R1861 VPWR.n309 VPWR.n4 1.69188
R1862 VPWR.n309 VPWR.n308 1.69188
R1863 VPWR.n131 VPWR.n130 1.69188
R1864 VPWR.n132 VPWR.n131 1.69188
R1865 VPWR.n469 VPWR.n310 1.69188
R1866 VPWR.n416 VPWR.n2 1.69188
R1867 VPWR.n401 VPWR.n2 1.69188
R1868 VPWR.n257 VPWR.n256 1.69188
R1869 VPWR.n256 VPWR.n255 1.69188
R1870 VPWR.n158 VPWR.n157 1.69188
R1871 VPWR.n159 VPWR.n158 1.69188
R1872 VPWR.n407 VPWR.n406 1.51082
R1873 VPWR.n382 VPWR.n379 1.4005
R1874 VPWR.n479 VPWR.n478 1.38219
R1875 VPWR.n276 VPWR.n274 1.2502
R1876 VPWR.n430 VPWR.n429 1.16414
R1877 VPWR.n502 VPWR.n496 1.143
R1878 VPWR.n519 VPWR.n513 1.143
R1879 VPWR.n481 VPWR.n479 1.13977
R1880 VPWR.n545 VPWR.n530 1.13675
R1881 VPWR.n144 VPWR.n143 1.12991
R1882 VPWR.n494 VPWR.n480 1.12991
R1883 VPWR.n511 VPWR.n497 1.12991
R1884 VPWR.n528 VPWR.n527 1.12991
R1885 VPWR.n381 VPWR.n338 1.07613
R1886 VPWR.n376 VPWR.n375 1.0005
R1887 VPWR.n513 VPWR.n512 0.862816
R1888 VPWR.n246 VPWR.n245 0.833988
R1889 VPWR.n495 VPWR.n479 0.823939
R1890 VPWR.n530 VPWR.n529 0.770881
R1891 VPWR.n371 VPWR.n370 0.753441
R1892 VPWR.n496 VPWR.n495 0.729231
R1893 VPWR.n472 VPWR 0.660687
R1894 VPWR.n395 VPWR.n394 0.635211
R1895 VPWR.n432 VPWR.n431 0.635211
R1896 VPWR.n250 VPWR.n249 0.595849
R1897 VPWR.n192 VPWR.n45 0.55065
R1898 VPWR.n243 VPWR.n242 0.529426
R1899 VPWR.n476 VPWR.n475 0.500125
R1900 VPWR.n195 VPWR.n194 0.500125
R1901 VPWR.n478 VPWR 0.467141
R1902 VPWR VPWR.n472 0.466259
R1903 VPWR.n131 VPWR.n103 0.431025
R1904 VPWR.n158 VPWR.n45 0.431025
R1905 VPWR.n423 VPWR.n422 0.42364
R1906 VPWR.n529 VPWR.n513 0.392323
R1907 VPWR.n193 VPWR.n3 0.3805
R1908 VPWR.n470 VPWR.n1 0.3805
R1909 VPWR.n194 VPWR.n23 0.3805
R1910 VPWR.n475 VPWR.n474 0.3805
R1911 VPWR.n139 VPWR.n138 0.376971
R1912 VPWR.n512 VPWR.n496 0.360318
R1913 VPWR.n389 VPWR.n337 0.323189
R1914 VPWR.n226 VPWR.n225 0.305262
R1915 VPWR.n232 VPWR.n35 0.305262
R1916 VPWR.n292 VPWR.n284 0.305262
R1917 VPWR.n433 VPWR.n325 0.305262
R1918 VPWR.n441 VPWR.n440 0.305262
R1919 VPWR.n489 VPWR.t171 0.27666
R1920 VPWR.n486 VPWR.t171 0.27666
R1921 VPWR.t85 VPWR.n507 0.27666
R1922 VPWR.n508 VPWR.t85 0.27666
R1923 VPWR.t172 VPWR.n524 0.27666
R1924 VPWR.n525 VPWR.t172 0.27666
R1925 VPWR.t163 VPWR.n538 0.27666
R1926 VPWR.n539 VPWR.t163 0.27666
R1927 VPWR.n293 VPWR.n283 0.239726
R1928 VPWR.n465 VPWR.n315 0.239726
R1929 VPWR.n268 VPWR.n267 0.227049
R1930 VPWR.n273 VPWR.n14 0.227049
R1931 VPWR.n397 VPWR.n396 0.227049
R1932 VPWR.n408 VPWR.n407 0.227049
R1933 VPWR.n124 VPWR 0.217591
R1934 VPWR.n226 VPWR.n224 0.209973
R1935 VPWR.n472 VPWR 0.168795
R1936 VPWR.n217 VPWR.n0 0.1603
R1937 VPWR.n469 VPWR.n309 0.1603
R1938 VPWR.n256 VPWR.n2 0.1603
R1939 VPWR VPWR.n12 0.145148
R1940 VPWR.n195 VPWR.n192 0.14385
R1941 VPWR.n131 VPWR.n3 0.14385
R1942 VPWR.n158 VPWR.n23 0.14385
R1943 VPWR.n124 VPWR 0.141725
R1944 VPWR.n283 VPWR 0.141725
R1945 VPWR.n315 VPWR 0.141725
R1946 VPWR.n277 VPWR.n10 0.140696
R1947 VPWR.n177 VPWR.n176 0.120292
R1948 VPWR.n176 VPWR.n60 0.120292
R1949 VPWR.n171 VPWR.n60 0.120292
R1950 VPWR.n169 VPWR.n64 0.120292
R1951 VPWR.n67 VPWR.n66 0.120292
R1952 VPWR.n163 VPWR.n67 0.120292
R1953 VPWR.n154 VPWR.n76 0.120292
R1954 VPWR.n149 VPWR.n91 0.120292
R1955 VPWR.n149 VPWR.n148 0.120292
R1956 VPWR.n147 VPWR.n93 0.120292
R1957 VPWR.n142 VPWR.n93 0.120292
R1958 VPWR.n141 VPWR.n97 0.120292
R1959 VPWR.n229 VPWR.n37 0.120292
R1960 VPWR.n234 VPWR.n37 0.120292
R1961 VPWR.n236 VPWR.n235 0.120292
R1962 VPWR.n261 VPWR.n260 0.120292
R1963 VPWR.n261 VPWR.n17 0.120292
R1964 VPWR.n265 VPWR.n17 0.120292
R1965 VPWR.n271 VPWR.n15 0.120292
R1966 VPWR.n272 VPWR.n271 0.120292
R1967 VPWR.n272 VPWR.n13 0.120292
R1968 VPWR.n373 VPWR.n372 0.120292
R1969 VPWR.n373 VPWR.n339 0.120292
R1970 VPWR.n383 VPWR.n339 0.120292
R1971 VPWR.n384 VPWR.n383 0.120292
R1972 VPWR.n385 VPWR.n384 0.120292
R1973 VPWR.n392 VPWR.n391 0.120292
R1974 VPWR.n393 VPWR.n392 0.120292
R1975 VPWR.n420 VPWR.n329 0.120292
R1976 VPWR.n426 VPWR.n329 0.120292
R1977 VPWR.n427 VPWR.n426 0.120292
R1978 VPWR.n428 VPWR.n427 0.120292
R1979 VPWR.n428 VPWR.n326 0.120292
R1980 VPWR.n434 VPWR.n326 0.120292
R1981 VPWR.n435 VPWR.n323 0.120292
R1982 VPWR.n442 VPWR.n323 0.120292
R1983 VPWR.n475 VPWR.n1 0.120125
R1984 VPWR.n194 VPWR.n193 0.120125
R1985 VPWR.n103 VPWR.n45 0.120125
R1986 VPWR.n242 VPWR.n241 0.106285
R1987 VPWR.n221 VPWR 0.104667
R1988 VPWR.n229 VPWR 0.104667
R1989 VPWR.n239 VPWR 0.104667
R1990 VPWR.n12 VPWR 0.098273
R1991 VPWR VPWR.n170 0.0981562
R1992 VPWR.n66 VPWR 0.0981562
R1993 VPWR VPWR.n162 0.0981562
R1994 VPWR VPWR.n147 0.0981562
R1995 VPWR VPWR.n141 0.0981562
R1996 VPWR.n227 VPWR 0.0981562
R1997 VPWR.n228 VPWR 0.0981562
R1998 VPWR.n235 VPWR 0.0981562
R1999 VPWR.n240 VPWR 0.0981562
R2000 VPWR.n266 VPWR 0.0981562
R2001 VPWR VPWR.n15 0.0981562
R2002 VPWR.n372 VPWR 0.0981562
R2003 VPWR.n391 VPWR 0.0981562
R2004 VPWR.n398 VPWR 0.0981562
R2005 VPWR.n399 VPWR 0.0981562
R2006 VPWR.n435 VPWR 0.0981562
R2007 VPWR.n91 VPWR 0.0968542
R2008 VPWR.n135 VPWR 0.0968542
R2009 VPWR.n222 VPWR 0.0968542
R2010 VPWR.n160 VPWR.n72 0.0950946
R2011 VPWR.n156 VPWR.n75 0.0950946
R2012 VPWR.n133 VPWR.n101 0.0950946
R2013 VPWR.n129 VPWR.n105 0.0950946
R2014 VPWR.n190 VPWR.n189 0.0950946
R2015 VPWR.n182 VPWR.n181 0.0950946
R2016 VPWR.n254 VPWR.n253 0.0950946
R2017 VPWR.n258 VPWR.n21 0.0950946
R2018 VPWR.n307 VPWR.n306 0.0950946
R2019 VPWR.n299 VPWR.n298 0.0950946
R2020 VPWR.n215 VPWR.n214 0.0950946
R2021 VPWR.n219 VPWR.n43 0.0950946
R2022 VPWR.n357 VPWR.n356 0.0950946
R2023 VPWR.n366 VPWR.n351 0.0950946
R2024 VPWR.n451 VPWR.n445 0.0950946
R2025 VPWR.n467 VPWR.n313 0.0950946
R2026 VPWR.n402 VPWR.n400 0.0950946
R2027 VPWR.n417 VPWR.n332 0.0950946
R2028 VPWR.n443 VPWR 0.0916458
R2029 VPWR VPWR.n177 0.0851354
R2030 VPWR VPWR.n169 0.0851354
R2031 VPWR.n188 VPWR.n48 0.0838333
R2032 VPWR.n213 VPWR.n197 0.0838333
R2033 VPWR.n31 VPWR.n28 0.0838333
R2034 VPWR.n300 VPWR.n294 0.0838333
R2035 VPWR.n358 VPWR.n354 0.0838333
R2036 VPWR.n412 VPWR.n411 0.0838333
R2037 VPWR.n466 VPWR.n314 0.0838333
R2038 VPWR.n187 VPWR.n50 0.0812292
R2039 VPWR.n82 VPWR.n81 0.0812292
R2040 VPWR.n108 VPWR.n100 0.0812292
R2041 VPWR.n212 VPWR.n201 0.0812292
R2042 VPWR.n252 VPWR.n251 0.0812292
R2043 VPWR.n361 VPWR.n359 0.0812292
R2044 VPWR.n409 VPWR.n335 0.0812292
R2045 VPWR VPWR.n134 0.0799271
R2046 VPWR VPWR.n6 0.0799271
R2047 VPWR.n444 VPWR 0.0799271
R2048 VPWR.n184 VPWR.n59 0.0760208
R2049 VPWR.n162 VPWR.n161 0.0760208
R2050 VPWR.n115 VPWR.n113 0.0760208
R2051 VPWR.n205 VPWR.n42 0.0760208
R2052 VPWR.n301 VPWR.n282 0.0760208
R2053 VPWR.n368 VPWR.n350 0.0760208
R2054 VPWR.n403 VPWR.n399 0.0760208
R2055 VPWR.n447 VPWR.n321 0.0760208
R2056 VPWR.n155 VPWR.n154 0.0708125
R2057 VPWR.n260 VPWR.n259 0.0708125
R2058 VPWR.n420 VPWR.n419 0.0708125
R2059 VPWR.n128 VPWR 0.0695104
R2060 VPWR.n85 VPWR.n83 0.0680676
R2061 VPWR.n85 VPWR.n84 0.0680676
R2062 VPWR.n112 VPWR.n110 0.0680676
R2063 VPWR.n112 VPWR.n111 0.0680676
R2064 VPWR.n178 VPWR.n49 0.0680676
R2065 VPWR.n180 VPWR.n178 0.0680676
R2066 VPWR.n30 VPWR.n26 0.0680676
R2067 VPWR.n30 VPWR.n29 0.0680676
R2068 VPWR.n295 VPWR.n7 0.0680676
R2069 VPWR.n297 VPWR.n295 0.0680676
R2070 VPWR.n200 VPWR.n198 0.0680676
R2071 VPWR.n200 VPWR.n199 0.0680676
R2072 VPWR.n362 VPWR.n353 0.0680676
R2073 VPWR.n363 VPWR.n362 0.0680676
R2074 VPWR.n450 VPWR.n448 0.0680676
R2075 VPWR.n448 VPWR.n446 0.0680676
R2076 VPWR.n413 VPWR.n334 0.0680676
R2077 VPWR.n414 VPWR.n413 0.0680676
R2078 VPWR.n87 VPWR 0.0643021
R2079 VPWR.n481 VPWR 0.06425
R2080 VPWR.n502 VPWR 0.06425
R2081 VPWR.n519 VPWR 0.06425
R2082 VPWR VPWR.n545 0.06425
R2083 VPWR.n305 VPWR 0.0590938
R2084 VPWR VPWR.n452 0.0590938
R2085 VPWR.n74 VPWR.n73 0.0574697
R2086 VPWR.n104 VPWR.n102 0.0574697
R2087 VPWR.n179 VPWR.n47 0.0574697
R2088 VPWR.n24 VPWR.n22 0.0574697
R2089 VPWR.n296 VPWR.n5 0.0574697
R2090 VPWR.n196 VPWR.n44 0.0574697
R2091 VPWR.n364 VPWR.n352 0.0574697
R2092 VPWR.n449 VPWR.n311 0.0574697
R2093 VPWR.n468 VPWR.n312 0.0574697
R2094 VPWR.n415 VPWR.n333 0.0574697
R2095 VPWR VPWR.n25 0.0538854
R2096 VPWR.n259 VPWR.n20 0.0499792
R2097 VPWR.n1 VPWR 0.047625
R2098 VPWR.n193 VPWR 0.047625
R2099 VPWR.n103 VPWR 0.047625
R2100 VPWR.n477 VPWR 0.0472062
R2101 VPWR.n471 VPWR 0.0472062
R2102 VPWR.n473 VPWR 0.0472062
R2103 VPWR VPWR.n477 0.0469161
R2104 VPWR VPWR.n471 0.0469161
R2105 VPWR.n473 VPWR 0.0469161
R2106 VPWR.n59 VPWR.n54 0.0447708
R2107 VPWR.n161 VPWR.n71 0.0447708
R2108 VPWR.n113 VPWR.n109 0.0447708
R2109 VPWR.n206 VPWR.n205 0.0447708
R2110 VPWR.n27 VPWR.n25 0.0447708
R2111 VPWR.n360 VPWR.n350 0.0447708
R2112 VPWR.n404 VPWR.n403 0.0447708
R2113 VPWR.n447 VPWR.n322 0.0447708
R2114 VPWR.n83 VPWR.n72 0.0410405
R2115 VPWR.n84 VPWR.n75 0.0410405
R2116 VPWR.n110 VPWR.n101 0.0410405
R2117 VPWR.n111 VPWR.n105 0.0410405
R2118 VPWR.n189 VPWR.n49 0.0410405
R2119 VPWR.n181 VPWR.n180 0.0410405
R2120 VPWR.n253 VPWR.n26 0.0410405
R2121 VPWR.n29 VPWR.n21 0.0410405
R2122 VPWR.n306 VPWR.n7 0.0410405
R2123 VPWR.n299 VPWR.n297 0.0410405
R2124 VPWR.n214 VPWR.n198 0.0410405
R2125 VPWR.n199 VPWR.n43 0.0410405
R2126 VPWR.n357 VPWR.n353 0.0410405
R2127 VPWR.n363 VPWR.n351 0.0410405
R2128 VPWR.n451 VPWR.n450 0.0410405
R2129 VPWR.n446 VPWR.n313 0.0410405
R2130 VPWR.n400 VPWR.n334 0.0410405
R2131 VPWR.n414 VPWR.n332 0.0410405
R2132 VPWR.n54 VPWR.n50 0.0395625
R2133 VPWR.n81 VPWR.n71 0.0395625
R2134 VPWR.n109 VPWR.n108 0.0395625
R2135 VPWR.n206 VPWR.n201 0.0395625
R2136 VPWR.n252 VPWR.n27 0.0395625
R2137 VPWR.n305 VPWR.n304 0.0395625
R2138 VPWR.n361 VPWR.n360 0.0395625
R2139 VPWR.n404 VPWR.n335 0.0395625
R2140 VPWR.n452 VPWR.n322 0.0395625
R2141 VPWR.n135 VPWR 0.0382604
R2142 VPWR VPWR.n443 0.0382604
R2143 VPWR.n88 VPWR 0.0356562
R2144 VPWR.n13 VPWR 0.0356562
R2145 VPWR.n88 VPWR.n87 0.0343542
R2146 VPWR.n28 VPWR.n20 0.0343542
R2147 VPWR.n411 VPWR.n410 0.0343542
R2148 VPWR.n419 VPWR 0.0343542
R2149 VPWR.n355 VPWR.n352 0.0292489
R2150 VPWR.n365 VPWR.n364 0.0292489
R2151 VPWR.n216 VPWR.n196 0.0292489
R2152 VPWR.n218 VPWR.n44 0.0292489
R2153 VPWR.n191 VPWR.n47 0.0292489
R2154 VPWR.n179 VPWR.n46 0.0292489
R2155 VPWR.n308 VPWR.n5 0.0292489
R2156 VPWR.n296 VPWR.n4 0.0292489
R2157 VPWR.n132 VPWR.n102 0.0292489
R2158 VPWR.n130 VPWR.n104 0.0292489
R2159 VPWR.n312 VPWR.n310 0.0292489
R2160 VPWR.n449 VPWR.n310 0.0292489
R2161 VPWR.n401 VPWR.n333 0.0292489
R2162 VPWR.n416 VPWR.n415 0.0292489
R2163 VPWR.n255 VPWR.n24 0.0292489
R2164 VPWR.n257 VPWR.n22 0.0292489
R2165 VPWR.n159 VPWR.n73 0.0292489
R2166 VPWR.n157 VPWR.n74 0.0292489
R2167 VPWR.n128 VPWR.n127 0.0291458
R2168 VPWR.n294 VPWR.n293 0.0291458
R2169 VPWR VPWR.n442 0.0291458
R2170 VPWR.n466 VPWR.n465 0.0291458
R2171 VPWR.n170 VPWR 0.0239375
R2172 VPWR VPWR.n76 0.0239375
R2173 VPWR VPWR.n97 0.0239375
R2174 VPWR VPWR.n221 0.0239375
R2175 VPWR.n478 VPWR 0.0231242
R2176 VPWR.n477 VPWR.n476 0.0231188
R2177 VPWR.n471 VPWR.n470 0.0231188
R2178 VPWR.n474 VPWR.n473 0.0231188
R2179 VPWR.n171 VPWR 0.0226354
R2180 VPWR VPWR.n64 0.0226354
R2181 VPWR.n163 VPWR 0.0226354
R2182 VPWR.n148 VPWR 0.0226354
R2183 VPWR.n142 VPWR 0.0226354
R2184 VPWR.n222 VPWR 0.0226354
R2185 VPWR VPWR.n227 0.0226354
R2186 VPWR VPWR.n234 0.0226354
R2187 VPWR VPWR.n239 0.0226354
R2188 VPWR.n240 VPWR 0.0226354
R2189 VPWR VPWR.n265 0.0226354
R2190 VPWR.n266 VPWR 0.0226354
R2191 VPWR.n11 VPWR 0.0226354
R2192 VPWR.n304 VPWR 0.0226354
R2193 VPWR.n282 VPWR 0.0226354
R2194 VPWR.n385 VPWR 0.0226354
R2195 VPWR.n393 VPWR 0.0226354
R2196 VPWR VPWR.n398 0.0226354
R2197 VPWR VPWR.n434 0.0226354
R2198 VPWR.n453 VPWR 0.0226354
R2199 VPWR VPWR.n86 0.0200312
R2200 VPWR.n476 VPWR.n0 0.018125
R2201 VPWR.n470 VPWR.n469 0.018125
R2202 VPWR.n474 VPWR.n2 0.018125
R2203 VPWR.n217 VPWR.n195 0.01695
R2204 VPWR.n309 VPWR.n3 0.01695
R2205 VPWR.n256 VPWR.n23 0.01695
R2206 VPWR.n127 VPWR 0.016125
R2207 VPWR VPWR.n228 0.016125
R2208 VPWR.n236 VPWR 0.016125
R2209 VPWR.n410 VPWR 0.016125
R2210 VPWR.n183 VPWR 0.0148229
R2211 VPWR.n155 VPWR 0.0148229
R2212 VPWR.n114 VPWR 0.0148229
R2213 VPWR.n418 VPWR.n417 0.0140135
R2214 VPWR.n418 VPWR 0.0140135
R2215 VPWR VPWR.n48 0.0122188
R2216 VPWR VPWR.n197 0.0122188
R2217 VPWR.n354 VPWR 0.0122188
R2218 VPWR.n184 VPWR.n183 0.0083125
R2219 VPWR.n115 VPWR.n114 0.0083125
R2220 VPWR.n220 VPWR.n42 0.0083125
R2221 VPWR VPWR.n220 0.0083125
R2222 VPWR.n301 VPWR.n300 0.0083125
R2223 VPWR.n368 VPWR.n367 0.0083125
R2224 VPWR.n367 VPWR 0.0083125
R2225 VPWR.n321 VPWR.n314 0.0083125
R2226 VPWR.n188 VPWR.n187 0.00310417
R2227 VPWR.n86 VPWR.n82 0.00310417
R2228 VPWR.n134 VPWR.n100 0.00310417
R2229 VPWR.n213 VPWR.n212 0.00310417
R2230 VPWR.n251 VPWR.n31 0.00310417
R2231 VPWR.n11 VPWR.n6 0.00310417
R2232 VPWR.n359 VPWR.n358 0.00310417
R2233 VPWR.n412 VPWR.n409 0.00310417
R2234 VPWR.n453 VPWR.n444 0.00310417
R2235 select1.n0 select1.t1 323.55
R2236 select1.n0 select1.t0 195.017
R2237 select1.n1 select1.n0 152
R2238 select1.n3 select1 18.8151
R2239 select1 select1.n2 10.2766
R2240 select1.n2 select1 6.7304
R2241 select1.n1 select1 1.45205
R2242 select1.n2 select1.n1 0.792253
R2243 select1.n3 select1 0.0384464
R2244 select1 select1.n3 0.0128547
R2245 passgatesCtrl_0.net10.n1 passgatesCtrl_0.net10.t4 260.322
R2246 passgatesCtrl_0.net10.n3 passgatesCtrl_0.net10.n0 207.22
R2247 passgatesCtrl_0.net10.n1 passgatesCtrl_0.net10.t3 175.169
R2248 passgatesCtrl_0.net10.n2 passgatesCtrl_0.net10.n1 153.13
R2249 passgatesCtrl_0.net10 passgatesCtrl_0.net10.t2 132.067
R2250 passgatesCtrl_0.net10.n0 passgatesCtrl_0.net10.t1 26.5955
R2251 passgatesCtrl_0.net10.n0 passgatesCtrl_0.net10.t0 26.5955
R2252 passgatesCtrl_0.net10 passgatesCtrl_0.net10.n3 17.4717
R2253 passgatesCtrl_0.net10.n3 passgatesCtrl_0.net10 12.2141
R2254 passgatesCtrl_0.net10 passgatesCtrl_0.net10.n2 9.39918
R2255 passgatesCtrl_0.net10.n2 passgatesCtrl_0.net10 3.2005
R2256 passgatesCtrl_0.net1.n12 passgatesCtrl_0.net1.t17 562.236
R2257 passgatesCtrl_0.net1.t17 passgatesCtrl_0.net1.t9 392.027
R2258 passgatesCtrl_0.net1.n20 passgatesCtrl_0.net1.t6 327.99
R2259 passgatesCtrl_0.net1.n3 passgatesCtrl_0.net1.t11 323.55
R2260 passgatesCtrl_0.net1.n1 passgatesCtrl_0.net1.t1 319.171
R2261 passgatesCtrl_0.net1.n24 passgatesCtrl_0.net1.t7 293.969
R2262 passgatesCtrl_0.net1.n8 passgatesCtrl_0.net1.t13 256.07
R2263 passgatesCtrl_0.net1.n17 passgatesCtrl_0.net1.t19 231.835
R2264 passgatesCtrl_0.net1.n6 passgatesCtrl_0.net1.t8 230.155
R2265 passgatesCtrl_0.net1 passgatesCtrl_0.net1.t0 209.923
R2266 passgatesCtrl_0.net1.n16 passgatesCtrl_0.net1.t18 206.19
R2267 passgatesCtrl_0.net1.n20 passgatesCtrl_0.net1.t15 199.457
R2268 passgatesCtrl_0.net1.n3 passgatesCtrl_0.net1.t2 195.017
R2269 passgatesCtrl_0.net1.n14 passgatesCtrl_0.net1.t5 185.376
R2270 passgatesCtrl_0.net1.n6 passgatesCtrl_0.net1.t3 157.856
R2271 passgatesCtrl_0.net1.n17 passgatesCtrl_0.net1.t14 157.07
R2272 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n16 154.657
R2273 passgatesCtrl_0.net1.n18 passgatesCtrl_0.net1.n17 154.048
R2274 passgatesCtrl_0.net1.n7 passgatesCtrl_0.net1.n6 153.147
R2275 passgatesCtrl_0.net1.n25 passgatesCtrl_0.net1.n24 152
R2276 passgatesCtrl_0.net1.n21 passgatesCtrl_0.net1.n20 152
R2277 passgatesCtrl_0.net1.n15 passgatesCtrl_0.net1.n14 152
R2278 passgatesCtrl_0.net1.n9 passgatesCtrl_0.net1.n8 152
R2279 passgatesCtrl_0.net1.n4 passgatesCtrl_0.net1.n3 152
R2280 passgatesCtrl_0.net1.n8 passgatesCtrl_0.net1.t12 150.03
R2281 passgatesCtrl_0.net1.n16 passgatesCtrl_0.net1.t16 148.35
R2282 passgatesCtrl_0.net1.n24 passgatesCtrl_0.net1.t4 138.338
R2283 passgatesCtrl_0.net1.n14 passgatesCtrl_0.net1.t10 137.177
R2284 passgatesCtrl_0.net1.n5 passgatesCtrl_0.net1 28.0894
R2285 passgatesCtrl_0.net1.n11 passgatesCtrl_0.net1.n10 25.2401
R2286 passgatesCtrl_0.net1.n13 passgatesCtrl_0.net1.n12 22.4834
R2287 passgatesCtrl_0.net1.n0 passgatesCtrl_0.net1 21.6175
R2288 passgatesCtrl_0.net1.n11 passgatesCtrl_0.net1.n7 20.5972
R2289 passgatesCtrl_0.net1.n23 passgatesCtrl_0.net1.n22 16.5589
R2290 passgatesCtrl_0.net1.n9 passgatesCtrl_0.net1 16.3845
R2291 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n25 15.2457
R2292 passgatesCtrl_0.net1.n26 passgatesCtrl_0.net1 14.6453
R2293 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n26 13.9801
R2294 passgatesCtrl_0.net1.n21 passgatesCtrl_0.net1 12.1605
R2295 passgatesCtrl_0.net1.n19 passgatesCtrl_0.net1.n0 11.55
R2296 passgatesCtrl_0.net1.n22 passgatesCtrl_0.net1 10.8805
R2297 passgatesCtrl_0.net1.n0 passgatesCtrl_0.net1.n15 10.8365
R2298 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n2 10.6976
R2299 passgatesCtrl_0.net1.n19 passgatesCtrl_0.net1.n18 9.3005
R2300 passgatesCtrl_0.net1.n12 passgatesCtrl_0.net1 8.92171
R2301 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n1 7.73474
R2302 passgatesCtrl_0.net1.n23 passgatesCtrl_0.net1.n19 7.40435
R2303 passgatesCtrl_0.net1.n5 passgatesCtrl_0.net1.n4 7.1685
R2304 passgatesCtrl_0.net1.n0 passgatesCtrl_0.net1.n13 6.03757
R2305 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n5 4.62272
R2306 passgatesCtrl_0.net1.n10 passgatesCtrl_0.net1.n9 4.6085
R2307 passgatesCtrl_0.net1.n10 passgatesCtrl_0.net1 4.58918
R2308 passgatesCtrl_0.net1.n18 passgatesCtrl_0.net1 4.3525
R2309 passgatesCtrl_0.net1.n26 passgatesCtrl_0.net1 4.26717
R2310 passgatesCtrl_0.net1.n22 passgatesCtrl_0.net1 3.62717
R2311 passgatesCtrl_0.net1.n13 passgatesCtrl_0.net1.n11 3.29171
R2312 passgatesCtrl_0.net1.n7 passgatesCtrl_0.net1 3.24826
R2313 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n23 3.14198
R2314 passgatesCtrl_0.net1.n15 passgatesCtrl_0.net1 3.0725
R2315 passgatesCtrl_0.net1.n4 passgatesCtrl_0.net1 2.9445
R2316 passgatesCtrl_0.net1.n1 passgatesCtrl_0.net1 2.48634
R2317 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n21 2.34717
R2318 passgatesCtrl_0.net1.n2 passgatesCtrl_0.net1 2.19479
R2319 passgatesCtrl_0.net1.n25 passgatesCtrl_0.net1 2.06502
R2320 passgatesCtrl_0.net1.n2 passgatesCtrl_0.net1 1.80756
R2321 passgatesCtrl_0.net1.n5 passgatesCtrl_0.net1 1.6645
R2322 A3.n1 A3.t3 26.3998
R2323 A3.n1 A3.t2 23.5483
R2324 A3.n0 A3.t0 12.7127
R2325 A3.n0 A3.t1 10.8578
R2326 A3.n2 A3.n1 3.12177
R2327 A3.n2 A3.n0 1.81453
R2328 A3.n3 A3.n2 1.1255
R2329 A3.n3 A3 0.210543
R2330 A3 A3.n3 0.0655
R2331 Z3.n1 Z3.t3 23.6581
R2332 Z3.n3 Z3.t2 23.3739
R2333 Z3.n1 Z3.t1 10.7528
R2334 Z3.n0 Z3.t0 10.6417
R2335 Z3.n2 Z3.n1 1.30064
R2336 Z3.n5 Z3.n4 0.924585
R2337 Z3.n3 Z3.n2 0.726502
R2338 Z3.n2 Z3.n0 0.512491
R2339 Z3.n4 Z3.n0 0.359663
R2340 Z3.n4 Z3.n3 0.216071
R2341 Z3.n5 Z3 0.0656042
R2342 Z3 Z3.n5 0.0376287
R2343 select0.n0 select0.t1 323.55
R2344 select0.n0 select0.t0 195.017
R2345 select0.n1 select0.n0 152
R2346 select0 select0.n2 14.4176
R2347 select0.n2 select0 6.7304
R2348 select0.n3 select0 2.87104
R2349 select0.n1 select0 1.45205
R2350 select0.n2 select0.n1 0.792253
R2351 select0.n3 select0 0.0696964
R2352 select0 select0.n3 0.0230291
R2353 Z2.n1 Z2.t0 23.6581
R2354 Z2.n3 Z2.t1 23.3739
R2355 Z2.n1 Z2.t3 10.7528
R2356 Z2.n0 Z2.t2 10.6417
R2357 Z2.n2 Z2.n1 1.30064
R2358 Z2.n5 Z2.n4 0.936641
R2359 Z2.n3 Z2.n2 0.726502
R2360 Z2.n2 Z2.n0 0.512491
R2361 Z2.n4 Z2.n0 0.359663
R2362 Z2.n4 Z2.n3 0.216071
R2363 Z2.n5 Z2 0.0776605
R2364 Z2 Z2.n5 0.0561931
R2365 A2.n1 A2.t0 26.3998
R2366 A2.n1 A2.t1 23.5483
R2367 A2.n0 A2.t3 12.7127
R2368 A2.n0 A2.t2 10.8578
R2369 A2.n2 A2.n1 3.12177
R2370 A2.n2 A2.n0 1.81453
R2371 A2.n3 A2.n2 1.1255
R2372 A2.n3 A2 0.219402
R2373 A2 A2.n3 0.0655
R2374 Z4.n1 Z4.t3 23.6581
R2375 Z4.n3 Z4.t2 23.3739
R2376 Z4.n1 Z4.t0 10.7528
R2377 Z4.n0 Z4.t1 10.6417
R2378 Z4.n2 Z4.n1 1.30064
R2379 Z4 Z4.n4 0.983856
R2380 Z4.n3 Z4.n2 0.726502
R2381 Z4.n2 Z4.n0 0.512491
R2382 Z4.n4 Z4.n0 0.359663
R2383 Z4.n4 Z4.n3 0.216071
R2384 A4.n1 A4.t3 26.3998
R2385 A4.n1 A4.t2 23.5483
R2386 A4.n0 A4.t0 12.7127
R2387 A4.n0 A4.t1 10.8578
R2388 A4.n2 A4.n1 3.12177
R2389 A4.n2 A4.n0 1.81453
R2390 A4.n3 A4.n2 1.1255
R2391 A4 A4.n3 0.134513
R2392 A4.n3 A4 0.0655
R2393 Z1.n1 Z1.t2 23.6581
R2394 Z1.n3 Z1.t3 23.3739
R2395 Z1.n1 Z1.t0 10.7528
R2396 Z1.n0 Z1.t1 10.6417
R2397 Z1.n2 Z1.n1 1.30064
R2398 Z1 Z1.n4 0.983856
R2399 Z1.n3 Z1.n2 0.726502
R2400 Z1.n2 Z1.n0 0.512491
R2401 Z1.n4 Z1.n0 0.359663
R2402 Z1.n4 Z1.n3 0.216071
R2403 A1.n1 A1.t2 26.3998
R2404 A1.n1 A1.t3 23.5483
R2405 A1.n0 A1.t0 12.7127
R2406 A1.n0 A1.t1 10.8578
R2407 A1.n2 A1.n1 3.12177
R2408 A1.n2 A1.n0 1.81453
R2409 A1.n3 A1.n2 1.1255
R2410 A1.n3 A1 0.21549
R2411 A1 A1.n3 0.0655
C0 passgatesCtrl_0.net6 a_n2057_n1942# 0.001427f
C1 passgatex4_0.GN1 passgatesCtrl_0.net1 0.055547f
C2 passgatesCtrl_0.net7 a_n1459_n3306# 1.39e-19
C3 passgatex4_0.GP4 a_n2883_n1648# 0.033357f
C4 A1 passgatesCtrl_0._02_ 2.53e-20
C5 passgatex4_0.GN4 Z4 0.443709f
C6 passgatex4_0.GN3 passgatex4_0.GN1 5.26e-19
C7 a_n491_n3280# a_n539_n3518# 5.96e-19
C8 passgatesCtrl_0.net3 passgatesCtrl_0._02_ 6.01e-20
C9 a_n1878_n4368# a_n1984_n4368# 0.313533f
C10 a_n801_n4216# passgatesCtrl_0._04_ 5.33e-19
C11 passgatesCtrl_0.net8 passgatesCtrl_0.net3 8.71e-21
C12 a_n1503_n2192# a_n1459_n3306# 6.43e-21
C13 passgatesCtrl_0.net6 a_n2639_n2040# 0.046149f
C14 passgatesCtrl_0._05_ passgatesCtrl_0.net2 0.019534f
C15 passgatesCtrl_0._03_ passgatex4_0.GP1 4.32e-20
C16 passgatesCtrl_0.net1 a_n2015_n2040# 0.134894f
C17 passgatesCtrl_0.net9 a_n1913_n1429# 0.031948f
C18 passgatex4_0.GP4 passgatesCtrl_0.net7 3.05e-20
C19 a_n2429_n1328# passgatesCtrl_0.net9 2.52e-19
C20 passgatesCtrl_0.net4 passgatesCtrl_0.net5 0.024789f
C21 passgatesCtrl_0.net5 a_n1003_n2040# 6.98e-19
C22 passgatex4_0.GN1 a_n995_n3605# 3.14e-19
C23 passgatex4_0.GN1 a_n1173_n2218# 1.7e-19
C24 passgatex4_0.GN3 a_n2015_n2040# 7.19e-21
C25 passgatesCtrl_0.net1 passgatex4_0.GN2 0.117828f
C26 passgatesCtrl_0.net2 a_n2975_n2192# 0.006018f
C27 passgatex4_0.GP2 A1 0.002086f
C28 passgatesCtrl_0.net4 a_n715_n3850# 8.15e-19
C29 select0 a_n1878_n4368# 3.96e-19
C30 VPWR a_n1637_n1429# 0.221714f
C31 passgatex4_0.GN3 passgatex4_0.GN2 0.051202f
C32 passgatex4_0.GP2 passgatesCtrl_0.net3 3.9e-21
C33 a_n1361_n1429# passgatesCtrl_0.net10 5.14e-19
C34 passgatesCtrl_0.net5 a_n1913_n1429# 0.038008f
C35 passgatesCtrl_0.net1 a_n2883_n1648# -6.59e-36
C36 passgatex4_0.GP4 passgatex4_0.GN4 3.44232f
C37 a_n1085_n1429# passgatesCtrl_0._00_ 4.99e-20
C38 a_n2429_n1328# passgatesCtrl_0.net5 8.98e-21
C39 select1 a_n1084_n4216# 0.005547f
C40 a_n1963_n3280# passgatesCtrl_0.net1 2.5e-19
C41 VPWR a_n491_n3280# 0.291441f
C42 a_n1635_n3306# a_n1459_n3306# 0.185422f
C43 a_n1173_n2218# passgatex4_0.GN2 0.001025f
C44 select0 a_n1984_n4368# 1.65e-19
C45 passgatesCtrl_0.net7 passgatesCtrl_0.net1 0.492308f
C46 passgatesCtrl_0.net2 passgatesCtrl_0._00_ 0.181488f
C47 a_n482_n4216# a_n715_n3850# 0.001428f
C48 passgatesCtrl_0._01_ a_n1045_n1942# 3.51e-19
C49 a_n597_n2040# a_n675_n1648# 0.003066f
C50 passgatex4_0.GN1 passgatesCtrl_0.net5 0.002166f
C51 passgatex4_0.GN3 passgatesCtrl_0.net7 1.52e-19
C52 passgatesCtrl_0.net1 a_n587_n3458# 0.002306f
C53 Z3 passgatex4_0.GN2 2.12e-20
C54 passgatesCtrl_0.net6 a_n1003_n2040# 2.87e-20
C55 passgatesCtrl_0._01_ a_n2185_n2218# 0.001002f
C56 passgatex4_0.GN4 passgatesCtrl_0.net1 5.43e-19
C57 passgatex4_0.GN1 a_n715_n3850# 0.001005f
C58 a_n1503_n2192# passgatesCtrl_0.net1 0.040031f
C59 a_n1459_n3306# passgatesCtrl_0.net2 0.096716f
C60 select1 passgatesCtrl_0.net2 0.026514f
C61 passgatex4_0.GN3 passgatex4_0.GN4 0.155269f
C62 passgatesCtrl_0.net6 a_n1913_n1429# 0.008072f
C63 a_n1503_n2192# passgatex4_0.GN3 1.78e-19
C64 a_n2015_n2040# passgatesCtrl_0.net5 0.012287f
C65 passgatesCtrl_0.net9 a_n2883_n1648# 0.123724f
C66 passgatesCtrl_0.net10 a_n675_n1648# 7.12e-20
C67 a_n597_n2040# passgatex4_0.GP1 9.87e-19
C68 passgatex4_0.GN1 A2 3.14e-19
C69 a_n539_n3518# passgatesCtrl_0._04_ 0.001297f
C70 passgatesCtrl_0.net5 passgatex4_0.GN2 0.011028f
C71 a_n2015_n2040# a_n2057_n1942# 3.5e-20
C72 a_n1503_n2192# a_n1173_n2218# 0.018393f
C73 passgatex4_0.GN3 Z2 0.00126f
C74 VPWR a_n1361_n1429# 0.211763f
C75 passgatesCtrl_0.net5 a_n2883_n1648# 4.81e-20
C76 passgatex4_0.GP4 passgatesCtrl_0.net2 0.005696f
C77 passgatesCtrl_0.net1 a_n1084_n4216# 0.004309f
C78 passgatesCtrl_0.net4 a_n1003_n2040# 0.001809f
C79 a_n1635_n3306# passgatesCtrl_0.net1 0.001693f
C80 passgatesCtrl_0.net7 passgatesCtrl_0.net9 1.77e-20
C81 VPWR a_n951_n2736# 0.193152f
C82 a_n1963_n3280# passgatesCtrl_0.net5 0.115837f
C83 a_n1637_n1429# passgatesCtrl_0.net8 0.001796f
C84 passgatex4_0.GP3 passgatex4_0.GP1 5.06e-19
C85 passgatex4_0.GN4 Z3 0.00128f
C86 A2 passgatex4_0.GN2 3.8137f
C87 passgatesCtrl_0.net1 a_n1085_n1429# 1.87e-20
C88 a_n1459_n3306# passgatesCtrl_0.net3 2.01e-19
C89 VPWR Z1 2.98463f
C90 a_n482_n4216# select0 0.266581f
C91 passgatex4_0.GN4 passgatesCtrl_0.net9 4.06e-19
C92 passgatesCtrl_0.net7 passgatesCtrl_0.net5 0.002751f
C93 passgatex4_0.GN3 a_n1085_n1429# 6.29e-19
C94 a_n1135_n4368# VPWR 0.162421f
C95 a_n1084_n4216# a_n995_n3605# 1.65e-19
C96 passgatesCtrl_0.net6 a_n2015_n2040# 0.013011f
C97 VPWR passgatesCtrl_0._04_ 0.211525f
C98 passgatesCtrl_0.net7 a_n715_n3850# 0.00214f
C99 passgatex4_0.GP2 a_n1637_n1429# 0.002575f
C100 Z3 Z2 7.67e-19
C101 passgatex4_0.GN1 select0 0.005832f
C102 passgatex4_0.GP4 A1 1.34e-19
C103 passgatesCtrl_0.net6 passgatex4_0.GN2 5.41e-20
C104 passgatesCtrl_0.net1 passgatesCtrl_0.net2 1.72543f
C105 passgatex4_0.GN4 passgatesCtrl_0.net5 0.05537f
C106 a_n1503_n2192# passgatesCtrl_0.net5 0.003576f
C107 a_n715_n3850# a_n587_n3458# 0.004764f
C108 a_n1173_n2218# a_n1085_n1429# 4.77e-20
C109 passgatex4_0.GN3 passgatesCtrl_0.net2 0.006039f
C110 passgatesCtrl_0.net6 a_n2883_n1648# 4.16e-19
C111 VPWR a_n2161_n4368# 0.173581f
C112 passgatex4_0.GN1 passgatesCtrl_0.net4 0.083575f
C113 passgatex4_0.GN1 a_n1003_n2040# 4.06e-19
C114 VPWR a_n675_n1648# 0.230164f
C115 passgatesCtrl_0.net2 a_n995_n3605# 0.043831f
C116 passgatesCtrl_0.net2 a_n1173_n2218# 0.177825f
C117 passgatex4_0.GN4 A2 1.95e-19
C118 a_n1085_n1429# passgatesCtrl_0.net9 4.15e-21
C119 passgatesCtrl_0.net6 passgatesCtrl_0.net7 5.12e-20
C120 passgatex4_0.GN4 a_n2639_n2040# 3.33e-20
C121 passgatesCtrl_0.net1 A1 0.049065f
C122 a_n1635_n3306# passgatesCtrl_0.net5 0.0036f
C123 VPWR passgatesCtrl_0._03_ 0.196287f
C124 passgatesCtrl_0.net4 passgatex4_0.GN2 0.005352f
C125 a_n1003_n2040# passgatex4_0.GN2 0.003895f
C126 VPWR passgatex4_0.GP1 2.34735f
C127 passgatesCtrl_0.net1 passgatesCtrl_0.net3 0.178768f
C128 passgatex4_0.GN3 A1 4.37e-19
C129 passgatesCtrl_0.net2 a_n2480_n4368# 0.162398f
C130 a_n2015_n2040# a_n1913_n1429# 1.05e-19
C131 passgatex4_0.GN1 a_n482_n4216# 0.00164f
C132 A2 Z2 4.51569f
C133 passgatesCtrl_0.net5 a_n1085_n1429# 0.032876f
C134 a_n1361_n1429# passgatesCtrl_0.net8 0.004727f
C135 passgatex4_0.GN4 passgatesCtrl_0.net6 0.043823f
C136 VPWR a_n1227_n2736# 0.241578f
C137 a_n1503_n2192# passgatesCtrl_0.net6 0.001672f
C138 VPWR a_n2465_n2164# 3.98e-19
C139 a_n1913_n1429# passgatex4_0.GN2 5.52e-20
C140 passgatesCtrl_0.net2 passgatesCtrl_0.net9 0.086587f
C141 a_n1135_n4368# a_n988_n4394# 0.003683f
C142 passgatesCtrl_0.net4 a_n1963_n3280# 0.001365f
C143 a_n1637_n1429# passgatesCtrl_0._00_ 1.44e-19
C144 VPWR a_n1045_n1942# 6.29e-19
C145 a_n988_n4394# passgatesCtrl_0._04_ 0.001033f
C146 VPWR passgatesCtrl_0._01_ 0.225859f
C147 passgatesCtrl_0._03_ a_n1507_n3280# 8.17e-20
C148 a_n995_n3605# passgatesCtrl_0.net3 1.28e-21
C149 a_n1173_n2218# passgatesCtrl_0.net3 0.010683f
C150 passgatesCtrl_0.net2 passgatesCtrl_0.net5 0.544042f
C151 passgatex4_0.GP2 a_n1361_n1429# 0.134077f
C152 VPWR a_n2185_n2218# 0.130016f
C153 passgatex4_0.GP3 passgatesCtrl_0.net10 0.234131f
C154 passgatesCtrl_0.net4 passgatesCtrl_0.net7 3.73e-19
C155 passgatesCtrl_0.net2 a_n715_n3850# 0.067356f
C156 Z3 A1 4.74e-21
C157 VPWR a_n801_n4216# 0.191329f
C158 a_n1084_n4216# a_n1984_n4368# 1.1e-19
C159 passgatesCtrl_0.net4 a_n587_n3458# 4.09e-19
C160 passgatex4_0.GN1 passgatex4_0.GN2 0.033541f
C161 passgatesCtrl_0.net7 a_n1913_n1429# 6.2e-20
C162 passgatex4_0.GP2 Z1 3.73e-21
C163 a_n1503_n2192# a_n1003_n2040# 4.74e-20
C164 passgatesCtrl_0.net2 a_n1878_n4368# 0.010759f
C165 passgatesCtrl_0.net6 a_n1085_n1429# 0.001258f
C166 passgatesCtrl_0._02_ a_n675_n1648# 0.194553f
C167 passgatex4_0.GN4 a_n1913_n1429# 0.112321f
C168 passgatesCtrl_0.net8 a_n675_n1648# 6.36e-19
C169 passgatesCtrl_0.net2 a_n2639_n2040# 0.180659f
C170 a_n2015_n2040# passgatex4_0.GN2 1.39e-19
C171 passgatesCtrl_0.net5 A1 5.61e-21
C172 select0 a_n1084_n4216# 0.001575f
C173 a_n482_n4216# passgatesCtrl_0.net7 6.47e-19
C174 passgatex4_0.GN4 a_n2429_n1328# 2.79e-21
C175 a_n715_n3850# A1 0.001233f
C176 passgatesCtrl_0.net5 passgatesCtrl_0.net3 0.001999f
C177 VPWR a_n597_n2040# 0.179575f
C178 a_n434_n1942# passgatex4_0.GP1 2.65e-19
C179 passgatesCtrl_0.net6 passgatesCtrl_0.net2 0.0936f
C180 passgatex4_0.GN1 passgatesCtrl_0.net7 0.028089f
C181 passgatesCtrl_0.net2 a_n1984_n4368# 0.051248f
C182 passgatesCtrl_0.net4 a_n1084_n4216# 0.00141f
C183 passgatex4_0.GP1 passgatesCtrl_0._02_ 6.66e-20
C184 passgatex4_0.GP2 a_n675_n1648# 5.94e-19
C185 passgatesCtrl_0.net4 a_n1635_n3306# 0.007618f
C186 A4 passgatex4_0.GP3 0.16204f
C187 passgatex4_0.GN1 a_n587_n3458# 1.58e-19
C188 A1 A2 1.81909f
C189 passgatex4_0.GN1 passgatex4_0.GN4 2.04e-19
C190 a_n1227_n2736# passgatesCtrl_0.net8 1.26e-20
C191 passgatesCtrl_0.net4 a_n1085_n1429# 2.63e-19
C192 a_n1361_n1429# passgatesCtrl_0._00_ 8.1e-20
C193 VPWR passgatesCtrl_0.net10 0.395163f
C194 A3 passgatex4_0.GP1 2.46e-21
C195 VPWR passgatex4_0.GP3 1.84344f
C196 select0 passgatesCtrl_0.net2 0.002824f
C197 passgatesCtrl_0.net7 passgatex4_0.GN2 0.34798f
C198 a_n1637_n1429# passgatesCtrl_0.net1 1.96e-19
C199 passgatex4_0.GP2 passgatex4_0.GP1 0.008406f
C200 passgatesCtrl_0.net8 a_n1045_n1942# 9.1e-19
C201 passgatesCtrl_0._01_ passgatesCtrl_0.net8 0.208131f
C202 a_n801_n4216# a_n988_n4394# 0.159555f
C203 passgatex4_0.GN1 Z2 4.77e-21
C204 passgatex4_0.GN3 a_n1637_n1429# 0.14217f
C205 a_n1503_n2192# a_n2015_n2040# 0.014264f
C206 passgatesCtrl_0.net8 a_n2185_n2218# 1.99e-21
C207 VPWR a_n1701_n4368# 0.143966f
C208 passgatex4_0.GP2 a_n1227_n2736# 4.59e-20
C209 passgatesCtrl_0.net4 passgatesCtrl_0.net2 0.097522f
C210 a_n1459_n3306# a_n1361_n1429# 8.17e-21
C211 passgatesCtrl_0.net2 a_n1003_n2040# 0.166925f
C212 passgatex4_0.GN4 passgatex4_0.GN2 5.8e-19
C213 a_n1503_n2192# passgatex4_0.GN2 4.62e-19
C214 a_n2189_n1429# a_n2185_n2218# 0.011493f
C215 a_n491_n3280# passgatesCtrl_0.net1 0.007927f
C216 VPWR a_n539_n3518# 0.259999f
C217 passgatex4_0.GN1 a_n1084_n4216# 4.22e-19
C218 passgatesCtrl_0.net7 a_n1963_n3280# 3.8e-20
C219 passgatesCtrl_0.net2 a_n1913_n1429# 3.2e-19
C220 passgatex4_0.GN4 a_n2883_n1648# 2.19e-19
C221 passgatesCtrl_0.net2 a_n2429_n1328# 1.42e-19
C222 passgatesCtrl_0._01_ passgatex4_0.GP2 4.67e-20
C223 select1 Z1 2.26e-19
C224 select0 A1 0.040389f
C225 passgatex4_0.GN1 a_n1085_n1429# 3.8e-19
C226 passgatesCtrl_0._05_ a_n2465_n2164# 5.76e-19
C227 Z2 passgatex4_0.GN2 0.427031f
C228 select0 passgatesCtrl_0.net3 1.33e-20
C229 a_n1135_n4368# select1 0.004485f
C230 a_n597_n2040# a_n434_n1942# 0.004767f
C231 a_n482_n4216# passgatesCtrl_0.net2 0.001264f
C232 select1 passgatesCtrl_0._04_ 3.6e-20
C233 passgatesCtrl_0.net4 A1 6.83e-21
C234 a_n597_n2040# passgatesCtrl_0._02_ 0.106303f
C235 VPWR A4 1.54289f
C236 passgatex4_0.GN4 passgatesCtrl_0.net7 4.64e-20
C237 a_n1503_n2192# passgatesCtrl_0.net7 2.69e-21
C238 passgatesCtrl_0._01_ passgatesCtrl_0._05_ 6.19e-21
C239 a_n1637_n1429# passgatesCtrl_0.net9 1.63e-19
C240 passgatesCtrl_0.net4 passgatesCtrl_0.net3 0.130377f
C241 a_n1003_n2040# passgatesCtrl_0.net3 7.73e-20
C242 passgatex4_0.GN1 passgatesCtrl_0.net2 0.068323f
C243 a_n1085_n1429# passgatex4_0.GN2 0.002397f
C244 select1 a_n2161_n4368# 0.002569f
C245 passgatesCtrl_0._01_ a_n2975_n2192# 3.25e-21
C246 a_n2975_n2192# a_n2185_n2218# 1.06e-20
C247 a_n1637_n1429# passgatesCtrl_0.net5 0.033814f
C248 passgatesCtrl_0.net10 passgatesCtrl_0._02_ 5.35e-20
C249 a_n1963_n3280# a_n1635_n3306# 0.017591f
C250 passgatesCtrl_0.net1 a_n1361_n1429# 2.44e-20
C251 passgatesCtrl_0.net2 a_n2015_n2040# 0.185322f
C252 passgatesCtrl_0.net8 passgatesCtrl_0.net10 1.06e-19
C253 a_n482_n4216# A1 0.001912f
C254 passgatex4_0.GN3 a_n1361_n1429# 0.109673f
C255 a_n1701_n4368# a_n988_n4394# 1.09e-19
C256 passgatesCtrl_0.net2 passgatex4_0.GN2 0.06846f
C257 a_n2189_n1429# passgatesCtrl_0.net10 0.041816f
C258 passgatesCtrl_0.net7 a_n1635_n3306# 1.83e-19
C259 a_n951_n2736# passgatesCtrl_0.net1 0.02864f
C260 a_n491_n3280# passgatesCtrl_0.net5 6.09e-20
C261 passgatex4_0.GP3 a_n2189_n1429# 0.110988f
C262 passgatesCtrl_0._03_ a_n1459_n3306# 9.63e-19
C263 select1 passgatesCtrl_0._03_ 4.71e-19
C264 passgatex4_0.GN1 A1 4.96968f
C265 a_n1459_n3306# passgatex4_0.GP1 1.14e-19
C266 VPWR a_n1507_n3280# 0.003544f
C267 passgatesCtrl_0.net1 Z1 3.3e-21
C268 passgatesCtrl_0.net2 a_n2883_n1648# 0.012477f
C269 A3 passgatex4_0.GP3 3.97267f
C270 passgatesCtrl_0.net7 a_n1085_n1429# 4.02e-19
C271 passgatesCtrl_0._01_ passgatesCtrl_0._00_ 5.18e-20
C272 passgatex4_0.GN1 passgatesCtrl_0.net3 0.357097f
C273 a_n2185_n2218# passgatesCtrl_0._00_ 0.0957f
C274 passgatex4_0.GP2 passgatesCtrl_0.net10 9.63e-20
C275 a_n1135_n4368# passgatesCtrl_0.net1 0.001335f
C276 passgatex4_0.GP2 passgatex4_0.GP3 0.007549f
C277 passgatesCtrl_0.net1 passgatesCtrl_0._04_ 0.050056f
C278 a_n1963_n3280# passgatesCtrl_0.net2 0.04096f
C279 passgatex4_0.GP4 passgatex4_0.GP1 2.41e-19
C280 a_n1637_n1429# passgatesCtrl_0.net6 0.218518f
C281 passgatesCtrl_0.net7 passgatesCtrl_0.net2 0.090257f
C282 A1 passgatex4_0.GN2 0.151745f
C283 passgatesCtrl_0._05_ passgatex4_0.GP3 6.13e-19
C284 passgatesCtrl_0.net3 passgatex4_0.GN2 0.069726f
C285 passgatesCtrl_0.net2 a_n587_n3458# 0.001719f
C286 a_n1361_n1429# passgatesCtrl_0.net9 7.62e-20
C287 passgatesCtrl_0.net1 a_n675_n1648# 8.22e-19
C288 a_n995_n3605# passgatesCtrl_0._04_ 0.294104f
C289 VPWR a_n988_n4394# 0.211037f
C290 a_n801_n4216# select1 0.001678f
C291 passgatex4_0.GN4 passgatesCtrl_0.net2 7.43e-19
C292 a_n1503_n2192# passgatesCtrl_0.net2 0.03779f
C293 passgatex4_0.GN1 a_n485_n2736# 0.003892f
C294 VPWR a_n434_n1942# 0.002344f
C295 passgatex4_0.GN3 a_n675_n1648# 1.89e-19
C296 VPWR passgatesCtrl_0._02_ 0.450634f
C297 a_n1361_n1429# passgatesCtrl_0.net5 0.230704f
C298 passgatex4_0.GP4 a_n2185_n2218# 2.89e-21
C299 VPWR passgatesCtrl_0.net8 0.561328f
C300 A3 A4 2.08862f
C301 passgatesCtrl_0._03_ passgatesCtrl_0.net1 9.6e-19
C302 passgatesCtrl_0.net7 A1 0.012018f
C303 passgatesCtrl_0.net1 passgatex4_0.GP1 0.003098f
C304 VPWR a_n2189_n1429# 0.195044f
C305 a_n951_n2736# passgatesCtrl_0.net5 6.35e-19
C306 passgatex4_0.GP2 A4 2.48e-20
C307 select0 a_n491_n3280# 4.9e-19
C308 passgatesCtrl_0.net7 passgatesCtrl_0.net3 0.034004f
C309 VPWR A3 1.61205f
C310 a_n1227_n2736# passgatesCtrl_0.net1 8.11e-19
C311 passgatex4_0.GN3 passgatex4_0.GP1 8.28e-19
C312 a_n587_n3458# A1 4.82e-20
C313 passgatesCtrl_0.net2 a_n1084_n4216# 0.001027f
C314 passgatesCtrl_0.net10 passgatesCtrl_0._00_ 0.005756f
C315 passgatex4_0.GN4 A1 1.92e-19
C316 a_n1635_n3306# passgatesCtrl_0.net2 0.200956f
C317 VPWR passgatex4_0.GP2 1.61055f
C318 passgatex4_0.GP3 passgatesCtrl_0._00_ 0.098299f
C319 a_n1637_n1429# a_n1913_n1429# 5.3e-19
C320 passgatesCtrl_0.net1 a_n1045_n1942# 0.001768f
C321 passgatesCtrl_0.net2 a_n1085_n1429# 0.006979f
C322 passgatesCtrl_0._01_ passgatesCtrl_0.net1 0.173572f
C323 a_n715_n3850# passgatesCtrl_0._04_ 0.099459f
C324 passgatesCtrl_0.net1 a_n2185_n2218# 0.184986f
C325 Z4 passgatex4_0.GP3 0.071646f
C326 a_n1227_n2736# a_n1173_n2218# 3.06e-19
C327 passgatesCtrl_0._01_ passgatex4_0.GN3 1.44e-19
C328 A1 Z2 0.004942f
C329 passgatex4_0.GN3 a_n2185_n2218# 4.42e-19
C330 passgatesCtrl_0.net6 a_n1361_n1429# 0.033794f
C331 VPWR passgatesCtrl_0._05_ 0.358831f
C332 a_n801_n4216# passgatesCtrl_0.net1 0.329151f
C333 passgatesCtrl_0.net7 a_n485_n2736# 0.002755f
C334 Z3 passgatex4_0.GP1 1.86e-21
C335 passgatesCtrl_0.net5 a_n675_n1648# 2.48e-19
C336 a_n1173_n2218# a_n1045_n1942# 0.005162f
C337 a_n1084_n4216# A1 7.64e-21
C338 VPWR a_n2975_n2192# 0.310075f
C339 passgatesCtrl_0._01_ a_n1173_n2218# 0.101852f
C340 a_n482_n4216# a_n491_n3280# 1.73e-21
C341 a_n1084_n4216# passgatesCtrl_0.net3 9.59e-22
C342 a_n1701_n4368# select1 0.004749f
C343 passgatex4_0.GP4 passgatesCtrl_0.net10 0.076097f
C344 a_n434_n1942# passgatesCtrl_0._02_ 4.96e-19
C345 passgatex4_0.GP4 passgatex4_0.GP3 0.057096f
C346 passgatex4_0.GN1 a_n491_n3280# 0.001658f
C347 a_n1135_n4368# a_n1984_n4368# 1.09e-19
C348 passgatesCtrl_0._03_ passgatesCtrl_0.net5 0.19429f
C349 passgatesCtrl_0.net5 passgatex4_0.GP1 0.0014f
C350 passgatesCtrl_0.net1 a_n597_n2040# 0.215616f
C351 passgatesCtrl_0.net8 passgatesCtrl_0._02_ 0.096563f
C352 a_n1637_n1429# passgatex4_0.GN2 2.05e-19
C353 a_n1227_n2736# passgatesCtrl_0.net5 0.002913f
C354 passgatesCtrl_0.net9 a_n2185_n2218# 6.62e-20
C355 select0 Z1 0.003513f
C356 VPWR passgatesCtrl_0._00_ 0.89146f
C357 passgatesCtrl_0.net2 A1 0.002113f
C358 A4 Z4 4.51497f
C359 a_n2161_n4368# a_n1984_n4368# 0.159555f
C360 a_n951_n2736# passgatesCtrl_0.net4 0.194653f
C361 passgatesCtrl_0.net2 passgatesCtrl_0.net3 0.095367f
C362 a_n951_n2736# a_n1003_n2040# 3.63e-19
C363 a_n1135_n4368# select0 5.8e-19
C364 passgatesCtrl_0.net5 a_n1045_n1942# 3.13e-20
C365 passgatex4_0.GP1 A2 0.122954f
C366 passgatesCtrl_0._01_ passgatesCtrl_0.net5 0.003676f
C367 passgatex4_0.GP2 passgatesCtrl_0._02_ 2.58e-19
C368 passgatesCtrl_0.net1 passgatesCtrl_0.net10 0.160369f
C369 a_n1173_n2218# a_n597_n2040# 8.8e-19
C370 passgatesCtrl_0.net5 a_n2185_n2218# 0.00379f
C371 VPWR Z4 2.81307f
C372 passgatesCtrl_0.net1 passgatex4_0.GP3 0.058232f
C373 passgatex4_0.GP2 passgatesCtrl_0.net8 0.008913f
C374 VPWR a_n1459_n3306# 0.260783f
C375 VPWR select1 1.30675f
C376 passgatex4_0.GN3 passgatesCtrl_0.net10 0.152678f
C377 passgatex4_0.GN3 passgatex4_0.GP3 2.37902f
C378 passgatesCtrl_0.net4 passgatesCtrl_0._04_ 0.00489f
C379 a_n1637_n1429# passgatesCtrl_0.net7 9.8e-20
C380 a_n2465_n2164# a_n2639_n2040# 0.006584f
C381 a_n2057_n1942# a_n2185_n2218# 0.005162f
C382 passgatesCtrl_0.net6 passgatesCtrl_0._03_ 2.14e-19
C383 passgatex4_0.GP2 A3 0.145029f
C384 passgatex4_0.GP4 A4 3.97306f
C385 a_n1701_n4368# passgatesCtrl_0.net1 3.89e-19
C386 a_n801_n4216# a_n715_n3850# 3.21e-19
C387 passgatex4_0.GN1 a_n1361_n1429# 2e-20
C388 passgatesCtrl_0.net1 a_n539_n3518# 0.107968f
C389 A1 passgatesCtrl_0.net3 1.84e-20
C390 passgatex4_0.GN4 a_n1637_n1429# 0.111188f
C391 passgatesCtrl_0._01_ a_n2639_n2040# 5.79e-21
C392 VPWR passgatex4_0.GP4 1.50532f
C393 passgatesCtrl_0.net7 a_n491_n3280# 0.200958f
C394 a_n2639_n2040# a_n2185_n2218# 0.002367f
C395 a_n951_n2736# passgatex4_0.GN1 0.135217f
C396 passgatesCtrl_0.net6 a_n1045_n1942# 2.07e-20
C397 passgatex4_0.GN1 Z1 0.428012f
C398 passgatesCtrl_0._01_ passgatesCtrl_0.net6 0.002059f
C399 select0 passgatex4_0.GP1 7.71e-19
C400 passgatesCtrl_0.net6 a_n2185_n2218# 0.029048f
C401 Z3 passgatex4_0.GP3 0.278332f
C402 a_n1135_n4368# passgatex4_0.GN1 1.78e-19
C403 passgatesCtrl_0.net9 passgatesCtrl_0.net10 0.181065f
C404 a_n1361_n1429# passgatex4_0.GN2 6.44e-19
C405 passgatex4_0.GP3 passgatesCtrl_0.net9 0.117574f
C406 passgatesCtrl_0.net4 passgatesCtrl_0._03_ 0.002493f
C407 passgatex4_0.GN1 passgatesCtrl_0._04_ 0.004444f
C408 passgatesCtrl_0.net4 passgatex4_0.GP1 3.09e-20
C409 passgatex4_0.GN3 A4 0.007063f
C410 a_n951_n2736# passgatex4_0.GN2 0.110403f
C411 a_n1227_n2736# passgatesCtrl_0.net4 0.041847f
C412 passgatesCtrl_0.net5 passgatesCtrl_0.net10 0.099696f
C413 VPWR passgatesCtrl_0.net1 2.63744f
C414 passgatesCtrl_0.net8 passgatesCtrl_0._00_ 1.17e-19
C415 Z1 passgatex4_0.GN2 6.82e-19
C416 passgatesCtrl_0.net3 a_n485_n2736# 0.011812f
C417 passgatex4_0.GP3 passgatesCtrl_0.net5 0.001185f
C418 VPWR passgatex4_0.GN3 0.518775f
C419 a_n2189_n1429# passgatesCtrl_0._00_ 6.88e-19
C420 passgatex4_0.GN1 a_n675_n1648# 8.62e-19
C421 select1 a_n988_n4394# 5.9e-19
C422 passgatesCtrl_0.net4 a_n1045_n1942# 2.33e-19
C423 a_n1003_n2040# a_n1045_n1942# 3.5e-20
C424 passgatesCtrl_0._05_ a_n2975_n2192# 0.225698f
C425 a_n801_n4216# select0 0.004124f
C426 passgatesCtrl_0._01_ a_n1003_n2040# 2.42e-19
C427 passgatesCtrl_0.net7 a_n1361_n1429# 1.77e-19
C428 passgatex4_0.GP2 passgatesCtrl_0._00_ 3.42e-20
C429 VPWR a_n995_n3605# 0.218874f
C430 VPWR a_n1173_n2218# 0.118575f
C431 a_n1637_n1429# passgatesCtrl_0.net2 6.58e-20
C432 passgatex4_0.GP3 A2 0.001646f
C433 a_n951_n2736# passgatesCtrl_0.net7 0.001413f
C434 A3 Z4 0.005563f
C435 passgatex4_0.GN4 a_n1361_n1429# 5.36e-19
C436 a_n1503_n2192# a_n1361_n1429# 0.010239f
C437 passgatex4_0.GN1 passgatex4_0.GP1 1.11922f
C438 a_n715_n3850# a_n539_n3518# 0.185422f
C439 passgatex4_0.GP3 a_n2639_n2040# 0.002737f
C440 passgatex4_0.GN2 a_n675_n1648# 0.021336f
C441 passgatex4_0.GP2 Z4 6e-21
C442 a_n1701_n4368# a_n1878_n4368# 0.134298f
C443 VPWR a_n2480_n4368# 0.27871f
C444 passgatex4_0.GN1 a_n1227_n2736# 0.109645f
C445 VPWR Z3 2.85844f
C446 passgatesCtrl_0._05_ passgatesCtrl_0._00_ 0.005299f
C447 a_n491_n3280# passgatesCtrl_0.net2 0.013113f
C448 passgatesCtrl_0.net6 passgatesCtrl_0.net10 0.043833f
C449 passgatesCtrl_0.net6 passgatex4_0.GP3 2.34e-19
C450 VPWR passgatesCtrl_0.net9 0.312028f
C451 passgatex4_0.GP4 a_n2189_n1429# 0.130626f
C452 passgatex4_0.GN1 a_n1045_n1942# 3.88e-20
C453 a_n587_n3458# passgatesCtrl_0._04_ 8.17e-20
C454 a_n2975_n2192# passgatesCtrl_0._00_ 0.012253f
C455 passgatesCtrl_0._01_ passgatex4_0.GN1 4.4e-20
C456 passgatex4_0.GP4 A3 0.001593f
C457 passgatex4_0.GP1 passgatex4_0.GN2 1.62948f
C458 a_n597_n2040# a_n1003_n2040# 4.09e-20
C459 a_n1701_n4368# a_n1984_n4368# 0.003683f
C460 VPWR passgatesCtrl_0.net5 0.609808f
C461 passgatex4_0.GP2 passgatex4_0.GP4 3.49e-19
C462 passgatesCtrl_0.net1 a_n988_n4394# 0.019707f
C463 passgatesCtrl_0.net7 a_n675_n1648# 0.109167f
C464 a_n1227_n2736# passgatex4_0.GN2 9.69e-19
C465 passgatesCtrl_0.net1 a_n434_n1942# 3.05e-19
C466 passgatex4_0.GN1 a_n801_n4216# 6.45e-19
C467 VPWR a_n715_n3850# 0.182247f
C468 passgatesCtrl_0._01_ a_n2015_n2040# 0.002311f
C469 passgatesCtrl_0.net1 passgatesCtrl_0._02_ 0.079473f
C470 a_n1361_n1429# a_n1085_n1429# 5.3e-19
C471 a_n491_n3280# A1 0.001919f
C472 passgatesCtrl_0._03_ a_n1963_n3280# 0.225915f
C473 A4 A2 2.39e-19
C474 VPWR a_n2057_n1942# 4.1e-19
C475 a_n2015_n2040# a_n2185_n2218# 0.101254f
C476 passgatesCtrl_0.net1 passgatesCtrl_0.net8 0.194974f
C477 a_n491_n3280# passgatesCtrl_0.net3 1.85e-19
C478 passgatesCtrl_0._01_ passgatex4_0.GN2 6.19e-19
C479 passgatex4_0.GN3 passgatesCtrl_0._02_ 1.13e-19
C480 VPWR a_n1878_n4368# 0.211692f
C481 a_n1701_n4368# select0 2.23e-19
C482 a_n1135_n4368# a_n1084_n4216# 0.134298f
C483 passgatex4_0.GP4 passgatesCtrl_0._05_ 6.86e-20
C484 passgatesCtrl_0.net1 a_n2189_n1429# 0.030465f
C485 passgatesCtrl_0.net7 passgatesCtrl_0._03_ 0.001559f
C486 passgatex4_0.GN3 passgatesCtrl_0.net8 0.002415f
C487 VPWR A2 1.62685f
C488 a_n988_n4394# a_n995_n3605# 0.011149f
C489 a_n1084_n4216# passgatesCtrl_0._04_ 2.48e-19
C490 passgatesCtrl_0.net7 passgatex4_0.GP1 0.068983f
C491 a_n1913_n1429# passgatesCtrl_0.net10 0.219762f
C492 passgatex4_0.GN3 a_n2189_n1429# 0.011181f
C493 select0 a_n539_n3518# 8.27e-19
C494 passgatesCtrl_0.net2 a_n1361_n1429# 1.59e-20
C495 VPWR a_n2639_n2040# 0.20743f
C496 a_n2429_n1328# passgatesCtrl_0.net10 0.009374f
C497 a_n1227_n2736# passgatesCtrl_0.net7 6.38e-19
C498 passgatex4_0.GP2 passgatesCtrl_0.net1 7.04e-20
C499 passgatex4_0.GN1 a_n597_n2040# 6.11e-19
C500 passgatex4_0.GN3 A3 3.80702f
C501 a_n2429_n1328# passgatex4_0.GP3 1.66e-19
C502 a_n1173_n2218# passgatesCtrl_0.net8 0.015061f
C503 passgatex4_0.GN4 passgatex4_0.GP1 3.45e-19
C504 a_n1503_n2192# passgatex4_0.GP1 3.01e-21
C505 a_n951_n2736# passgatesCtrl_0.net2 1.46e-19
C506 passgatesCtrl_0.net4 a_n539_n3518# 1.79e-19
C507 VPWR passgatesCtrl_0.net6 0.615644f
C508 passgatex4_0.GN3 passgatex4_0.GP2 2.40528f
C509 VPWR a_n1984_n4368# 0.222008f
C510 passgatesCtrl_0.net2 Z1 2.55e-19
C511 a_n1135_n4368# passgatesCtrl_0.net2 6.62e-19
C512 passgatesCtrl_0._05_ passgatesCtrl_0.net1 0.001365f
C513 passgatex4_0.GP1 Z2 0.065749f
C514 passgatex4_0.GP2 a_n1173_n2218# 5.22e-19
C515 passgatesCtrl_0.net2 passgatesCtrl_0._04_ 0.096582f
C516 select1 a_n1459_n3306# 3.4e-19
C517 a_n1085_n1429# a_n675_n1648# 0.031466f
C518 passgatex4_0.GN1 passgatex4_0.GP3 3.37e-19
C519 a_n597_n2040# passgatex4_0.GN2 0.009622f
C520 passgatex4_0.GP4 passgatesCtrl_0._00_ 0.039155f
C521 passgatesCtrl_0._01_ a_n1503_n2192# 0.213841f
C522 VPWR select0 0.625418f
C523 passgatesCtrl_0.net1 a_n2975_n2192# 7.01e-19
C524 passgatex4_0.GN4 a_n2185_n2218# 2.2e-21
C525 a_n1361_n1429# passgatesCtrl_0.net3 6.41e-20
C526 A3 Z3 4.51555f
C527 passgatesCtrl_0._03_ a_n1635_n3306# 0.074703f
C528 a_n2189_n1429# passgatesCtrl_0.net9 0.219432f
C529 a_n482_n4216# a_n539_n3518# 0.003312f
C530 a_n1635_n3306# passgatex4_0.GP1 6.97e-20
C531 a_n951_n2736# A1 1.79e-20
C532 passgatesCtrl_0.net5 passgatesCtrl_0._02_ 4.38e-19
C533 passgatesCtrl_0.net2 a_n2161_n4368# 0.383661f
C534 passgatex4_0.GP2 Z3 0.063817f
C535 a_n1227_n2736# a_n1084_n4216# 4.03e-19
C536 passgatex4_0.GP4 Z4 0.278468f
C537 passgatesCtrl_0.net5 passgatesCtrl_0.net8 0.012208f
C538 passgatesCtrl_0.net2 a_n675_n1648# 1.87e-20
C539 A1 Z1 4.51541f
C540 a_n951_n2736# passgatesCtrl_0.net3 0.037807f
C541 VPWR passgatesCtrl_0.net4 0.442407f
C542 VPWR a_n1003_n2040# 0.076471f
C543 passgatex4_0.GN1 a_n539_n3518# 0.001234f
C544 passgatesCtrl_0.net10 passgatex4_0.GN2 4.61e-20
C545 passgatex4_0.GP2 passgatesCtrl_0.net9 8.22e-21
C546 passgatesCtrl_0.net5 a_n2189_n1429# 0.002712f
C547 a_n1135_n4368# A1 2.48e-21
C548 passgatex4_0.GP3 passgatex4_0.GN2 0.001327f
C549 a_n1878_n4368# a_n988_n4394# 1.1e-19
C550 passgatesCtrl_0._04_ A1 2.11e-20
C551 a_n1227_n2736# a_n1085_n1429# 2.57e-19
C552 passgatesCtrl_0.net7 a_n597_n2040# 0.010689f
C553 VPWR a_n1913_n1429# 0.196943f
C554 passgatesCtrl_0.net10 a_n2883_n1648# 5.56e-19
C555 VPWR a_n2429_n1328# 1.96e-19
C556 passgatex4_0.GP3 a_n2883_n1648# 0.008642f
C557 passgatesCtrl_0.net1 passgatesCtrl_0._00_ 0.110008f
C558 passgatex4_0.GP2 passgatesCtrl_0.net5 0.125101f
C559 passgatesCtrl_0._03_ passgatesCtrl_0.net2 0.265291f
C560 passgatesCtrl_0.net2 passgatex4_0.GP1 0.078988f
C561 passgatex4_0.GN3 passgatesCtrl_0._00_ 6.68e-20
C562 passgatesCtrl_0.net4 a_n1507_n3280# 5.55e-19
C563 a_n1503_n2192# a_n597_n2040# 1.1e-19
C564 VPWR a_n482_n4216# 0.290651f
C565 a_n1227_n2736# passgatesCtrl_0.net2 0.006314f
C566 passgatesCtrl_0.net2 a_n2465_n2164# 0.001995f
C567 a_n988_n4394# a_n1984_n4368# 0.002297f
C568 A1 a_n675_n1648# 2.71e-20
C569 passgatesCtrl_0.net7 passgatesCtrl_0.net10 4.64e-20
C570 A3 A2 1.81997f
C571 a_n1459_n3306# passgatesCtrl_0.net1 0.20481f
C572 passgatex4_0.GN3 Z4 1.95e-20
C573 select1 passgatesCtrl_0.net1 0.002895f
C574 a_n1173_n2218# passgatesCtrl_0._00_ 1.7e-21
C575 VPWR passgatex4_0.GN1 0.938241f
C576 passgatesCtrl_0.net6 passgatesCtrl_0.net8 0.02671f
C577 passgatesCtrl_0.net2 a_n1045_n1942# 0.001911f
C578 passgatex4_0.GP2 A2 3.97567f
C579 passgatesCtrl_0._01_ passgatesCtrl_0.net2 0.218705f
C580 passgatesCtrl_0.net6 a_n2189_n1429# 1.92e-20
C581 passgatex4_0.GN4 passgatesCtrl_0.net10 0.039325f
C582 passgatesCtrl_0.net2 a_n2185_n2218# 0.042928f
C583 select0 a_n988_n4394# 0.001977f
C584 passgatex4_0.GN4 passgatex4_0.GP3 3.23503f
C585 A1 passgatex4_0.GP1 4.03203f
C586 VPWR a_n2015_n2040# 0.097823f
C587 passgatex4_0.GP4 passgatesCtrl_0.net1 0.00512f
C588 passgatesCtrl_0.net7 a_n539_n3518# 0.004605f
C589 a_n801_n4216# passgatesCtrl_0.net2 6.52e-19
C590 select1 a_n995_n3605# 2.55e-19
C591 passgatesCtrl_0.net3 passgatex4_0.GP1 0.001814f
C592 passgatex4_0.GP2 passgatesCtrl_0.net6 0.001965f
C593 passgatesCtrl_0.net9 passgatesCtrl_0._00_ 0.099215f
C594 VPWR passgatex4_0.GN2 0.389408f
C595 passgatex4_0.GN3 passgatex4_0.GP4 0.048689f
C596 a_n1227_n2736# passgatesCtrl_0.net3 0.23425f
C597 passgatex4_0.GP3 Z2 1.03e-20
C598 passgatesCtrl_0._05_ a_n2639_n2040# 0.114102f
C599 Z3 Z4 0.002331f
C600 a_n1003_n2040# passgatesCtrl_0._02_ 0.054258f
C601 VPWR a_n2883_n1648# 0.258847f
C602 select1 a_n2480_n4368# 0.270124f
C603 passgatesCtrl_0.net4 passgatesCtrl_0.net8 5.72e-20
C604 passgatesCtrl_0.net5 passgatesCtrl_0._00_ 0.002004f
C605 a_n1003_n2040# passgatesCtrl_0.net8 0.002587f
C606 a_n2975_n2192# a_n2639_n2040# 0.015664f
C607 passgatesCtrl_0.net6 passgatesCtrl_0._05_ 0.289483f
C608 a_n1637_n1429# a_n1361_n1429# 5.3e-19
C609 passgatesCtrl_0._01_ passgatesCtrl_0.net3 6.43e-19
C610 VPWR a_n1963_n3280# 0.266692f
C611 passgatesCtrl_0.net2 a_n597_n2040# 0.154638f
C612 a_n801_n4216# A1 1.16e-20
C613 passgatesCtrl_0.net8 a_n1913_n1429# 3.98e-20
C614 a_n1085_n1429# passgatesCtrl_0.net10 2.12e-19
C615 a_n2057_n1942# passgatesCtrl_0._00_ 3.51e-19
C616 passgatesCtrl_0.net6 a_n2975_n2192# 0.108594f
C617 passgatex4_0.GP1 a_n485_n2736# 2.46e-19
C618 a_n2189_n1429# a_n1913_n1429# 5.3e-19
C619 VPWR passgatesCtrl_0.net7 0.589224f
C620 passgatex4_0.GN4 A4 3.8425f
C621 passgatex4_0.GP4 Z3 1.58e-20
C622 a_n1459_n3306# passgatesCtrl_0.net5 7.33e-19
C623 passgatex4_0.GN3 passgatesCtrl_0.net1 0.027691f
C624 select1 passgatesCtrl_0.net5 2.72e-19
C625 passgatex4_0.GN1 a_n988_n4394# 4.16e-19
C626 VPWR a_n587_n3458# 2.56e-19
C627 passgatex4_0.GP4 passgatesCtrl_0.net9 0.376983f
C628 select1 a_n715_n3850# 1.42e-19
C629 passgatex4_0.GN1 a_n434_n1942# 1.09e-19
C630 a_n2639_n2040# passgatesCtrl_0._00_ 0.054291f
C631 VPWR passgatex4_0.GN4 0.255383f
C632 passgatesCtrl_0.net2 passgatesCtrl_0.net10 0.082322f
C633 VPWR a_n1503_n2192# 0.26412f
C634 passgatesCtrl_0.net2 passgatex4_0.GP3 0.137787f
C635 passgatex4_0.GN1 passgatesCtrl_0._02_ 0.005251f
C636 passgatesCtrl_0.net1 a_n995_n3605# 0.008453f
C637 passgatesCtrl_0.net1 a_n1173_n2218# 0.059436f
C638 a_n491_n3280# Z1 1.26e-20
C639 passgatex4_0.GN1 passgatesCtrl_0.net8 1.87e-19
C640 passgatex4_0.GP4 passgatesCtrl_0.net5 0.005756f
C641 select1 a_n1878_n4368# 0.009355f
C642 passgatesCtrl_0.net6 passgatesCtrl_0._00_ 0.194746f
C643 a_n597_n2040# passgatesCtrl_0.net3 7.1e-21
C644 a_n1701_n4368# passgatesCtrl_0.net2 0.003464f
C645 VPWR Z2 2.84785f
C646 passgatesCtrl_0.net2 a_n539_n3518# 0.242957f
C647 passgatex4_0.GP2 passgatex4_0.GN1 0.002408f
C648 passgatex4_0.GN2 passgatesCtrl_0._02_ 0.237149f
C649 VPWR a_n1084_n4216# 0.201932f
C650 passgatex4_0.GN3 Z3 0.427101f
C651 passgatesCtrl_0.net1 passgatesCtrl_0.net9 0.061468f
C652 VPWR a_n1635_n3306# 0.225849f
C653 select1 a_n1984_n4368# 0.00809f
C654 passgatex4_0.GP4 A2 1.28e-19
C655 passgatesCtrl_0.net8 passgatex4_0.GN2 0.00108f
C656 passgatex4_0.GP3 A1 2.76e-19
C657 passgatex4_0.GN3 passgatesCtrl_0.net9 0.015603f
C658 passgatex4_0.GP4 a_n2639_n2040# 1.28e-20
C659 VPWR a_n1085_n1429# 0.219592f
C660 passgatesCtrl_0.net1 passgatesCtrl_0.net5 0.088832f
C661 A3 passgatex4_0.GN2 0.00661f
C662 a_n2189_n1429# a_n2883_n1648# 0.002068f
C663 passgatesCtrl_0.net1 a_n715_n3850# 0.224224f
C664 passgatex4_0.GN3 passgatesCtrl_0.net5 0.188564f
C665 passgatex4_0.GP4 passgatesCtrl_0.net6 2.47e-20
C666 passgatex4_0.GP2 passgatex4_0.GN2 1.51461f
C667 passgatesCtrl_0.net7 a_n434_n1942# 5.23e-19
C668 select1 select0 0.083731f
C669 a_n539_n3518# A1 0.002355f
C670 passgatesCtrl_0.net1 a_n2057_n1942# 0.00235f
C671 passgatesCtrl_0._03_ a_n491_n3280# 7.41e-20
C672 a_n491_n3280# passgatex4_0.GP1 0.109714f
C673 a_n1635_n3306# a_n1507_n3280# 0.004764f
C674 passgatesCtrl_0.net7 passgatesCtrl_0._02_ 0.003983f
C675 a_n1913_n1429# passgatesCtrl_0._00_ 2.75e-19
C676 a_n539_n3518# passgatesCtrl_0.net3 6.41e-21
C677 VPWR passgatesCtrl_0.net2 3.00507f
C678 passgatesCtrl_0.net7 passgatesCtrl_0.net8 2.52e-19
C679 passgatesCtrl_0.net1 a_n1878_n4368# 6.03e-19
C680 a_n1173_n2218# passgatesCtrl_0.net5 0.001684f
C681 a_n951_n2736# Z1 1e-20
C682 passgatesCtrl_0.net4 a_n1459_n3306# 0.010474f
C683 passgatesCtrl_0._01_ a_n1637_n1429# 2.78e-19
C684 passgatesCtrl_0.net4 select1 0.003108f
C685 passgatesCtrl_0.net7 a_n2189_n1429# 2.69e-20
C686 a_n715_n3850# a_n995_n3605# 3.02e-19
C687 passgatesCtrl_0.net1 a_n2639_n2040# 0.084866f
C688 a_n1503_n2192# passgatesCtrl_0._02_ 4.67e-20
C689 passgatex4_0.GN3 A2 0.161523f
C690 passgatex4_0.GN4 passgatesCtrl_0.net8 5.26e-19
C691 a_n1503_n2192# passgatesCtrl_0.net8 0.107924f
C692 passgatesCtrl_0._05_ a_n2883_n1648# 6.71e-20
C693 passgatex4_0.GN4 a_n2189_n1429# 2.84e-19
C694 passgatex4_0.GP2 passgatesCtrl_0.net7 3.18e-19
C695 passgatesCtrl_0.net6 passgatesCtrl_0.net1 0.502444f
C696 passgatesCtrl_0.net2 a_n1507_n3280# 5.53e-19
C697 passgatesCtrl_0.net1 a_n1984_n4368# 2.27e-19
C698 passgatex4_0.GN4 A3 0.183073f
C699 passgatesCtrl_0.net5 passgatesCtrl_0.net9 0.011574f
C700 a_n1084_n4216# a_n988_n4394# 0.313533f
C701 VPWR A1 1.84639f
C702 a_n2975_n2192# a_n2883_n1648# 1.44e-19
C703 passgatex4_0.GN3 passgatesCtrl_0.net6 0.151115f
C704 passgatex4_0.GP2 passgatex4_0.GN4 0.041571f
C705 a_n1503_n2192# passgatex4_0.GP2 3.34e-21
C706 VPWR passgatesCtrl_0.net3 0.348944f
C707 passgatex4_0.GP4 a_n1913_n1429# 0.109546f
C708 Z1 a_n675_n1648# 3.24e-20
C709 passgatex4_0.GP4 a_n2429_n1328# 5.08e-19
C710 a_n2015_n2040# passgatesCtrl_0._00_ 1.34e-19
C711 passgatex4_0.GN1 a_n1459_n3306# 4.47e-21
C712 Z3 A2 0.004565f
C713 passgatex4_0.GN1 select1 1.61e-19
C714 A3 Z2 1.49e-20
C715 passgatesCtrl_0.net6 a_n1173_n2218# 2.62e-19
C716 select0 passgatesCtrl_0.net1 0.025769f
C717 a_n1085_n1429# passgatesCtrl_0._02_ 7.02e-19
C718 passgatex4_0.GP2 Z2 0.278333f
C719 passgatex4_0.GN4 passgatesCtrl_0._05_ 3.95e-20
C720 passgatesCtrl_0.net5 a_n2057_n1942# 2.64e-19
C721 a_n1085_n1429# passgatesCtrl_0.net8 0.201804f
C722 passgatesCtrl_0.net9 a_n2639_n2040# 2.03e-19
C723 a_n951_n2736# passgatex4_0.GP1 9.85e-21
C724 passgatesCtrl_0.net4 passgatesCtrl_0.net1 0.142351f
C725 passgatesCtrl_0._00_ a_n2883_n1648# 0.229802f
C726 passgatesCtrl_0.net1 a_n1003_n2040# 0.158092f
C727 passgatesCtrl_0.net2 a_n988_n4394# 7.27e-19
C728 Z1 passgatex4_0.GP1 0.278495f
C729 passgatesCtrl_0.net5 a_n1878_n4368# 3.52e-19
C730 passgatesCtrl_0.net2 a_n434_n1942# 9.54e-19
C731 a_n951_n2736# a_n1227_n2736# 5.3e-19
C732 passgatex4_0.GN1 passgatex4_0.GP4 1.4e-19
C733 a_n1637_n1429# passgatesCtrl_0.net10 0.030972f
C734 VPWR a_n485_n2736# 0.00616f
C735 passgatesCtrl_0._01_ a_n1361_n1429# 1.94e-20
C736 passgatesCtrl_0.net6 passgatesCtrl_0.net9 5.48e-19
C737 passgatesCtrl_0.net2 passgatesCtrl_0._02_ 0.092244f
C738 passgatesCtrl_0.net1 a_n1913_n1429# 0.006122f
C739 passgatex4_0.GP2 a_n1085_n1429# 0.11066f
C740 passgatesCtrl_0.net2 passgatesCtrl_0.net8 0.129f
C741 passgatex4_0.GN3 a_n1913_n1429# 0.034066f
C742 a_n1135_n4368# a_n1227_n2736# 1.17e-20
C743 passgatesCtrl_0.net2 a_n2189_n1429# 3.62e-20
C744 passgatesCtrl_0.net4 a_n995_n3605# 0.110271f
C745 passgatesCtrl_0.net4 a_n1173_n2218# 0.001325f
C746 passgatex4_0.GN3 a_n2429_n1328# 9.54e-20
C747 a_n1003_n2040# a_n995_n3605# 4.27e-20
C748 a_n1173_n2218# a_n1003_n2040# 0.101254f
C749 passgatesCtrl_0.net6 passgatesCtrl_0.net5 0.372649f
C750 passgatesCtrl_0.net5 a_n1984_n4368# 1.71e-19
C751 select1 a_n1963_n3280# 3.96e-19
C752 a_n482_n4216# passgatesCtrl_0.net1 0.167305f
C753 passgatex4_0.GP4 passgatex4_0.GN2 3.27e-19
C754 passgatex4_0.GN4 passgatesCtrl_0._00_ 3.91e-19
C755 a_n988_n4394# A1 1.54e-20
C756 passgatex4_0.GP1 a_n675_n1648# 0.001422f
C757 passgatex4_0.GP2 passgatesCtrl_0.net2 3.91e-20
C758 a_n1503_n2192# passgatesCtrl_0._00_ 5.79e-21
C759 Z4 VGND 2.706298f
C760 A4 VGND 3.775201f
C761 Z3 VGND 2.493104f
C762 A3 VGND 3.16981f
C763 Z2 VGND 2.453408f
C764 A2 VGND 3.285328f
C765 Z1 VGND 2.856037f
C766 A1 VGND 3.713512f
C767 select0 VGND 0.611662f
C768 select1 VGND 1.92417f
C769 VPWR VGND 0.101815p
C770 a_n1135_n4368# VGND 0.171495f
C771 a_n1701_n4368# VGND 0.108493f
C772 a_n482_n4216# VGND 0.309602f
C773 a_n801_n4216# VGND 0.268985f
C774 a_n988_n4394# VGND 0.277513f
C775 a_n1084_n4216# VGND 0.27241f
C776 a_n1878_n4368# VGND 0.260674f
C777 a_n1984_n4368# VGND 0.250918f
C778 a_n2161_n4368# VGND 0.286148f
C779 a_n2480_n4368# VGND 0.328097f
C780 a_n587_n3458# VGND 0.005492f
C781 a_n539_n3518# VGND 0.241098f
C782 a_n715_n3850# VGND 0.229487f
C783 passgatesCtrl_0._04_ VGND 0.264876f
C784 a_n995_n3605# VGND 0.260858f
C785 a_n1507_n3280# VGND 0.005035f
C786 passgatex4_0.GP1 VGND 2.27865f
C787 a_n491_n3280# VGND 0.274026f
C788 a_n1459_n3306# VGND 0.254131f
C789 a_n1635_n3306# VGND 0.235093f
C790 a_n1963_n3280# VGND 0.277418f
C791 passgatesCtrl_0._03_ VGND 0.368268f
C792 a_n485_n2736# VGND 2.19e-19
C793 passgatex4_0.GN2 VGND 4.32804f
C794 passgatex4_0.GN1 VGND 3.99205f
C795 a_n951_n2736# VGND 0.268527f
C796 passgatesCtrl_0.net4 VGND 0.647109f
C797 a_n1227_n2736# VGND 0.2678f
C798 passgatesCtrl_0.net3 VGND 0.42716f
C799 a_n434_n1942# VGND 5.62e-19
C800 a_n1045_n1942# VGND 7.49e-19
C801 a_n1003_n2040# VGND 0.298899f
C802 a_n2465_n2164# VGND 0.005723f
C803 a_n2057_n1942# VGND 8.59e-19
C804 a_n2015_n2040# VGND 0.295323f
C805 a_n597_n2040# VGND 0.234177f
C806 a_n1173_n2218# VGND 0.254047f
C807 a_n1503_n2192# VGND 0.224474f
C808 passgatesCtrl_0._01_ VGND 0.199048f
C809 a_n2185_n2218# VGND 0.267196f
C810 a_n2639_n2040# VGND 0.257089f
C811 a_n2975_n2192# VGND 0.252788f
C812 passgatesCtrl_0._05_ VGND 0.341727f
C813 passgatesCtrl_0.net7 VGND 0.453064f
C814 passgatex4_0.GP2 VGND 2.23556f
C815 passgatex4_0.GN3 VGND 3.82555f
C816 passgatex4_0.GN4 VGND 5.2369f
C817 passgatex4_0.GP4 VGND 5.2081f
C818 passgatex4_0.GP3 VGND 2.17467f
C819 a_n2429_n1328# VGND 0.001779f
C820 a_n675_n1648# VGND 0.258431f
C821 passgatesCtrl_0._02_ VGND 0.366887f
C822 passgatesCtrl_0.net8 VGND 0.333624f
C823 a_n1085_n1429# VGND 0.250109f
C824 passgatesCtrl_0.net5 VGND 0.6309f
C825 a_n1361_n1429# VGND 0.21514f
C826 passgatesCtrl_0.net6 VGND 0.300978f
C827 a_n1637_n1429# VGND 0.2182f
C828 passgatesCtrl_0.net10 VGND -0.162684f
C829 a_n1913_n1429# VGND 0.220816f
C830 passgatesCtrl_0.net9 VGND 0.33083f
C831 a_n2189_n1429# VGND 0.238577f
C832 passgatesCtrl_0.net1 VGND 3.170257f
C833 passgatesCtrl_0.net2 VGND 4.630451f
C834 a_n2883_n1648# VGND 0.241645f
C835 passgatesCtrl_0._00_ VGND 0.297612f
C836 A1.t0 VGND 0.838615f
C837 A1.t1 VGND 0.481433f
C838 A1.n0 VGND 4.66276f
C839 A1.t2 VGND 0.867976f
C840 A1.t3 VGND 0.614013f
C841 A1.n1 VGND 4.76729f
C842 A1.n2 VGND 0.754061f
C843 A1.n3 VGND 0.235366f
C844 Z1.t1 VGND 0.368287f
C845 Z1.n0 VGND 0.549919f
C846 Z1.t0 VGND 0.37568f
C847 Z1.t2 VGND 0.498536f
C848 Z1.n1 VGND 2.51576f
C849 Z1.n2 VGND 0.851227f
C850 Z1.t3 VGND 0.485176f
C851 Z1.n3 VGND 0.603414f
C852 Z1.n4 VGND 0.766774f
C853 A4.t0 VGND 0.893471f
C854 A4.t1 VGND 0.512925f
C855 A4.n0 VGND 4.96776f
C856 A4.t3 VGND 0.924752f
C857 A4.t2 VGND 0.654177f
C858 A4.n1 VGND 5.07912f
C859 A4.n2 VGND 0.803386f
C860 A4.n3 VGND 0.175929f
C861 Z4.t1 VGND 0.356732f
C862 Z4.n0 VGND 0.532664f
C863 Z4.t0 VGND 0.363892f
C864 Z4.t3 VGND 0.482893f
C865 Z4.n1 VGND 2.43682f
C866 Z4.n2 VGND 0.824519f
C867 Z4.t2 VGND 0.469953f
C868 Z4.n3 VGND 0.584481f
C869 Z4.n4 VGND 0.742715f
C870 A2.t3 VGND 0.763965f
C871 A2.t2 VGND 0.438578f
C872 A2.n0 VGND 4.2477f
C873 A2.t0 VGND 0.790712f
C874 A2.t1 VGND 0.559356f
C875 A2.n1 VGND 4.34292f
C876 A2.n2 VGND 0.686937f
C877 A2.n3 VGND 0.222065f
C878 Z2.t2 VGND 0.358466f
C879 Z2.n0 VGND 0.535254f
C880 Z2.t3 VGND 0.365662f
C881 Z2.t0 VGND 0.485241f
C882 Z2.n1 VGND 2.44867f
C883 Z2.n2 VGND 0.828528f
C884 Z2.t1 VGND 0.472238f
C885 Z2.n3 VGND 0.587323f
C886 Z2.n4 VGND 0.723782f
C887 Z2.n5 VGND 0.319875f
C888 Z3.t0 VGND 0.361967f
C889 Z3.n0 VGND 0.540482f
C890 Z3.t1 VGND 0.369233f
C891 Z3.t3 VGND 0.48998f
C892 Z3.n1 VGND 2.47259f
C893 Z3.n2 VGND 0.83662f
C894 Z3.t2 VGND 0.47685f
C895 Z3.n3 VGND 0.593059f
C896 Z3.n4 VGND 0.728589f
C897 Z3.n5 VGND 0.33185f
C898 A3.t0 VGND 0.893706f
C899 A3.t1 VGND 0.51306f
C900 A3.n0 VGND 4.969069f
C901 A3.t3 VGND 0.924996f
C902 A3.t2 VGND 0.654349f
C903 A3.n1 VGND 5.08046f
C904 A3.n2 VGND 0.803598f
C905 A3.n3 VGND 0.264739f
C906 passgatesCtrl_0.net1.n0 VGND 0.226539f
C907 passgatesCtrl_0.net1.t1 VGND 0.053408f
C908 passgatesCtrl_0.net1.n1 VGND 0.014253f
C909 passgatesCtrl_0.net1.t0 VGND 0.033625f
C910 passgatesCtrl_0.net1.n2 VGND 0.02627f
C911 passgatesCtrl_0.net1.t11 VGND 0.01948f
C912 passgatesCtrl_0.net1.t2 VGND 0.013193f
C913 passgatesCtrl_0.net1.n3 VGND 0.052945f
C914 passgatesCtrl_0.net1.n4 VGND 0.021541f
C915 passgatesCtrl_0.net1.n5 VGND 0.027845f
C916 passgatesCtrl_0.net1.t3 VGND 0.015219f
C917 passgatesCtrl_0.net1.t8 VGND 0.024374f
C918 passgatesCtrl_0.net1.n6 VGND 0.046451f
C919 passgatesCtrl_0.net1.n7 VGND 0.05146f
C920 passgatesCtrl_0.net1.t13 VGND 0.016147f
C921 passgatesCtrl_0.net1.t12 VGND 0.011096f
C922 passgatesCtrl_0.net1.n8 VGND 0.046923f
C923 passgatesCtrl_0.net1.n9 VGND 0.01118f
C924 passgatesCtrl_0.net1.n10 VGND 0.021551f
C925 passgatesCtrl_0.net1.n11 VGND 0.171457f
C926 passgatesCtrl_0.net1.t9 VGND 0.022577f
C927 passgatesCtrl_0.net1.t17 VGND 0.052767f
C928 passgatesCtrl_0.net1.n12 VGND 0.058498f
C929 passgatesCtrl_0.net1.n13 VGND 0.193324f
C930 passgatesCtrl_0.net1.t10 VGND 0.010521f
C931 passgatesCtrl_0.net1.t5 VGND 0.012736f
C932 passgatesCtrl_0.net1.n14 VGND 0.042403f
C933 passgatesCtrl_0.net1.n15 VGND 0.009709f
C934 passgatesCtrl_0.net1.t16 VGND 0.010838f
C935 passgatesCtrl_0.net1.t18 VGND 0.013595f
C936 passgatesCtrl_0.net1.n16 VGND 0.030532f
C937 passgatesCtrl_0.net1.t14 VGND 0.015192f
C938 passgatesCtrl_0.net1.t19 VGND 0.024522f
C939 passgatesCtrl_0.net1.n17 VGND 0.049813f
C940 passgatesCtrl_0.net1.n18 VGND 0.013363f
C941 passgatesCtrl_0.net1.n19 VGND 0.13082f
C942 passgatesCtrl_0.net1.t6 VGND 0.019673f
C943 passgatesCtrl_0.net1.t15 VGND 0.013358f
C944 passgatesCtrl_0.net1.n20 VGND 0.046479f
C945 passgatesCtrl_0.net1.n21 VGND 0.011125f
C946 passgatesCtrl_0.net1.n22 VGND 0.054042f
C947 passgatesCtrl_0.net1.n23 VGND 0.220245f
C948 passgatesCtrl_0.net1.t7 VGND 0.022351f
C949 passgatesCtrl_0.net1.t4 VGND 0.010599f
C950 passgatesCtrl_0.net1.n24 VGND 0.080089f
C951 passgatesCtrl_0.net1.n25 VGND 0.01726f
C952 passgatesCtrl_0.net1.n26 VGND 0.016365f
C953 passgatesCtrl_0.net10.t2 VGND -0.055929f
C954 passgatesCtrl_0.net10.t1 VGND -0.028065f
C955 passgatesCtrl_0.net10.t0 VGND -0.028065f
C956 passgatesCtrl_0.net10.n0 VGND -0.063496f
C957 passgatesCtrl_0.net10.t3 VGND -0.027227f
C958 passgatesCtrl_0.net10.t4 VGND -0.043656f
C959 passgatesCtrl_0.net10.n1 VGND -0.087973f
C960 passgatesCtrl_0.net10.n2 VGND -0.035052f
C961 passgatesCtrl_0.net10.n3 VGND -0.16161f
C962 VPWR.n0 VGND 0.115638f
C963 VPWR.n1 VGND 0.176137f
C964 VPWR.n2 VGND 0.115638f
C965 VPWR.n3 VGND 0.104151f
C966 VPWR.n4 VGND 0.003054f
C967 VPWR.n5 VGND 0.003159f
C968 VPWR.n6 VGND 0.001813f
C969 VPWR.n7 VGND 0.001417f
C970 VPWR.t103 VGND 0.278603f
C971 VPWR.t31 VGND 0.021284f
C972 VPWR.t99 VGND 0.029392f
C973 VPWR.t127 VGND 0.28885f
C974 VPWR.t13 VGND 0.021284f
C975 VPWR.t0 VGND 0.045608f
C976 VPWR.t104 VGND 0.110472f
C977 VPWR.n8 VGND 0.135354f
C978 VPWR.n9 VGND 0.015324f
C979 VPWR.t63 VGND 0.004539f
C980 VPWR.n10 VGND 0.01112f
C981 VPWR.n11 VGND 5.46e-19
C982 VPWR.n12 VGND 0.00398f
C983 VPWR.n13 VGND 0.003417f
C984 VPWR.t35 VGND 0.004921f
C985 VPWR.n14 VGND 0.009822f
C986 VPWR.n15 VGND 0.004796f
C987 VPWR.t180 VGND 0.065381f
C988 VPWR.n16 VGND 0.029387f
C989 VPWR.n17 VGND 0.005284f
C990 VPWR.t1 VGND 0.001371f
C991 VPWR.t2 VGND 0.001371f
C992 VPWR.n18 VGND 0.002981f
C993 VPWR.n19 VGND 0.006462f
C994 VPWR.n20 VGND 0.001838f
C995 VPWR.n21 VGND 0.001771f
C996 VPWR.n22 VGND 0.003159f
C997 VPWR.n23 VGND 0.104151f
C998 VPWR.n24 VGND 0.003159f
C999 VPWR.n25 VGND 0.002158f
C1000 VPWR.n26 VGND 0.001417f
C1001 VPWR.n27 VGND 0.001838f
C1002 VPWR.n28 VGND 0.002585f
C1003 VPWR.n29 VGND 0.001417f
C1004 VPWR.n30 VGND 0.001771f
C1005 VPWR.n31 VGND 0.001895f
C1006 VPWR.t155 VGND 6.78e-19
C1007 VPWR.t175 VGND 0.00103f
C1008 VPWR.n32 VGND 0.00172f
C1009 VPWR.n33 VGND 0.002685f
C1010 VPWR.n34 VGND 0.001801f
C1011 VPWR.n35 VGND 0.004842f
C1012 VPWR.t159 VGND 0.001371f
C1013 VPWR.t151 VGND 0.001371f
C1014 VPWR.n36 VGND 0.003045f
C1015 VPWR.n37 VGND 0.005284f
C1016 VPWR.t192 VGND 0.026295f
C1017 VPWR.t100 VGND 0.001371f
C1018 VPWR.t158 VGND 0.001371f
C1019 VPWR.n38 VGND 0.002981f
C1020 VPWR.n39 VGND 0.013419f
C1021 VPWR.t154 VGND 0.001371f
C1022 VPWR.t126 VGND 0.001371f
C1023 VPWR.n40 VGND 0.003045f
C1024 VPWR.n41 VGND 0.008241f
C1025 VPWR.n42 VGND 0.001838f
C1026 VPWR.n43 VGND 0.001771f
C1027 VPWR.n44 VGND 0.003159f
C1028 VPWR.n45 VGND 0.40558f
C1029 VPWR.n46 VGND 0.003054f
C1030 VPWR.n47 VGND 0.003159f
C1031 VPWR.n48 VGND 0.0021f
C1032 VPWR.n49 VGND 0.001417f
C1033 VPWR.n50 VGND 0.002642f
C1034 VPWR.t44 VGND 0.004509f
C1035 VPWR.t193 VGND 0.009569f
C1036 VPWR.n52 VGND 0.024536f
C1037 VPWR.t45 VGND 0.004509f
C1038 VPWR.n53 VGND 0.013365f
C1039 VPWR.n54 VGND 0.001838f
C1040 VPWR.t29 VGND 0.004509f
C1041 VPWR.t189 VGND 0.009569f
C1042 VPWR.n56 VGND 0.024536f
C1043 VPWR.t30 VGND 0.004509f
C1044 VPWR.n57 VGND 0.013365f
C1045 VPWR.n58 VGND 0.001871f
C1046 VPWR.n59 VGND 0.002642f
C1047 VPWR.n60 VGND 0.005284f
C1048 VPWR.t167 VGND 0.00103f
C1049 VPWR.t12 VGND 0.001556f
C1050 VPWR.n61 VGND 0.004648f
C1051 VPWR.t121 VGND 0.001371f
C1052 VPWR.t165 VGND 0.001371f
C1053 VPWR.n62 VGND 0.002981f
C1054 VPWR.t102 VGND 0.00276f
C1055 VPWR.n63 VGND 0.0092f
C1056 VPWR.n64 VGND 0.00313f
C1057 VPWR.t84 VGND 0.001371f
C1058 VPWR.t98 VGND 0.001371f
C1059 VPWR.n65 VGND 0.003045f
C1060 VPWR.n66 VGND 0.004796f
C1061 VPWR.n67 VGND 0.005284f
C1062 VPWR.t109 VGND 0.001055f
C1063 VPWR.t146 VGND 0.001556f
C1064 VPWR.n68 VGND 0.004775f
C1065 VPWR.t10 VGND 0.001371f
C1066 VPWR.t80 VGND 0.001371f
C1067 VPWR.n69 VGND 0.003045f
C1068 VPWR.n70 VGND 0.007905f
C1069 VPWR.n71 VGND 0.001838f
C1070 VPWR.n72 VGND 0.001771f
C1071 VPWR.n73 VGND 0.003159f
C1072 VPWR.n74 VGND 0.003159f
C1073 VPWR.n75 VGND 0.001771f
C1074 VPWR.n76 VGND 0.003159f
C1075 VPWR.t70 VGND 0.001371f
C1076 VPWR.t6 VGND 0.001371f
C1077 VPWR.n77 VGND 0.003045f
C1078 VPWR.n78 VGND 0.007905f
C1079 VPWR.n79 VGND 0.0012f
C1080 VPWR.t148 VGND 0.001371f
C1081 VPWR.t125 VGND 0.001371f
C1082 VPWR.n80 VGND 0.003045f
C1083 VPWR.n81 VGND 0.002642f
C1084 VPWR.n82 VGND 0.001838f
C1085 VPWR.n83 VGND 0.001417f
C1086 VPWR.n84 VGND 0.001417f
C1087 VPWR.n85 VGND 0.001771f
C1088 VPWR.n86 VGND 4.88e-19
C1089 VPWR.n87 VGND 0.002154f
C1090 VPWR.n88 VGND 0.001522f
C1091 VPWR.n89 VGND 0.008241f
C1092 VPWR.t106 VGND 0.002717f
C1093 VPWR.t72 VGND 0.001371f
C1094 VPWR.t68 VGND 0.001371f
C1095 VPWR.n90 VGND 0.003045f
C1096 VPWR.n91 VGND 0.004767f
C1097 VPWR.n92 VGND 0.001536f
C1098 VPWR.n93 VGND 0.005284f
C1099 VPWR.t134 VGND 0.001371f
C1100 VPWR.t92 VGND 0.001371f
C1101 VPWR.n94 VGND 0.003045f
C1102 VPWR.t88 VGND 0.001055f
C1103 VPWR.t119 VGND 0.001556f
C1104 VPWR.n95 VGND 0.004765f
C1105 VPWR.t123 VGND 0.006321f
C1106 VPWR.t90 VGND 0.002709f
C1107 VPWR.n96 VGND 0.005531f
C1108 VPWR.n97 VGND 0.003159f
C1109 VPWR.t115 VGND 0.006322f
C1110 VPWR.t82 VGND 5.06e-19
C1111 VPWR.t113 VGND 0.001358f
C1112 VPWR.n98 VGND 0.006196f
C1113 VPWR.t28 VGND 0.046562f
C1114 VPWR.t107 VGND 0.024382f
C1115 VPWR.t166 VGND 0.024212f
C1116 VPWR.t120 VGND 0.016424f
C1117 VPWR.t11 VGND 0.0149f
C1118 VPWR.t164 VGND 0.021503f
C1119 VPWR.t101 VGND 0.030985f
C1120 VPWR.t83 VGND 0.006603f
C1121 VPWR.t86 VGND 0.013545f
C1122 VPWR.t108 VGND 0.013545f
C1123 VPWR.t97 VGND 0.016593f
C1124 VPWR.t145 VGND 0.026583f
C1125 VPWR.t9 VGND 0.020149f
C1126 VPWR.t79 VGND 0.015577f
C1127 VPWR.t69 VGND 0.015577f
C1128 VPWR.t5 VGND 0.025905f
C1129 VPWR.t147 VGND 0.015408f
C1130 VPWR.t124 VGND 0.031324f
C1131 VPWR.t71 VGND 0.019979f
C1132 VPWR.t67 VGND 0.032509f
C1133 VPWR.t170 VGND 0.026583f
C1134 VPWR.t87 VGND 0.005249f
C1135 VPWR.t133 VGND 0.016593f
C1136 VPWR.t118 VGND 0.0149f
C1137 VPWR.t91 VGND 0.026921f
C1138 VPWR.t122 VGND 0.011344f
C1139 VPWR.t89 VGND 0.014223f
C1140 VPWR.t114 VGND 0.014223f
C1141 VPWR.t112 VGND 0.011852f
C1142 VPWR.t16 VGND 0.046731f
C1143 VPWR.t139 VGND 0.013545f
C1144 VPWR.t77 VGND 0.011006f
C1145 VPWR.t73 VGND 0.015577f
C1146 VPWR.t143 VGND 0.038604f
C1147 VPWR.t81 VGND 0.038991f
C1148 VPWR.n99 VGND 0.001536f
C1149 VPWR.n100 VGND 0.001838f
C1150 VPWR.n101 VGND 0.001771f
C1151 VPWR.n102 VGND 0.003159f
C1152 VPWR.n103 VGND 0.185574f
C1153 VPWR.n104 VGND 0.003159f
C1154 VPWR.n105 VGND 0.001771f
C1155 VPWR.t144 VGND 0.001371f
C1156 VPWR.t74 VGND 0.001371f
C1157 VPWR.n106 VGND 0.003045f
C1158 VPWR.n107 VGND 0.007905f
C1159 VPWR.n108 VGND 0.002642f
C1160 VPWR.n109 VGND 0.001838f
C1161 VPWR.n110 VGND 0.001417f
C1162 VPWR.n111 VGND 0.001417f
C1163 VPWR.n112 VGND 0.001771f
C1164 VPWR.n113 VGND 0.002642f
C1165 VPWR.n114 VGND 4.88e-19
C1166 VPWR.n115 VGND 0.001838f
C1167 VPWR.t78 VGND 0.001371f
C1168 VPWR.t140 VGND 0.001371f
C1169 VPWR.n116 VGND 0.003045f
C1170 VPWR.n117 VGND 0.007905f
C1171 VPWR.t17 VGND 0.004509f
C1172 VPWR.t181 VGND 0.009569f
C1173 VPWR.n119 VGND 0.024536f
C1174 VPWR.t18 VGND 0.004509f
C1175 VPWR.n120 VGND 0.013365f
C1176 VPWR.t53 VGND 0.004509f
C1177 VPWR.t177 VGND 0.009569f
C1178 VPWR.n122 VGND 0.024536f
C1179 VPWR.t54 VGND 0.004509f
C1180 VPWR.n123 VGND 0.013365f
C1181 VPWR.n124 VGND 0.005481f
C1182 VPWR.n125 VGND 0.011299f
C1183 VPWR.n126 VGND 0.001241f
C1184 VPWR.n127 VGND 9.76e-19
C1185 VPWR.n128 VGND 0.002158f
C1186 VPWR.n129 VGND 0.002767f
C1187 VPWR.n130 VGND 0.003054f
C1188 VPWR.n131 VGND 0.197333f
C1189 VPWR.n132 VGND 0.003054f
C1190 VPWR.n133 VGND 0.002767f
C1191 VPWR.n134 VGND 0.001813f
C1192 VPWR.n135 VGND 0.002958f
C1193 VPWR.n136 VGND 0.010251f
C1194 VPWR.n137 VGND 0.006524f
C1195 VPWR.n138 VGND 0.008048f
C1196 VPWR.n139 VGND 9.46e-19
C1197 VPWR.n140 VGND 0.001475f
C1198 VPWR.n141 VGND 0.004796f
C1199 VPWR.n142 VGND 0.00313f
C1200 VPWR.n143 VGND 4.27e-19
C1201 VPWR.n144 VGND 0.007931f
C1202 VPWR.n145 VGND 0.001505f
C1203 VPWR.n146 VGND 0.013321f
C1204 VPWR.n147 VGND 0.004796f
C1205 VPWR.n148 VGND 0.00313f
C1206 VPWR.n149 VGND 0.005284f
C1207 VPWR.n150 VGND 0.001536f
C1208 VPWR.n151 VGND 0.008007f
C1209 VPWR.n152 VGND 0.001795f
C1210 VPWR.n153 VGND 0.001251f
C1211 VPWR.n154 VGND 0.004193f
C1212 VPWR.n155 VGND 0.001871f
C1213 VPWR.n156 VGND 0.002767f
C1214 VPWR.n157 VGND 0.003054f
C1215 VPWR.n158 VGND 0.197333f
C1216 VPWR.n159 VGND 0.003054f
C1217 VPWR.n160 VGND 0.002767f
C1218 VPWR.n161 VGND 0.002646f
C1219 VPWR.n162 VGND 0.003819f
C1220 VPWR.n163 VGND 0.00313f
C1221 VPWR.n164 VGND 0.001282f
C1222 VPWR.n165 VGND 0.007176f
C1223 VPWR.n166 VGND 0.007926f
C1224 VPWR.n167 VGND 0.001536f
C1225 VPWR.n168 VGND 0.001638f
C1226 VPWR.n169 VGND 0.004509f
C1227 VPWR.n170 VGND 0.002671f
C1228 VPWR.n171 VGND 0.00313f
C1229 VPWR.n172 VGND 0.001587f
C1230 VPWR.n173 VGND 0.007309f
C1231 VPWR.n174 VGND 0.006996f
C1232 VPWR.n175 VGND 0.001261f
C1233 VPWR.n176 VGND 0.005284f
C1234 VPWR.n177 VGND 0.004509f
C1235 VPWR.n178 VGND 0.001771f
C1236 VPWR.n179 VGND 0.003159f
C1237 VPWR.n180 VGND 0.001417f
C1238 VPWR.n181 VGND 0.001771f
C1239 VPWR.n182 VGND 0.002767f
C1240 VPWR.n183 VGND 4.92e-19
C1241 VPWR.n184 VGND 0.001838f
C1242 VPWR.n185 VGND 0.001577f
C1243 VPWR.n186 VGND 0.011306f
C1244 VPWR.n187 VGND 0.001838f
C1245 VPWR.n188 VGND 0.001895f
C1246 VPWR.n189 VGND 0.001771f
C1247 VPWR.n190 VGND 0.002767f
C1248 VPWR.n191 VGND 0.003054f
C1249 VPWR.n192 VGND 0.237185f
C1250 VPWR.n193 VGND 0.176137f
C1251 VPWR.n194 VGND 0.384936f
C1252 VPWR.n195 VGND 0.145773f
C1253 VPWR.n196 VGND 0.003159f
C1254 VPWR.n197 VGND 0.0021f
C1255 VPWR.n198 VGND 0.001417f
C1256 VPWR.n199 VGND 0.001417f
C1257 VPWR.n200 VGND 0.001771f
C1258 VPWR.n201 VGND 0.002642f
C1259 VPWR.t32 VGND 0.004509f
C1260 VPWR.t182 VGND 0.009569f
C1261 VPWR.n203 VGND 0.024536f
C1262 VPWR.t33 VGND 0.004509f
C1263 VPWR.n204 VGND 0.013365f
C1264 VPWR.n205 VGND 0.002642f
C1265 VPWR.n206 VGND 0.001838f
C1266 VPWR.t61 VGND 0.004509f
C1267 VPWR.t188 VGND 0.009569f
C1268 VPWR.n208 VGND 0.024536f
C1269 VPWR.t62 VGND 0.004509f
C1270 VPWR.n209 VGND 0.013365f
C1271 VPWR.n210 VGND 0.001241f
C1272 VPWR.n211 VGND 0.011306f
C1273 VPWR.n212 VGND 0.001838f
C1274 VPWR.n213 VGND 0.001895f
C1275 VPWR.n214 VGND 0.001771f
C1276 VPWR.n215 VGND 0.002767f
C1277 VPWR.n216 VGND 0.003054f
C1278 VPWR.n217 VGND 0.114872f
C1279 VPWR.n218 VGND 0.003054f
C1280 VPWR.n219 VGND 0.002767f
C1281 VPWR.n220 VGND 3.49e-19
C1282 VPWR.n221 VGND 0.002814f
C1283 VPWR.n222 VGND 0.002613f
C1284 VPWR.n223 VGND 0.001333f
C1285 VPWR.t160 VGND 0.006334f
C1286 VPWR.n224 VGND 0.010785f
C1287 VPWR.t55 VGND 0.004472f
C1288 VPWR.n225 VGND 0.007877f
C1289 VPWR.n226 VGND 0.00348f
C1290 VPWR.n227 VGND 0.002642f
C1291 VPWR.n228 VGND 0.002498f
C1292 VPWR.n229 VGND 0.004939f
C1293 VPWR.n230 VGND 0.013871f
C1294 VPWR.n231 VGND 0.019633f
C1295 VPWR.t56 VGND 0.004472f
C1296 VPWR.n232 VGND 0.007877f
C1297 VPWR.n233 VGND 0.035693f
C1298 VPWR.n234 VGND 0.00313f
C1299 VPWR.n235 VGND 0.004796f
C1300 VPWR.n236 VGND 0.002987f
C1301 VPWR.n237 VGND 0.008233f
C1302 VPWR.n238 VGND 0.00118f
C1303 VPWR.n239 VGND 0.002786f
C1304 VPWR.n240 VGND 0.002642f
C1305 VPWR.n241 VGND 0.001085f
C1306 VPWR.n242 VGND 0.001024f
C1307 VPWR.t34 VGND 0.004921f
C1308 VPWR.n243 VGND 0.003786f
C1309 VPWR.n244 VGND 0.006238f
C1310 VPWR.n245 VGND 0.005553f
C1311 VPWR.n246 VGND 0.005274f
C1312 VPWR.t105 VGND 9.3e-19
C1313 VPWR.t128 VGND 0.003822f
C1314 VPWR.n247 VGND 0.003518f
C1315 VPWR.n248 VGND 0.002638f
C1316 VPWR.n249 VGND 0.005017f
C1317 VPWR.n250 VGND 0.005583f
C1318 VPWR.n251 VGND 0.001838f
C1319 VPWR.n252 VGND 0.002642f
C1320 VPWR.n253 VGND 0.001771f
C1321 VPWR.n254 VGND 0.002767f
C1322 VPWR.n255 VGND 0.003054f
C1323 VPWR.n256 VGND 0.114872f
C1324 VPWR.n257 VGND 0.003054f
C1325 VPWR.n258 VGND 0.002767f
C1326 VPWR.n259 VGND 0.002646f
C1327 VPWR.n260 VGND 0.004193f
C1328 VPWR.n261 VGND 0.005284f
C1329 VPWR.n262 VGND 0.00666f
C1330 VPWR.n263 VGND 0.012423f
C1331 VPWR.n264 VGND 0.005301f
C1332 VPWR.n265 VGND 0.00313f
C1333 VPWR.n266 VGND 0.002642f
C1334 VPWR.n267 VGND 0.006595f
C1335 VPWR.t14 VGND 0.004472f
C1336 VPWR.n268 VGND 0.010271f
C1337 VPWR.n269 VGND 0.018051f
C1338 VPWR.n270 VGND 0.018051f
C1339 VPWR.n271 VGND 0.005284f
C1340 VPWR.n272 VGND 0.005284f
C1341 VPWR.n273 VGND 0.006545f
C1342 VPWR.n274 VGND 0.01473f
C1343 VPWR.t186 VGND 0.033554f
C1344 VPWR.n275 VGND 0.056186f
C1345 VPWR.t15 VGND 0.004472f
C1346 VPWR.n276 VGND 0.011514f
C1347 VPWR.n277 VGND 0.019201f
C1348 VPWR.t46 VGND 0.004509f
C1349 VPWR.t196 VGND 0.009569f
C1350 VPWR.n279 VGND 0.024536f
C1351 VPWR.t47 VGND 0.004509f
C1352 VPWR.n280 VGND 0.012134f
C1353 VPWR.t191 VGND 0.018664f
C1354 VPWR.n281 VGND 0.016882f
C1355 VPWR.n282 VGND 0.002154f
C1356 VPWR.n283 VGND 0.006059f
C1357 VPWR.t64 VGND 0.004472f
C1358 VPWR.n284 VGND 0.004409f
C1359 VPWR.t57 VGND 0.004509f
C1360 VPWR.t194 VGND 0.009569f
C1361 VPWR.n286 VGND 0.024536f
C1362 VPWR.t58 VGND 0.004509f
C1363 VPWR.n287 VGND 0.013365f
C1364 VPWR.t39 VGND 0.004509f
C1365 VPWR.t176 VGND 0.009569f
C1366 VPWR.n289 VGND 0.024536f
C1367 VPWR.t40 VGND 0.004509f
C1368 VPWR.n290 VGND 0.013365f
C1369 VPWR.n291 VGND 0.011265f
C1370 VPWR.n292 VGND 0.004909f
C1371 VPWR.n293 VGND 0.006786f
C1372 VPWR.n294 VGND 0.002474f
C1373 VPWR.n295 VGND 0.001771f
C1374 VPWR.n296 VGND 0.003159f
C1375 VPWR.n297 VGND 0.001417f
C1376 VPWR.n298 VGND 0.002767f
C1377 VPWR.n299 VGND 0.001771f
C1378 VPWR.n300 VGND 0.00201f
C1379 VPWR.n301 VGND 0.001838f
C1380 VPWR.n302 VGND 0.014674f
C1381 VPWR.n303 VGND 0.011685f
C1382 VPWR.n304 VGND 0.00135f
C1383 VPWR.n305 VGND 0.002154f
C1384 VPWR.n306 VGND 0.001771f
C1385 VPWR.n307 VGND 0.002767f
C1386 VPWR.n308 VGND 0.003054f
C1387 VPWR.n309 VGND 0.114872f
C1388 VPWR.n311 VGND 0.00308f
C1389 VPWR.n312 VGND 0.003159f
C1390 VPWR.n313 VGND 0.001771f
C1391 VPWR.n314 VGND 0.00201f
C1392 VPWR.n315 VGND 0.006059f
C1393 VPWR.t36 VGND 0.045885f
C1394 VPWR.t110 VGND 0.011175f
C1395 VPWR.t161 VGND 0.016593f
C1396 VPWR.t152 VGND 0.016085f
C1397 VPWR.t141 VGND 0.0149f
C1398 VPWR.t7 VGND 0.037927f
C1399 VPWR.t173 VGND 0.030138f
C1400 VPWR.t137 VGND 0.016085f
C1401 VPWR.t75 VGND 0.026583f
C1402 VPWR.t95 VGND 0.019641f
C1403 VPWR.t131 VGND 0.0149f
C1404 VPWR.t3 VGND 0.016085f
C1405 VPWR.t156 VGND 0.026583f
C1406 VPWR.t50 VGND 0.060277f
C1407 VPWR.t22 VGND 0.022858f
C1408 VPWR.t168 VGND 0.032001f
C1409 VPWR.t93 VGND 0.047917f
C1410 VPWR.t129 VGND 0.047917f
C1411 VPWR.t116 VGND 0.040297f
C1412 VPWR.t149 VGND 0.020487f
C1413 VPWR.t25 VGND 0.016085f
C1414 VPWR.t135 VGND 0.027091f
C1415 VPWR.t41 VGND 0.072976f
C1416 VPWR.t19 VGND 0.075007f
C1417 VPWR.n316 VGND 0.036145f
C1418 VPWR.n317 VGND 0.019586f
C1419 VPWR.t48 VGND 0.004472f
C1420 VPWR.t197 VGND 0.018829f
C1421 VPWR.n319 VGND 0.032712f
C1422 VPWR.t49 VGND 0.004472f
C1423 VPWR.n320 VGND 0.01877f
C1424 VPWR.n321 VGND 0.001838f
C1425 VPWR.n322 VGND 0.001838f
C1426 VPWR.n323 VGND 0.005284f
C1427 VPWR.t184 VGND 0.018664f
C1428 VPWR.t150 VGND 0.002858f
C1429 VPWR.t136 VGND 8.29e-19
C1430 VPWR.n324 VGND 0.00309f
C1431 VPWR.t26 VGND 0.004472f
C1432 VPWR.n325 VGND 0.007877f
C1433 VPWR.n326 VGND 0.005284f
C1434 VPWR.t130 VGND 0.002858f
C1435 VPWR.t117 VGND 8.29e-19
C1436 VPWR.n327 VGND 0.00309f
C1437 VPWR.n328 VGND 0.00666f
C1438 VPWR.n329 VGND 0.005284f
C1439 VPWR.t185 VGND 0.065173f
C1440 VPWR.t169 VGND 0.002858f
C1441 VPWR.t94 VGND 8.29e-19
C1442 VPWR.n330 VGND 0.00309f
C1443 VPWR.n331 VGND 0.006347f
C1444 VPWR.n332 VGND 0.001771f
C1445 VPWR.n333 VGND 0.003159f
C1446 VPWR.n334 VGND 0.001417f
C1447 VPWR.n335 VGND 0.002642f
C1448 VPWR.t187 VGND 0.018664f
C1449 VPWR.n336 VGND 0.018051f
C1450 VPWR.n337 VGND 0.002787f
C1451 VPWR.n338 VGND 0.002817f
C1452 VPWR.n339 VGND 0.005284f
C1453 VPWR.t162 VGND 8.29e-19
C1454 VPWR.t142 VGND 0.002858f
C1455 VPWR.n340 VGND 0.00309f
C1456 VPWR.n341 VGND 0.00481f
C1457 VPWR.t111 VGND 6.78e-19
C1458 VPWR.t153 VGND 0.00103f
C1459 VPWR.n342 VGND 0.001759f
C1460 VPWR.t65 VGND 0.004509f
C1461 VPWR.t190 VGND 0.009569f
C1462 VPWR.n344 VGND 0.024536f
C1463 VPWR.t66 VGND 0.004509f
C1464 VPWR.n345 VGND 0.013365f
C1465 VPWR.t37 VGND 0.004509f
C1466 VPWR.t195 VGND 0.009569f
C1467 VPWR.n347 VGND 0.024536f
C1468 VPWR.t38 VGND 0.004509f
C1469 VPWR.n348 VGND 0.013365f
C1470 VPWR.n349 VGND 0.011306f
C1471 VPWR.n350 VGND 0.002642f
C1472 VPWR.n351 VGND 0.001771f
C1473 VPWR.n352 VGND 0.003159f
C1474 VPWR.n353 VGND 0.001417f
C1475 VPWR.n354 VGND 0.0021f
C1476 VPWR.n355 VGND 0.003054f
C1477 VPWR.n356 VGND 0.002767f
C1478 VPWR.n357 VGND 0.001771f
C1479 VPWR.n358 VGND 0.001895f
C1480 VPWR.n359 VGND 0.001838f
C1481 VPWR.n360 VGND 0.001838f
C1482 VPWR.n361 VGND 0.002642f
C1483 VPWR.n362 VGND 0.001771f
C1484 VPWR.n363 VGND 0.001417f
C1485 VPWR.n364 VGND 0.003159f
C1486 VPWR.n365 VGND 0.003054f
C1487 VPWR.n366 VGND 0.002767f
C1488 VPWR.n367 VGND 3.49e-19
C1489 VPWR.n368 VGND 0.001838f
C1490 VPWR.n369 VGND 0.001556f
C1491 VPWR.n370 VGND 0.00444f
C1492 VPWR.n371 VGND 4.17e-19
C1493 VPWR.n372 VGND 0.004796f
C1494 VPWR.n373 VGND 0.005284f
C1495 VPWR.n374 VGND 0.001368f
C1496 VPWR.n375 VGND 0.002831f
C1497 VPWR.n376 VGND 0.002987f
C1498 VPWR.t8 VGND 9.3e-19
C1499 VPWR.n377 VGND 0.002638f
C1500 VPWR.t138 VGND 0.003822f
C1501 VPWR.n378 VGND 0.003518f
C1502 VPWR.n379 VGND 0.00314f
C1503 VPWR.t174 VGND 8.29e-19
C1504 VPWR.t76 VGND 0.002858f
C1505 VPWR.n380 VGND 0.003049f
C1506 VPWR.n381 VGND 0.003043f
C1507 VPWR.n382 VGND 0.002625f
C1508 VPWR.n383 VGND 0.005284f
C1509 VPWR.n384 VGND 0.005284f
C1510 VPWR.n385 VGND 0.00313f
C1511 VPWR.n386 VGND 0.001434f
C1512 VPWR.t96 VGND 0.001371f
C1513 VPWR.t4 VGND 0.001371f
C1514 VPWR.n387 VGND 0.003045f
C1515 VPWR.t132 VGND 8.29e-19
C1516 VPWR.t157 VGND 0.002858f
C1517 VPWR.n388 VGND 0.003049f
C1518 VPWR.n389 VGND 0.002437f
C1519 VPWR.n390 VGND 0.008432f
C1520 VPWR.n391 VGND 0.004796f
C1521 VPWR.n392 VGND 0.005284f
C1522 VPWR.n393 VGND 0.00313f
C1523 VPWR.n394 VGND 0.002697f
C1524 VPWR.t23 VGND 0.004921f
C1525 VPWR.n395 VGND 0.003542f
C1526 VPWR.t51 VGND 0.004472f
C1527 VPWR.n396 VGND 0.010271f
C1528 VPWR.n397 VGND 0.007784f
C1529 VPWR.n398 VGND 0.002642f
C1530 VPWR.n399 VGND 0.003819f
C1531 VPWR.n400 VGND 0.001771f
C1532 VPWR.n401 VGND 0.003054f
C1533 VPWR.n402 VGND 0.002767f
C1534 VPWR.n403 VGND 0.002646f
C1535 VPWR.n404 VGND 0.001838f
C1536 VPWR.n405 VGND 0.013995f
C1537 VPWR.n406 VGND 0.01912f
C1538 VPWR.t52 VGND 0.004472f
C1539 VPWR.n407 VGND 0.005606f
C1540 VPWR.n408 VGND 0.008033f
C1541 VPWR.n409 VGND 0.001838f
C1542 VPWR.n410 VGND 0.001091f
C1543 VPWR.n411 VGND 0.002585f
C1544 VPWR.n412 VGND 0.001895f
C1545 VPWR.n413 VGND 0.001771f
C1546 VPWR.n414 VGND 0.001417f
C1547 VPWR.n415 VGND 0.003159f
C1548 VPWR.n416 VGND 0.003054f
C1549 VPWR.n417 VGND 0.001443f
C1550 VPWR.n418 VGND 3.54e-19
C1551 VPWR.n419 VGND 0.002297f
C1552 VPWR.n420 VGND 0.004193f
C1553 VPWR.n421 VGND 0.00666f
C1554 VPWR.n422 VGND 0.003475f
C1555 VPWR.n423 VGND 0.005431f
C1556 VPWR.n424 VGND 0.030297f
C1557 VPWR.n425 VGND 0.005103f
C1558 VPWR.n426 VGND 0.005284f
C1559 VPWR.n427 VGND 0.005284f
C1560 VPWR.n428 VGND 0.005284f
C1561 VPWR.n429 VGND 0.003728f
C1562 VPWR.n430 VGND 0.006987f
C1563 VPWR.t24 VGND 0.004921f
C1564 VPWR.n431 VGND 0.003424f
C1565 VPWR.n432 VGND 0.002582f
C1566 VPWR.n433 VGND 0.005198f
C1567 VPWR.n434 VGND 0.00313f
C1568 VPWR.n435 VGND 0.004796f
C1569 VPWR.n436 VGND 0.010554f
C1570 VPWR.n437 VGND 0.01081f
C1571 VPWR.n438 VGND 0.006332f
C1572 VPWR.n439 VGND 0.016882f
C1573 VPWR.t27 VGND 0.004472f
C1574 VPWR.n440 VGND 0.004409f
C1575 VPWR.n441 VGND 0.004909f
C1576 VPWR.n442 VGND 0.003274f
C1577 VPWR.n443 VGND 0.002843f
C1578 VPWR.n444 VGND 0.001813f
C1579 VPWR.n445 VGND 0.002741f
C1580 VPWR.n446 VGND 0.001417f
C1581 VPWR.n447 VGND 0.002642f
C1582 VPWR.n448 VGND 0.001771f
C1583 VPWR.n449 VGND 0.003159f
C1584 VPWR.n450 VGND 0.001417f
C1585 VPWR.n451 VGND 0.001771f
C1586 VPWR.n452 VGND 0.002154f
C1587 VPWR.n453 VGND 5.46e-19
C1588 VPWR.t20 VGND 0.004472f
C1589 VPWR.t179 VGND 0.018829f
C1590 VPWR.n455 VGND 0.032712f
C1591 VPWR.t21 VGND 0.004472f
C1592 VPWR.n456 VGND 0.01877f
C1593 VPWR.t42 VGND 0.004509f
C1594 VPWR.t178 VGND 0.009569f
C1595 VPWR.n458 VGND 0.024536f
C1596 VPWR.t43 VGND 0.004509f
C1597 VPWR.n459 VGND 0.013365f
C1598 VPWR.t59 VGND 0.004509f
C1599 VPWR.t183 VGND 0.009569f
C1600 VPWR.n461 VGND 0.024536f
C1601 VPWR.t60 VGND 0.004509f
C1602 VPWR.n462 VGND 0.013365f
C1603 VPWR.n463 VGND 0.011004f
C1604 VPWR.n464 VGND 0.015879f
C1605 VPWR.n465 VGND 0.006786f
C1606 VPWR.n466 VGND 0.002474f
C1607 VPWR.n467 VGND 0.002741f
C1608 VPWR.n468 VGND 0.00308f
C1609 VPWR.n469 VGND 0.115638f
C1610 VPWR.n470 VGND 0.026229f
C1611 VPWR.n471 VGND 0.075814f
C1612 VPWR.n472 VGND 0.360185f
C1613 VPWR.n473 VGND 0.075814f
C1614 VPWR.n474 VGND 0.026229f
C1615 VPWR.n475 VGND 0.384936f
C1616 VPWR.n476 VGND 0.067851f
C1617 VPWR.n477 VGND 0.075814f
C1618 VPWR.n478 VGND 0.122169f
C1619 VPWR.n479 VGND 0.100437f
C1620 VPWR.n480 VGND 1.93e-19
C1621 VPWR.n481 VGND 0.032316f
C1622 VPWR.n482 VGND 0.060473f
C1623 VPWR.n483 VGND 0.068782f
C1624 VPWR.n484 VGND 0.050377f
C1625 VPWR.t171 VGND 0.555684f
C1626 VPWR.n485 VGND 0.102743f
C1627 VPWR.n487 VGND 0.417917f
C1628 VPWR.n488 VGND 0.050377f
C1629 VPWR.n490 VGND 0.417917f
C1630 VPWR.n491 VGND 0.049622f
C1631 VPWR.n492 VGND 0.030592f
C1632 VPWR.n493 VGND 0.005583f
C1633 VPWR.n494 VGND 0.005464f
C1634 VPWR.n495 VGND 0.082022f
C1635 VPWR.n496 VGND 0.050682f
C1636 VPWR.n497 VGND 0.030459f
C1637 VPWR.n498 VGND 0.005613f
C1638 VPWR.n499 VGND 0.417917f
C1639 VPWR.n500 VGND 0.417917f
C1640 VPWR.n501 VGND 0.049622f
C1641 VPWR.n502 VGND 0.032078f
C1642 VPWR.n503 VGND 0.060473f
C1643 VPWR.n504 VGND 0.102743f
C1644 VPWR.n505 VGND 0.068782f
C1645 VPWR.n506 VGND 0.050377f
C1646 VPWR.t85 VGND 0.555684f
C1647 VPWR.n509 VGND 0.050377f
C1648 VPWR.n510 VGND 0.00177f
C1649 VPWR.n511 VGND 0.004f
C1650 VPWR.n512 VGND 0.074678f
C1651 VPWR.n513 VGND 0.051989f
C1652 VPWR.n514 VGND 0.030561f
C1653 VPWR.n515 VGND 0.005613f
C1654 VPWR.n516 VGND 0.417917f
C1655 VPWR.n517 VGND 0.417917f
C1656 VPWR.n518 VGND 0.049622f
C1657 VPWR.n519 VGND 0.032078f
C1658 VPWR.n520 VGND 0.060473f
C1659 VPWR.n521 VGND 0.102743f
C1660 VPWR.n522 VGND 0.068782f
C1661 VPWR.n523 VGND 0.050377f
C1662 VPWR.t172 VGND 0.555684f
C1663 VPWR.n526 VGND 0.050377f
C1664 VPWR.n527 VGND 0.001668f
C1665 VPWR.n528 VGND 0.003994f
C1666 VPWR.n529 VGND 0.076174f
C1667 VPWR.n530 VGND 0.06566f
C1668 VPWR.n531 VGND 0.102743f
C1669 VPWR.n532 VGND 0.023085f
C1670 VPWR.n533 VGND 0.049622f
C1671 VPWR.n534 VGND 0.417917f
C1672 VPWR.n535 VGND 0.417917f
C1673 VPWR.n536 VGND 0.068782f
C1674 VPWR.n537 VGND 0.050377f
C1675 VPWR.t163 VGND 0.555684f
C1676 VPWR.n540 VGND 0.050377f
C1677 VPWR.n541 VGND 2.14e-19
C1678 VPWR.n542 VGND 0.030592f
C1679 VPWR.n543 VGND 0.005562f
C1680 VPWR.n544 VGND 0.060473f
C1681 VPWR.n545 VGND 0.032334f
C1682 passgatesCtrl_0.net2.n0 VGND 0.241262f
C1683 passgatesCtrl_0.net2.t0 VGND 0.052358f
C1684 passgatesCtrl_0.net2.n1 VGND 0.013973f
C1685 passgatesCtrl_0.net2.t3 VGND 0.019097f
C1686 passgatesCtrl_0.net2.t7 VGND 0.012934f
C1687 passgatesCtrl_0.net2.n2 VGND 0.052064f
C1688 passgatesCtrl_0.net2.t1 VGND 0.032964f
C1689 passgatesCtrl_0.net2.n3 VGND 0.011845f
C1690 passgatesCtrl_0.net2.n4 VGND 0.031329f
C1691 passgatesCtrl_0.net2.t6 VGND 0.022133f
C1692 passgatesCtrl_0.net2.t15 VGND 0.05173f
C1693 passgatesCtrl_0.net2.n5 VGND 0.062148f
C1694 passgatesCtrl_0.net2.t10 VGND 0.014926f
C1695 passgatesCtrl_0.net2.t19 VGND 0.023903f
C1696 passgatesCtrl_0.net2.n6 VGND 0.04516f
C1697 passgatesCtrl_0.net2.n7 VGND 0.063372f
C1698 passgatesCtrl_0.net2.t16 VGND 0.010242f
C1699 passgatesCtrl_0.net2.t2 VGND 0.012844f
C1700 passgatesCtrl_0.net2.n8 VGND 0.047082f
C1701 passgatesCtrl_0.net2.n9 VGND 0.216971f
C1702 passgatesCtrl_0.net2.n10 VGND 0.157732f
C1703 passgatesCtrl_0.net2.t17 VGND 0.010314f
C1704 passgatesCtrl_0.net2.t9 VGND 0.012486f
C1705 passgatesCtrl_0.net2.n11 VGND 0.041569f
C1706 passgatesCtrl_0.net2.n12 VGND 0.009518f
C1707 passgatesCtrl_0.net2.t12 VGND 0.016063f
C1708 passgatesCtrl_0.net2.t8 VGND 0.011059f
C1709 passgatesCtrl_0.net2.n13 VGND 0.038188f
C1710 passgatesCtrl_0.net2.n14 VGND 0.010881f
C1711 passgatesCtrl_0.net2.t4 VGND 0.014893f
C1712 passgatesCtrl_0.net2.t11 VGND 0.023864f
C1713 passgatesCtrl_0.net2.n15 VGND 0.047068f
C1714 passgatesCtrl_0.net2.n16 VGND 0.061051f
C1715 passgatesCtrl_0.net2.n17 VGND 0.168444f
C1716 passgatesCtrl_0.net2.t18 VGND 0.01039f
C1717 passgatesCtrl_0.net2.t14 VGND 0.021912f
C1718 passgatesCtrl_0.net2.n18 VGND 0.078683f
C1719 passgatesCtrl_0.net2.n19 VGND 0.017108f
C1720 passgatesCtrl_0.net2.n20 VGND 0.16814f
C1721 passgatesCtrl_0.net2.t5 VGND 0.013096f
C1722 passgatesCtrl_0.net2.t13 VGND 0.019286f
C1723 passgatesCtrl_0.net2.n21 VGND 0.045566f
C1724 passgatesCtrl_0.net2.n22 VGND 0.010906f
C1725 passgatesCtrl_0.net2.n23 VGND 0.364405f
C1726 passgatesCtrl_0.net2.n24 VGND 0.041229f
.ends

