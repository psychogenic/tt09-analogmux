magic
tech sky130A
magscale 1 2
timestamp 1728289486
<< locali >>
rect 1344 -3944 1452 -3942
<< viali >>
rect 1520 -3138 1566 -3096
rect 1526 -3246 1562 -3138
rect 1790 -3252 1836 -3108
rect 1140 -3340 1204 -3296
rect 1250 -3344 1296 -3284
rect 1418 -3342 1480 -3294
rect 1690 -3342 1756 -3294
rect 1812 -3342 1862 -3294
rect 1239 -3677 1273 -3643
rect 768 -3906 816 -3678
rect 1786 -3712 1832 -3652
rect 952 -3820 1006 -3774
rect 1080 -3822 1190 -3778
rect 1680 -3834 1732 -3718
rect 2232 -3874 2284 -3734
rect 2426 -3832 2474 -3656
rect 2608 -3820 2662 -3776
rect 2724 -3838 2846 -3774
rect 1344 -3942 1452 -3890
rect 1898 -3934 2006 -3890
rect 1148 -4328 1184 -4204
rect 1324 -4334 1380 -4194
rect 1598 -4334 1650 -4196
rect 1966 -4336 2022 -4214
rect 1234 -4426 1298 -4382
rect 1516 -4428 1568 -4384
rect 1880 -4430 1940 -4382
rect 2148 -4430 2206 -4382
rect 1146 -4564 1186 -4484
rect 1968 -4558 2022 -4492
rect 2254 -4542 2302 -4388
<< metal1 >>
rect 792 -3050 802 -2984
rect 2046 -3050 2056 -2984
rect 2134 -3048 2144 -2972
rect 2214 -3048 2224 -2972
rect 2326 -2980 2576 -2966
rect 2326 -3060 2526 -2980
rect 2590 -3060 2600 -2980
rect 1508 -3096 1578 -3090
rect 1508 -3138 1520 -3096
rect 1566 -3138 1578 -3096
rect 1784 -3102 1842 -3096
rect 1784 -3108 2610 -3102
rect 1784 -3120 1790 -3108
rect 1508 -3144 1526 -3138
rect 828 -3156 898 -3154
rect 674 -3162 1481 -3156
rect 674 -3214 787 -3162
rect 839 -3214 1481 -3162
rect 674 -3222 1481 -3214
rect 1246 -3272 1290 -3260
rect 1244 -3284 1302 -3272
rect 670 -3290 1212 -3286
rect 670 -3292 1216 -3290
rect 670 -3350 942 -3292
rect 1000 -3296 1216 -3292
rect 1000 -3340 1140 -3296
rect 1204 -3340 1216 -3296
rect 1000 -3346 1216 -3340
rect 1244 -3344 1250 -3284
rect 1000 -3350 1212 -3346
rect 670 -3352 1212 -3350
rect 1244 -3352 1254 -3344
rect 1322 -3352 1332 -3284
rect 1415 -3288 1481 -3222
rect 1520 -3246 1526 -3144
rect 1562 -3144 1578 -3138
rect 1562 -3186 1574 -3144
rect 1520 -3258 1532 -3246
rect 1406 -3294 1492 -3288
rect 1406 -3342 1418 -3294
rect 1480 -3342 1492 -3294
rect 1406 -3348 1492 -3342
rect 1522 -3348 1532 -3258
rect 1592 -3348 1602 -3186
rect 1776 -3252 1790 -3120
rect 1836 -3144 2610 -3108
rect 1836 -3252 1880 -3144
rect 1776 -3254 1880 -3252
rect 1784 -3264 1874 -3254
rect 1678 -3294 1768 -3288
rect 1678 -3342 1690 -3294
rect 1756 -3342 1768 -3294
rect 1678 -3348 1768 -3342
rect 1800 -3294 1874 -3264
rect 1800 -3342 1812 -3294
rect 1862 -3342 1874 -3294
rect 1800 -3348 1874 -3342
rect 1244 -3356 1302 -3352
rect 1246 -3362 1290 -3356
rect 1685 -3400 1751 -3348
rect 666 -3466 1751 -3400
rect 1126 -3592 1136 -3522
rect 1198 -3592 1208 -3522
rect 1610 -3590 1620 -3524
rect 2108 -3590 2118 -3524
rect 2246 -3592 2256 -3526
rect 2490 -3592 2500 -3526
rect 2694 -3590 2704 -3528
rect 2762 -3590 2772 -3528
rect 1227 -3640 1285 -3637
rect 1226 -3642 1285 -3640
rect 1392 -3642 1398 -3634
rect 1226 -3643 1398 -3642
rect 762 -3678 822 -3666
rect 762 -3680 768 -3678
rect 740 -3686 768 -3680
rect 702 -3904 712 -3686
rect 766 -3904 768 -3686
rect 762 -3906 768 -3904
rect 816 -3906 822 -3678
rect 1226 -3677 1239 -3643
rect 1273 -3677 1398 -3643
rect 1226 -3678 1398 -3677
rect 1226 -3680 1285 -3678
rect 1227 -3683 1285 -3680
rect 1392 -3686 1398 -3678
rect 1450 -3686 1456 -3634
rect 1780 -3652 1838 -3640
rect 1520 -3668 1530 -3664
rect 1518 -3714 1530 -3668
rect 956 -3720 1530 -3714
rect 1594 -3720 1604 -3664
rect 1670 -3718 1682 -3698
rect 956 -3742 1602 -3720
rect 956 -3768 1018 -3742
rect 940 -3774 1018 -3768
rect 940 -3820 952 -3774
rect 1006 -3820 1018 -3774
rect 1060 -3772 1200 -3770
rect 1060 -3777 1202 -3772
rect 1233 -3777 1239 -3776
rect 940 -3826 1018 -3820
rect 1057 -3778 1239 -3777
rect 1057 -3822 1080 -3778
rect 1190 -3822 1239 -3778
rect 1057 -3827 1239 -3822
rect 1060 -3828 1202 -3827
rect 1233 -3828 1239 -3827
rect 1291 -3828 1297 -3776
rect 1670 -3834 1680 -3718
rect 1734 -3750 1742 -3698
rect 1780 -3712 1786 -3652
rect 1832 -3668 1838 -3652
rect 2420 -3656 2480 -3644
rect 2420 -3660 2426 -3656
rect 2474 -3660 2480 -3656
rect 1832 -3712 1870 -3668
rect 1780 -3720 1870 -3712
rect 1922 -3720 1948 -3668
rect 1780 -3724 1838 -3720
rect 2226 -3726 2290 -3722
rect 1732 -3834 1742 -3750
rect 2222 -3734 2298 -3726
rect 1772 -3814 1778 -3762
rect 1830 -3767 1836 -3762
rect 2222 -3767 2232 -3734
rect 1830 -3809 2232 -3767
rect 1830 -3814 1836 -3809
rect 1670 -3838 1742 -3834
rect 1674 -3846 1738 -3838
rect 1332 -3888 1466 -3882
rect 1908 -3884 1996 -3864
rect 2222 -3874 2232 -3809
rect 2284 -3874 2298 -3734
rect 2418 -3832 2426 -3660
rect 2418 -3836 2428 -3832
rect 2496 -3836 2506 -3660
rect 2596 -3772 2674 -3770
rect 2594 -3776 2674 -3772
rect 2712 -3774 2858 -3768
rect 2712 -3775 2724 -3774
rect 2594 -3820 2608 -3776
rect 2662 -3820 2674 -3776
rect 2594 -3826 2674 -3820
rect 2711 -3825 2724 -3775
rect 2420 -3844 2480 -3836
rect 2222 -3880 2298 -3874
rect 2598 -3880 2662 -3826
rect 2712 -3838 2724 -3825
rect 2846 -3838 2858 -3774
rect 2712 -3844 2858 -3838
rect 1886 -3888 2018 -3884
rect 762 -3918 822 -3906
rect 932 -3952 942 -3888
rect 1006 -3890 1838 -3888
rect 1006 -3942 1344 -3890
rect 1452 -3894 1838 -3890
rect 1452 -3942 1778 -3894
rect 1006 -3952 1032 -3942
rect 1334 -3950 1468 -3942
rect 1766 -3946 1778 -3942
rect 1830 -3946 1838 -3894
rect 1882 -3890 2020 -3888
rect 1882 -3934 1898 -3890
rect 2006 -3934 2020 -3890
rect 2218 -3932 2668 -3880
rect 1882 -3944 2020 -3934
rect 1766 -3952 1838 -3946
rect 778 -4014 788 -3960
rect 844 -3982 854 -3960
rect 1922 -3973 1984 -3944
rect 1676 -3982 1682 -3973
rect 844 -4014 1682 -3982
rect 796 -4016 1682 -4014
rect 1676 -4025 1682 -4016
rect 1734 -3982 1740 -3973
rect 1922 -3982 1986 -3973
rect 2795 -3982 2845 -3844
rect 1734 -4001 2845 -3982
rect 1734 -4016 2837 -4001
rect 1734 -4025 1740 -4016
rect 1922 -4025 1986 -4016
rect 1488 -4138 1498 -4072
rect 1824 -4138 1834 -4072
rect 2144 -4138 2150 -4078
rect 2210 -4138 2216 -4078
rect 2518 -4144 2528 -4056
rect 2608 -4144 2618 -4056
rect 1130 -4204 1204 -4144
rect 1318 -4194 1386 -4182
rect 1130 -4328 1148 -4204
rect 1184 -4328 1204 -4204
rect 1130 -4342 1204 -4328
rect 1314 -4334 1324 -4194
rect 1380 -4334 1390 -4194
rect 1592 -4196 1656 -4184
rect 1588 -4334 1598 -4196
rect 1650 -4334 1660 -4196
rect 1960 -4214 2028 -4202
rect 1960 -4216 1966 -4214
rect 2022 -4216 2028 -4214
rect 1318 -4346 1386 -4334
rect 1592 -4346 1656 -4334
rect 1958 -4336 1966 -4216
rect 1958 -4338 1968 -4336
rect 2026 -4338 2036 -4216
rect 2154 -4262 2160 -4210
rect 2212 -4215 2218 -4210
rect 2422 -4215 2428 -4210
rect 2212 -4257 2428 -4215
rect 2212 -4262 2218 -4257
rect 2422 -4262 2428 -4257
rect 2480 -4262 2486 -4210
rect 1960 -4348 2028 -4338
rect 1222 -4382 1310 -4376
rect 703 -4450 709 -4398
rect 761 -4409 767 -4398
rect 1222 -4409 1234 -4382
rect 761 -4426 1234 -4409
rect 1298 -4426 1310 -4382
rect 761 -4432 1310 -4426
rect 761 -4439 1295 -4432
rect 1394 -4434 1400 -4382
rect 1452 -4390 1458 -4382
rect 1504 -4384 1580 -4378
rect 1868 -4382 1952 -4376
rect 1504 -4390 1516 -4384
rect 1452 -4425 1516 -4390
rect 1452 -4434 1458 -4425
rect 1504 -4428 1516 -4425
rect 1568 -4428 1580 -4384
rect 1504 -4434 1580 -4428
rect 761 -4450 767 -4439
rect 1864 -4442 1874 -4382
rect 1940 -4436 1952 -4382
rect 1940 -4442 1950 -4436
rect 1128 -4570 1138 -4470
rect 1192 -4570 1202 -4470
rect 1980 -4480 2028 -4348
rect 2136 -4382 2218 -4376
rect 2136 -4430 2148 -4382
rect 2136 -4434 2160 -4430
rect 2212 -4434 2218 -4382
rect 2136 -4436 2218 -4434
rect 2248 -4388 2308 -4376
rect 1962 -4492 2028 -4480
rect 1962 -4558 1968 -4492
rect 2022 -4558 2028 -4492
rect 2248 -4542 2254 -4388
rect 2302 -4390 2308 -4388
rect 2320 -4542 2330 -4390
rect 2248 -4554 2308 -4542
rect 1962 -4570 2028 -4558
rect 778 -4680 788 -4614
rect 1102 -4680 1112 -4614
rect 1128 -4628 1202 -4570
rect 1128 -4634 1136 -4628
rect 1130 -4688 1136 -4634
rect 1196 -4688 1202 -4628
rect 2332 -4680 2342 -4614
rect 2656 -4680 2666 -4614
rect 2696 -4684 2702 -4624
rect 2762 -4684 2768 -4624
<< via1 >>
rect 802 -3050 2046 -2984
rect 2144 -3048 2214 -2972
rect 2526 -3060 2590 -2980
rect 787 -3214 839 -3162
rect 942 -3350 1000 -3292
rect 1254 -3344 1296 -3284
rect 1296 -3344 1322 -3284
rect 1254 -3352 1322 -3344
rect 1532 -3246 1562 -3186
rect 1562 -3246 1592 -3186
rect 1532 -3348 1592 -3246
rect 1136 -3592 1198 -3522
rect 1620 -3590 2108 -3524
rect 2256 -3592 2490 -3526
rect 2704 -3590 2762 -3528
rect 712 -3904 766 -3686
rect 1398 -3686 1450 -3634
rect 1530 -3720 1594 -3664
rect 1682 -3718 1734 -3698
rect 1239 -3828 1291 -3776
rect 1682 -3750 1732 -3718
rect 1732 -3750 1734 -3718
rect 1870 -3720 1922 -3668
rect 1778 -3814 1830 -3762
rect 2428 -3832 2474 -3660
rect 2474 -3832 2496 -3660
rect 2428 -3836 2496 -3832
rect 942 -3952 1006 -3888
rect 1778 -3946 1830 -3894
rect 788 -4014 844 -3960
rect 1682 -4025 1734 -3973
rect 1498 -4138 1824 -4072
rect 2150 -4138 2210 -4078
rect 2528 -4144 2608 -4056
rect 1324 -4334 1380 -4194
rect 1598 -4334 1650 -4196
rect 1968 -4336 2022 -4216
rect 2022 -4336 2026 -4216
rect 1968 -4338 2026 -4336
rect 2160 -4262 2212 -4210
rect 2428 -4262 2480 -4210
rect 709 -4450 761 -4398
rect 1400 -4434 1452 -4382
rect 1874 -4430 1880 -4382
rect 1880 -4430 1940 -4382
rect 1874 -4442 1940 -4430
rect 1138 -4484 1192 -4470
rect 1138 -4564 1146 -4484
rect 1146 -4564 1186 -4484
rect 1186 -4564 1192 -4484
rect 1138 -4570 1192 -4564
rect 2160 -4430 2206 -4382
rect 2206 -4430 2212 -4382
rect 2160 -4434 2212 -4430
rect 2258 -4542 2302 -4390
rect 2302 -4542 2320 -4390
rect 788 -4680 1102 -4614
rect 1136 -4688 1196 -4628
rect 2342 -4680 2656 -4614
rect 2702 -4684 2762 -4624
<< metal2 >>
rect 2144 -2972 2214 -2962
rect 802 -2984 2046 -2974
rect 802 -3060 2046 -3050
rect 2144 -3058 2214 -3048
rect 2526 -2980 2596 -2970
rect 787 -3162 839 -3156
rect 787 -3220 839 -3214
rect 1526 -3176 1562 -3132
rect 1526 -3186 1592 -3176
rect 712 -3686 766 -3676
rect 712 -3914 766 -3904
rect 720 -4392 750 -3914
rect 794 -3950 833 -3220
rect 1526 -3246 1532 -3186
rect 926 -3292 1006 -3282
rect 1254 -3284 1322 -3274
rect 926 -3350 942 -3292
rect 1000 -3350 1006 -3292
rect 926 -3370 1006 -3350
rect 788 -3960 844 -3950
rect 788 -4024 844 -4014
rect 876 -4234 910 -3710
rect 958 -3878 1006 -3370
rect 1240 -3352 1254 -3286
rect 1240 -3362 1322 -3352
rect 1532 -3358 1592 -3348
rect 942 -3888 1006 -3878
rect 942 -3966 1006 -3952
rect 1136 -3522 1198 -3512
rect 1136 -3602 1198 -3592
rect 709 -4398 761 -4392
rect 709 -4456 761 -4450
rect 720 -4798 750 -4456
rect 1136 -4470 1196 -3602
rect 1240 -3770 1290 -3362
rect 1398 -3634 1450 -3628
rect 1538 -3654 1588 -3358
rect 1620 -3524 2108 -3514
rect 1620 -3600 2108 -3590
rect 1398 -3692 1450 -3686
rect 1530 -3664 1594 -3654
rect 1239 -3776 1291 -3770
rect 1239 -3834 1291 -3828
rect 1324 -4194 1380 -4184
rect 1324 -4344 1380 -4334
rect 1136 -4570 1138 -4470
rect 1192 -4570 1196 -4470
rect 788 -4614 1102 -4604
rect 788 -4690 1102 -4680
rect 1136 -4628 1196 -4570
rect 1136 -4694 1196 -4688
rect 1332 -4798 1362 -4344
rect 1411 -4376 1441 -3692
rect 1870 -3668 1922 -3662
rect 1530 -3730 1594 -3720
rect 1682 -3698 1734 -3692
rect 1870 -3726 1922 -3720
rect 1682 -3756 1734 -3750
rect 1691 -3967 1725 -3756
rect 1778 -3762 1830 -3756
rect 1778 -3820 1830 -3814
rect 1783 -3894 1825 -3820
rect 1772 -3946 1778 -3894
rect 1830 -3946 1836 -3894
rect 1682 -3973 1734 -3967
rect 1682 -4031 1734 -4025
rect 1498 -4072 1824 -4062
rect 1498 -4148 1824 -4138
rect 1598 -4196 1650 -4186
rect 1598 -4344 1650 -4334
rect 1400 -4382 1452 -4376
rect 1400 -4440 1452 -4434
rect 1411 -4798 1441 -4440
rect 1610 -4798 1640 -4344
rect 1874 -4372 1918 -3726
rect 2150 -4078 2210 -3058
rect 2590 -3060 2596 -2980
rect 2526 -3070 2596 -3060
rect 2256 -3526 2490 -3516
rect 2256 -3602 2490 -3592
rect 2150 -4144 2210 -4138
rect 2428 -3660 2496 -3650
rect 2428 -3846 2496 -3836
rect 1968 -4216 2026 -4206
rect 2160 -4210 2212 -4204
rect 2160 -4268 2212 -4262
rect 2428 -4210 2480 -3846
rect 2536 -3988 2596 -3070
rect 2704 -3528 2762 -3518
rect 2702 -3590 2704 -3528
rect 2528 -4056 2608 -3988
rect 2528 -4156 2608 -4144
rect 2428 -4268 2480 -4262
rect 1968 -4348 2026 -4338
rect 1874 -4382 1940 -4372
rect 1874 -4452 1940 -4442
rect 1879 -4798 1913 -4452
rect 1980 -4798 2010 -4348
rect 2165 -4376 2207 -4268
rect 2160 -4382 2212 -4376
rect 2160 -4440 2212 -4434
rect 2258 -4390 2320 -4380
rect 2170 -4798 2203 -4440
rect 2258 -4552 2320 -4542
rect 2262 -4798 2295 -4552
rect 2342 -4614 2656 -4604
rect 2342 -4690 2656 -4680
rect 2702 -4624 2762 -3590
rect 2702 -4690 2762 -4684
<< via2 >>
rect 802 -3050 2046 -2984
rect 1620 -3590 2108 -3524
rect 788 -4680 1102 -4614
rect 1498 -4138 1824 -4072
rect 2256 -3592 2490 -3526
rect 2342 -4680 2656 -4614
<< metal3 >>
rect 750 -2984 2774 -2966
rect 750 -3050 802 -2984
rect 2046 -3050 2774 -2984
rect 750 -3062 2774 -3050
rect 750 -3524 2774 -3510
rect 750 -3590 1620 -3524
rect 2108 -3526 2774 -3524
rect 2108 -3590 2256 -3526
rect 750 -3592 2256 -3590
rect 2490 -3592 2774 -3526
rect 750 -3606 2774 -3592
rect 752 -4072 2776 -4054
rect 752 -4138 1498 -4072
rect 1824 -4138 2776 -4072
rect 752 -4150 2776 -4138
rect 752 -4614 2776 -4598
rect 752 -4680 788 -4614
rect 1102 -4680 2342 -4614
rect 2656 -4680 2776 -4614
rect 752 -4694 2776 -4680
use sky130_fd_sc_hd__inv_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1120 0 1 -3558
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  x2
timestamp 1704896540
transform 1 0 1396 0 1 -3558
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1948 0 1 -3558
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  x4
timestamp 1704896540
transform -1 0 2408 0 -1 -3558
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  x5
timestamp 1704896540
transform 1 0 1120 0 1 -4646
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  x6
timestamp 1704896540
transform 1 0 1764 0 1 -4646
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1212 0 -1 -3558
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1764 0 -1 -3558
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  x9
timestamp 1704896540
transform -1 0 2316 0 -1 -3558
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  x10
timestamp 1704896540
transform -1 0 2868 0 -1 -3558
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  x11
timestamp 1704896540
transform 1 0 1212 0 1 -4646
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  x12
timestamp 1704896540
transform 1 0 1488 0 1 -4646
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  x13
timestamp 1704896540
transform 1 0 1856 0 1 -4646
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  x14
timestamp 1704896540
transform 1 0 2132 0 1 -4646
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2040 0 1 -3558
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  x16
timestamp 1704896540
transform 1 0 2408 0 1 -4646
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  x17
timestamp 1704896540
transform 1 0 752 0 1 -4646
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  x18
timestamp 1704896540
transform 1 0 1672 0 1 -3558
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  x19
timestamp 1704896540
transform 1 0 752 0 1 -3558
box -38 -48 406 592
<< labels >>
flabel metal1 676 -3352 742 -3290 0 FreeSans 800 0 0 0 SEL0
port 0 nsew
flabel metal1 682 -3218 748 -3156 0 FreeSans 800 0 0 0 SEL1
port 1 nsew
flabel metal1 674 -3464 740 -3402 0 FreeSans 800 0 0 0 SEL2
port 2 nsew
flabel metal2 722 -4794 748 -4720 0 FreeSans 480 0 0 0 gno0
port 3 nsew
flabel metal2 1334 -4794 1360 -4720 0 FreeSans 480 0 0 0 gpo0
port 4 nsew
flabel metal2 1412 -4792 1438 -4718 0 FreeSans 480 0 0 0 gno1
port 5 nsew
flabel metal2 1612 -4794 1638 -4720 0 FreeSans 480 0 0 0 gpo1
port 6 nsew
flabel metal2 1884 -4792 1910 -4718 0 FreeSans 480 0 0 0 gno2
port 7 nsew
flabel metal2 1982 -4792 2008 -4718 0 FreeSans 480 0 0 0 gpo2
port 8 nsew
flabel metal2 2172 -4792 2198 -4718 0 FreeSans 480 0 0 0 gno3
port 9 nsew
flabel metal2 2266 -4792 2292 -4718 0 FreeSans 480 0 0 0 gpo3
port 10 nsew
flabel metal1 2466 -3142 2602 -3104 0 FreeSans 480 0 0 0 nSEL2
port 11 nsew
flabel metal3 2642 -3054 2766 -2980 0 FreeSans 640 0 0 0 VPWR
port 12 nsew
flabel metal3 2600 -4146 2768 -4058 0 FreeSans 640 0 0 0 VPWR
port 12 nsew
flabel metal3 780 -3604 948 -3516 0 FreeSans 640 0 0 0 VGND
port 13 nsew
flabel metal3 766 -4690 934 -4602 0 FreeSans 640 0 0 0 VGND
port 13 nsew
flabel metal2 1246 -3348 1310 -3294 0 FreeSans 320 0 0 0 nSEL0
flabel metal2 1534 -3350 1592 -3302 0 FreeSans 320 0 0 0 nSEL1
<< end >>
