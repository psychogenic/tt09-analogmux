magic
tech sky130A
magscale 1 2
timestamp 1728339728
<< viali >>
rect 2697 9537 2731 9571
rect 2513 9333 2547 9367
rect 2053 8449 2087 8483
rect 2145 8381 2179 8415
rect 2421 8313 2455 8347
rect 3249 7837 3283 7871
rect 2982 7769 3016 7803
rect 1869 7701 1903 7735
rect 1678 7497 1712 7531
rect 1501 7361 1535 7395
rect 1593 7361 1627 7395
rect 1777 7361 1811 7395
rect 2982 7361 3016 7395
rect 3249 7293 3283 7327
rect 1869 7225 1903 7259
rect 2421 6953 2455 6987
rect 3065 6953 3099 6987
rect 2973 6817 3007 6851
rect 3065 6749 3099 6783
rect 3249 6749 3283 6783
rect 2237 6681 2271 6715
rect 2789 6681 2823 6715
rect 2437 6613 2471 6647
rect 2605 6613 2639 6647
rect 2237 5865 2271 5899
rect 6009 5661 6043 5695
rect 3525 5593 3559 5627
rect 4721 5525 4755 5559
rect 4353 5321 4387 5355
rect 6561 5321 6595 5355
rect 5488 5253 5522 5287
rect 6009 5185 6043 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7757 5185 7791 5219
rect 3801 5117 3835 5151
rect 4261 5117 4295 5151
rect 5733 5117 5767 5151
rect 7021 5117 7055 5151
rect 7481 5117 7515 5151
rect 4169 5049 4203 5083
rect 5825 5049 5859 5083
rect 6377 5049 6411 5083
rect 7389 5049 7423 5083
rect 6929 4981 6963 5015
rect 7573 4981 7607 5015
rect 3617 4709 3651 4743
rect 2237 4641 2271 4675
rect 5089 4641 5123 4675
rect 1961 4573 1995 4607
rect 2145 4573 2179 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 4997 4573 5031 4607
rect 5460 4573 5494 4607
rect 5733 4573 5767 4607
rect 2504 4505 2538 4539
rect 2053 4437 2087 4471
rect 4905 4437 4939 4471
rect 5457 4437 5491 4471
rect 5641 4437 5675 4471
rect 7021 4437 7055 4471
rect 3065 4233 3099 4267
rect 5058 4165 5092 4199
rect 6920 4165 6954 4199
rect 1409 4097 1443 4131
rect 1593 4097 1627 4131
rect 1685 4097 1719 4131
rect 1941 4097 1975 4131
rect 3525 4097 3559 4131
rect 4629 4097 4663 4131
rect 6653 4097 6687 4131
rect 1501 4029 1535 4063
rect 3157 4029 3191 4063
rect 3617 4029 3651 4063
rect 4169 4029 4203 4063
rect 4353 4029 4387 4063
rect 4445 4029 4479 4063
rect 4537 4029 4571 4063
rect 4813 4029 4847 4063
rect 6193 3893 6227 3927
rect 8033 3893 8067 3927
rect 4445 3689 4479 3723
rect 4629 3689 4663 3723
rect 4905 3689 4939 3723
rect 4169 3621 4203 3655
rect 4721 3621 4755 3655
rect 3801 3553 3835 3587
rect 1961 3485 1995 3519
rect 3985 3485 4019 3519
rect 5181 3485 5215 3519
rect 6653 3485 6687 3519
rect 4491 3451 4525 3485
rect 2228 3417 2262 3451
rect 4261 3417 4295 3451
rect 4884 3417 4918 3451
rect 5089 3417 5123 3451
rect 5448 3417 5482 3451
rect 6920 3417 6954 3451
rect 3341 3349 3375 3383
rect 6561 3349 6595 3383
rect 8033 3349 8067 3383
rect 2421 3145 2455 3179
rect 4169 3145 4203 3179
rect 5549 3145 5583 3179
rect 6561 3145 6595 3179
rect 6653 3145 6687 3179
rect 7573 3145 7607 3179
rect 5733 3077 5767 3111
rect 6929 3077 6963 3111
rect 2605 3009 2639 3043
rect 2881 3009 2915 3043
rect 3065 3009 3099 3043
rect 3341 3009 3375 3043
rect 3985 3009 4019 3043
rect 5825 3009 5859 3043
rect 5917 3009 5951 3043
rect 6745 3009 6779 3043
rect 7113 3009 7147 3043
rect 8033 3009 8067 3043
rect 3157 2941 3191 2975
rect 3525 2941 3559 2975
rect 3801 2941 3835 2975
rect 7205 2941 7239 2975
rect 7297 2941 7331 2975
rect 7389 2941 7423 2975
rect 7665 2941 7699 2975
rect 7941 2941 7975 2975
rect 6101 2873 6135 2907
rect 6377 2805 6411 2839
rect 8125 2533 8159 2567
rect 1593 2397 1627 2431
rect 1961 2397 1995 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5641 2397 5675 2431
rect 6561 2397 6595 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 8401 2397 8435 2431
rect 1409 2261 1443 2295
rect 1777 2261 1811 2295
rect 2697 2261 2731 2295
rect 3801 2261 3835 2295
rect 4537 2261 4571 2295
rect 5457 2261 5491 2295
rect 6377 2261 6411 2295
rect 7297 2261 7331 2295
rect 8217 2261 8251 2295
<< metal1 >>
rect 1104 9818 8740 9840
rect 1104 9766 1810 9818
rect 1862 9766 1874 9818
rect 1926 9766 1938 9818
rect 1990 9766 2002 9818
rect 2054 9766 2066 9818
rect 2118 9766 3130 9818
rect 3182 9766 3194 9818
rect 3246 9766 3258 9818
rect 3310 9766 3322 9818
rect 3374 9766 3386 9818
rect 3438 9766 4450 9818
rect 4502 9766 4514 9818
rect 4566 9766 4578 9818
rect 4630 9766 4642 9818
rect 4694 9766 4706 9818
rect 4758 9766 5770 9818
rect 5822 9766 5834 9818
rect 5886 9766 5898 9818
rect 5950 9766 5962 9818
rect 6014 9766 6026 9818
rect 6078 9766 7090 9818
rect 7142 9766 7154 9818
rect 7206 9766 7218 9818
rect 7270 9766 7282 9818
rect 7334 9766 7346 9818
rect 7398 9766 8410 9818
rect 8462 9766 8474 9818
rect 8526 9766 8538 9818
rect 8590 9766 8602 9818
rect 8654 9766 8666 9818
rect 8718 9766 8740 9818
rect 1104 9744 8740 9766
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2464 9540 2697 9568
rect 2464 9528 2470 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2501 9367 2559 9373
rect 2501 9364 2513 9367
rect 2188 9336 2513 9364
rect 2188 9324 2194 9336
rect 2501 9333 2513 9336
rect 2547 9333 2559 9367
rect 2501 9327 2559 9333
rect 1104 9274 8740 9296
rect 1104 9222 1150 9274
rect 1202 9222 1214 9274
rect 1266 9222 1278 9274
rect 1330 9222 1342 9274
rect 1394 9222 1406 9274
rect 1458 9222 2470 9274
rect 2522 9222 2534 9274
rect 2586 9222 2598 9274
rect 2650 9222 2662 9274
rect 2714 9222 2726 9274
rect 2778 9222 3790 9274
rect 3842 9222 3854 9274
rect 3906 9222 3918 9274
rect 3970 9222 3982 9274
rect 4034 9222 4046 9274
rect 4098 9222 5110 9274
rect 5162 9222 5174 9274
rect 5226 9222 5238 9274
rect 5290 9222 5302 9274
rect 5354 9222 5366 9274
rect 5418 9222 6430 9274
rect 6482 9222 6494 9274
rect 6546 9222 6558 9274
rect 6610 9222 6622 9274
rect 6674 9222 6686 9274
rect 6738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 7942 9274
rect 7994 9222 8006 9274
rect 8058 9222 8740 9274
rect 1104 9200 8740 9222
rect 1104 8730 8740 8752
rect 1104 8678 1810 8730
rect 1862 8678 1874 8730
rect 1926 8678 1938 8730
rect 1990 8678 2002 8730
rect 2054 8678 2066 8730
rect 2118 8678 3130 8730
rect 3182 8678 3194 8730
rect 3246 8678 3258 8730
rect 3310 8678 3322 8730
rect 3374 8678 3386 8730
rect 3438 8678 4450 8730
rect 4502 8678 4514 8730
rect 4566 8678 4578 8730
rect 4630 8678 4642 8730
rect 4694 8678 4706 8730
rect 4758 8678 5770 8730
rect 5822 8678 5834 8730
rect 5886 8678 5898 8730
rect 5950 8678 5962 8730
rect 6014 8678 6026 8730
rect 6078 8678 7090 8730
rect 7142 8678 7154 8730
rect 7206 8678 7218 8730
rect 7270 8678 7282 8730
rect 7334 8678 7346 8730
rect 7398 8678 8410 8730
rect 8462 8678 8474 8730
rect 8526 8678 8538 8730
rect 8590 8678 8602 8730
rect 8654 8678 8666 8730
rect 8718 8678 8740 8730
rect 1104 8656 8740 8678
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1636 8452 2053 8480
rect 1636 8440 1642 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2130 8372 2136 8424
rect 2188 8372 2194 8424
rect 2409 8347 2467 8353
rect 2409 8313 2421 8347
rect 2455 8344 2467 8347
rect 2866 8344 2872 8356
rect 2455 8316 2872 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 1104 8186 8740 8208
rect 1104 8134 1150 8186
rect 1202 8134 1214 8186
rect 1266 8134 1278 8186
rect 1330 8134 1342 8186
rect 1394 8134 1406 8186
rect 1458 8134 2470 8186
rect 2522 8134 2534 8186
rect 2586 8134 2598 8186
rect 2650 8134 2662 8186
rect 2714 8134 2726 8186
rect 2778 8134 3790 8186
rect 3842 8134 3854 8186
rect 3906 8134 3918 8186
rect 3970 8134 3982 8186
rect 4034 8134 4046 8186
rect 4098 8134 5110 8186
rect 5162 8134 5174 8186
rect 5226 8134 5238 8186
rect 5290 8134 5302 8186
rect 5354 8134 5366 8186
rect 5418 8134 6430 8186
rect 6482 8134 6494 8186
rect 6546 8134 6558 8186
rect 6610 8134 6622 8186
rect 6674 8134 6686 8186
rect 6738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 7942 8186
rect 7994 8134 8006 8186
rect 8058 8134 8740 8186
rect 1104 8112 8740 8134
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 2280 7840 3249 7868
rect 2280 7828 2286 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 2866 7760 2872 7812
rect 2924 7800 2930 7812
rect 2970 7803 3028 7809
rect 2970 7800 2982 7803
rect 2924 7772 2982 7800
rect 2924 7760 2930 7772
rect 2970 7769 2982 7772
rect 3016 7769 3028 7803
rect 2970 7763 3028 7769
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1636 7704 1869 7732
rect 1636 7692 1642 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 1104 7642 8740 7664
rect 1104 7590 1810 7642
rect 1862 7590 1874 7642
rect 1926 7590 1938 7642
rect 1990 7590 2002 7642
rect 2054 7590 2066 7642
rect 2118 7590 3130 7642
rect 3182 7590 3194 7642
rect 3246 7590 3258 7642
rect 3310 7590 3322 7642
rect 3374 7590 3386 7642
rect 3438 7590 4450 7642
rect 4502 7590 4514 7642
rect 4566 7590 4578 7642
rect 4630 7590 4642 7642
rect 4694 7590 4706 7642
rect 4758 7590 5770 7642
rect 5822 7590 5834 7642
rect 5886 7590 5898 7642
rect 5950 7590 5962 7642
rect 6014 7590 6026 7642
rect 6078 7590 7090 7642
rect 7142 7590 7154 7642
rect 7206 7590 7218 7642
rect 7270 7590 7282 7642
rect 7334 7590 7346 7642
rect 7398 7590 8410 7642
rect 8462 7590 8474 7642
rect 8526 7590 8538 7642
rect 8590 7590 8602 7642
rect 8654 7590 8666 7642
rect 8718 7590 8740 7642
rect 1104 7568 8740 7590
rect 1666 7531 1724 7537
rect 1666 7497 1678 7531
rect 1712 7528 1724 7531
rect 3050 7528 3056 7540
rect 1712 7500 3056 7528
rect 1712 7497 1724 7500
rect 1666 7491 1724 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 2130 7460 2136 7472
rect 1504 7432 2136 7460
rect 1504 7401 1532 7432
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 1578 7352 1584 7404
rect 1636 7352 1642 7404
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 1670 7216 1676 7268
rect 1728 7256 1734 7268
rect 1780 7256 1808 7355
rect 2958 7352 2964 7404
rect 3016 7401 3022 7404
rect 3016 7355 3028 7401
rect 3016 7352 3022 7355
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7293 3295 7327
rect 3237 7287 3295 7293
rect 1857 7259 1915 7265
rect 1857 7256 1869 7259
rect 1728 7228 1869 7256
rect 1728 7216 1734 7228
rect 1857 7225 1869 7228
rect 1903 7225 1915 7259
rect 1857 7219 1915 7225
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 3252 7188 3280 7287
rect 2280 7160 3280 7188
rect 2280 7148 2286 7160
rect 1104 7098 8740 7120
rect 1104 7046 1150 7098
rect 1202 7046 1214 7098
rect 1266 7046 1278 7098
rect 1330 7046 1342 7098
rect 1394 7046 1406 7098
rect 1458 7046 2470 7098
rect 2522 7046 2534 7098
rect 2586 7046 2598 7098
rect 2650 7046 2662 7098
rect 2714 7046 2726 7098
rect 2778 7046 3790 7098
rect 3842 7046 3854 7098
rect 3906 7046 3918 7098
rect 3970 7046 3982 7098
rect 4034 7046 4046 7098
rect 4098 7046 5110 7098
rect 5162 7046 5174 7098
rect 5226 7046 5238 7098
rect 5290 7046 5302 7098
rect 5354 7046 5366 7098
rect 5418 7046 6430 7098
rect 6482 7046 6494 7098
rect 6546 7046 6558 7098
rect 6610 7046 6622 7098
rect 6674 7046 6686 7098
rect 6738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 7942 7098
rect 7994 7046 8006 7098
rect 8058 7046 8740 7098
rect 1104 7024 8740 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 1728 6956 2421 6984
rect 1728 6944 1734 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 3053 6987 3111 6993
rect 3053 6984 3065 6987
rect 3016 6956 3065 6984
rect 3016 6944 3022 6956
rect 3053 6953 3065 6956
rect 3099 6953 3111 6987
rect 3053 6947 3111 6953
rect 2866 6808 2872 6860
rect 2924 6848 2930 6860
rect 2961 6851 3019 6857
rect 2961 6848 2973 6851
rect 2924 6820 2973 6848
rect 2924 6808 2930 6820
rect 2961 6817 2973 6820
rect 3007 6848 3019 6851
rect 3007 6820 3280 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 3252 6789 3280 6820
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 1486 6672 1492 6724
rect 1544 6712 1550 6724
rect 2225 6715 2283 6721
rect 2225 6712 2237 6715
rect 1544 6684 2237 6712
rect 1544 6672 1550 6684
rect 2225 6681 2237 6684
rect 2271 6681 2283 6715
rect 2777 6715 2835 6721
rect 2777 6712 2789 6715
rect 2225 6675 2283 6681
rect 2608 6684 2789 6712
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2608 6653 2636 6684
rect 2777 6681 2789 6684
rect 2823 6681 2835 6715
rect 2777 6675 2835 6681
rect 2425 6647 2483 6653
rect 2425 6644 2437 6647
rect 2188 6616 2437 6644
rect 2188 6604 2194 6616
rect 2425 6613 2437 6616
rect 2471 6613 2483 6647
rect 2425 6607 2483 6613
rect 2593 6647 2651 6653
rect 2593 6613 2605 6647
rect 2639 6613 2651 6647
rect 2593 6607 2651 6613
rect 1104 6554 8740 6576
rect 1104 6502 1810 6554
rect 1862 6502 1874 6554
rect 1926 6502 1938 6554
rect 1990 6502 2002 6554
rect 2054 6502 2066 6554
rect 2118 6502 3130 6554
rect 3182 6502 3194 6554
rect 3246 6502 3258 6554
rect 3310 6502 3322 6554
rect 3374 6502 3386 6554
rect 3438 6502 4450 6554
rect 4502 6502 4514 6554
rect 4566 6502 4578 6554
rect 4630 6502 4642 6554
rect 4694 6502 4706 6554
rect 4758 6502 5770 6554
rect 5822 6502 5834 6554
rect 5886 6502 5898 6554
rect 5950 6502 5962 6554
rect 6014 6502 6026 6554
rect 6078 6502 7090 6554
rect 7142 6502 7154 6554
rect 7206 6502 7218 6554
rect 7270 6502 7282 6554
rect 7334 6502 7346 6554
rect 7398 6502 8410 6554
rect 8462 6502 8474 6554
rect 8526 6502 8538 6554
rect 8590 6502 8602 6554
rect 8654 6502 8666 6554
rect 8718 6502 8740 6554
rect 1104 6480 8740 6502
rect 1104 6010 8740 6032
rect 1104 5958 1150 6010
rect 1202 5958 1214 6010
rect 1266 5958 1278 6010
rect 1330 5958 1342 6010
rect 1394 5958 1406 6010
rect 1458 5958 2470 6010
rect 2522 5958 2534 6010
rect 2586 5958 2598 6010
rect 2650 5958 2662 6010
rect 2714 5958 2726 6010
rect 2778 5958 3790 6010
rect 3842 5958 3854 6010
rect 3906 5958 3918 6010
rect 3970 5958 3982 6010
rect 4034 5958 4046 6010
rect 4098 5958 5110 6010
rect 5162 5958 5174 6010
rect 5226 5958 5238 6010
rect 5290 5958 5302 6010
rect 5354 5958 5366 6010
rect 5418 5958 6430 6010
rect 6482 5958 6494 6010
rect 6546 5958 6558 6010
rect 6610 5958 6622 6010
rect 6674 5958 6686 6010
rect 6738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 7942 6010
rect 7994 5958 8006 6010
rect 8058 5958 8740 6010
rect 1104 5936 8740 5958
rect 2222 5856 2228 5908
rect 2280 5856 2286 5908
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5692 6055 5695
rect 6822 5692 6828 5704
rect 6043 5664 6828 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 3513 5627 3571 5633
rect 3513 5593 3525 5627
rect 3559 5593 3571 5627
rect 3513 5587 3571 5593
rect 3528 5556 3556 5587
rect 4709 5559 4767 5565
rect 4709 5556 4721 5559
rect 3528 5528 4721 5556
rect 4709 5525 4721 5528
rect 4755 5556 4767 5559
rect 5442 5556 5448 5568
rect 4755 5528 5448 5556
rect 4755 5525 4767 5528
rect 4709 5519 4767 5525
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 1104 5466 8740 5488
rect 1104 5414 1810 5466
rect 1862 5414 1874 5466
rect 1926 5414 1938 5466
rect 1990 5414 2002 5466
rect 2054 5414 2066 5466
rect 2118 5414 3130 5466
rect 3182 5414 3194 5466
rect 3246 5414 3258 5466
rect 3310 5414 3322 5466
rect 3374 5414 3386 5466
rect 3438 5414 4450 5466
rect 4502 5414 4514 5466
rect 4566 5414 4578 5466
rect 4630 5414 4642 5466
rect 4694 5414 4706 5466
rect 4758 5414 5770 5466
rect 5822 5414 5834 5466
rect 5886 5414 5898 5466
rect 5950 5414 5962 5466
rect 6014 5414 6026 5466
rect 6078 5414 7090 5466
rect 7142 5414 7154 5466
rect 7206 5414 7218 5466
rect 7270 5414 7282 5466
rect 7334 5414 7346 5466
rect 7398 5414 8410 5466
rect 8462 5414 8474 5466
rect 8526 5414 8538 5466
rect 8590 5414 8602 5466
rect 8654 5414 8666 5466
rect 8718 5414 8740 5466
rect 1104 5392 8740 5414
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 6270 5352 6276 5364
rect 4387 5324 6276 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 6270 5312 6276 5324
rect 6328 5352 6334 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6328 5324 6561 5352
rect 6328 5312 6334 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 5476 5287 5534 5293
rect 5476 5253 5488 5287
rect 5522 5284 5534 5287
rect 5810 5284 5816 5296
rect 5522 5256 5816 5284
rect 5522 5253 5534 5256
rect 5476 5247 5534 5253
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 4264 5188 6009 5216
rect 4264 5157 4292 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6144 5188 6653 5216
rect 6144 5176 6150 5188
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 6822 5216 6828 5228
rect 6779 5188 6828 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7484 5188 7757 5216
rect 3789 5151 3847 5157
rect 3789 5117 3801 5151
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5117 4307 5151
rect 4249 5111 4307 5117
rect 3804 5012 3832 5111
rect 5718 5108 5724 5160
rect 5776 5108 5782 5160
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7484 5157 7512 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 4154 5040 4160 5092
rect 4212 5040 4218 5092
rect 4264 5052 4476 5080
rect 4264 5012 4292 5052
rect 4448 5024 4476 5052
rect 5810 5040 5816 5092
rect 5868 5040 5874 5092
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 6365 5083 6423 5089
rect 6365 5080 6377 5083
rect 6052 5052 6377 5080
rect 6052 5040 6058 5052
rect 6365 5049 6377 5052
rect 6411 5049 6423 5083
rect 6365 5043 6423 5049
rect 7377 5083 7435 5089
rect 7377 5049 7389 5083
rect 7423 5080 7435 5083
rect 7423 5052 7512 5080
rect 7423 5049 7435 5052
rect 7377 5043 7435 5049
rect 7484 5024 7512 5052
rect 3804 4984 4292 5012
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 6917 5015 6975 5021
rect 6917 5012 6929 5015
rect 4488 4984 6929 5012
rect 4488 4972 4494 4984
rect 6917 4981 6929 4984
rect 6963 4981 6975 5015
rect 6917 4975 6975 4981
rect 7466 4972 7472 5024
rect 7524 4972 7530 5024
rect 7558 4972 7564 5024
rect 7616 4972 7622 5024
rect 1104 4922 8740 4944
rect 1104 4870 1150 4922
rect 1202 4870 1214 4922
rect 1266 4870 1278 4922
rect 1330 4870 1342 4922
rect 1394 4870 1406 4922
rect 1458 4870 2470 4922
rect 2522 4870 2534 4922
rect 2586 4870 2598 4922
rect 2650 4870 2662 4922
rect 2714 4870 2726 4922
rect 2778 4870 3790 4922
rect 3842 4870 3854 4922
rect 3906 4870 3918 4922
rect 3970 4870 3982 4922
rect 4034 4870 4046 4922
rect 4098 4870 5110 4922
rect 5162 4870 5174 4922
rect 5226 4870 5238 4922
rect 5290 4870 5302 4922
rect 5354 4870 5366 4922
rect 5418 4870 6430 4922
rect 6482 4870 6494 4922
rect 6546 4870 6558 4922
rect 6610 4870 6622 4922
rect 6674 4870 6686 4922
rect 6738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 7942 4922
rect 7994 4870 8006 4922
rect 8058 4870 8740 4922
rect 1104 4848 8740 4870
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 6086 4808 6092 4820
rect 2924 4780 6092 4808
rect 2924 4768 2930 4780
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 3510 4700 3516 4752
rect 3568 4740 3574 4752
rect 3605 4743 3663 4749
rect 3605 4740 3617 4743
rect 3568 4712 3617 4740
rect 3568 4700 3574 4712
rect 3605 4709 3617 4712
rect 3651 4740 3663 4743
rect 5442 4740 5448 4752
rect 3651 4712 5448 4740
rect 3651 4709 3663 4712
rect 3605 4703 3663 4709
rect 5442 4700 5448 4712
rect 5500 4740 5506 4752
rect 5994 4740 6000 4752
rect 5500 4712 6000 4740
rect 5500 4700 5506 4712
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 2222 4632 2228 4684
rect 2280 4632 2286 4684
rect 4890 4672 4896 4684
rect 4264 4644 4896 4672
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4604 2191 4607
rect 2958 4604 2964 4616
rect 2179 4576 2964 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 1964 4536 1992 4567
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 4264 4613 4292 4644
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 6178 4672 6184 4684
rect 5123 4644 6184 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4430 4564 4436 4616
rect 4488 4564 4494 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4798 4604 4804 4616
rect 4755 4576 4804 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 4798 4564 4804 4576
rect 4856 4604 4862 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4856 4576 4997 4604
rect 4856 4564 4862 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 5448 4607 5506 4613
rect 5448 4604 5460 4607
rect 4985 4567 5043 4573
rect 5092 4576 5460 4604
rect 2492 4539 2550 4545
rect 1964 4508 2176 4536
rect 1394 4428 1400 4480
rect 1452 4468 1458 4480
rect 2041 4471 2099 4477
rect 2041 4468 2053 4471
rect 1452 4440 2053 4468
rect 1452 4428 1458 4440
rect 2041 4437 2053 4440
rect 2087 4437 2099 4471
rect 2148 4468 2176 4508
rect 2492 4505 2504 4539
rect 2538 4536 2550 4539
rect 3050 4536 3056 4548
rect 2538 4508 3056 4536
rect 2538 4505 2550 4508
rect 2492 4499 2550 4505
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 5092 4536 5120 4576
rect 5448 4573 5460 4576
rect 5494 4573 5506 4607
rect 5448 4567 5506 4573
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5684 4576 5733 4604
rect 5684 4564 5690 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 4264 4508 5120 4536
rect 4264 4480 4292 4508
rect 2866 4468 2872 4480
rect 2148 4440 2872 4468
rect 2041 4431 2099 4437
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 4246 4428 4252 4480
rect 4304 4428 4310 4480
rect 4890 4428 4896 4480
rect 4948 4428 4954 4480
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5534 4468 5540 4480
rect 5491 4440 5540 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5626 4428 5632 4480
rect 5684 4428 5690 4480
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 6638 4468 6644 4480
rect 5776 4440 6644 4468
rect 5776 4428 5782 4440
rect 6638 4428 6644 4440
rect 6696 4468 6702 4480
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6696 4440 7021 4468
rect 6696 4428 6702 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7009 4431 7067 4437
rect 1104 4378 8740 4400
rect 1104 4326 1810 4378
rect 1862 4326 1874 4378
rect 1926 4326 1938 4378
rect 1990 4326 2002 4378
rect 2054 4326 2066 4378
rect 2118 4326 3130 4378
rect 3182 4326 3194 4378
rect 3246 4326 3258 4378
rect 3310 4326 3322 4378
rect 3374 4326 3386 4378
rect 3438 4326 4450 4378
rect 4502 4326 4514 4378
rect 4566 4326 4578 4378
rect 4630 4326 4642 4378
rect 4694 4326 4706 4378
rect 4758 4326 5770 4378
rect 5822 4326 5834 4378
rect 5886 4326 5898 4378
rect 5950 4326 5962 4378
rect 6014 4326 6026 4378
rect 6078 4326 7090 4378
rect 7142 4326 7154 4378
rect 7206 4326 7218 4378
rect 7270 4326 7282 4378
rect 7334 4326 7346 4378
rect 7398 4326 8410 4378
rect 8462 4326 8474 4378
rect 8526 4326 8538 4378
rect 8590 4326 8602 4378
rect 8654 4326 8666 4378
rect 8718 4326 8740 4378
rect 1104 4304 8740 4326
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3053 4267 3111 4273
rect 3053 4264 3065 4267
rect 3016 4236 3065 4264
rect 3016 4224 3022 4236
rect 3053 4233 3065 4236
rect 3099 4233 3111 4267
rect 3053 4227 3111 4233
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 6822 4264 6828 4276
rect 4488 4236 6828 4264
rect 4488 4224 4494 4236
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 2038 4196 2044 4208
rect 1688 4168 2044 4196
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 1578 4088 1584 4140
rect 1636 4088 1642 4140
rect 1688 4137 1716 4168
rect 2038 4156 2044 4168
rect 2096 4196 2102 4208
rect 2222 4196 2228 4208
rect 2096 4168 2228 4196
rect 2096 4156 2102 4168
rect 2222 4156 2228 4168
rect 2280 4156 2286 4208
rect 4448 4196 4476 4224
rect 4264 4168 4476 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1929 4131 1987 4137
rect 1929 4128 1941 4131
rect 1673 4091 1731 4097
rect 1780 4100 1941 4128
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 1780 4060 1808 4100
rect 1929 4097 1941 4100
rect 1975 4097 1987 4131
rect 1929 4091 1987 4097
rect 3510 4088 3516 4140
rect 3568 4088 3574 4140
rect 1535 4032 1808 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 3145 4063 3203 4069
rect 3145 4060 3157 4063
rect 3108 4032 3157 4060
rect 3108 4020 3114 4032
rect 3145 4029 3157 4032
rect 3191 4029 3203 4063
rect 3145 4023 3203 4029
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 3620 3992 3648 4023
rect 4154 4020 4160 4072
rect 4212 4020 4218 4072
rect 4264 4060 4292 4168
rect 4890 4156 4896 4208
rect 4948 4196 4954 4208
rect 5046 4199 5104 4205
rect 5046 4196 5058 4199
rect 4948 4168 5058 4196
rect 4948 4156 4954 4168
rect 5046 4165 5058 4168
rect 5092 4165 5104 4199
rect 5046 4159 5104 4165
rect 6908 4199 6966 4205
rect 6908 4165 6920 4199
rect 6954 4196 6966 4199
rect 7558 4196 7564 4208
rect 6954 4168 7564 4196
rect 6954 4165 6966 4168
rect 6908 4159 6966 4165
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4706 4128 4712 4140
rect 4663 4100 4712 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4706 4088 4712 4100
rect 4764 4128 4770 4140
rect 6086 4128 6092 4140
rect 4764 4100 6092 4128
rect 4764 4088 4770 4100
rect 6086 4088 6092 4100
rect 6144 4128 6150 4140
rect 6270 4128 6276 4140
rect 6144 4100 6276 4128
rect 6144 4088 6150 4100
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6638 4088 6644 4140
rect 6696 4088 6702 4140
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 4264 4032 4353 4060
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 4246 3992 4252 4004
rect 3620 3964 4252 3992
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 4448 3992 4476 4023
rect 4522 4020 4528 4072
rect 4580 4020 4586 4072
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 4614 3992 4620 4004
rect 4448 3964 4620 3992
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 4816 3924 4844 4023
rect 5718 3924 5724 3936
rect 4816 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6270 3924 6276 3936
rect 6227 3896 6276 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8294 3924 8300 3936
rect 8067 3896 8300 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 1104 3834 8740 3856
rect 1104 3782 1150 3834
rect 1202 3782 1214 3834
rect 1266 3782 1278 3834
rect 1330 3782 1342 3834
rect 1394 3782 1406 3834
rect 1458 3782 2470 3834
rect 2522 3782 2534 3834
rect 2586 3782 2598 3834
rect 2650 3782 2662 3834
rect 2714 3782 2726 3834
rect 2778 3782 3790 3834
rect 3842 3782 3854 3834
rect 3906 3782 3918 3834
rect 3970 3782 3982 3834
rect 4034 3782 4046 3834
rect 4098 3782 5110 3834
rect 5162 3782 5174 3834
rect 5226 3782 5238 3834
rect 5290 3782 5302 3834
rect 5354 3782 5366 3834
rect 5418 3782 6430 3834
rect 6482 3782 6494 3834
rect 6546 3782 6558 3834
rect 6610 3782 6622 3834
rect 6674 3782 6686 3834
rect 6738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 7942 3834
rect 7994 3782 8006 3834
rect 8058 3782 8740 3834
rect 1104 3760 8740 3782
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 3602 3720 3608 3732
rect 2924 3692 3608 3720
rect 2924 3680 2930 3692
rect 3602 3680 3608 3692
rect 3660 3720 3666 3732
rect 4430 3720 4436 3732
rect 3660 3692 3832 3720
rect 3660 3680 3666 3692
rect 3804 3593 3832 3692
rect 3988 3692 4436 3720
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2038 3516 2044 3528
rect 1995 3488 2044 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 2216 3451 2274 3457
rect 2216 3417 2228 3451
rect 2262 3448 2274 3451
rect 2406 3448 2412 3460
rect 2262 3420 2412 3448
rect 2262 3417 2274 3420
rect 2216 3411 2274 3417
rect 2406 3408 2412 3420
rect 2464 3408 2470 3460
rect 3804 3448 3832 3547
rect 3988 3525 4016 3692
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 4798 3720 4804 3732
rect 4663 3692 4804 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 4890 3680 4896 3732
rect 4948 3680 4954 3732
rect 6086 3680 6092 3732
rect 6144 3720 6150 3732
rect 6454 3720 6460 3732
rect 6144 3692 6460 3720
rect 6144 3680 6150 3692
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 4157 3655 4215 3661
rect 4157 3621 4169 3655
rect 4203 3652 4215 3655
rect 4246 3652 4252 3664
rect 4203 3624 4252 3652
rect 4203 3621 4215 3624
rect 4157 3615 4215 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 4709 3655 4767 3661
rect 4709 3621 4721 3655
rect 4755 3621 4767 3655
rect 4709 3615 4767 3621
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4154 3516 4160 3528
rect 4019 3488 4160 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4724 3516 4752 3615
rect 4480 3491 4752 3516
rect 4479 3488 4752 3491
rect 5169 3519 5227 3525
rect 4479 3485 4537 3488
rect 4249 3451 4307 3457
rect 4249 3448 4261 3451
rect 3804 3420 4261 3448
rect 4249 3417 4261 3420
rect 4295 3417 4307 3451
rect 4479 3451 4491 3485
rect 4525 3451 4537 3485
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5718 3516 5724 3528
rect 5215 3488 5724 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5718 3476 5724 3488
rect 5776 3516 5782 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 5776 3488 6653 3516
rect 5776 3476 5782 3488
rect 6641 3485 6653 3488
rect 6687 3516 6699 3519
rect 6730 3516 6736 3528
rect 6687 3488 6736 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 4479 3445 4537 3451
rect 4872 3451 4930 3457
rect 4249 3411 4307 3417
rect 4872 3417 4884 3451
rect 4918 3448 4930 3451
rect 4982 3448 4988 3460
rect 4918 3420 4988 3448
rect 4918 3417 4930 3420
rect 4872 3411 4930 3417
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 3329 3383 3387 3389
rect 3329 3380 3341 3383
rect 3108 3352 3341 3380
rect 3108 3340 3114 3352
rect 3329 3349 3341 3352
rect 3375 3349 3387 3383
rect 4264 3380 4292 3411
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 5077 3451 5135 3457
rect 5077 3417 5089 3451
rect 5123 3448 5135 3451
rect 5258 3448 5264 3460
rect 5123 3420 5264 3448
rect 5123 3417 5135 3420
rect 5077 3411 5135 3417
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 5436 3451 5494 3457
rect 5436 3417 5448 3451
rect 5482 3448 5494 3451
rect 5626 3448 5632 3460
rect 5482 3420 5632 3448
rect 5482 3417 5494 3420
rect 5436 3411 5494 3417
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 6362 3448 6368 3460
rect 6104 3420 6368 3448
rect 4614 3380 4620 3392
rect 4264 3352 4620 3380
rect 3329 3343 3387 3349
rect 4614 3340 4620 3352
rect 4672 3380 4678 3392
rect 6104 3380 6132 3420
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 6908 3451 6966 3457
rect 6908 3417 6920 3451
rect 6954 3448 6966 3451
rect 7650 3448 7656 3460
rect 6954 3420 7656 3448
rect 6954 3417 6966 3420
rect 6908 3411 6966 3417
rect 7650 3408 7656 3420
rect 7708 3408 7714 3460
rect 4672 3352 6132 3380
rect 4672 3340 4678 3352
rect 6178 3340 6184 3392
rect 6236 3380 6242 3392
rect 6549 3383 6607 3389
rect 6549 3380 6561 3383
rect 6236 3352 6561 3380
rect 6236 3340 6242 3352
rect 6549 3349 6561 3352
rect 6595 3380 6607 3383
rect 7558 3380 7564 3392
rect 6595 3352 7564 3380
rect 6595 3349 6607 3352
rect 6549 3343 6607 3349
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8018 3340 8024 3392
rect 8076 3340 8082 3392
rect 1104 3290 8740 3312
rect 1104 3238 1810 3290
rect 1862 3238 1874 3290
rect 1926 3238 1938 3290
rect 1990 3238 2002 3290
rect 2054 3238 2066 3290
rect 2118 3238 3130 3290
rect 3182 3238 3194 3290
rect 3246 3238 3258 3290
rect 3310 3238 3322 3290
rect 3374 3238 3386 3290
rect 3438 3238 4450 3290
rect 4502 3238 4514 3290
rect 4566 3238 4578 3290
rect 4630 3238 4642 3290
rect 4694 3238 4706 3290
rect 4758 3238 5770 3290
rect 5822 3238 5834 3290
rect 5886 3238 5898 3290
rect 5950 3238 5962 3290
rect 6014 3238 6026 3290
rect 6078 3238 7090 3290
rect 7142 3238 7154 3290
rect 7206 3238 7218 3290
rect 7270 3238 7282 3290
rect 7334 3238 7346 3290
rect 7398 3238 8410 3290
rect 8462 3238 8474 3290
rect 8526 3238 8538 3290
rect 8590 3238 8602 3290
rect 8654 3238 8666 3290
rect 8718 3238 8740 3290
rect 1104 3216 8740 3238
rect 2406 3136 2412 3188
rect 2464 3136 2470 3188
rect 4154 3136 4160 3188
rect 4212 3136 4218 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 5592 3148 6561 3176
rect 5592 3136 5598 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 6822 3176 6828 3188
rect 6687 3148 6828 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 1578 3068 1584 3120
rect 1636 3108 1642 3120
rect 3694 3108 3700 3120
rect 1636 3080 2912 3108
rect 1636 3068 1642 3080
rect 2884 3049 2912 3080
rect 3068 3080 3700 3108
rect 3068 3052 3096 3080
rect 3694 3068 3700 3080
rect 3752 3108 3758 3120
rect 5721 3111 5779 3117
rect 3752 3080 4016 3108
rect 3752 3068 3758 3080
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2869 3043 2927 3049
rect 2639 3012 2774 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2746 2836 2774 3012
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 2884 2972 2912 3003
rect 3050 3000 3056 3052
rect 3108 3000 3114 3052
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3602 3040 3608 3052
rect 3375 3012 3608 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 3988 3049 4016 3080
rect 5721 3077 5733 3111
rect 5767 3108 5779 3111
rect 6178 3108 6184 3120
rect 5767 3080 6184 3108
rect 5767 3077 5779 3080
rect 5721 3071 5779 3077
rect 6178 3068 6184 3080
rect 6236 3068 6242 3120
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5810 3040 5816 3052
rect 5040 3012 5816 3040
rect 5040 3000 5046 3012
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6454 3040 6460 3052
rect 5960 3012 6460 3040
rect 5960 3000 5966 3012
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 3145 2975 3203 2981
rect 3145 2972 3157 2975
rect 2884 2944 3157 2972
rect 3145 2941 3157 2944
rect 3191 2941 3203 2975
rect 3145 2935 3203 2941
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 3559 2944 3801 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 5828 2972 5856 3000
rect 6270 2972 6276 2984
rect 5828 2944 6276 2972
rect 3789 2935 3847 2941
rect 2958 2864 2964 2916
rect 3016 2904 3022 2916
rect 3528 2904 3556 2935
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 3016 2876 3556 2904
rect 3016 2864 3022 2876
rect 5626 2864 5632 2916
rect 5684 2904 5690 2916
rect 5902 2904 5908 2916
rect 5684 2876 5908 2904
rect 5684 2864 5690 2876
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6089 2907 6147 2913
rect 6089 2873 6101 2907
rect 6135 2873 6147 2907
rect 6564 2904 6592 3139
rect 6822 3136 6828 3148
rect 6880 3176 6886 3188
rect 7282 3176 7288 3188
rect 6880 3148 7288 3176
rect 6880 3136 6886 3148
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7561 3179 7619 3185
rect 7561 3176 7573 3179
rect 7524 3148 7573 3176
rect 7524 3136 7530 3148
rect 7561 3145 7573 3148
rect 7607 3145 7619 3179
rect 7561 3139 7619 3145
rect 6917 3111 6975 3117
rect 6917 3077 6929 3111
rect 6963 3108 6975 3111
rect 8294 3108 8300 3120
rect 6963 3080 8300 3108
rect 6963 3077 6975 3080
rect 6917 3071 6975 3077
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 7116 3049 7144 3080
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6696 3012 6745 3040
rect 6696 3000 6702 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 6748 2972 6776 3003
rect 8018 3000 8024 3052
rect 8076 3000 8082 3052
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 6748 2944 7205 2972
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 7282 2932 7288 2984
rect 7340 2932 7346 2984
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 7392 2904 7420 2935
rect 7650 2932 7656 2984
rect 7708 2932 7714 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7760 2944 7941 2972
rect 6564 2876 7420 2904
rect 6089 2867 6147 2873
rect 4246 2836 4252 2848
rect 2746 2808 4252 2836
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 6104 2836 6132 2867
rect 5500 2808 6132 2836
rect 6365 2839 6423 2845
rect 5500 2796 5506 2808
rect 6365 2805 6377 2839
rect 6411 2836 6423 2839
rect 7006 2836 7012 2848
rect 6411 2808 7012 2836
rect 6411 2805 6423 2808
rect 6365 2799 6423 2805
rect 7006 2796 7012 2808
rect 7064 2836 7070 2848
rect 7760 2836 7788 2944
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 7064 2808 7788 2836
rect 7064 2796 7070 2808
rect 1104 2746 8740 2768
rect 1104 2694 1150 2746
rect 1202 2694 1214 2746
rect 1266 2694 1278 2746
rect 1330 2694 1342 2746
rect 1394 2694 1406 2746
rect 1458 2694 2470 2746
rect 2522 2694 2534 2746
rect 2586 2694 2598 2746
rect 2650 2694 2662 2746
rect 2714 2694 2726 2746
rect 2778 2694 3790 2746
rect 3842 2694 3854 2746
rect 3906 2694 3918 2746
rect 3970 2694 3982 2746
rect 4034 2694 4046 2746
rect 4098 2694 5110 2746
rect 5162 2694 5174 2746
rect 5226 2694 5238 2746
rect 5290 2694 5302 2746
rect 5354 2694 5366 2746
rect 5418 2694 6430 2746
rect 6482 2694 6494 2746
rect 6546 2694 6558 2746
rect 6610 2694 6622 2746
rect 6674 2694 6686 2746
rect 6738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 7942 2746
rect 7994 2694 8006 2746
rect 8058 2694 8740 2746
rect 1104 2672 8740 2694
rect 8113 2567 8171 2573
rect 8113 2533 8125 2567
rect 8159 2564 8171 2567
rect 9030 2564 9036 2576
rect 8159 2536 9036 2564
rect 8159 2533 8171 2536
rect 8113 2527 8171 2533
rect 9030 2524 9036 2536
rect 9088 2524 9094 2576
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1544 2400 1593 2428
rect 1544 2388 1550 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 1728 2400 1961 2428
rect 1728 2388 1734 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 2958 2428 2964 2440
rect 2915 2400 2964 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3694 2388 3700 2440
rect 3752 2428 3758 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3752 2400 3985 2428
rect 3752 2388 3758 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5442 2428 5448 2440
rect 4755 2400 5448 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5626 2388 5632 2440
rect 5684 2388 5690 2440
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5868 2400 6561 2428
rect 5868 2388 5874 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7558 2428 7564 2440
rect 7515 2400 7564 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8110 2428 8116 2440
rect 7975 2400 8116 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8352 2400 8401 2428
rect 8352 2388 8358 2400
rect 8389 2397 8401 2400
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 750 2252 756 2304
rect 808 2292 814 2304
rect 1397 2295 1455 2301
rect 1397 2292 1409 2295
rect 808 2264 1409 2292
rect 808 2252 814 2264
rect 1397 2261 1409 2264
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 1670 2252 1676 2304
rect 1728 2292 1734 2304
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 1728 2264 1777 2292
rect 1728 2252 1734 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 1765 2255 1823 2261
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 2685 2295 2743 2301
rect 2685 2292 2697 2295
rect 2648 2264 2697 2292
rect 2648 2252 2654 2264
rect 2685 2261 2697 2264
rect 2731 2261 2743 2295
rect 2685 2255 2743 2261
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3568 2264 3801 2292
rect 3568 2252 3574 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 4338 2252 4344 2304
rect 4396 2292 4402 2304
rect 4525 2295 4583 2301
rect 4525 2292 4537 2295
rect 4396 2264 4537 2292
rect 4396 2252 4402 2264
rect 4525 2261 4537 2264
rect 4571 2261 4583 2295
rect 4525 2255 4583 2261
rect 5350 2252 5356 2304
rect 5408 2292 5414 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5408 2264 5457 2292
rect 5408 2252 5414 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6270 2252 6276 2304
rect 6328 2292 6334 2304
rect 6365 2295 6423 2301
rect 6365 2292 6377 2295
rect 6328 2264 6377 2292
rect 6328 2252 6334 2264
rect 6365 2261 6377 2264
rect 6411 2261 6423 2295
rect 6365 2255 6423 2261
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7064 2264 7297 2292
rect 7064 2252 7070 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 8202 2252 8208 2304
rect 8260 2252 8266 2304
rect 1104 2202 8740 2224
rect 1104 2150 1810 2202
rect 1862 2150 1874 2202
rect 1926 2150 1938 2202
rect 1990 2150 2002 2202
rect 2054 2150 2066 2202
rect 2118 2150 3130 2202
rect 3182 2150 3194 2202
rect 3246 2150 3258 2202
rect 3310 2150 3322 2202
rect 3374 2150 3386 2202
rect 3438 2150 4450 2202
rect 4502 2150 4514 2202
rect 4566 2150 4578 2202
rect 4630 2150 4642 2202
rect 4694 2150 4706 2202
rect 4758 2150 5770 2202
rect 5822 2150 5834 2202
rect 5886 2150 5898 2202
rect 5950 2150 5962 2202
rect 6014 2150 6026 2202
rect 6078 2150 7090 2202
rect 7142 2150 7154 2202
rect 7206 2150 7218 2202
rect 7270 2150 7282 2202
rect 7334 2150 7346 2202
rect 7398 2150 8410 2202
rect 8462 2150 8474 2202
rect 8526 2150 8538 2202
rect 8590 2150 8602 2202
rect 8654 2150 8666 2202
rect 8718 2150 8740 2202
rect 1104 2128 8740 2150
<< via1 >>
rect 1810 9766 1862 9818
rect 1874 9766 1926 9818
rect 1938 9766 1990 9818
rect 2002 9766 2054 9818
rect 2066 9766 2118 9818
rect 3130 9766 3182 9818
rect 3194 9766 3246 9818
rect 3258 9766 3310 9818
rect 3322 9766 3374 9818
rect 3386 9766 3438 9818
rect 4450 9766 4502 9818
rect 4514 9766 4566 9818
rect 4578 9766 4630 9818
rect 4642 9766 4694 9818
rect 4706 9766 4758 9818
rect 5770 9766 5822 9818
rect 5834 9766 5886 9818
rect 5898 9766 5950 9818
rect 5962 9766 6014 9818
rect 6026 9766 6078 9818
rect 7090 9766 7142 9818
rect 7154 9766 7206 9818
rect 7218 9766 7270 9818
rect 7282 9766 7334 9818
rect 7346 9766 7398 9818
rect 8410 9766 8462 9818
rect 8474 9766 8526 9818
rect 8538 9766 8590 9818
rect 8602 9766 8654 9818
rect 8666 9766 8718 9818
rect 2412 9528 2464 9580
rect 2136 9324 2188 9376
rect 1150 9222 1202 9274
rect 1214 9222 1266 9274
rect 1278 9222 1330 9274
rect 1342 9222 1394 9274
rect 1406 9222 1458 9274
rect 2470 9222 2522 9274
rect 2534 9222 2586 9274
rect 2598 9222 2650 9274
rect 2662 9222 2714 9274
rect 2726 9222 2778 9274
rect 3790 9222 3842 9274
rect 3854 9222 3906 9274
rect 3918 9222 3970 9274
rect 3982 9222 4034 9274
rect 4046 9222 4098 9274
rect 5110 9222 5162 9274
rect 5174 9222 5226 9274
rect 5238 9222 5290 9274
rect 5302 9222 5354 9274
rect 5366 9222 5418 9274
rect 6430 9222 6482 9274
rect 6494 9222 6546 9274
rect 6558 9222 6610 9274
rect 6622 9222 6674 9274
rect 6686 9222 6738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 7942 9222 7994 9274
rect 8006 9222 8058 9274
rect 1810 8678 1862 8730
rect 1874 8678 1926 8730
rect 1938 8678 1990 8730
rect 2002 8678 2054 8730
rect 2066 8678 2118 8730
rect 3130 8678 3182 8730
rect 3194 8678 3246 8730
rect 3258 8678 3310 8730
rect 3322 8678 3374 8730
rect 3386 8678 3438 8730
rect 4450 8678 4502 8730
rect 4514 8678 4566 8730
rect 4578 8678 4630 8730
rect 4642 8678 4694 8730
rect 4706 8678 4758 8730
rect 5770 8678 5822 8730
rect 5834 8678 5886 8730
rect 5898 8678 5950 8730
rect 5962 8678 6014 8730
rect 6026 8678 6078 8730
rect 7090 8678 7142 8730
rect 7154 8678 7206 8730
rect 7218 8678 7270 8730
rect 7282 8678 7334 8730
rect 7346 8678 7398 8730
rect 8410 8678 8462 8730
rect 8474 8678 8526 8730
rect 8538 8678 8590 8730
rect 8602 8678 8654 8730
rect 8666 8678 8718 8730
rect 1584 8440 1636 8492
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2872 8304 2924 8356
rect 1150 8134 1202 8186
rect 1214 8134 1266 8186
rect 1278 8134 1330 8186
rect 1342 8134 1394 8186
rect 1406 8134 1458 8186
rect 2470 8134 2522 8186
rect 2534 8134 2586 8186
rect 2598 8134 2650 8186
rect 2662 8134 2714 8186
rect 2726 8134 2778 8186
rect 3790 8134 3842 8186
rect 3854 8134 3906 8186
rect 3918 8134 3970 8186
rect 3982 8134 4034 8186
rect 4046 8134 4098 8186
rect 5110 8134 5162 8186
rect 5174 8134 5226 8186
rect 5238 8134 5290 8186
rect 5302 8134 5354 8186
rect 5366 8134 5418 8186
rect 6430 8134 6482 8186
rect 6494 8134 6546 8186
rect 6558 8134 6610 8186
rect 6622 8134 6674 8186
rect 6686 8134 6738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 7942 8134 7994 8186
rect 8006 8134 8058 8186
rect 2228 7828 2280 7880
rect 2872 7760 2924 7812
rect 1584 7692 1636 7744
rect 1810 7590 1862 7642
rect 1874 7590 1926 7642
rect 1938 7590 1990 7642
rect 2002 7590 2054 7642
rect 2066 7590 2118 7642
rect 3130 7590 3182 7642
rect 3194 7590 3246 7642
rect 3258 7590 3310 7642
rect 3322 7590 3374 7642
rect 3386 7590 3438 7642
rect 4450 7590 4502 7642
rect 4514 7590 4566 7642
rect 4578 7590 4630 7642
rect 4642 7590 4694 7642
rect 4706 7590 4758 7642
rect 5770 7590 5822 7642
rect 5834 7590 5886 7642
rect 5898 7590 5950 7642
rect 5962 7590 6014 7642
rect 6026 7590 6078 7642
rect 7090 7590 7142 7642
rect 7154 7590 7206 7642
rect 7218 7590 7270 7642
rect 7282 7590 7334 7642
rect 7346 7590 7398 7642
rect 8410 7590 8462 7642
rect 8474 7590 8526 7642
rect 8538 7590 8590 7642
rect 8602 7590 8654 7642
rect 8666 7590 8718 7642
rect 3056 7488 3108 7540
rect 2136 7420 2188 7472
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 1676 7216 1728 7268
rect 2964 7395 3016 7404
rect 2964 7361 2982 7395
rect 2982 7361 3016 7395
rect 2964 7352 3016 7361
rect 2228 7148 2280 7200
rect 1150 7046 1202 7098
rect 1214 7046 1266 7098
rect 1278 7046 1330 7098
rect 1342 7046 1394 7098
rect 1406 7046 1458 7098
rect 2470 7046 2522 7098
rect 2534 7046 2586 7098
rect 2598 7046 2650 7098
rect 2662 7046 2714 7098
rect 2726 7046 2778 7098
rect 3790 7046 3842 7098
rect 3854 7046 3906 7098
rect 3918 7046 3970 7098
rect 3982 7046 4034 7098
rect 4046 7046 4098 7098
rect 5110 7046 5162 7098
rect 5174 7046 5226 7098
rect 5238 7046 5290 7098
rect 5302 7046 5354 7098
rect 5366 7046 5418 7098
rect 6430 7046 6482 7098
rect 6494 7046 6546 7098
rect 6558 7046 6610 7098
rect 6622 7046 6674 7098
rect 6686 7046 6738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 7942 7046 7994 7098
rect 8006 7046 8058 7098
rect 1676 6944 1728 6996
rect 2964 6944 3016 6996
rect 2872 6808 2924 6860
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 1492 6672 1544 6724
rect 2136 6604 2188 6656
rect 1810 6502 1862 6554
rect 1874 6502 1926 6554
rect 1938 6502 1990 6554
rect 2002 6502 2054 6554
rect 2066 6502 2118 6554
rect 3130 6502 3182 6554
rect 3194 6502 3246 6554
rect 3258 6502 3310 6554
rect 3322 6502 3374 6554
rect 3386 6502 3438 6554
rect 4450 6502 4502 6554
rect 4514 6502 4566 6554
rect 4578 6502 4630 6554
rect 4642 6502 4694 6554
rect 4706 6502 4758 6554
rect 5770 6502 5822 6554
rect 5834 6502 5886 6554
rect 5898 6502 5950 6554
rect 5962 6502 6014 6554
rect 6026 6502 6078 6554
rect 7090 6502 7142 6554
rect 7154 6502 7206 6554
rect 7218 6502 7270 6554
rect 7282 6502 7334 6554
rect 7346 6502 7398 6554
rect 8410 6502 8462 6554
rect 8474 6502 8526 6554
rect 8538 6502 8590 6554
rect 8602 6502 8654 6554
rect 8666 6502 8718 6554
rect 1150 5958 1202 6010
rect 1214 5958 1266 6010
rect 1278 5958 1330 6010
rect 1342 5958 1394 6010
rect 1406 5958 1458 6010
rect 2470 5958 2522 6010
rect 2534 5958 2586 6010
rect 2598 5958 2650 6010
rect 2662 5958 2714 6010
rect 2726 5958 2778 6010
rect 3790 5958 3842 6010
rect 3854 5958 3906 6010
rect 3918 5958 3970 6010
rect 3982 5958 4034 6010
rect 4046 5958 4098 6010
rect 5110 5958 5162 6010
rect 5174 5958 5226 6010
rect 5238 5958 5290 6010
rect 5302 5958 5354 6010
rect 5366 5958 5418 6010
rect 6430 5958 6482 6010
rect 6494 5958 6546 6010
rect 6558 5958 6610 6010
rect 6622 5958 6674 6010
rect 6686 5958 6738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 7942 5958 7994 6010
rect 8006 5958 8058 6010
rect 2228 5899 2280 5908
rect 2228 5865 2237 5899
rect 2237 5865 2271 5899
rect 2271 5865 2280 5899
rect 2228 5856 2280 5865
rect 6828 5652 6880 5704
rect 5448 5516 5500 5568
rect 1810 5414 1862 5466
rect 1874 5414 1926 5466
rect 1938 5414 1990 5466
rect 2002 5414 2054 5466
rect 2066 5414 2118 5466
rect 3130 5414 3182 5466
rect 3194 5414 3246 5466
rect 3258 5414 3310 5466
rect 3322 5414 3374 5466
rect 3386 5414 3438 5466
rect 4450 5414 4502 5466
rect 4514 5414 4566 5466
rect 4578 5414 4630 5466
rect 4642 5414 4694 5466
rect 4706 5414 4758 5466
rect 5770 5414 5822 5466
rect 5834 5414 5886 5466
rect 5898 5414 5950 5466
rect 5962 5414 6014 5466
rect 6026 5414 6078 5466
rect 7090 5414 7142 5466
rect 7154 5414 7206 5466
rect 7218 5414 7270 5466
rect 7282 5414 7334 5466
rect 7346 5414 7398 5466
rect 8410 5414 8462 5466
rect 8474 5414 8526 5466
rect 8538 5414 8590 5466
rect 8602 5414 8654 5466
rect 8666 5414 8718 5466
rect 6276 5312 6328 5364
rect 5816 5244 5868 5296
rect 6092 5176 6144 5228
rect 6828 5176 6880 5228
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 4160 5083 4212 5092
rect 4160 5049 4169 5083
rect 4169 5049 4203 5083
rect 4203 5049 4212 5083
rect 4160 5040 4212 5049
rect 5816 5083 5868 5092
rect 5816 5049 5825 5083
rect 5825 5049 5859 5083
rect 5859 5049 5868 5083
rect 5816 5040 5868 5049
rect 6000 5040 6052 5092
rect 4436 4972 4488 5024
rect 7472 4972 7524 5024
rect 7564 5015 7616 5024
rect 7564 4981 7573 5015
rect 7573 4981 7607 5015
rect 7607 4981 7616 5015
rect 7564 4972 7616 4981
rect 1150 4870 1202 4922
rect 1214 4870 1266 4922
rect 1278 4870 1330 4922
rect 1342 4870 1394 4922
rect 1406 4870 1458 4922
rect 2470 4870 2522 4922
rect 2534 4870 2586 4922
rect 2598 4870 2650 4922
rect 2662 4870 2714 4922
rect 2726 4870 2778 4922
rect 3790 4870 3842 4922
rect 3854 4870 3906 4922
rect 3918 4870 3970 4922
rect 3982 4870 4034 4922
rect 4046 4870 4098 4922
rect 5110 4870 5162 4922
rect 5174 4870 5226 4922
rect 5238 4870 5290 4922
rect 5302 4870 5354 4922
rect 5366 4870 5418 4922
rect 6430 4870 6482 4922
rect 6494 4870 6546 4922
rect 6558 4870 6610 4922
rect 6622 4870 6674 4922
rect 6686 4870 6738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 7942 4870 7994 4922
rect 8006 4870 8058 4922
rect 2872 4768 2924 4820
rect 6092 4768 6144 4820
rect 3516 4700 3568 4752
rect 5448 4700 5500 4752
rect 6000 4700 6052 4752
rect 2228 4675 2280 4684
rect 2228 4641 2237 4675
rect 2237 4641 2271 4675
rect 2271 4641 2280 4675
rect 2228 4632 2280 4641
rect 2964 4564 3016 4616
rect 4896 4632 4948 4684
rect 6184 4632 6236 4684
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 4804 4564 4856 4616
rect 1400 4428 1452 4480
rect 3056 4496 3108 4548
rect 5632 4564 5684 4616
rect 2872 4428 2924 4480
rect 4252 4428 4304 4480
rect 4896 4471 4948 4480
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 4896 4428 4948 4437
rect 5540 4428 5592 4480
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 5724 4428 5776 4480
rect 6644 4428 6696 4480
rect 1810 4326 1862 4378
rect 1874 4326 1926 4378
rect 1938 4326 1990 4378
rect 2002 4326 2054 4378
rect 2066 4326 2118 4378
rect 3130 4326 3182 4378
rect 3194 4326 3246 4378
rect 3258 4326 3310 4378
rect 3322 4326 3374 4378
rect 3386 4326 3438 4378
rect 4450 4326 4502 4378
rect 4514 4326 4566 4378
rect 4578 4326 4630 4378
rect 4642 4326 4694 4378
rect 4706 4326 4758 4378
rect 5770 4326 5822 4378
rect 5834 4326 5886 4378
rect 5898 4326 5950 4378
rect 5962 4326 6014 4378
rect 6026 4326 6078 4378
rect 7090 4326 7142 4378
rect 7154 4326 7206 4378
rect 7218 4326 7270 4378
rect 7282 4326 7334 4378
rect 7346 4326 7398 4378
rect 8410 4326 8462 4378
rect 8474 4326 8526 4378
rect 8538 4326 8590 4378
rect 8602 4326 8654 4378
rect 8666 4326 8718 4378
rect 2964 4224 3016 4276
rect 4436 4224 4488 4276
rect 6828 4224 6880 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 2044 4156 2096 4208
rect 2228 4156 2280 4208
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 3056 4020 3108 4072
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 4896 4156 4948 4208
rect 7564 4156 7616 4208
rect 4712 4088 4764 4140
rect 6092 4088 6144 4140
rect 6276 4088 6328 4140
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 4252 3952 4304 4004
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 4620 3952 4672 4004
rect 5724 3884 5776 3936
rect 6276 3884 6328 3936
rect 8300 3884 8352 3936
rect 1150 3782 1202 3834
rect 1214 3782 1266 3834
rect 1278 3782 1330 3834
rect 1342 3782 1394 3834
rect 1406 3782 1458 3834
rect 2470 3782 2522 3834
rect 2534 3782 2586 3834
rect 2598 3782 2650 3834
rect 2662 3782 2714 3834
rect 2726 3782 2778 3834
rect 3790 3782 3842 3834
rect 3854 3782 3906 3834
rect 3918 3782 3970 3834
rect 3982 3782 4034 3834
rect 4046 3782 4098 3834
rect 5110 3782 5162 3834
rect 5174 3782 5226 3834
rect 5238 3782 5290 3834
rect 5302 3782 5354 3834
rect 5366 3782 5418 3834
rect 6430 3782 6482 3834
rect 6494 3782 6546 3834
rect 6558 3782 6610 3834
rect 6622 3782 6674 3834
rect 6686 3782 6738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 7942 3782 7994 3834
rect 8006 3782 8058 3834
rect 2872 3680 2924 3732
rect 3608 3680 3660 3732
rect 4436 3723 4488 3732
rect 2044 3476 2096 3528
rect 2412 3408 2464 3460
rect 4436 3689 4445 3723
rect 4445 3689 4479 3723
rect 4479 3689 4488 3723
rect 4436 3680 4488 3689
rect 4804 3680 4856 3732
rect 4896 3723 4948 3732
rect 4896 3689 4905 3723
rect 4905 3689 4939 3723
rect 4939 3689 4948 3723
rect 4896 3680 4948 3689
rect 6092 3680 6144 3732
rect 6460 3680 6512 3732
rect 4252 3612 4304 3664
rect 4160 3476 4212 3528
rect 5724 3476 5776 3528
rect 6736 3476 6788 3528
rect 3056 3340 3108 3392
rect 4988 3408 5040 3460
rect 5264 3408 5316 3460
rect 5632 3408 5684 3460
rect 4620 3340 4672 3392
rect 6368 3408 6420 3460
rect 7656 3408 7708 3460
rect 6184 3340 6236 3392
rect 7564 3340 7616 3392
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 1810 3238 1862 3290
rect 1874 3238 1926 3290
rect 1938 3238 1990 3290
rect 2002 3238 2054 3290
rect 2066 3238 2118 3290
rect 3130 3238 3182 3290
rect 3194 3238 3246 3290
rect 3258 3238 3310 3290
rect 3322 3238 3374 3290
rect 3386 3238 3438 3290
rect 4450 3238 4502 3290
rect 4514 3238 4566 3290
rect 4578 3238 4630 3290
rect 4642 3238 4694 3290
rect 4706 3238 4758 3290
rect 5770 3238 5822 3290
rect 5834 3238 5886 3290
rect 5898 3238 5950 3290
rect 5962 3238 6014 3290
rect 6026 3238 6078 3290
rect 7090 3238 7142 3290
rect 7154 3238 7206 3290
rect 7218 3238 7270 3290
rect 7282 3238 7334 3290
rect 7346 3238 7398 3290
rect 8410 3238 8462 3290
rect 8474 3238 8526 3290
rect 8538 3238 8590 3290
rect 8602 3238 8654 3290
rect 8666 3238 8718 3290
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 4160 3179 4212 3188
rect 4160 3145 4169 3179
rect 4169 3145 4203 3179
rect 4203 3145 4212 3179
rect 4160 3136 4212 3145
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 1584 3068 1636 3120
rect 3700 3068 3752 3120
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3608 3000 3660 3052
rect 6184 3068 6236 3120
rect 4988 3000 5040 3052
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 6460 3000 6512 3052
rect 2964 2864 3016 2916
rect 6276 2932 6328 2984
rect 5632 2864 5684 2916
rect 5908 2864 5960 2916
rect 6828 3136 6880 3188
rect 7288 3136 7340 3188
rect 7472 3136 7524 3188
rect 6644 3000 6696 3052
rect 8300 3068 8352 3120
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 7656 2975 7708 2984
rect 7656 2941 7665 2975
rect 7665 2941 7699 2975
rect 7699 2941 7708 2975
rect 7656 2932 7708 2941
rect 4252 2796 4304 2848
rect 5448 2796 5500 2848
rect 7012 2796 7064 2848
rect 1150 2694 1202 2746
rect 1214 2694 1266 2746
rect 1278 2694 1330 2746
rect 1342 2694 1394 2746
rect 1406 2694 1458 2746
rect 2470 2694 2522 2746
rect 2534 2694 2586 2746
rect 2598 2694 2650 2746
rect 2662 2694 2714 2746
rect 2726 2694 2778 2746
rect 3790 2694 3842 2746
rect 3854 2694 3906 2746
rect 3918 2694 3970 2746
rect 3982 2694 4034 2746
rect 4046 2694 4098 2746
rect 5110 2694 5162 2746
rect 5174 2694 5226 2746
rect 5238 2694 5290 2746
rect 5302 2694 5354 2746
rect 5366 2694 5418 2746
rect 6430 2694 6482 2746
rect 6494 2694 6546 2746
rect 6558 2694 6610 2746
rect 6622 2694 6674 2746
rect 6686 2694 6738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 7942 2694 7994 2746
rect 8006 2694 8058 2746
rect 9036 2524 9088 2576
rect 1492 2388 1544 2440
rect 1676 2388 1728 2440
rect 2964 2388 3016 2440
rect 3700 2388 3752 2440
rect 5448 2388 5500 2440
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 5816 2388 5868 2440
rect 7564 2388 7616 2440
rect 8116 2388 8168 2440
rect 8300 2388 8352 2440
rect 756 2252 808 2304
rect 1676 2252 1728 2304
rect 2596 2252 2648 2304
rect 3516 2252 3568 2304
rect 4344 2252 4396 2304
rect 5356 2252 5408 2304
rect 6276 2252 6328 2304
rect 7012 2252 7064 2304
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 1810 2150 1862 2202
rect 1874 2150 1926 2202
rect 1938 2150 1990 2202
rect 2002 2150 2054 2202
rect 2066 2150 2118 2202
rect 3130 2150 3182 2202
rect 3194 2150 3246 2202
rect 3258 2150 3310 2202
rect 3322 2150 3374 2202
rect 3386 2150 3438 2202
rect 4450 2150 4502 2202
rect 4514 2150 4566 2202
rect 4578 2150 4630 2202
rect 4642 2150 4694 2202
rect 4706 2150 4758 2202
rect 5770 2150 5822 2202
rect 5834 2150 5886 2202
rect 5898 2150 5950 2202
rect 5962 2150 6014 2202
rect 6026 2150 6078 2202
rect 7090 2150 7142 2202
rect 7154 2150 7206 2202
rect 7218 2150 7270 2202
rect 7282 2150 7334 2202
rect 7346 2150 7398 2202
rect 8410 2150 8462 2202
rect 8474 2150 8526 2202
rect 8538 2150 8590 2202
rect 8602 2150 8654 2202
rect 8666 2150 8718 2202
<< metal2 >>
rect 2410 10086 2466 10886
rect 1810 9820 2118 9829
rect 1810 9818 1816 9820
rect 1872 9818 1896 9820
rect 1952 9818 1976 9820
rect 2032 9818 2056 9820
rect 2112 9818 2118 9820
rect 1872 9766 1874 9818
rect 2054 9766 2056 9818
rect 1810 9764 1816 9766
rect 1872 9764 1896 9766
rect 1952 9764 1976 9766
rect 2032 9764 2056 9766
rect 2112 9764 2118 9766
rect 1810 9755 2118 9764
rect 2424 9586 2452 10086
rect 6918 9990 6974 10790
rect 6918 9976 6960 9990
rect 3130 9820 3438 9829
rect 3130 9818 3136 9820
rect 3192 9818 3216 9820
rect 3272 9818 3296 9820
rect 3352 9818 3376 9820
rect 3432 9818 3438 9820
rect 3192 9766 3194 9818
rect 3374 9766 3376 9818
rect 3130 9764 3136 9766
rect 3192 9764 3216 9766
rect 3272 9764 3296 9766
rect 3352 9764 3376 9766
rect 3432 9764 3438 9766
rect 3130 9755 3438 9764
rect 4450 9820 4758 9829
rect 4450 9818 4456 9820
rect 4512 9818 4536 9820
rect 4592 9818 4616 9820
rect 4672 9818 4696 9820
rect 4752 9818 4758 9820
rect 4512 9766 4514 9818
rect 4694 9766 4696 9818
rect 4450 9764 4456 9766
rect 4512 9764 4536 9766
rect 4592 9764 4616 9766
rect 4672 9764 4696 9766
rect 4752 9764 4758 9766
rect 4450 9755 4758 9764
rect 5770 9820 6078 9829
rect 5770 9818 5776 9820
rect 5832 9818 5856 9820
rect 5912 9818 5936 9820
rect 5992 9818 6016 9820
rect 6072 9818 6078 9820
rect 5832 9766 5834 9818
rect 6014 9766 6016 9818
rect 5770 9764 5776 9766
rect 5832 9764 5856 9766
rect 5912 9764 5936 9766
rect 5992 9764 6016 9766
rect 6072 9764 6078 9766
rect 5770 9755 6078 9764
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1150 9276 1458 9285
rect 1150 9274 1156 9276
rect 1212 9274 1236 9276
rect 1292 9274 1316 9276
rect 1372 9274 1396 9276
rect 1452 9274 1458 9276
rect 1212 9222 1214 9274
rect 1394 9222 1396 9274
rect 1150 9220 1156 9222
rect 1212 9220 1236 9222
rect 1292 9220 1316 9222
rect 1372 9220 1396 9222
rect 1452 9220 1458 9222
rect 1150 9211 1458 9220
rect 1810 8732 2118 8741
rect 1810 8730 1816 8732
rect 1872 8730 1896 8732
rect 1952 8730 1976 8732
rect 2032 8730 2056 8732
rect 2112 8730 2118 8732
rect 1872 8678 1874 8730
rect 2054 8678 2056 8730
rect 1810 8676 1816 8678
rect 1872 8676 1896 8678
rect 1952 8676 1976 8678
rect 2032 8676 2056 8678
rect 2112 8676 2118 8678
rect 1810 8667 2118 8676
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1150 8188 1458 8197
rect 1150 8186 1156 8188
rect 1212 8186 1236 8188
rect 1292 8186 1316 8188
rect 1372 8186 1396 8188
rect 1452 8186 1458 8188
rect 1212 8134 1214 8186
rect 1394 8134 1396 8186
rect 1150 8132 1156 8134
rect 1212 8132 1236 8134
rect 1292 8132 1316 8134
rect 1372 8132 1396 8134
rect 1452 8132 1458 8134
rect 1150 8123 1458 8132
rect 1596 7750 1624 8434
rect 2148 8430 2176 9318
rect 2470 9276 2778 9285
rect 2470 9274 2476 9276
rect 2532 9274 2556 9276
rect 2612 9274 2636 9276
rect 2692 9274 2716 9276
rect 2772 9274 2778 9276
rect 2532 9222 2534 9274
rect 2714 9222 2716 9274
rect 2470 9220 2476 9222
rect 2532 9220 2556 9222
rect 2612 9220 2636 9222
rect 2692 9220 2716 9222
rect 2772 9220 2778 9222
rect 2470 9211 2778 9220
rect 3790 9276 4098 9285
rect 3790 9274 3796 9276
rect 3852 9274 3876 9276
rect 3932 9274 3956 9276
rect 4012 9274 4036 9276
rect 4092 9274 4098 9276
rect 3852 9222 3854 9274
rect 4034 9222 4036 9274
rect 3790 9220 3796 9222
rect 3852 9220 3876 9222
rect 3932 9220 3956 9222
rect 4012 9220 4036 9222
rect 4092 9220 4098 9222
rect 3790 9211 4098 9220
rect 5110 9276 5418 9285
rect 5110 9274 5116 9276
rect 5172 9274 5196 9276
rect 5252 9274 5276 9276
rect 5332 9274 5356 9276
rect 5412 9274 5418 9276
rect 5172 9222 5174 9274
rect 5354 9222 5356 9274
rect 5110 9220 5116 9222
rect 5172 9220 5196 9222
rect 5252 9220 5276 9222
rect 5332 9220 5356 9222
rect 5412 9220 5418 9222
rect 5110 9211 5418 9220
rect 6430 9276 6738 9285
rect 6430 9274 6436 9276
rect 6492 9274 6516 9276
rect 6572 9274 6596 9276
rect 6652 9274 6676 9276
rect 6732 9274 6738 9276
rect 6492 9222 6494 9274
rect 6674 9222 6676 9274
rect 6430 9220 6436 9222
rect 6492 9220 6516 9222
rect 6572 9220 6596 9222
rect 6652 9220 6676 9222
rect 6732 9220 6738 9222
rect 6430 9211 6738 9220
rect 3130 8732 3438 8741
rect 3130 8730 3136 8732
rect 3192 8730 3216 8732
rect 3272 8730 3296 8732
rect 3352 8730 3376 8732
rect 3432 8730 3438 8732
rect 3192 8678 3194 8730
rect 3374 8678 3376 8730
rect 3130 8676 3136 8678
rect 3192 8676 3216 8678
rect 3272 8676 3296 8678
rect 3352 8676 3376 8678
rect 3432 8676 3438 8678
rect 3130 8667 3438 8676
rect 4450 8732 4758 8741
rect 4450 8730 4456 8732
rect 4512 8730 4536 8732
rect 4592 8730 4616 8732
rect 4672 8730 4696 8732
rect 4752 8730 4758 8732
rect 4512 8678 4514 8730
rect 4694 8678 4696 8730
rect 4450 8676 4456 8678
rect 4512 8676 4536 8678
rect 4592 8676 4616 8678
rect 4672 8676 4696 8678
rect 4752 8676 4758 8678
rect 4450 8667 4758 8676
rect 5770 8732 6078 8741
rect 5770 8730 5776 8732
rect 5832 8730 5856 8732
rect 5912 8730 5936 8732
rect 5992 8730 6016 8732
rect 6072 8730 6078 8732
rect 5832 8678 5834 8730
rect 6014 8678 6016 8730
rect 5770 8676 5776 8678
rect 5832 8676 5856 8678
rect 5912 8676 5936 8678
rect 5992 8676 6016 8678
rect 6072 8676 6078 8678
rect 5770 8667 6078 8676
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7410 1624 7686
rect 1810 7644 2118 7653
rect 1810 7642 1816 7644
rect 1872 7642 1896 7644
rect 1952 7642 1976 7644
rect 2032 7642 2056 7644
rect 2112 7642 2118 7644
rect 1872 7590 1874 7642
rect 2054 7590 2056 7642
rect 1810 7588 1816 7590
rect 1872 7588 1896 7590
rect 1952 7588 1976 7590
rect 2032 7588 2056 7590
rect 2112 7588 2118 7590
rect 1810 7579 2118 7588
rect 2148 7478 2176 8366
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2470 8188 2778 8197
rect 2470 8186 2476 8188
rect 2532 8186 2556 8188
rect 2612 8186 2636 8188
rect 2692 8186 2716 8188
rect 2772 8186 2778 8188
rect 2532 8134 2534 8186
rect 2714 8134 2716 8186
rect 2470 8132 2476 8134
rect 2532 8132 2556 8134
rect 2612 8132 2636 8134
rect 2692 8132 2716 8134
rect 2772 8132 2778 8134
rect 2470 8123 2778 8132
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1150 7100 1458 7109
rect 1150 7098 1156 7100
rect 1212 7098 1236 7100
rect 1292 7098 1316 7100
rect 1372 7098 1396 7100
rect 1452 7098 1458 7100
rect 1212 7046 1214 7098
rect 1394 7046 1396 7098
rect 1150 7044 1156 7046
rect 1212 7044 1236 7046
rect 1292 7044 1316 7046
rect 1372 7044 1396 7046
rect 1452 7044 1458 7046
rect 1150 7035 1458 7044
rect 1596 6914 1624 7346
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1688 7002 1716 7210
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1504 6886 1624 6914
rect 1504 6730 1532 6886
rect 1492 6724 1544 6730
rect 1492 6666 1544 6672
rect 1150 6012 1458 6021
rect 1150 6010 1156 6012
rect 1212 6010 1236 6012
rect 1292 6010 1316 6012
rect 1372 6010 1396 6012
rect 1452 6010 1458 6012
rect 1212 5958 1214 6010
rect 1394 5958 1396 6010
rect 1150 5956 1156 5958
rect 1212 5956 1236 5958
rect 1292 5956 1316 5958
rect 1372 5956 1396 5958
rect 1452 5956 1458 5958
rect 1150 5947 1458 5956
rect 1150 4924 1458 4933
rect 1150 4922 1156 4924
rect 1212 4922 1236 4924
rect 1292 4922 1316 4924
rect 1372 4922 1396 4924
rect 1452 4922 1458 4924
rect 1212 4870 1214 4922
rect 1394 4870 1396 4922
rect 1150 4868 1156 4870
rect 1212 4868 1236 4870
rect 1292 4868 1316 4870
rect 1372 4868 1396 4870
rect 1452 4868 1458 4870
rect 1150 4859 1458 4868
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1412 4146 1440 4422
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1150 3836 1458 3845
rect 1150 3834 1156 3836
rect 1212 3834 1236 3836
rect 1292 3834 1316 3836
rect 1372 3834 1396 3836
rect 1452 3834 1458 3836
rect 1212 3782 1214 3834
rect 1394 3782 1396 3834
rect 1150 3780 1156 3782
rect 1212 3780 1236 3782
rect 1292 3780 1316 3782
rect 1372 3780 1396 3782
rect 1452 3780 1458 3782
rect 1150 3771 1458 3780
rect 1150 2748 1458 2757
rect 1150 2746 1156 2748
rect 1212 2746 1236 2748
rect 1292 2746 1316 2748
rect 1372 2746 1396 2748
rect 1452 2746 1458 2748
rect 1212 2694 1214 2746
rect 1394 2694 1396 2746
rect 1150 2692 1156 2694
rect 1212 2692 1236 2694
rect 1292 2692 1316 2694
rect 1372 2692 1396 2694
rect 1452 2692 1458 2694
rect 1150 2683 1458 2692
rect 1504 2446 1532 6666
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1596 3126 1624 4082
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1688 2446 1716 6938
rect 2148 6662 2176 7414
rect 2240 7206 2268 7822
rect 2884 7818 2912 8298
rect 3790 8188 4098 8197
rect 3790 8186 3796 8188
rect 3852 8186 3876 8188
rect 3932 8186 3956 8188
rect 4012 8186 4036 8188
rect 4092 8186 4098 8188
rect 3852 8134 3854 8186
rect 4034 8134 4036 8186
rect 3790 8132 3796 8134
rect 3852 8132 3876 8134
rect 3932 8132 3956 8134
rect 4012 8132 4036 8134
rect 4092 8132 4098 8134
rect 3790 8123 4098 8132
rect 5110 8188 5418 8197
rect 5110 8186 5116 8188
rect 5172 8186 5196 8188
rect 5252 8186 5276 8188
rect 5332 8186 5356 8188
rect 5412 8186 5418 8188
rect 5172 8134 5174 8186
rect 5354 8134 5356 8186
rect 5110 8132 5116 8134
rect 5172 8132 5196 8134
rect 5252 8132 5276 8134
rect 5332 8132 5356 8134
rect 5412 8132 5418 8134
rect 5110 8123 5418 8132
rect 6430 8188 6738 8197
rect 6430 8186 6436 8188
rect 6492 8186 6516 8188
rect 6572 8186 6596 8188
rect 6652 8186 6676 8188
rect 6732 8186 6738 8188
rect 6492 8134 6494 8186
rect 6674 8134 6676 8186
rect 6430 8132 6436 8134
rect 6492 8132 6516 8134
rect 6572 8132 6596 8134
rect 6652 8132 6676 8134
rect 6732 8132 6738 8134
rect 6430 8123 6738 8132
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 3130 7644 3438 7653
rect 3130 7642 3136 7644
rect 3192 7642 3216 7644
rect 3272 7642 3296 7644
rect 3352 7642 3376 7644
rect 3432 7642 3438 7644
rect 3192 7590 3194 7642
rect 3374 7590 3376 7642
rect 3130 7588 3136 7590
rect 3192 7588 3216 7590
rect 3272 7588 3296 7590
rect 3352 7588 3376 7590
rect 3432 7588 3438 7590
rect 3130 7579 3438 7588
rect 4450 7644 4758 7653
rect 4450 7642 4456 7644
rect 4512 7642 4536 7644
rect 4592 7642 4616 7644
rect 4672 7642 4696 7644
rect 4752 7642 4758 7644
rect 4512 7590 4514 7642
rect 4694 7590 4696 7642
rect 4450 7588 4456 7590
rect 4512 7588 4536 7590
rect 4592 7588 4616 7590
rect 4672 7588 4696 7590
rect 4752 7588 4758 7590
rect 4450 7579 4758 7588
rect 5770 7644 6078 7653
rect 5770 7642 5776 7644
rect 5832 7642 5856 7644
rect 5912 7642 5936 7644
rect 5992 7642 6016 7644
rect 6072 7642 6078 7644
rect 5832 7590 5834 7642
rect 6014 7590 6016 7642
rect 5770 7588 5776 7590
rect 5832 7588 5856 7590
rect 5912 7588 5936 7590
rect 5992 7588 6016 7590
rect 6072 7588 6078 7590
rect 5770 7579 6078 7588
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1810 6556 2118 6565
rect 1810 6554 1816 6556
rect 1872 6554 1896 6556
rect 1952 6554 1976 6556
rect 2032 6554 2056 6556
rect 2112 6554 2118 6556
rect 1872 6502 1874 6554
rect 2054 6502 2056 6554
rect 1810 6500 1816 6502
rect 1872 6500 1896 6502
rect 1952 6500 1976 6502
rect 2032 6500 2056 6502
rect 2112 6500 2118 6502
rect 1810 6491 2118 6500
rect 2240 5914 2268 7142
rect 2470 7100 2778 7109
rect 2470 7098 2476 7100
rect 2532 7098 2556 7100
rect 2612 7098 2636 7100
rect 2692 7098 2716 7100
rect 2772 7098 2778 7100
rect 2532 7046 2534 7098
rect 2714 7046 2716 7098
rect 2470 7044 2476 7046
rect 2532 7044 2556 7046
rect 2612 7044 2636 7046
rect 2692 7044 2716 7046
rect 2772 7044 2778 7046
rect 2470 7035 2778 7044
rect 2976 7002 3004 7346
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2470 6012 2778 6021
rect 2470 6010 2476 6012
rect 2532 6010 2556 6012
rect 2612 6010 2636 6012
rect 2692 6010 2716 6012
rect 2772 6010 2778 6012
rect 2532 5958 2534 6010
rect 2714 5958 2716 6010
rect 2470 5956 2476 5958
rect 2532 5956 2556 5958
rect 2612 5956 2636 5958
rect 2692 5956 2716 5958
rect 2772 5956 2778 5958
rect 2470 5947 2778 5956
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 1810 5468 2118 5477
rect 1810 5466 1816 5468
rect 1872 5466 1896 5468
rect 1952 5466 1976 5468
rect 2032 5466 2056 5468
rect 2112 5466 2118 5468
rect 1872 5414 1874 5466
rect 2054 5414 2056 5466
rect 1810 5412 1816 5414
rect 1872 5412 1896 5414
rect 1952 5412 1976 5414
rect 2032 5412 2056 5414
rect 2112 5412 2118 5414
rect 1810 5403 2118 5412
rect 2240 4690 2268 5850
rect 2470 4924 2778 4933
rect 2470 4922 2476 4924
rect 2532 4922 2556 4924
rect 2612 4922 2636 4924
rect 2692 4922 2716 4924
rect 2772 4922 2778 4924
rect 2532 4870 2534 4922
rect 2714 4870 2716 4922
rect 2470 4868 2476 4870
rect 2532 4868 2556 4870
rect 2612 4868 2636 4870
rect 2692 4868 2716 4870
rect 2772 4868 2778 4870
rect 2470 4859 2778 4868
rect 2884 4826 2912 6802
rect 3068 6798 3096 7482
rect 3790 7100 4098 7109
rect 3790 7098 3796 7100
rect 3852 7098 3876 7100
rect 3932 7098 3956 7100
rect 4012 7098 4036 7100
rect 4092 7098 4098 7100
rect 3852 7046 3854 7098
rect 4034 7046 4036 7098
rect 3790 7044 3796 7046
rect 3852 7044 3876 7046
rect 3932 7044 3956 7046
rect 4012 7044 4036 7046
rect 4092 7044 4098 7046
rect 3790 7035 4098 7044
rect 5110 7100 5418 7109
rect 5110 7098 5116 7100
rect 5172 7098 5196 7100
rect 5252 7098 5276 7100
rect 5332 7098 5356 7100
rect 5412 7098 5418 7100
rect 5172 7046 5174 7098
rect 5354 7046 5356 7098
rect 5110 7044 5116 7046
rect 5172 7044 5196 7046
rect 5252 7044 5276 7046
rect 5332 7044 5356 7046
rect 5412 7044 5418 7046
rect 5110 7035 5418 7044
rect 6430 7100 6738 7109
rect 6430 7098 6436 7100
rect 6492 7098 6516 7100
rect 6572 7098 6596 7100
rect 6652 7098 6676 7100
rect 6732 7098 6738 7100
rect 6492 7046 6494 7098
rect 6674 7046 6676 7098
rect 6430 7044 6436 7046
rect 6492 7044 6516 7046
rect 6572 7044 6596 7046
rect 6652 7044 6676 7046
rect 6732 7044 6738 7046
rect 6430 7035 6738 7044
rect 6932 6882 6960 9976
rect 7090 9820 7398 9829
rect 7090 9818 7096 9820
rect 7152 9818 7176 9820
rect 7232 9818 7256 9820
rect 7312 9818 7336 9820
rect 7392 9818 7398 9820
rect 7152 9766 7154 9818
rect 7334 9766 7336 9818
rect 7090 9764 7096 9766
rect 7152 9764 7176 9766
rect 7232 9764 7256 9766
rect 7312 9764 7336 9766
rect 7392 9764 7398 9766
rect 7090 9755 7398 9764
rect 8410 9820 8718 9829
rect 8410 9818 8416 9820
rect 8472 9818 8496 9820
rect 8552 9818 8576 9820
rect 8632 9818 8656 9820
rect 8712 9818 8718 9820
rect 8472 9766 8474 9818
rect 8654 9766 8656 9818
rect 8410 9764 8416 9766
rect 8472 9764 8496 9766
rect 8552 9764 8576 9766
rect 8632 9764 8656 9766
rect 8712 9764 8718 9766
rect 8410 9755 8718 9764
rect 7750 9276 8058 9285
rect 7750 9274 7756 9276
rect 7812 9274 7836 9276
rect 7892 9274 7916 9276
rect 7972 9274 7996 9276
rect 8052 9274 8058 9276
rect 7812 9222 7814 9274
rect 7994 9222 7996 9274
rect 7750 9220 7756 9222
rect 7812 9220 7836 9222
rect 7892 9220 7916 9222
rect 7972 9220 7996 9222
rect 8052 9220 8058 9222
rect 7750 9211 8058 9220
rect 7090 8732 7398 8741
rect 7090 8730 7096 8732
rect 7152 8730 7176 8732
rect 7232 8730 7256 8732
rect 7312 8730 7336 8732
rect 7392 8730 7398 8732
rect 7152 8678 7154 8730
rect 7334 8678 7336 8730
rect 7090 8676 7096 8678
rect 7152 8676 7176 8678
rect 7232 8676 7256 8678
rect 7312 8676 7336 8678
rect 7392 8676 7398 8678
rect 7090 8667 7398 8676
rect 8410 8732 8718 8741
rect 8410 8730 8416 8732
rect 8472 8730 8496 8732
rect 8552 8730 8576 8732
rect 8632 8730 8656 8732
rect 8712 8730 8718 8732
rect 8472 8678 8474 8730
rect 8654 8678 8656 8730
rect 8410 8676 8416 8678
rect 8472 8676 8496 8678
rect 8552 8676 8576 8678
rect 8632 8676 8656 8678
rect 8712 8676 8718 8678
rect 8410 8667 8718 8676
rect 7750 8188 8058 8197
rect 7750 8186 7756 8188
rect 7812 8186 7836 8188
rect 7892 8186 7916 8188
rect 7972 8186 7996 8188
rect 8052 8186 8058 8188
rect 7812 8134 7814 8186
rect 7994 8134 7996 8186
rect 7750 8132 7756 8134
rect 7812 8132 7836 8134
rect 7892 8132 7916 8134
rect 7972 8132 7996 8134
rect 8052 8132 8058 8134
rect 7750 8123 8058 8132
rect 7090 7644 7398 7653
rect 7090 7642 7096 7644
rect 7152 7642 7176 7644
rect 7232 7642 7256 7644
rect 7312 7642 7336 7644
rect 7392 7642 7398 7644
rect 7152 7590 7154 7642
rect 7334 7590 7336 7642
rect 7090 7588 7096 7590
rect 7152 7588 7176 7590
rect 7232 7588 7256 7590
rect 7312 7588 7336 7590
rect 7392 7588 7398 7590
rect 7090 7579 7398 7588
rect 8410 7644 8718 7653
rect 8410 7642 8416 7644
rect 8472 7642 8496 7644
rect 8552 7642 8576 7644
rect 8632 7642 8656 7644
rect 8712 7642 8718 7644
rect 8472 7590 8474 7642
rect 8654 7590 8656 7642
rect 8410 7588 8416 7590
rect 8472 7588 8496 7590
rect 8552 7588 8576 7590
rect 8632 7588 8656 7590
rect 8712 7588 8718 7590
rect 8410 7579 8718 7588
rect 7750 7100 8058 7109
rect 7750 7098 7756 7100
rect 7812 7098 7836 7100
rect 7892 7098 7916 7100
rect 7972 7098 7996 7100
rect 8052 7098 8058 7100
rect 7812 7046 7814 7098
rect 7994 7046 7996 7098
rect 7750 7044 7756 7046
rect 7812 7044 7836 7046
rect 7892 7044 7916 7046
rect 7972 7044 7996 7046
rect 8052 7044 8058 7046
rect 7750 7035 8058 7044
rect 6840 6854 6960 6882
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3130 6556 3438 6565
rect 3130 6554 3136 6556
rect 3192 6554 3216 6556
rect 3272 6554 3296 6556
rect 3352 6554 3376 6556
rect 3432 6554 3438 6556
rect 3192 6502 3194 6554
rect 3374 6502 3376 6554
rect 3130 6500 3136 6502
rect 3192 6500 3216 6502
rect 3272 6500 3296 6502
rect 3352 6500 3376 6502
rect 3432 6500 3438 6502
rect 3130 6491 3438 6500
rect 4450 6556 4758 6565
rect 4450 6554 4456 6556
rect 4512 6554 4536 6556
rect 4592 6554 4616 6556
rect 4672 6554 4696 6556
rect 4752 6554 4758 6556
rect 4512 6502 4514 6554
rect 4694 6502 4696 6554
rect 4450 6500 4456 6502
rect 4512 6500 4536 6502
rect 4592 6500 4616 6502
rect 4672 6500 4696 6502
rect 4752 6500 4758 6502
rect 4450 6491 4758 6500
rect 5770 6556 6078 6565
rect 5770 6554 5776 6556
rect 5832 6554 5856 6556
rect 5912 6554 5936 6556
rect 5992 6554 6016 6556
rect 6072 6554 6078 6556
rect 5832 6502 5834 6554
rect 6014 6502 6016 6554
rect 5770 6500 5776 6502
rect 5832 6500 5856 6502
rect 5912 6500 5936 6502
rect 5992 6500 6016 6502
rect 6072 6500 6078 6502
rect 5770 6491 6078 6500
rect 3790 6012 4098 6021
rect 3790 6010 3796 6012
rect 3852 6010 3876 6012
rect 3932 6010 3956 6012
rect 4012 6010 4036 6012
rect 4092 6010 4098 6012
rect 3852 5958 3854 6010
rect 4034 5958 4036 6010
rect 3790 5956 3796 5958
rect 3852 5956 3876 5958
rect 3932 5956 3956 5958
rect 4012 5956 4036 5958
rect 4092 5956 4098 5958
rect 3790 5947 4098 5956
rect 5110 6012 5418 6021
rect 5110 6010 5116 6012
rect 5172 6010 5196 6012
rect 5252 6010 5276 6012
rect 5332 6010 5356 6012
rect 5412 6010 5418 6012
rect 5172 5958 5174 6010
rect 5354 5958 5356 6010
rect 5110 5956 5116 5958
rect 5172 5956 5196 5958
rect 5252 5956 5276 5958
rect 5332 5956 5356 5958
rect 5412 5956 5418 5958
rect 5110 5947 5418 5956
rect 6430 6012 6738 6021
rect 6430 6010 6436 6012
rect 6492 6010 6516 6012
rect 6572 6010 6596 6012
rect 6652 6010 6676 6012
rect 6732 6010 6738 6012
rect 6492 5958 6494 6010
rect 6674 5958 6676 6010
rect 6430 5956 6436 5958
rect 6492 5956 6516 5958
rect 6572 5956 6596 5958
rect 6652 5956 6676 5958
rect 6732 5956 6738 5958
rect 6430 5947 6738 5956
rect 6840 5710 6868 6854
rect 7090 6556 7398 6565
rect 7090 6554 7096 6556
rect 7152 6554 7176 6556
rect 7232 6554 7256 6556
rect 7312 6554 7336 6556
rect 7392 6554 7398 6556
rect 7152 6502 7154 6554
rect 7334 6502 7336 6554
rect 7090 6500 7096 6502
rect 7152 6500 7176 6502
rect 7232 6500 7256 6502
rect 7312 6500 7336 6502
rect 7392 6500 7398 6502
rect 7090 6491 7398 6500
rect 8410 6556 8718 6565
rect 8410 6554 8416 6556
rect 8472 6554 8496 6556
rect 8552 6554 8576 6556
rect 8632 6554 8656 6556
rect 8712 6554 8718 6556
rect 8472 6502 8474 6554
rect 8654 6502 8656 6554
rect 8410 6500 8416 6502
rect 8472 6500 8496 6502
rect 8552 6500 8576 6502
rect 8632 6500 8656 6502
rect 8712 6500 8718 6502
rect 8410 6491 8718 6500
rect 7750 6012 8058 6021
rect 7750 6010 7756 6012
rect 7812 6010 7836 6012
rect 7892 6010 7916 6012
rect 7972 6010 7996 6012
rect 8052 6010 8058 6012
rect 7812 5958 7814 6010
rect 7994 5958 7996 6010
rect 7750 5956 7756 5958
rect 7812 5956 7836 5958
rect 7892 5956 7916 5958
rect 7972 5956 7996 5958
rect 8052 5956 8058 5958
rect 7750 5947 8058 5956
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 5448 5568 5500 5574
rect 5500 5516 5580 5522
rect 5448 5510 5580 5516
rect 5460 5494 5580 5510
rect 3130 5468 3438 5477
rect 3130 5466 3136 5468
rect 3192 5466 3216 5468
rect 3272 5466 3296 5468
rect 3352 5466 3376 5468
rect 3432 5466 3438 5468
rect 3192 5414 3194 5466
rect 3374 5414 3376 5466
rect 3130 5412 3136 5414
rect 3192 5412 3216 5414
rect 3272 5412 3296 5414
rect 3352 5412 3376 5414
rect 3432 5412 3438 5414
rect 3130 5403 3438 5412
rect 4450 5468 4758 5477
rect 4450 5466 4456 5468
rect 4512 5466 4536 5468
rect 4592 5466 4616 5468
rect 4672 5466 4696 5468
rect 4752 5466 4758 5468
rect 4512 5414 4514 5466
rect 4694 5414 4696 5466
rect 4450 5412 4456 5414
rect 4512 5412 4536 5414
rect 4592 5412 4616 5414
rect 4672 5412 4696 5414
rect 4752 5412 4758 5414
rect 4450 5403 4758 5412
rect 5552 5386 5580 5494
rect 5770 5468 6078 5477
rect 5770 5466 5776 5468
rect 5832 5466 5856 5468
rect 5912 5466 5936 5468
rect 5992 5466 6016 5468
rect 6072 5466 6078 5468
rect 5832 5414 5834 5466
rect 6014 5414 6016 5466
rect 5770 5412 5776 5414
rect 5832 5412 5856 5414
rect 5912 5412 5936 5414
rect 5992 5412 6016 5414
rect 6072 5412 6078 5414
rect 5770 5403 6078 5412
rect 7090 5468 7398 5477
rect 7090 5466 7096 5468
rect 7152 5466 7176 5468
rect 7232 5466 7256 5468
rect 7312 5466 7336 5468
rect 7392 5466 7398 5468
rect 7152 5414 7154 5466
rect 7334 5414 7336 5466
rect 7090 5412 7096 5414
rect 7152 5412 7176 5414
rect 7232 5412 7256 5414
rect 7312 5412 7336 5414
rect 7392 5412 7398 5414
rect 7090 5403 7398 5412
rect 8410 5468 8718 5477
rect 8410 5466 8416 5468
rect 8472 5466 8496 5468
rect 8552 5466 8576 5468
rect 8632 5466 8656 5468
rect 8712 5466 8718 5468
rect 8472 5414 8474 5466
rect 8654 5414 8656 5466
rect 8410 5412 8416 5414
rect 8472 5412 8496 5414
rect 8552 5412 8576 5414
rect 8632 5412 8656 5414
rect 8712 5412 8718 5414
rect 8410 5403 8718 5412
rect 5552 5358 5672 5386
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3790 4924 4098 4933
rect 3790 4922 3796 4924
rect 3852 4922 3876 4924
rect 3932 4922 3956 4924
rect 4012 4922 4036 4924
rect 4092 4922 4098 4924
rect 3852 4870 3854 4922
rect 4034 4870 4036 4922
rect 3790 4868 3796 4870
rect 3852 4868 3876 4870
rect 3932 4868 3956 4870
rect 4012 4868 4036 4870
rect 4092 4868 4098 4870
rect 3790 4859 4098 4868
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 1810 4380 2118 4389
rect 1810 4378 1816 4380
rect 1872 4378 1896 4380
rect 1952 4378 1976 4380
rect 2032 4378 2056 4380
rect 2112 4378 2118 4380
rect 1872 4326 1874 4378
rect 2054 4326 2056 4378
rect 1810 4324 1816 4326
rect 1872 4324 1896 4326
rect 1952 4324 1976 4326
rect 2032 4324 2056 4326
rect 2112 4324 2118 4326
rect 1810 4315 2118 4324
rect 2240 4214 2268 4626
rect 2884 4486 2912 4762
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2044 4208 2096 4214
rect 2044 4150 2096 4156
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 2056 3534 2084 4150
rect 2470 3836 2778 3845
rect 2470 3834 2476 3836
rect 2532 3834 2556 3836
rect 2612 3834 2636 3836
rect 2692 3834 2716 3836
rect 2772 3834 2778 3836
rect 2532 3782 2534 3834
rect 2714 3782 2716 3834
rect 2470 3780 2476 3782
rect 2532 3780 2556 3782
rect 2612 3780 2636 3782
rect 2692 3780 2716 3782
rect 2772 3780 2778 3782
rect 2470 3771 2778 3780
rect 2884 3738 2912 4422
rect 2976 4282 3004 4558
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 1810 3292 2118 3301
rect 1810 3290 1816 3292
rect 1872 3290 1896 3292
rect 1952 3290 1976 3292
rect 2032 3290 2056 3292
rect 2112 3290 2118 3292
rect 1872 3238 1874 3290
rect 2054 3238 2056 3290
rect 1810 3236 1816 3238
rect 1872 3236 1896 3238
rect 1952 3236 1976 3238
rect 2032 3236 2056 3238
rect 2112 3236 2118 3238
rect 1810 3227 2118 3236
rect 2424 3194 2452 3402
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2976 2922 3004 4218
rect 3068 4078 3096 4490
rect 3130 4380 3438 4389
rect 3130 4378 3136 4380
rect 3192 4378 3216 4380
rect 3272 4378 3296 4380
rect 3352 4378 3376 4380
rect 3432 4378 3438 4380
rect 3192 4326 3194 4378
rect 3374 4326 3376 4378
rect 3130 4324 3136 4326
rect 3192 4324 3216 4326
rect 3272 4324 3296 4326
rect 3352 4324 3376 4326
rect 3432 4324 3438 4326
rect 3130 4315 3438 4324
rect 3528 4146 3556 4694
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 4172 4078 4200 5034
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4622 4476 4966
rect 5110 4924 5418 4933
rect 5110 4922 5116 4924
rect 5172 4922 5196 4924
rect 5252 4922 5276 4924
rect 5332 4922 5356 4924
rect 5412 4922 5418 4924
rect 5172 4870 5174 4922
rect 5354 4870 5356 4922
rect 5110 4868 5116 4870
rect 5172 4868 5196 4870
rect 5252 4868 5276 4870
rect 5332 4868 5356 4870
rect 5412 4868 5418 4870
rect 5110 4859 5418 4868
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4908 4570 4936 4626
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4264 4010 4292 4422
rect 4450 4380 4758 4389
rect 4450 4378 4456 4380
rect 4512 4378 4536 4380
rect 4592 4378 4616 4380
rect 4672 4378 4696 4380
rect 4752 4378 4758 4380
rect 4512 4326 4514 4378
rect 4694 4326 4696 4378
rect 4450 4324 4456 4326
rect 4512 4324 4536 4326
rect 4592 4324 4616 4326
rect 4672 4324 4696 4326
rect 4752 4324 4758 4326
rect 4450 4315 4758 4324
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 3790 3836 4098 3845
rect 3790 3834 3796 3836
rect 3852 3834 3876 3836
rect 3932 3834 3956 3836
rect 4012 3834 4036 3836
rect 4092 3834 4098 3836
rect 3852 3782 3854 3834
rect 4034 3782 4036 3834
rect 3790 3780 3796 3782
rect 3852 3780 3876 3782
rect 3932 3780 3956 3782
rect 4012 3780 4036 3782
rect 4092 3780 4098 3782
rect 3790 3771 4098 3780
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3068 3058 3096 3334
rect 3130 3292 3438 3301
rect 3130 3290 3136 3292
rect 3192 3290 3216 3292
rect 3272 3290 3296 3292
rect 3352 3290 3376 3292
rect 3432 3290 3438 3292
rect 3192 3238 3194 3290
rect 3374 3238 3376 3290
rect 3130 3236 3136 3238
rect 3192 3236 3216 3238
rect 3272 3236 3296 3238
rect 3352 3236 3376 3238
rect 3432 3236 3438 3238
rect 3130 3227 3438 3236
rect 3620 3058 3648 3674
rect 4264 3670 4292 3946
rect 4448 3738 4476 4218
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4528 4072 4580 4078
rect 4526 4040 4528 4049
rect 4580 4040 4582 4049
rect 4526 3975 4582 3984
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 3194 4200 3470
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2470 2748 2778 2757
rect 2470 2746 2476 2748
rect 2532 2746 2556 2748
rect 2612 2746 2636 2748
rect 2692 2746 2716 2748
rect 2772 2746 2778 2748
rect 2532 2694 2534 2746
rect 2714 2694 2716 2746
rect 2470 2692 2476 2694
rect 2532 2692 2556 2694
rect 2612 2692 2636 2694
rect 2692 2692 2716 2694
rect 2772 2692 2778 2694
rect 2470 2683 2778 2692
rect 2976 2446 3004 2858
rect 3712 2446 3740 3062
rect 4264 2854 4292 3606
rect 4632 3398 4660 3946
rect 4724 3618 4752 4082
rect 4816 3738 4844 4558
rect 4908 4542 5028 4570
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4214 4936 4422
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4908 3618 4936 3674
rect 4724 3590 4936 3618
rect 5000 3466 5028 4542
rect 5460 4049 5488 4694
rect 5644 4622 5672 5358
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5736 4486 5764 5102
rect 5828 5098 5856 5238
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6012 4758 6040 5034
rect 6104 4826 6132 5170
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5446 4040 5502 4049
rect 5446 3975 5502 3984
rect 5110 3836 5418 3845
rect 5110 3834 5116 3836
rect 5172 3834 5196 3836
rect 5252 3834 5276 3836
rect 5332 3834 5356 3836
rect 5412 3834 5418 3836
rect 5172 3782 5174 3834
rect 5354 3782 5356 3834
rect 5110 3780 5116 3782
rect 5172 3780 5196 3782
rect 5252 3780 5276 3782
rect 5332 3780 5356 3782
rect 5412 3780 5418 3782
rect 5110 3771 5418 3780
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 5264 3460 5316 3466
rect 5460 3448 5488 3975
rect 5316 3420 5488 3448
rect 5264 3402 5316 3408
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4450 3292 4758 3301
rect 4450 3290 4456 3292
rect 4512 3290 4536 3292
rect 4592 3290 4616 3292
rect 4672 3290 4696 3292
rect 4752 3290 4758 3292
rect 4512 3238 4514 3290
rect 4694 3238 4696 3290
rect 4450 3236 4456 3238
rect 4512 3236 4536 3238
rect 4592 3236 4616 3238
rect 4672 3236 4696 3238
rect 4752 3236 4758 3238
rect 4450 3227 4758 3236
rect 5000 3058 5028 3402
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5460 2854 5488 3420
rect 5552 3194 5580 4422
rect 5644 3466 5672 4422
rect 5770 4380 6078 4389
rect 5770 4378 5776 4380
rect 5832 4378 5856 4380
rect 5912 4378 5936 4380
rect 5992 4378 6016 4380
rect 6072 4378 6078 4380
rect 5832 4326 5834 4378
rect 6014 4326 6016 4378
rect 5770 4324 5776 4326
rect 5832 4324 5856 4326
rect 5912 4324 5936 4326
rect 5992 4324 6016 4326
rect 6072 4324 6078 4326
rect 5770 4315 6078 4324
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3534 5764 3878
rect 6104 3738 6132 4082
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 6196 3398 6224 4626
rect 6288 4146 6316 5306
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6430 4924 6738 4933
rect 6430 4922 6436 4924
rect 6492 4922 6516 4924
rect 6572 4922 6596 4924
rect 6652 4922 6676 4924
rect 6732 4922 6738 4924
rect 6492 4870 6494 4922
rect 6674 4870 6676 4922
rect 6430 4868 6436 4870
rect 6492 4868 6516 4870
rect 6572 4868 6596 4870
rect 6652 4868 6676 4870
rect 6732 4868 6738 4870
rect 6430 4859 6738 4868
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6656 4146 6684 4422
rect 6840 4282 6868 5170
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6840 4162 6868 4218
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6644 4140 6696 4146
rect 6840 4134 6960 4162
rect 6644 4082 6696 4088
rect 6656 4026 6684 4082
rect 6656 3998 6868 4026
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 5770 3292 6078 3301
rect 5770 3290 5776 3292
rect 5832 3290 5856 3292
rect 5912 3290 5936 3292
rect 5992 3290 6016 3292
rect 6072 3290 6078 3292
rect 5832 3238 5834 3290
rect 6014 3238 6016 3290
rect 5770 3236 5776 3238
rect 5832 3236 5856 3238
rect 5912 3236 5936 3238
rect 5992 3236 6016 3238
rect 6072 3236 6078 3238
rect 5770 3227 6078 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6196 3126 6224 3334
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 3790 2748 4098 2757
rect 3790 2746 3796 2748
rect 3852 2746 3876 2748
rect 3932 2746 3956 2748
rect 4012 2746 4036 2748
rect 4092 2746 4098 2748
rect 3852 2694 3854 2746
rect 4034 2694 4036 2746
rect 3790 2692 3796 2694
rect 3852 2692 3876 2694
rect 3932 2692 3956 2694
rect 4012 2692 4036 2694
rect 4092 2692 4098 2694
rect 3790 2683 4098 2692
rect 5110 2748 5418 2757
rect 5110 2746 5116 2748
rect 5172 2746 5196 2748
rect 5252 2746 5276 2748
rect 5332 2746 5356 2748
rect 5412 2746 5418 2748
rect 5172 2694 5174 2746
rect 5354 2694 5356 2746
rect 5110 2692 5116 2694
rect 5172 2692 5196 2694
rect 5252 2692 5276 2694
rect 5332 2692 5356 2694
rect 5412 2692 5418 2694
rect 5110 2683 5418 2692
rect 5460 2446 5488 2790
rect 5644 2446 5672 2858
rect 5828 2446 5856 2994
rect 5920 2922 5948 2994
rect 6288 2990 6316 3878
rect 6430 3836 6738 3845
rect 6430 3834 6436 3836
rect 6492 3834 6516 3836
rect 6572 3834 6596 3836
rect 6652 3834 6676 3836
rect 6732 3834 6738 3836
rect 6492 3782 6494 3834
rect 6674 3782 6676 3834
rect 6430 3780 6436 3782
rect 6492 3780 6516 3782
rect 6572 3780 6596 3782
rect 6652 3780 6676 3782
rect 6732 3780 6738 3782
rect 6430 3771 6738 3780
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6380 2938 6408 3402
rect 6472 3058 6500 3674
rect 6840 3618 6868 3998
rect 6748 3590 6868 3618
rect 6748 3534 6776 3590
rect 6736 3528 6788 3534
rect 6932 3482 6960 4134
rect 6736 3470 6788 3476
rect 6840 3454 6960 3482
rect 6840 3194 6868 3454
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6656 2938 6684 2994
rect 5908 2916 5960 2922
rect 6380 2910 6684 2938
rect 5908 2858 5960 2864
rect 7024 2854 7052 5102
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7090 4380 7398 4389
rect 7090 4378 7096 4380
rect 7152 4378 7176 4380
rect 7232 4378 7256 4380
rect 7312 4378 7336 4380
rect 7392 4378 7398 4380
rect 7152 4326 7154 4378
rect 7334 4326 7336 4378
rect 7090 4324 7096 4326
rect 7152 4324 7176 4326
rect 7232 4324 7256 4326
rect 7312 4324 7336 4326
rect 7392 4324 7398 4326
rect 7090 4315 7398 4324
rect 7090 3292 7398 3301
rect 7090 3290 7096 3292
rect 7152 3290 7176 3292
rect 7232 3290 7256 3292
rect 7312 3290 7336 3292
rect 7392 3290 7398 3292
rect 7152 3238 7154 3290
rect 7334 3238 7336 3290
rect 7090 3236 7096 3238
rect 7152 3236 7176 3238
rect 7232 3236 7256 3238
rect 7312 3236 7336 3238
rect 7392 3236 7398 3238
rect 7090 3227 7398 3236
rect 7484 3194 7512 4966
rect 7576 4214 7604 4966
rect 7750 4924 8058 4933
rect 7750 4922 7756 4924
rect 7812 4922 7836 4924
rect 7892 4922 7916 4924
rect 7972 4922 7996 4924
rect 8052 4922 8058 4924
rect 7812 4870 7814 4922
rect 7994 4870 7996 4922
rect 7750 4868 7756 4870
rect 7812 4868 7836 4870
rect 7892 4868 7916 4870
rect 7972 4868 7996 4870
rect 8052 4868 8058 4870
rect 7750 4859 8058 4868
rect 8410 4380 8718 4389
rect 8410 4378 8416 4380
rect 8472 4378 8496 4380
rect 8552 4378 8576 4380
rect 8632 4378 8656 4380
rect 8712 4378 8718 4380
rect 8472 4326 8474 4378
rect 8654 4326 8656 4378
rect 8410 4324 8416 4326
rect 8472 4324 8496 4326
rect 8552 4324 8576 4326
rect 8632 4324 8656 4326
rect 8712 4324 8718 4326
rect 8410 4315 8718 4324
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 7750 3836 8058 3845
rect 7750 3834 7756 3836
rect 7812 3834 7836 3836
rect 7892 3834 7916 3836
rect 7972 3834 7996 3836
rect 8052 3834 8058 3836
rect 7812 3782 7814 3834
rect 7994 3782 7996 3834
rect 7750 3780 7756 3782
rect 7812 3780 7836 3782
rect 7892 3780 7916 3782
rect 7972 3780 7996 3782
rect 8052 3780 8058 3782
rect 7750 3771 8058 3780
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7300 2990 7328 3130
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6430 2748 6738 2757
rect 6430 2746 6436 2748
rect 6492 2746 6516 2748
rect 6572 2746 6596 2748
rect 6652 2746 6676 2748
rect 6732 2746 6738 2748
rect 6492 2694 6494 2746
rect 6674 2694 6676 2746
rect 6430 2692 6436 2694
rect 6492 2692 6516 2694
rect 6572 2692 6596 2694
rect 6652 2692 6676 2694
rect 6732 2692 6738 2694
rect 6430 2683 6738 2692
rect 7576 2446 7604 3334
rect 7668 2990 7696 3402
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8036 3058 8064 3334
rect 8312 3126 8340 3878
rect 8410 3292 8718 3301
rect 8410 3290 8416 3292
rect 8472 3290 8496 3292
rect 8552 3290 8576 3292
rect 8632 3290 8656 3292
rect 8712 3290 8718 3292
rect 8472 3238 8474 3290
rect 8654 3238 8656 3290
rect 8410 3236 8416 3238
rect 8472 3236 8496 3238
rect 8552 3236 8576 3238
rect 8632 3236 8656 3238
rect 8712 3236 8718 3238
rect 8410 3227 8718 3236
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 8036 2938 8064 2994
rect 8036 2910 8156 2938
rect 7750 2748 8058 2757
rect 7750 2746 7756 2748
rect 7812 2746 7836 2748
rect 7892 2746 7916 2748
rect 7972 2746 7996 2748
rect 8052 2746 8058 2748
rect 7812 2694 7814 2746
rect 7994 2694 7996 2746
rect 7750 2692 7756 2694
rect 7812 2692 7836 2694
rect 7892 2692 7916 2694
rect 7972 2692 7996 2694
rect 8052 2692 8058 2694
rect 7750 2683 8058 2692
rect 8128 2446 8156 2910
rect 8312 2446 8340 3062
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 756 2304 808 2310
rect 756 2246 808 2252
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 7012 2304 7064 2310
rect 8208 2304 8260 2310
rect 7012 2246 7064 2252
rect 8128 2264 8208 2292
rect 768 1782 796 2246
rect 1688 1782 1716 2246
rect 1810 2204 2118 2213
rect 1810 2202 1816 2204
rect 1872 2202 1896 2204
rect 1952 2202 1976 2204
rect 2032 2202 2056 2204
rect 2112 2202 2118 2204
rect 1872 2150 1874 2202
rect 2054 2150 2056 2202
rect 1810 2148 1816 2150
rect 1872 2148 1896 2150
rect 1952 2148 1976 2150
rect 2032 2148 2056 2150
rect 2112 2148 2118 2150
rect 1810 2139 2118 2148
rect 2608 1782 2636 2246
rect 3130 2204 3438 2213
rect 3130 2202 3136 2204
rect 3192 2202 3216 2204
rect 3272 2202 3296 2204
rect 3352 2202 3376 2204
rect 3432 2202 3438 2204
rect 3192 2150 3194 2202
rect 3374 2150 3376 2202
rect 3130 2148 3136 2150
rect 3192 2148 3216 2150
rect 3272 2148 3296 2150
rect 3352 2148 3376 2150
rect 3432 2148 3438 2150
rect 3130 2139 3438 2148
rect 3528 1782 3556 2246
rect 4356 1992 4384 2246
rect 4450 2204 4758 2213
rect 4450 2202 4456 2204
rect 4512 2202 4536 2204
rect 4592 2202 4616 2204
rect 4672 2202 4696 2204
rect 4752 2202 4758 2204
rect 4512 2150 4514 2202
rect 4694 2150 4696 2202
rect 4450 2148 4456 2150
rect 4512 2148 4536 2150
rect 4592 2148 4616 2150
rect 4672 2148 4696 2150
rect 4752 2148 4758 2150
rect 4450 2139 4758 2148
rect 4356 1964 4476 1992
rect 4356 1962 4384 1964
rect 4448 1782 4476 1964
rect 5368 1782 5396 2246
rect 5770 2204 6078 2213
rect 5770 2202 5776 2204
rect 5832 2202 5856 2204
rect 5912 2202 5936 2204
rect 5992 2202 6016 2204
rect 6072 2202 6078 2204
rect 5832 2150 5834 2202
rect 6014 2150 6016 2202
rect 5770 2148 5776 2150
rect 5832 2148 5856 2150
rect 5912 2148 5936 2150
rect 5992 2148 6016 2150
rect 6072 2148 6078 2150
rect 5770 2139 6078 2148
rect 6288 1782 6316 2246
rect 7024 1952 7052 2246
rect 7090 2204 7398 2213
rect 7090 2202 7096 2204
rect 7152 2202 7176 2204
rect 7232 2202 7256 2204
rect 7312 2202 7336 2204
rect 7392 2202 7398 2204
rect 7152 2150 7154 2202
rect 7334 2150 7336 2202
rect 7090 2148 7096 2150
rect 7152 2148 7176 2150
rect 7232 2148 7256 2150
rect 7312 2148 7336 2150
rect 7392 2148 7398 2150
rect 7090 2139 7398 2148
rect 7024 1924 7236 1952
rect 7208 1782 7236 1924
rect 8128 1782 8156 2264
rect 8208 2246 8260 2252
rect 8410 2204 8718 2213
rect 8410 2202 8416 2204
rect 8472 2202 8496 2204
rect 8552 2202 8576 2204
rect 8632 2202 8656 2204
rect 8712 2202 8718 2204
rect 8472 2150 8474 2202
rect 8654 2150 8656 2202
rect 8410 2148 8416 2150
rect 8472 2148 8496 2150
rect 8552 2148 8576 2150
rect 8632 2148 8656 2150
rect 8712 2148 8718 2150
rect 8410 2139 8718 2148
rect 9048 1782 9076 2518
rect 754 982 810 1782
rect 1674 982 1730 1782
rect 2594 982 2650 1782
rect 3514 982 3570 1782
rect 4434 982 4490 1782
rect 5354 982 5410 1782
rect 6274 982 6330 1782
rect 7194 982 7250 1782
rect 8114 982 8170 1782
rect 9034 982 9090 1782
<< via2 >>
rect 1816 9818 1872 9820
rect 1896 9818 1952 9820
rect 1976 9818 2032 9820
rect 2056 9818 2112 9820
rect 1816 9766 1862 9818
rect 1862 9766 1872 9818
rect 1896 9766 1926 9818
rect 1926 9766 1938 9818
rect 1938 9766 1952 9818
rect 1976 9766 1990 9818
rect 1990 9766 2002 9818
rect 2002 9766 2032 9818
rect 2056 9766 2066 9818
rect 2066 9766 2112 9818
rect 1816 9764 1872 9766
rect 1896 9764 1952 9766
rect 1976 9764 2032 9766
rect 2056 9764 2112 9766
rect 3136 9818 3192 9820
rect 3216 9818 3272 9820
rect 3296 9818 3352 9820
rect 3376 9818 3432 9820
rect 3136 9766 3182 9818
rect 3182 9766 3192 9818
rect 3216 9766 3246 9818
rect 3246 9766 3258 9818
rect 3258 9766 3272 9818
rect 3296 9766 3310 9818
rect 3310 9766 3322 9818
rect 3322 9766 3352 9818
rect 3376 9766 3386 9818
rect 3386 9766 3432 9818
rect 3136 9764 3192 9766
rect 3216 9764 3272 9766
rect 3296 9764 3352 9766
rect 3376 9764 3432 9766
rect 4456 9818 4512 9820
rect 4536 9818 4592 9820
rect 4616 9818 4672 9820
rect 4696 9818 4752 9820
rect 4456 9766 4502 9818
rect 4502 9766 4512 9818
rect 4536 9766 4566 9818
rect 4566 9766 4578 9818
rect 4578 9766 4592 9818
rect 4616 9766 4630 9818
rect 4630 9766 4642 9818
rect 4642 9766 4672 9818
rect 4696 9766 4706 9818
rect 4706 9766 4752 9818
rect 4456 9764 4512 9766
rect 4536 9764 4592 9766
rect 4616 9764 4672 9766
rect 4696 9764 4752 9766
rect 5776 9818 5832 9820
rect 5856 9818 5912 9820
rect 5936 9818 5992 9820
rect 6016 9818 6072 9820
rect 5776 9766 5822 9818
rect 5822 9766 5832 9818
rect 5856 9766 5886 9818
rect 5886 9766 5898 9818
rect 5898 9766 5912 9818
rect 5936 9766 5950 9818
rect 5950 9766 5962 9818
rect 5962 9766 5992 9818
rect 6016 9766 6026 9818
rect 6026 9766 6072 9818
rect 5776 9764 5832 9766
rect 5856 9764 5912 9766
rect 5936 9764 5992 9766
rect 6016 9764 6072 9766
rect 1156 9274 1212 9276
rect 1236 9274 1292 9276
rect 1316 9274 1372 9276
rect 1396 9274 1452 9276
rect 1156 9222 1202 9274
rect 1202 9222 1212 9274
rect 1236 9222 1266 9274
rect 1266 9222 1278 9274
rect 1278 9222 1292 9274
rect 1316 9222 1330 9274
rect 1330 9222 1342 9274
rect 1342 9222 1372 9274
rect 1396 9222 1406 9274
rect 1406 9222 1452 9274
rect 1156 9220 1212 9222
rect 1236 9220 1292 9222
rect 1316 9220 1372 9222
rect 1396 9220 1452 9222
rect 1816 8730 1872 8732
rect 1896 8730 1952 8732
rect 1976 8730 2032 8732
rect 2056 8730 2112 8732
rect 1816 8678 1862 8730
rect 1862 8678 1872 8730
rect 1896 8678 1926 8730
rect 1926 8678 1938 8730
rect 1938 8678 1952 8730
rect 1976 8678 1990 8730
rect 1990 8678 2002 8730
rect 2002 8678 2032 8730
rect 2056 8678 2066 8730
rect 2066 8678 2112 8730
rect 1816 8676 1872 8678
rect 1896 8676 1952 8678
rect 1976 8676 2032 8678
rect 2056 8676 2112 8678
rect 1156 8186 1212 8188
rect 1236 8186 1292 8188
rect 1316 8186 1372 8188
rect 1396 8186 1452 8188
rect 1156 8134 1202 8186
rect 1202 8134 1212 8186
rect 1236 8134 1266 8186
rect 1266 8134 1278 8186
rect 1278 8134 1292 8186
rect 1316 8134 1330 8186
rect 1330 8134 1342 8186
rect 1342 8134 1372 8186
rect 1396 8134 1406 8186
rect 1406 8134 1452 8186
rect 1156 8132 1212 8134
rect 1236 8132 1292 8134
rect 1316 8132 1372 8134
rect 1396 8132 1452 8134
rect 2476 9274 2532 9276
rect 2556 9274 2612 9276
rect 2636 9274 2692 9276
rect 2716 9274 2772 9276
rect 2476 9222 2522 9274
rect 2522 9222 2532 9274
rect 2556 9222 2586 9274
rect 2586 9222 2598 9274
rect 2598 9222 2612 9274
rect 2636 9222 2650 9274
rect 2650 9222 2662 9274
rect 2662 9222 2692 9274
rect 2716 9222 2726 9274
rect 2726 9222 2772 9274
rect 2476 9220 2532 9222
rect 2556 9220 2612 9222
rect 2636 9220 2692 9222
rect 2716 9220 2772 9222
rect 3796 9274 3852 9276
rect 3876 9274 3932 9276
rect 3956 9274 4012 9276
rect 4036 9274 4092 9276
rect 3796 9222 3842 9274
rect 3842 9222 3852 9274
rect 3876 9222 3906 9274
rect 3906 9222 3918 9274
rect 3918 9222 3932 9274
rect 3956 9222 3970 9274
rect 3970 9222 3982 9274
rect 3982 9222 4012 9274
rect 4036 9222 4046 9274
rect 4046 9222 4092 9274
rect 3796 9220 3852 9222
rect 3876 9220 3932 9222
rect 3956 9220 4012 9222
rect 4036 9220 4092 9222
rect 5116 9274 5172 9276
rect 5196 9274 5252 9276
rect 5276 9274 5332 9276
rect 5356 9274 5412 9276
rect 5116 9222 5162 9274
rect 5162 9222 5172 9274
rect 5196 9222 5226 9274
rect 5226 9222 5238 9274
rect 5238 9222 5252 9274
rect 5276 9222 5290 9274
rect 5290 9222 5302 9274
rect 5302 9222 5332 9274
rect 5356 9222 5366 9274
rect 5366 9222 5412 9274
rect 5116 9220 5172 9222
rect 5196 9220 5252 9222
rect 5276 9220 5332 9222
rect 5356 9220 5412 9222
rect 6436 9274 6492 9276
rect 6516 9274 6572 9276
rect 6596 9274 6652 9276
rect 6676 9274 6732 9276
rect 6436 9222 6482 9274
rect 6482 9222 6492 9274
rect 6516 9222 6546 9274
rect 6546 9222 6558 9274
rect 6558 9222 6572 9274
rect 6596 9222 6610 9274
rect 6610 9222 6622 9274
rect 6622 9222 6652 9274
rect 6676 9222 6686 9274
rect 6686 9222 6732 9274
rect 6436 9220 6492 9222
rect 6516 9220 6572 9222
rect 6596 9220 6652 9222
rect 6676 9220 6732 9222
rect 3136 8730 3192 8732
rect 3216 8730 3272 8732
rect 3296 8730 3352 8732
rect 3376 8730 3432 8732
rect 3136 8678 3182 8730
rect 3182 8678 3192 8730
rect 3216 8678 3246 8730
rect 3246 8678 3258 8730
rect 3258 8678 3272 8730
rect 3296 8678 3310 8730
rect 3310 8678 3322 8730
rect 3322 8678 3352 8730
rect 3376 8678 3386 8730
rect 3386 8678 3432 8730
rect 3136 8676 3192 8678
rect 3216 8676 3272 8678
rect 3296 8676 3352 8678
rect 3376 8676 3432 8678
rect 4456 8730 4512 8732
rect 4536 8730 4592 8732
rect 4616 8730 4672 8732
rect 4696 8730 4752 8732
rect 4456 8678 4502 8730
rect 4502 8678 4512 8730
rect 4536 8678 4566 8730
rect 4566 8678 4578 8730
rect 4578 8678 4592 8730
rect 4616 8678 4630 8730
rect 4630 8678 4642 8730
rect 4642 8678 4672 8730
rect 4696 8678 4706 8730
rect 4706 8678 4752 8730
rect 4456 8676 4512 8678
rect 4536 8676 4592 8678
rect 4616 8676 4672 8678
rect 4696 8676 4752 8678
rect 5776 8730 5832 8732
rect 5856 8730 5912 8732
rect 5936 8730 5992 8732
rect 6016 8730 6072 8732
rect 5776 8678 5822 8730
rect 5822 8678 5832 8730
rect 5856 8678 5886 8730
rect 5886 8678 5898 8730
rect 5898 8678 5912 8730
rect 5936 8678 5950 8730
rect 5950 8678 5962 8730
rect 5962 8678 5992 8730
rect 6016 8678 6026 8730
rect 6026 8678 6072 8730
rect 5776 8676 5832 8678
rect 5856 8676 5912 8678
rect 5936 8676 5992 8678
rect 6016 8676 6072 8678
rect 1816 7642 1872 7644
rect 1896 7642 1952 7644
rect 1976 7642 2032 7644
rect 2056 7642 2112 7644
rect 1816 7590 1862 7642
rect 1862 7590 1872 7642
rect 1896 7590 1926 7642
rect 1926 7590 1938 7642
rect 1938 7590 1952 7642
rect 1976 7590 1990 7642
rect 1990 7590 2002 7642
rect 2002 7590 2032 7642
rect 2056 7590 2066 7642
rect 2066 7590 2112 7642
rect 1816 7588 1872 7590
rect 1896 7588 1952 7590
rect 1976 7588 2032 7590
rect 2056 7588 2112 7590
rect 2476 8186 2532 8188
rect 2556 8186 2612 8188
rect 2636 8186 2692 8188
rect 2716 8186 2772 8188
rect 2476 8134 2522 8186
rect 2522 8134 2532 8186
rect 2556 8134 2586 8186
rect 2586 8134 2598 8186
rect 2598 8134 2612 8186
rect 2636 8134 2650 8186
rect 2650 8134 2662 8186
rect 2662 8134 2692 8186
rect 2716 8134 2726 8186
rect 2726 8134 2772 8186
rect 2476 8132 2532 8134
rect 2556 8132 2612 8134
rect 2636 8132 2692 8134
rect 2716 8132 2772 8134
rect 1156 7098 1212 7100
rect 1236 7098 1292 7100
rect 1316 7098 1372 7100
rect 1396 7098 1452 7100
rect 1156 7046 1202 7098
rect 1202 7046 1212 7098
rect 1236 7046 1266 7098
rect 1266 7046 1278 7098
rect 1278 7046 1292 7098
rect 1316 7046 1330 7098
rect 1330 7046 1342 7098
rect 1342 7046 1372 7098
rect 1396 7046 1406 7098
rect 1406 7046 1452 7098
rect 1156 7044 1212 7046
rect 1236 7044 1292 7046
rect 1316 7044 1372 7046
rect 1396 7044 1452 7046
rect 1156 6010 1212 6012
rect 1236 6010 1292 6012
rect 1316 6010 1372 6012
rect 1396 6010 1452 6012
rect 1156 5958 1202 6010
rect 1202 5958 1212 6010
rect 1236 5958 1266 6010
rect 1266 5958 1278 6010
rect 1278 5958 1292 6010
rect 1316 5958 1330 6010
rect 1330 5958 1342 6010
rect 1342 5958 1372 6010
rect 1396 5958 1406 6010
rect 1406 5958 1452 6010
rect 1156 5956 1212 5958
rect 1236 5956 1292 5958
rect 1316 5956 1372 5958
rect 1396 5956 1452 5958
rect 1156 4922 1212 4924
rect 1236 4922 1292 4924
rect 1316 4922 1372 4924
rect 1396 4922 1452 4924
rect 1156 4870 1202 4922
rect 1202 4870 1212 4922
rect 1236 4870 1266 4922
rect 1266 4870 1278 4922
rect 1278 4870 1292 4922
rect 1316 4870 1330 4922
rect 1330 4870 1342 4922
rect 1342 4870 1372 4922
rect 1396 4870 1406 4922
rect 1406 4870 1452 4922
rect 1156 4868 1212 4870
rect 1236 4868 1292 4870
rect 1316 4868 1372 4870
rect 1396 4868 1452 4870
rect 1156 3834 1212 3836
rect 1236 3834 1292 3836
rect 1316 3834 1372 3836
rect 1396 3834 1452 3836
rect 1156 3782 1202 3834
rect 1202 3782 1212 3834
rect 1236 3782 1266 3834
rect 1266 3782 1278 3834
rect 1278 3782 1292 3834
rect 1316 3782 1330 3834
rect 1330 3782 1342 3834
rect 1342 3782 1372 3834
rect 1396 3782 1406 3834
rect 1406 3782 1452 3834
rect 1156 3780 1212 3782
rect 1236 3780 1292 3782
rect 1316 3780 1372 3782
rect 1396 3780 1452 3782
rect 1156 2746 1212 2748
rect 1236 2746 1292 2748
rect 1316 2746 1372 2748
rect 1396 2746 1452 2748
rect 1156 2694 1202 2746
rect 1202 2694 1212 2746
rect 1236 2694 1266 2746
rect 1266 2694 1278 2746
rect 1278 2694 1292 2746
rect 1316 2694 1330 2746
rect 1330 2694 1342 2746
rect 1342 2694 1372 2746
rect 1396 2694 1406 2746
rect 1406 2694 1452 2746
rect 1156 2692 1212 2694
rect 1236 2692 1292 2694
rect 1316 2692 1372 2694
rect 1396 2692 1452 2694
rect 3796 8186 3852 8188
rect 3876 8186 3932 8188
rect 3956 8186 4012 8188
rect 4036 8186 4092 8188
rect 3796 8134 3842 8186
rect 3842 8134 3852 8186
rect 3876 8134 3906 8186
rect 3906 8134 3918 8186
rect 3918 8134 3932 8186
rect 3956 8134 3970 8186
rect 3970 8134 3982 8186
rect 3982 8134 4012 8186
rect 4036 8134 4046 8186
rect 4046 8134 4092 8186
rect 3796 8132 3852 8134
rect 3876 8132 3932 8134
rect 3956 8132 4012 8134
rect 4036 8132 4092 8134
rect 5116 8186 5172 8188
rect 5196 8186 5252 8188
rect 5276 8186 5332 8188
rect 5356 8186 5412 8188
rect 5116 8134 5162 8186
rect 5162 8134 5172 8186
rect 5196 8134 5226 8186
rect 5226 8134 5238 8186
rect 5238 8134 5252 8186
rect 5276 8134 5290 8186
rect 5290 8134 5302 8186
rect 5302 8134 5332 8186
rect 5356 8134 5366 8186
rect 5366 8134 5412 8186
rect 5116 8132 5172 8134
rect 5196 8132 5252 8134
rect 5276 8132 5332 8134
rect 5356 8132 5412 8134
rect 6436 8186 6492 8188
rect 6516 8186 6572 8188
rect 6596 8186 6652 8188
rect 6676 8186 6732 8188
rect 6436 8134 6482 8186
rect 6482 8134 6492 8186
rect 6516 8134 6546 8186
rect 6546 8134 6558 8186
rect 6558 8134 6572 8186
rect 6596 8134 6610 8186
rect 6610 8134 6622 8186
rect 6622 8134 6652 8186
rect 6676 8134 6686 8186
rect 6686 8134 6732 8186
rect 6436 8132 6492 8134
rect 6516 8132 6572 8134
rect 6596 8132 6652 8134
rect 6676 8132 6732 8134
rect 3136 7642 3192 7644
rect 3216 7642 3272 7644
rect 3296 7642 3352 7644
rect 3376 7642 3432 7644
rect 3136 7590 3182 7642
rect 3182 7590 3192 7642
rect 3216 7590 3246 7642
rect 3246 7590 3258 7642
rect 3258 7590 3272 7642
rect 3296 7590 3310 7642
rect 3310 7590 3322 7642
rect 3322 7590 3352 7642
rect 3376 7590 3386 7642
rect 3386 7590 3432 7642
rect 3136 7588 3192 7590
rect 3216 7588 3272 7590
rect 3296 7588 3352 7590
rect 3376 7588 3432 7590
rect 4456 7642 4512 7644
rect 4536 7642 4592 7644
rect 4616 7642 4672 7644
rect 4696 7642 4752 7644
rect 4456 7590 4502 7642
rect 4502 7590 4512 7642
rect 4536 7590 4566 7642
rect 4566 7590 4578 7642
rect 4578 7590 4592 7642
rect 4616 7590 4630 7642
rect 4630 7590 4642 7642
rect 4642 7590 4672 7642
rect 4696 7590 4706 7642
rect 4706 7590 4752 7642
rect 4456 7588 4512 7590
rect 4536 7588 4592 7590
rect 4616 7588 4672 7590
rect 4696 7588 4752 7590
rect 5776 7642 5832 7644
rect 5856 7642 5912 7644
rect 5936 7642 5992 7644
rect 6016 7642 6072 7644
rect 5776 7590 5822 7642
rect 5822 7590 5832 7642
rect 5856 7590 5886 7642
rect 5886 7590 5898 7642
rect 5898 7590 5912 7642
rect 5936 7590 5950 7642
rect 5950 7590 5962 7642
rect 5962 7590 5992 7642
rect 6016 7590 6026 7642
rect 6026 7590 6072 7642
rect 5776 7588 5832 7590
rect 5856 7588 5912 7590
rect 5936 7588 5992 7590
rect 6016 7588 6072 7590
rect 1816 6554 1872 6556
rect 1896 6554 1952 6556
rect 1976 6554 2032 6556
rect 2056 6554 2112 6556
rect 1816 6502 1862 6554
rect 1862 6502 1872 6554
rect 1896 6502 1926 6554
rect 1926 6502 1938 6554
rect 1938 6502 1952 6554
rect 1976 6502 1990 6554
rect 1990 6502 2002 6554
rect 2002 6502 2032 6554
rect 2056 6502 2066 6554
rect 2066 6502 2112 6554
rect 1816 6500 1872 6502
rect 1896 6500 1952 6502
rect 1976 6500 2032 6502
rect 2056 6500 2112 6502
rect 2476 7098 2532 7100
rect 2556 7098 2612 7100
rect 2636 7098 2692 7100
rect 2716 7098 2772 7100
rect 2476 7046 2522 7098
rect 2522 7046 2532 7098
rect 2556 7046 2586 7098
rect 2586 7046 2598 7098
rect 2598 7046 2612 7098
rect 2636 7046 2650 7098
rect 2650 7046 2662 7098
rect 2662 7046 2692 7098
rect 2716 7046 2726 7098
rect 2726 7046 2772 7098
rect 2476 7044 2532 7046
rect 2556 7044 2612 7046
rect 2636 7044 2692 7046
rect 2716 7044 2772 7046
rect 2476 6010 2532 6012
rect 2556 6010 2612 6012
rect 2636 6010 2692 6012
rect 2716 6010 2772 6012
rect 2476 5958 2522 6010
rect 2522 5958 2532 6010
rect 2556 5958 2586 6010
rect 2586 5958 2598 6010
rect 2598 5958 2612 6010
rect 2636 5958 2650 6010
rect 2650 5958 2662 6010
rect 2662 5958 2692 6010
rect 2716 5958 2726 6010
rect 2726 5958 2772 6010
rect 2476 5956 2532 5958
rect 2556 5956 2612 5958
rect 2636 5956 2692 5958
rect 2716 5956 2772 5958
rect 1816 5466 1872 5468
rect 1896 5466 1952 5468
rect 1976 5466 2032 5468
rect 2056 5466 2112 5468
rect 1816 5414 1862 5466
rect 1862 5414 1872 5466
rect 1896 5414 1926 5466
rect 1926 5414 1938 5466
rect 1938 5414 1952 5466
rect 1976 5414 1990 5466
rect 1990 5414 2002 5466
rect 2002 5414 2032 5466
rect 2056 5414 2066 5466
rect 2066 5414 2112 5466
rect 1816 5412 1872 5414
rect 1896 5412 1952 5414
rect 1976 5412 2032 5414
rect 2056 5412 2112 5414
rect 2476 4922 2532 4924
rect 2556 4922 2612 4924
rect 2636 4922 2692 4924
rect 2716 4922 2772 4924
rect 2476 4870 2522 4922
rect 2522 4870 2532 4922
rect 2556 4870 2586 4922
rect 2586 4870 2598 4922
rect 2598 4870 2612 4922
rect 2636 4870 2650 4922
rect 2650 4870 2662 4922
rect 2662 4870 2692 4922
rect 2716 4870 2726 4922
rect 2726 4870 2772 4922
rect 2476 4868 2532 4870
rect 2556 4868 2612 4870
rect 2636 4868 2692 4870
rect 2716 4868 2772 4870
rect 3796 7098 3852 7100
rect 3876 7098 3932 7100
rect 3956 7098 4012 7100
rect 4036 7098 4092 7100
rect 3796 7046 3842 7098
rect 3842 7046 3852 7098
rect 3876 7046 3906 7098
rect 3906 7046 3918 7098
rect 3918 7046 3932 7098
rect 3956 7046 3970 7098
rect 3970 7046 3982 7098
rect 3982 7046 4012 7098
rect 4036 7046 4046 7098
rect 4046 7046 4092 7098
rect 3796 7044 3852 7046
rect 3876 7044 3932 7046
rect 3956 7044 4012 7046
rect 4036 7044 4092 7046
rect 5116 7098 5172 7100
rect 5196 7098 5252 7100
rect 5276 7098 5332 7100
rect 5356 7098 5412 7100
rect 5116 7046 5162 7098
rect 5162 7046 5172 7098
rect 5196 7046 5226 7098
rect 5226 7046 5238 7098
rect 5238 7046 5252 7098
rect 5276 7046 5290 7098
rect 5290 7046 5302 7098
rect 5302 7046 5332 7098
rect 5356 7046 5366 7098
rect 5366 7046 5412 7098
rect 5116 7044 5172 7046
rect 5196 7044 5252 7046
rect 5276 7044 5332 7046
rect 5356 7044 5412 7046
rect 6436 7098 6492 7100
rect 6516 7098 6572 7100
rect 6596 7098 6652 7100
rect 6676 7098 6732 7100
rect 6436 7046 6482 7098
rect 6482 7046 6492 7098
rect 6516 7046 6546 7098
rect 6546 7046 6558 7098
rect 6558 7046 6572 7098
rect 6596 7046 6610 7098
rect 6610 7046 6622 7098
rect 6622 7046 6652 7098
rect 6676 7046 6686 7098
rect 6686 7046 6732 7098
rect 6436 7044 6492 7046
rect 6516 7044 6572 7046
rect 6596 7044 6652 7046
rect 6676 7044 6732 7046
rect 7096 9818 7152 9820
rect 7176 9818 7232 9820
rect 7256 9818 7312 9820
rect 7336 9818 7392 9820
rect 7096 9766 7142 9818
rect 7142 9766 7152 9818
rect 7176 9766 7206 9818
rect 7206 9766 7218 9818
rect 7218 9766 7232 9818
rect 7256 9766 7270 9818
rect 7270 9766 7282 9818
rect 7282 9766 7312 9818
rect 7336 9766 7346 9818
rect 7346 9766 7392 9818
rect 7096 9764 7152 9766
rect 7176 9764 7232 9766
rect 7256 9764 7312 9766
rect 7336 9764 7392 9766
rect 8416 9818 8472 9820
rect 8496 9818 8552 9820
rect 8576 9818 8632 9820
rect 8656 9818 8712 9820
rect 8416 9766 8462 9818
rect 8462 9766 8472 9818
rect 8496 9766 8526 9818
rect 8526 9766 8538 9818
rect 8538 9766 8552 9818
rect 8576 9766 8590 9818
rect 8590 9766 8602 9818
rect 8602 9766 8632 9818
rect 8656 9766 8666 9818
rect 8666 9766 8712 9818
rect 8416 9764 8472 9766
rect 8496 9764 8552 9766
rect 8576 9764 8632 9766
rect 8656 9764 8712 9766
rect 7756 9274 7812 9276
rect 7836 9274 7892 9276
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 7756 9222 7802 9274
rect 7802 9222 7812 9274
rect 7836 9222 7866 9274
rect 7866 9222 7878 9274
rect 7878 9222 7892 9274
rect 7916 9222 7930 9274
rect 7930 9222 7942 9274
rect 7942 9222 7972 9274
rect 7996 9222 8006 9274
rect 8006 9222 8052 9274
rect 7756 9220 7812 9222
rect 7836 9220 7892 9222
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 7096 8730 7152 8732
rect 7176 8730 7232 8732
rect 7256 8730 7312 8732
rect 7336 8730 7392 8732
rect 7096 8678 7142 8730
rect 7142 8678 7152 8730
rect 7176 8678 7206 8730
rect 7206 8678 7218 8730
rect 7218 8678 7232 8730
rect 7256 8678 7270 8730
rect 7270 8678 7282 8730
rect 7282 8678 7312 8730
rect 7336 8678 7346 8730
rect 7346 8678 7392 8730
rect 7096 8676 7152 8678
rect 7176 8676 7232 8678
rect 7256 8676 7312 8678
rect 7336 8676 7392 8678
rect 8416 8730 8472 8732
rect 8496 8730 8552 8732
rect 8576 8730 8632 8732
rect 8656 8730 8712 8732
rect 8416 8678 8462 8730
rect 8462 8678 8472 8730
rect 8496 8678 8526 8730
rect 8526 8678 8538 8730
rect 8538 8678 8552 8730
rect 8576 8678 8590 8730
rect 8590 8678 8602 8730
rect 8602 8678 8632 8730
rect 8656 8678 8666 8730
rect 8666 8678 8712 8730
rect 8416 8676 8472 8678
rect 8496 8676 8552 8678
rect 8576 8676 8632 8678
rect 8656 8676 8712 8678
rect 7756 8186 7812 8188
rect 7836 8186 7892 8188
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 7756 8134 7802 8186
rect 7802 8134 7812 8186
rect 7836 8134 7866 8186
rect 7866 8134 7878 8186
rect 7878 8134 7892 8186
rect 7916 8134 7930 8186
rect 7930 8134 7942 8186
rect 7942 8134 7972 8186
rect 7996 8134 8006 8186
rect 8006 8134 8052 8186
rect 7756 8132 7812 8134
rect 7836 8132 7892 8134
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 7096 7642 7152 7644
rect 7176 7642 7232 7644
rect 7256 7642 7312 7644
rect 7336 7642 7392 7644
rect 7096 7590 7142 7642
rect 7142 7590 7152 7642
rect 7176 7590 7206 7642
rect 7206 7590 7218 7642
rect 7218 7590 7232 7642
rect 7256 7590 7270 7642
rect 7270 7590 7282 7642
rect 7282 7590 7312 7642
rect 7336 7590 7346 7642
rect 7346 7590 7392 7642
rect 7096 7588 7152 7590
rect 7176 7588 7232 7590
rect 7256 7588 7312 7590
rect 7336 7588 7392 7590
rect 8416 7642 8472 7644
rect 8496 7642 8552 7644
rect 8576 7642 8632 7644
rect 8656 7642 8712 7644
rect 8416 7590 8462 7642
rect 8462 7590 8472 7642
rect 8496 7590 8526 7642
rect 8526 7590 8538 7642
rect 8538 7590 8552 7642
rect 8576 7590 8590 7642
rect 8590 7590 8602 7642
rect 8602 7590 8632 7642
rect 8656 7590 8666 7642
rect 8666 7590 8712 7642
rect 8416 7588 8472 7590
rect 8496 7588 8552 7590
rect 8576 7588 8632 7590
rect 8656 7588 8712 7590
rect 7756 7098 7812 7100
rect 7836 7098 7892 7100
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 7756 7046 7802 7098
rect 7802 7046 7812 7098
rect 7836 7046 7866 7098
rect 7866 7046 7878 7098
rect 7878 7046 7892 7098
rect 7916 7046 7930 7098
rect 7930 7046 7942 7098
rect 7942 7046 7972 7098
rect 7996 7046 8006 7098
rect 8006 7046 8052 7098
rect 7756 7044 7812 7046
rect 7836 7044 7892 7046
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 3136 6554 3192 6556
rect 3216 6554 3272 6556
rect 3296 6554 3352 6556
rect 3376 6554 3432 6556
rect 3136 6502 3182 6554
rect 3182 6502 3192 6554
rect 3216 6502 3246 6554
rect 3246 6502 3258 6554
rect 3258 6502 3272 6554
rect 3296 6502 3310 6554
rect 3310 6502 3322 6554
rect 3322 6502 3352 6554
rect 3376 6502 3386 6554
rect 3386 6502 3432 6554
rect 3136 6500 3192 6502
rect 3216 6500 3272 6502
rect 3296 6500 3352 6502
rect 3376 6500 3432 6502
rect 4456 6554 4512 6556
rect 4536 6554 4592 6556
rect 4616 6554 4672 6556
rect 4696 6554 4752 6556
rect 4456 6502 4502 6554
rect 4502 6502 4512 6554
rect 4536 6502 4566 6554
rect 4566 6502 4578 6554
rect 4578 6502 4592 6554
rect 4616 6502 4630 6554
rect 4630 6502 4642 6554
rect 4642 6502 4672 6554
rect 4696 6502 4706 6554
rect 4706 6502 4752 6554
rect 4456 6500 4512 6502
rect 4536 6500 4592 6502
rect 4616 6500 4672 6502
rect 4696 6500 4752 6502
rect 5776 6554 5832 6556
rect 5856 6554 5912 6556
rect 5936 6554 5992 6556
rect 6016 6554 6072 6556
rect 5776 6502 5822 6554
rect 5822 6502 5832 6554
rect 5856 6502 5886 6554
rect 5886 6502 5898 6554
rect 5898 6502 5912 6554
rect 5936 6502 5950 6554
rect 5950 6502 5962 6554
rect 5962 6502 5992 6554
rect 6016 6502 6026 6554
rect 6026 6502 6072 6554
rect 5776 6500 5832 6502
rect 5856 6500 5912 6502
rect 5936 6500 5992 6502
rect 6016 6500 6072 6502
rect 3796 6010 3852 6012
rect 3876 6010 3932 6012
rect 3956 6010 4012 6012
rect 4036 6010 4092 6012
rect 3796 5958 3842 6010
rect 3842 5958 3852 6010
rect 3876 5958 3906 6010
rect 3906 5958 3918 6010
rect 3918 5958 3932 6010
rect 3956 5958 3970 6010
rect 3970 5958 3982 6010
rect 3982 5958 4012 6010
rect 4036 5958 4046 6010
rect 4046 5958 4092 6010
rect 3796 5956 3852 5958
rect 3876 5956 3932 5958
rect 3956 5956 4012 5958
rect 4036 5956 4092 5958
rect 5116 6010 5172 6012
rect 5196 6010 5252 6012
rect 5276 6010 5332 6012
rect 5356 6010 5412 6012
rect 5116 5958 5162 6010
rect 5162 5958 5172 6010
rect 5196 5958 5226 6010
rect 5226 5958 5238 6010
rect 5238 5958 5252 6010
rect 5276 5958 5290 6010
rect 5290 5958 5302 6010
rect 5302 5958 5332 6010
rect 5356 5958 5366 6010
rect 5366 5958 5412 6010
rect 5116 5956 5172 5958
rect 5196 5956 5252 5958
rect 5276 5956 5332 5958
rect 5356 5956 5412 5958
rect 6436 6010 6492 6012
rect 6516 6010 6572 6012
rect 6596 6010 6652 6012
rect 6676 6010 6732 6012
rect 6436 5958 6482 6010
rect 6482 5958 6492 6010
rect 6516 5958 6546 6010
rect 6546 5958 6558 6010
rect 6558 5958 6572 6010
rect 6596 5958 6610 6010
rect 6610 5958 6622 6010
rect 6622 5958 6652 6010
rect 6676 5958 6686 6010
rect 6686 5958 6732 6010
rect 6436 5956 6492 5958
rect 6516 5956 6572 5958
rect 6596 5956 6652 5958
rect 6676 5956 6732 5958
rect 7096 6554 7152 6556
rect 7176 6554 7232 6556
rect 7256 6554 7312 6556
rect 7336 6554 7392 6556
rect 7096 6502 7142 6554
rect 7142 6502 7152 6554
rect 7176 6502 7206 6554
rect 7206 6502 7218 6554
rect 7218 6502 7232 6554
rect 7256 6502 7270 6554
rect 7270 6502 7282 6554
rect 7282 6502 7312 6554
rect 7336 6502 7346 6554
rect 7346 6502 7392 6554
rect 7096 6500 7152 6502
rect 7176 6500 7232 6502
rect 7256 6500 7312 6502
rect 7336 6500 7392 6502
rect 8416 6554 8472 6556
rect 8496 6554 8552 6556
rect 8576 6554 8632 6556
rect 8656 6554 8712 6556
rect 8416 6502 8462 6554
rect 8462 6502 8472 6554
rect 8496 6502 8526 6554
rect 8526 6502 8538 6554
rect 8538 6502 8552 6554
rect 8576 6502 8590 6554
rect 8590 6502 8602 6554
rect 8602 6502 8632 6554
rect 8656 6502 8666 6554
rect 8666 6502 8712 6554
rect 8416 6500 8472 6502
rect 8496 6500 8552 6502
rect 8576 6500 8632 6502
rect 8656 6500 8712 6502
rect 7756 6010 7812 6012
rect 7836 6010 7892 6012
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 7756 5958 7802 6010
rect 7802 5958 7812 6010
rect 7836 5958 7866 6010
rect 7866 5958 7878 6010
rect 7878 5958 7892 6010
rect 7916 5958 7930 6010
rect 7930 5958 7942 6010
rect 7942 5958 7972 6010
rect 7996 5958 8006 6010
rect 8006 5958 8052 6010
rect 7756 5956 7812 5958
rect 7836 5956 7892 5958
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 3136 5466 3192 5468
rect 3216 5466 3272 5468
rect 3296 5466 3352 5468
rect 3376 5466 3432 5468
rect 3136 5414 3182 5466
rect 3182 5414 3192 5466
rect 3216 5414 3246 5466
rect 3246 5414 3258 5466
rect 3258 5414 3272 5466
rect 3296 5414 3310 5466
rect 3310 5414 3322 5466
rect 3322 5414 3352 5466
rect 3376 5414 3386 5466
rect 3386 5414 3432 5466
rect 3136 5412 3192 5414
rect 3216 5412 3272 5414
rect 3296 5412 3352 5414
rect 3376 5412 3432 5414
rect 4456 5466 4512 5468
rect 4536 5466 4592 5468
rect 4616 5466 4672 5468
rect 4696 5466 4752 5468
rect 4456 5414 4502 5466
rect 4502 5414 4512 5466
rect 4536 5414 4566 5466
rect 4566 5414 4578 5466
rect 4578 5414 4592 5466
rect 4616 5414 4630 5466
rect 4630 5414 4642 5466
rect 4642 5414 4672 5466
rect 4696 5414 4706 5466
rect 4706 5414 4752 5466
rect 4456 5412 4512 5414
rect 4536 5412 4592 5414
rect 4616 5412 4672 5414
rect 4696 5412 4752 5414
rect 5776 5466 5832 5468
rect 5856 5466 5912 5468
rect 5936 5466 5992 5468
rect 6016 5466 6072 5468
rect 5776 5414 5822 5466
rect 5822 5414 5832 5466
rect 5856 5414 5886 5466
rect 5886 5414 5898 5466
rect 5898 5414 5912 5466
rect 5936 5414 5950 5466
rect 5950 5414 5962 5466
rect 5962 5414 5992 5466
rect 6016 5414 6026 5466
rect 6026 5414 6072 5466
rect 5776 5412 5832 5414
rect 5856 5412 5912 5414
rect 5936 5412 5992 5414
rect 6016 5412 6072 5414
rect 7096 5466 7152 5468
rect 7176 5466 7232 5468
rect 7256 5466 7312 5468
rect 7336 5466 7392 5468
rect 7096 5414 7142 5466
rect 7142 5414 7152 5466
rect 7176 5414 7206 5466
rect 7206 5414 7218 5466
rect 7218 5414 7232 5466
rect 7256 5414 7270 5466
rect 7270 5414 7282 5466
rect 7282 5414 7312 5466
rect 7336 5414 7346 5466
rect 7346 5414 7392 5466
rect 7096 5412 7152 5414
rect 7176 5412 7232 5414
rect 7256 5412 7312 5414
rect 7336 5412 7392 5414
rect 8416 5466 8472 5468
rect 8496 5466 8552 5468
rect 8576 5466 8632 5468
rect 8656 5466 8712 5468
rect 8416 5414 8462 5466
rect 8462 5414 8472 5466
rect 8496 5414 8526 5466
rect 8526 5414 8538 5466
rect 8538 5414 8552 5466
rect 8576 5414 8590 5466
rect 8590 5414 8602 5466
rect 8602 5414 8632 5466
rect 8656 5414 8666 5466
rect 8666 5414 8712 5466
rect 8416 5412 8472 5414
rect 8496 5412 8552 5414
rect 8576 5412 8632 5414
rect 8656 5412 8712 5414
rect 3796 4922 3852 4924
rect 3876 4922 3932 4924
rect 3956 4922 4012 4924
rect 4036 4922 4092 4924
rect 3796 4870 3842 4922
rect 3842 4870 3852 4922
rect 3876 4870 3906 4922
rect 3906 4870 3918 4922
rect 3918 4870 3932 4922
rect 3956 4870 3970 4922
rect 3970 4870 3982 4922
rect 3982 4870 4012 4922
rect 4036 4870 4046 4922
rect 4046 4870 4092 4922
rect 3796 4868 3852 4870
rect 3876 4868 3932 4870
rect 3956 4868 4012 4870
rect 4036 4868 4092 4870
rect 1816 4378 1872 4380
rect 1896 4378 1952 4380
rect 1976 4378 2032 4380
rect 2056 4378 2112 4380
rect 1816 4326 1862 4378
rect 1862 4326 1872 4378
rect 1896 4326 1926 4378
rect 1926 4326 1938 4378
rect 1938 4326 1952 4378
rect 1976 4326 1990 4378
rect 1990 4326 2002 4378
rect 2002 4326 2032 4378
rect 2056 4326 2066 4378
rect 2066 4326 2112 4378
rect 1816 4324 1872 4326
rect 1896 4324 1952 4326
rect 1976 4324 2032 4326
rect 2056 4324 2112 4326
rect 2476 3834 2532 3836
rect 2556 3834 2612 3836
rect 2636 3834 2692 3836
rect 2716 3834 2772 3836
rect 2476 3782 2522 3834
rect 2522 3782 2532 3834
rect 2556 3782 2586 3834
rect 2586 3782 2598 3834
rect 2598 3782 2612 3834
rect 2636 3782 2650 3834
rect 2650 3782 2662 3834
rect 2662 3782 2692 3834
rect 2716 3782 2726 3834
rect 2726 3782 2772 3834
rect 2476 3780 2532 3782
rect 2556 3780 2612 3782
rect 2636 3780 2692 3782
rect 2716 3780 2772 3782
rect 1816 3290 1872 3292
rect 1896 3290 1952 3292
rect 1976 3290 2032 3292
rect 2056 3290 2112 3292
rect 1816 3238 1862 3290
rect 1862 3238 1872 3290
rect 1896 3238 1926 3290
rect 1926 3238 1938 3290
rect 1938 3238 1952 3290
rect 1976 3238 1990 3290
rect 1990 3238 2002 3290
rect 2002 3238 2032 3290
rect 2056 3238 2066 3290
rect 2066 3238 2112 3290
rect 1816 3236 1872 3238
rect 1896 3236 1952 3238
rect 1976 3236 2032 3238
rect 2056 3236 2112 3238
rect 3136 4378 3192 4380
rect 3216 4378 3272 4380
rect 3296 4378 3352 4380
rect 3376 4378 3432 4380
rect 3136 4326 3182 4378
rect 3182 4326 3192 4378
rect 3216 4326 3246 4378
rect 3246 4326 3258 4378
rect 3258 4326 3272 4378
rect 3296 4326 3310 4378
rect 3310 4326 3322 4378
rect 3322 4326 3352 4378
rect 3376 4326 3386 4378
rect 3386 4326 3432 4378
rect 3136 4324 3192 4326
rect 3216 4324 3272 4326
rect 3296 4324 3352 4326
rect 3376 4324 3432 4326
rect 5116 4922 5172 4924
rect 5196 4922 5252 4924
rect 5276 4922 5332 4924
rect 5356 4922 5412 4924
rect 5116 4870 5162 4922
rect 5162 4870 5172 4922
rect 5196 4870 5226 4922
rect 5226 4870 5238 4922
rect 5238 4870 5252 4922
rect 5276 4870 5290 4922
rect 5290 4870 5302 4922
rect 5302 4870 5332 4922
rect 5356 4870 5366 4922
rect 5366 4870 5412 4922
rect 5116 4868 5172 4870
rect 5196 4868 5252 4870
rect 5276 4868 5332 4870
rect 5356 4868 5412 4870
rect 4456 4378 4512 4380
rect 4536 4378 4592 4380
rect 4616 4378 4672 4380
rect 4696 4378 4752 4380
rect 4456 4326 4502 4378
rect 4502 4326 4512 4378
rect 4536 4326 4566 4378
rect 4566 4326 4578 4378
rect 4578 4326 4592 4378
rect 4616 4326 4630 4378
rect 4630 4326 4642 4378
rect 4642 4326 4672 4378
rect 4696 4326 4706 4378
rect 4706 4326 4752 4378
rect 4456 4324 4512 4326
rect 4536 4324 4592 4326
rect 4616 4324 4672 4326
rect 4696 4324 4752 4326
rect 3796 3834 3852 3836
rect 3876 3834 3932 3836
rect 3956 3834 4012 3836
rect 4036 3834 4092 3836
rect 3796 3782 3842 3834
rect 3842 3782 3852 3834
rect 3876 3782 3906 3834
rect 3906 3782 3918 3834
rect 3918 3782 3932 3834
rect 3956 3782 3970 3834
rect 3970 3782 3982 3834
rect 3982 3782 4012 3834
rect 4036 3782 4046 3834
rect 4046 3782 4092 3834
rect 3796 3780 3852 3782
rect 3876 3780 3932 3782
rect 3956 3780 4012 3782
rect 4036 3780 4092 3782
rect 3136 3290 3192 3292
rect 3216 3290 3272 3292
rect 3296 3290 3352 3292
rect 3376 3290 3432 3292
rect 3136 3238 3182 3290
rect 3182 3238 3192 3290
rect 3216 3238 3246 3290
rect 3246 3238 3258 3290
rect 3258 3238 3272 3290
rect 3296 3238 3310 3290
rect 3310 3238 3322 3290
rect 3322 3238 3352 3290
rect 3376 3238 3386 3290
rect 3386 3238 3432 3290
rect 3136 3236 3192 3238
rect 3216 3236 3272 3238
rect 3296 3236 3352 3238
rect 3376 3236 3432 3238
rect 4526 4020 4528 4040
rect 4528 4020 4580 4040
rect 4580 4020 4582 4040
rect 4526 3984 4582 4020
rect 2476 2746 2532 2748
rect 2556 2746 2612 2748
rect 2636 2746 2692 2748
rect 2716 2746 2772 2748
rect 2476 2694 2522 2746
rect 2522 2694 2532 2746
rect 2556 2694 2586 2746
rect 2586 2694 2598 2746
rect 2598 2694 2612 2746
rect 2636 2694 2650 2746
rect 2650 2694 2662 2746
rect 2662 2694 2692 2746
rect 2716 2694 2726 2746
rect 2726 2694 2772 2746
rect 2476 2692 2532 2694
rect 2556 2692 2612 2694
rect 2636 2692 2692 2694
rect 2716 2692 2772 2694
rect 5446 3984 5502 4040
rect 5116 3834 5172 3836
rect 5196 3834 5252 3836
rect 5276 3834 5332 3836
rect 5356 3834 5412 3836
rect 5116 3782 5162 3834
rect 5162 3782 5172 3834
rect 5196 3782 5226 3834
rect 5226 3782 5238 3834
rect 5238 3782 5252 3834
rect 5276 3782 5290 3834
rect 5290 3782 5302 3834
rect 5302 3782 5332 3834
rect 5356 3782 5366 3834
rect 5366 3782 5412 3834
rect 5116 3780 5172 3782
rect 5196 3780 5252 3782
rect 5276 3780 5332 3782
rect 5356 3780 5412 3782
rect 4456 3290 4512 3292
rect 4536 3290 4592 3292
rect 4616 3290 4672 3292
rect 4696 3290 4752 3292
rect 4456 3238 4502 3290
rect 4502 3238 4512 3290
rect 4536 3238 4566 3290
rect 4566 3238 4578 3290
rect 4578 3238 4592 3290
rect 4616 3238 4630 3290
rect 4630 3238 4642 3290
rect 4642 3238 4672 3290
rect 4696 3238 4706 3290
rect 4706 3238 4752 3290
rect 4456 3236 4512 3238
rect 4536 3236 4592 3238
rect 4616 3236 4672 3238
rect 4696 3236 4752 3238
rect 5776 4378 5832 4380
rect 5856 4378 5912 4380
rect 5936 4378 5992 4380
rect 6016 4378 6072 4380
rect 5776 4326 5822 4378
rect 5822 4326 5832 4378
rect 5856 4326 5886 4378
rect 5886 4326 5898 4378
rect 5898 4326 5912 4378
rect 5936 4326 5950 4378
rect 5950 4326 5962 4378
rect 5962 4326 5992 4378
rect 6016 4326 6026 4378
rect 6026 4326 6072 4378
rect 5776 4324 5832 4326
rect 5856 4324 5912 4326
rect 5936 4324 5992 4326
rect 6016 4324 6072 4326
rect 6436 4922 6492 4924
rect 6516 4922 6572 4924
rect 6596 4922 6652 4924
rect 6676 4922 6732 4924
rect 6436 4870 6482 4922
rect 6482 4870 6492 4922
rect 6516 4870 6546 4922
rect 6546 4870 6558 4922
rect 6558 4870 6572 4922
rect 6596 4870 6610 4922
rect 6610 4870 6622 4922
rect 6622 4870 6652 4922
rect 6676 4870 6686 4922
rect 6686 4870 6732 4922
rect 6436 4868 6492 4870
rect 6516 4868 6572 4870
rect 6596 4868 6652 4870
rect 6676 4868 6732 4870
rect 5776 3290 5832 3292
rect 5856 3290 5912 3292
rect 5936 3290 5992 3292
rect 6016 3290 6072 3292
rect 5776 3238 5822 3290
rect 5822 3238 5832 3290
rect 5856 3238 5886 3290
rect 5886 3238 5898 3290
rect 5898 3238 5912 3290
rect 5936 3238 5950 3290
rect 5950 3238 5962 3290
rect 5962 3238 5992 3290
rect 6016 3238 6026 3290
rect 6026 3238 6072 3290
rect 5776 3236 5832 3238
rect 5856 3236 5912 3238
rect 5936 3236 5992 3238
rect 6016 3236 6072 3238
rect 3796 2746 3852 2748
rect 3876 2746 3932 2748
rect 3956 2746 4012 2748
rect 4036 2746 4092 2748
rect 3796 2694 3842 2746
rect 3842 2694 3852 2746
rect 3876 2694 3906 2746
rect 3906 2694 3918 2746
rect 3918 2694 3932 2746
rect 3956 2694 3970 2746
rect 3970 2694 3982 2746
rect 3982 2694 4012 2746
rect 4036 2694 4046 2746
rect 4046 2694 4092 2746
rect 3796 2692 3852 2694
rect 3876 2692 3932 2694
rect 3956 2692 4012 2694
rect 4036 2692 4092 2694
rect 5116 2746 5172 2748
rect 5196 2746 5252 2748
rect 5276 2746 5332 2748
rect 5356 2746 5412 2748
rect 5116 2694 5162 2746
rect 5162 2694 5172 2746
rect 5196 2694 5226 2746
rect 5226 2694 5238 2746
rect 5238 2694 5252 2746
rect 5276 2694 5290 2746
rect 5290 2694 5302 2746
rect 5302 2694 5332 2746
rect 5356 2694 5366 2746
rect 5366 2694 5412 2746
rect 5116 2692 5172 2694
rect 5196 2692 5252 2694
rect 5276 2692 5332 2694
rect 5356 2692 5412 2694
rect 6436 3834 6492 3836
rect 6516 3834 6572 3836
rect 6596 3834 6652 3836
rect 6676 3834 6732 3836
rect 6436 3782 6482 3834
rect 6482 3782 6492 3834
rect 6516 3782 6546 3834
rect 6546 3782 6558 3834
rect 6558 3782 6572 3834
rect 6596 3782 6610 3834
rect 6610 3782 6622 3834
rect 6622 3782 6652 3834
rect 6676 3782 6686 3834
rect 6686 3782 6732 3834
rect 6436 3780 6492 3782
rect 6516 3780 6572 3782
rect 6596 3780 6652 3782
rect 6676 3780 6732 3782
rect 7096 4378 7152 4380
rect 7176 4378 7232 4380
rect 7256 4378 7312 4380
rect 7336 4378 7392 4380
rect 7096 4326 7142 4378
rect 7142 4326 7152 4378
rect 7176 4326 7206 4378
rect 7206 4326 7218 4378
rect 7218 4326 7232 4378
rect 7256 4326 7270 4378
rect 7270 4326 7282 4378
rect 7282 4326 7312 4378
rect 7336 4326 7346 4378
rect 7346 4326 7392 4378
rect 7096 4324 7152 4326
rect 7176 4324 7232 4326
rect 7256 4324 7312 4326
rect 7336 4324 7392 4326
rect 7096 3290 7152 3292
rect 7176 3290 7232 3292
rect 7256 3290 7312 3292
rect 7336 3290 7392 3292
rect 7096 3238 7142 3290
rect 7142 3238 7152 3290
rect 7176 3238 7206 3290
rect 7206 3238 7218 3290
rect 7218 3238 7232 3290
rect 7256 3238 7270 3290
rect 7270 3238 7282 3290
rect 7282 3238 7312 3290
rect 7336 3238 7346 3290
rect 7346 3238 7392 3290
rect 7096 3236 7152 3238
rect 7176 3236 7232 3238
rect 7256 3236 7312 3238
rect 7336 3236 7392 3238
rect 7756 4922 7812 4924
rect 7836 4922 7892 4924
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 7756 4870 7802 4922
rect 7802 4870 7812 4922
rect 7836 4870 7866 4922
rect 7866 4870 7878 4922
rect 7878 4870 7892 4922
rect 7916 4870 7930 4922
rect 7930 4870 7942 4922
rect 7942 4870 7972 4922
rect 7996 4870 8006 4922
rect 8006 4870 8052 4922
rect 7756 4868 7812 4870
rect 7836 4868 7892 4870
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8416 4378 8472 4380
rect 8496 4378 8552 4380
rect 8576 4378 8632 4380
rect 8656 4378 8712 4380
rect 8416 4326 8462 4378
rect 8462 4326 8472 4378
rect 8496 4326 8526 4378
rect 8526 4326 8538 4378
rect 8538 4326 8552 4378
rect 8576 4326 8590 4378
rect 8590 4326 8602 4378
rect 8602 4326 8632 4378
rect 8656 4326 8666 4378
rect 8666 4326 8712 4378
rect 8416 4324 8472 4326
rect 8496 4324 8552 4326
rect 8576 4324 8632 4326
rect 8656 4324 8712 4326
rect 7756 3834 7812 3836
rect 7836 3834 7892 3836
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 7756 3782 7802 3834
rect 7802 3782 7812 3834
rect 7836 3782 7866 3834
rect 7866 3782 7878 3834
rect 7878 3782 7892 3834
rect 7916 3782 7930 3834
rect 7930 3782 7942 3834
rect 7942 3782 7972 3834
rect 7996 3782 8006 3834
rect 8006 3782 8052 3834
rect 7756 3780 7812 3782
rect 7836 3780 7892 3782
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 6436 2746 6492 2748
rect 6516 2746 6572 2748
rect 6596 2746 6652 2748
rect 6676 2746 6732 2748
rect 6436 2694 6482 2746
rect 6482 2694 6492 2746
rect 6516 2694 6546 2746
rect 6546 2694 6558 2746
rect 6558 2694 6572 2746
rect 6596 2694 6610 2746
rect 6610 2694 6622 2746
rect 6622 2694 6652 2746
rect 6676 2694 6686 2746
rect 6686 2694 6732 2746
rect 6436 2692 6492 2694
rect 6516 2692 6572 2694
rect 6596 2692 6652 2694
rect 6676 2692 6732 2694
rect 8416 3290 8472 3292
rect 8496 3290 8552 3292
rect 8576 3290 8632 3292
rect 8656 3290 8712 3292
rect 8416 3238 8462 3290
rect 8462 3238 8472 3290
rect 8496 3238 8526 3290
rect 8526 3238 8538 3290
rect 8538 3238 8552 3290
rect 8576 3238 8590 3290
rect 8590 3238 8602 3290
rect 8602 3238 8632 3290
rect 8656 3238 8666 3290
rect 8666 3238 8712 3290
rect 8416 3236 8472 3238
rect 8496 3236 8552 3238
rect 8576 3236 8632 3238
rect 8656 3236 8712 3238
rect 7756 2746 7812 2748
rect 7836 2746 7892 2748
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 7756 2694 7802 2746
rect 7802 2694 7812 2746
rect 7836 2694 7866 2746
rect 7866 2694 7878 2746
rect 7878 2694 7892 2746
rect 7916 2694 7930 2746
rect 7930 2694 7942 2746
rect 7942 2694 7972 2746
rect 7996 2694 8006 2746
rect 8006 2694 8052 2746
rect 7756 2692 7812 2694
rect 7836 2692 7892 2694
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 1816 2202 1872 2204
rect 1896 2202 1952 2204
rect 1976 2202 2032 2204
rect 2056 2202 2112 2204
rect 1816 2150 1862 2202
rect 1862 2150 1872 2202
rect 1896 2150 1926 2202
rect 1926 2150 1938 2202
rect 1938 2150 1952 2202
rect 1976 2150 1990 2202
rect 1990 2150 2002 2202
rect 2002 2150 2032 2202
rect 2056 2150 2066 2202
rect 2066 2150 2112 2202
rect 1816 2148 1872 2150
rect 1896 2148 1952 2150
rect 1976 2148 2032 2150
rect 2056 2148 2112 2150
rect 3136 2202 3192 2204
rect 3216 2202 3272 2204
rect 3296 2202 3352 2204
rect 3376 2202 3432 2204
rect 3136 2150 3182 2202
rect 3182 2150 3192 2202
rect 3216 2150 3246 2202
rect 3246 2150 3258 2202
rect 3258 2150 3272 2202
rect 3296 2150 3310 2202
rect 3310 2150 3322 2202
rect 3322 2150 3352 2202
rect 3376 2150 3386 2202
rect 3386 2150 3432 2202
rect 3136 2148 3192 2150
rect 3216 2148 3272 2150
rect 3296 2148 3352 2150
rect 3376 2148 3432 2150
rect 4456 2202 4512 2204
rect 4536 2202 4592 2204
rect 4616 2202 4672 2204
rect 4696 2202 4752 2204
rect 4456 2150 4502 2202
rect 4502 2150 4512 2202
rect 4536 2150 4566 2202
rect 4566 2150 4578 2202
rect 4578 2150 4592 2202
rect 4616 2150 4630 2202
rect 4630 2150 4642 2202
rect 4642 2150 4672 2202
rect 4696 2150 4706 2202
rect 4706 2150 4752 2202
rect 4456 2148 4512 2150
rect 4536 2148 4592 2150
rect 4616 2148 4672 2150
rect 4696 2148 4752 2150
rect 5776 2202 5832 2204
rect 5856 2202 5912 2204
rect 5936 2202 5992 2204
rect 6016 2202 6072 2204
rect 5776 2150 5822 2202
rect 5822 2150 5832 2202
rect 5856 2150 5886 2202
rect 5886 2150 5898 2202
rect 5898 2150 5912 2202
rect 5936 2150 5950 2202
rect 5950 2150 5962 2202
rect 5962 2150 5992 2202
rect 6016 2150 6026 2202
rect 6026 2150 6072 2202
rect 5776 2148 5832 2150
rect 5856 2148 5912 2150
rect 5936 2148 5992 2150
rect 6016 2148 6072 2150
rect 7096 2202 7152 2204
rect 7176 2202 7232 2204
rect 7256 2202 7312 2204
rect 7336 2202 7392 2204
rect 7096 2150 7142 2202
rect 7142 2150 7152 2202
rect 7176 2150 7206 2202
rect 7206 2150 7218 2202
rect 7218 2150 7232 2202
rect 7256 2150 7270 2202
rect 7270 2150 7282 2202
rect 7282 2150 7312 2202
rect 7336 2150 7346 2202
rect 7346 2150 7392 2202
rect 7096 2148 7152 2150
rect 7176 2148 7232 2150
rect 7256 2148 7312 2150
rect 7336 2148 7392 2150
rect 8416 2202 8472 2204
rect 8496 2202 8552 2204
rect 8576 2202 8632 2204
rect 8656 2202 8712 2204
rect 8416 2150 8462 2202
rect 8462 2150 8472 2202
rect 8496 2150 8526 2202
rect 8526 2150 8538 2202
rect 8538 2150 8552 2202
rect 8576 2150 8590 2202
rect 8590 2150 8602 2202
rect 8602 2150 8632 2202
rect 8656 2150 8666 2202
rect 8666 2150 8712 2202
rect 8416 2148 8472 2150
rect 8496 2148 8552 2150
rect 8576 2148 8632 2150
rect 8656 2148 8712 2150
<< metal3 >>
rect 1800 10204 8722 10260
rect 1800 10006 2136 10204
rect 8522 10006 8722 10204
rect 1800 9944 8722 10006
rect 1800 9825 2084 9944
rect 1800 9824 2122 9825
rect 1800 9760 1812 9824
rect 1876 9760 1892 9824
rect 1956 9760 1972 9824
rect 2036 9760 2052 9824
rect 2116 9760 2122 9824
rect 1800 9759 2122 9760
rect 3122 9824 3458 9944
rect 4452 9825 4768 9944
rect 5772 9825 6088 9944
rect 7090 9825 7406 9944
rect 3122 9760 3132 9824
rect 3196 9760 3212 9824
rect 3276 9760 3292 9824
rect 3356 9760 3372 9824
rect 3436 9760 3458 9824
rect 1800 9710 2084 9759
rect 3122 9550 3458 9760
rect 4446 9824 4768 9825
rect 4446 9760 4452 9824
rect 4516 9760 4532 9824
rect 4596 9760 4612 9824
rect 4676 9760 4692 9824
rect 4756 9760 4768 9824
rect 4446 9759 4768 9760
rect 5766 9824 6088 9825
rect 5766 9760 5772 9824
rect 5836 9760 5852 9824
rect 5916 9760 5932 9824
rect 5996 9760 6012 9824
rect 6076 9760 6088 9824
rect 5766 9759 6088 9760
rect 7086 9824 7406 9825
rect 7086 9760 7092 9824
rect 7156 9760 7172 9824
rect 7236 9760 7252 9824
rect 7316 9760 7332 9824
rect 7396 9760 7406 9824
rect 7086 9759 7406 9760
rect 4452 9572 4768 9759
rect 5772 9586 6088 9759
rect 7090 9594 7406 9759
rect 8406 9824 8722 9944
rect 8406 9760 8412 9824
rect 8476 9760 8492 9824
rect 8556 9760 8572 9824
rect 8636 9760 8652 9824
rect 8716 9760 8722 9824
rect 8406 9600 8722 9760
rect 1146 9280 1462 9281
rect 1146 9216 1152 9280
rect 1216 9216 1232 9280
rect 1296 9216 1312 9280
rect 1376 9216 1392 9280
rect 1456 9216 1462 9280
rect 1146 9215 1462 9216
rect 2466 9280 2782 9281
rect 2466 9216 2472 9280
rect 2536 9216 2552 9280
rect 2616 9216 2632 9280
rect 2696 9216 2712 9280
rect 2776 9216 2782 9280
rect 2466 9215 2782 9216
rect 3786 9280 4102 9281
rect 3786 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4102 9280
rect 3786 9215 4102 9216
rect 5106 9280 5422 9281
rect 5106 9216 5112 9280
rect 5176 9216 5192 9280
rect 5256 9216 5272 9280
rect 5336 9216 5352 9280
rect 5416 9216 5422 9280
rect 5106 9215 5422 9216
rect 6426 9280 6742 9281
rect 6426 9216 6432 9280
rect 6496 9216 6512 9280
rect 6576 9216 6592 9280
rect 6656 9216 6672 9280
rect 6736 9216 6742 9280
rect 6426 9215 6742 9216
rect 7746 9280 8062 9281
rect 7746 9216 7752 9280
rect 7816 9216 7832 9280
rect 7896 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8062 9280
rect 7746 9215 8062 9216
rect 1806 8736 2122 8737
rect 1806 8672 1812 8736
rect 1876 8672 1892 8736
rect 1956 8672 1972 8736
rect 2036 8672 2052 8736
rect 2116 8672 2122 8736
rect 1806 8671 2122 8672
rect 3126 8736 3442 8737
rect 3126 8672 3132 8736
rect 3196 8672 3212 8736
rect 3276 8672 3292 8736
rect 3356 8672 3372 8736
rect 3436 8672 3442 8736
rect 3126 8671 3442 8672
rect 4446 8736 4762 8737
rect 4446 8672 4452 8736
rect 4516 8672 4532 8736
rect 4596 8672 4612 8736
rect 4676 8672 4692 8736
rect 4756 8672 4762 8736
rect 4446 8671 4762 8672
rect 5766 8736 6082 8737
rect 5766 8672 5772 8736
rect 5836 8672 5852 8736
rect 5916 8672 5932 8736
rect 5996 8672 6012 8736
rect 6076 8672 6082 8736
rect 5766 8671 6082 8672
rect 7086 8736 7402 8737
rect 7086 8672 7092 8736
rect 7156 8672 7172 8736
rect 7236 8672 7252 8736
rect 7316 8672 7332 8736
rect 7396 8672 7402 8736
rect 7086 8671 7402 8672
rect 8406 8736 8722 8737
rect 8406 8672 8412 8736
rect 8476 8672 8492 8736
rect 8556 8672 8572 8736
rect 8636 8672 8652 8736
rect 8716 8672 8722 8736
rect 8406 8671 8722 8672
rect 1146 8192 1462 8193
rect 1146 8128 1152 8192
rect 1216 8128 1232 8192
rect 1296 8128 1312 8192
rect 1376 8128 1392 8192
rect 1456 8128 1462 8192
rect 1146 8127 1462 8128
rect 2466 8192 2782 8193
rect 2466 8128 2472 8192
rect 2536 8128 2552 8192
rect 2616 8128 2632 8192
rect 2696 8128 2712 8192
rect 2776 8128 2782 8192
rect 2466 8127 2782 8128
rect 3786 8192 4102 8193
rect 3786 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4102 8192
rect 3786 8127 4102 8128
rect 5106 8192 5422 8193
rect 5106 8128 5112 8192
rect 5176 8128 5192 8192
rect 5256 8128 5272 8192
rect 5336 8128 5352 8192
rect 5416 8128 5422 8192
rect 5106 8127 5422 8128
rect 6426 8192 6742 8193
rect 6426 8128 6432 8192
rect 6496 8128 6512 8192
rect 6576 8128 6592 8192
rect 6656 8128 6672 8192
rect 6736 8128 6742 8192
rect 6426 8127 6742 8128
rect 7746 8192 8062 8193
rect 7746 8128 7752 8192
rect 7816 8128 7832 8192
rect 7896 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8062 8192
rect 7746 8127 8062 8128
rect 1806 7648 2122 7649
rect 1806 7584 1812 7648
rect 1876 7584 1892 7648
rect 1956 7584 1972 7648
rect 2036 7584 2052 7648
rect 2116 7584 2122 7648
rect 1806 7583 2122 7584
rect 3126 7648 3442 7649
rect 3126 7584 3132 7648
rect 3196 7584 3212 7648
rect 3276 7584 3292 7648
rect 3356 7584 3372 7648
rect 3436 7584 3442 7648
rect 3126 7583 3442 7584
rect 4446 7648 4762 7649
rect 4446 7584 4452 7648
rect 4516 7584 4532 7648
rect 4596 7584 4612 7648
rect 4676 7584 4692 7648
rect 4756 7584 4762 7648
rect 4446 7583 4762 7584
rect 5766 7648 6082 7649
rect 5766 7584 5772 7648
rect 5836 7584 5852 7648
rect 5916 7584 5932 7648
rect 5996 7584 6012 7648
rect 6076 7584 6082 7648
rect 5766 7583 6082 7584
rect 7086 7648 7402 7649
rect 7086 7584 7092 7648
rect 7156 7584 7172 7648
rect 7236 7584 7252 7648
rect 7316 7584 7332 7648
rect 7396 7584 7402 7648
rect 7086 7583 7402 7584
rect 8406 7648 8722 7649
rect 8406 7584 8412 7648
rect 8476 7584 8492 7648
rect 8556 7584 8572 7648
rect 8636 7584 8652 7648
rect 8716 7584 8722 7648
rect 8406 7583 8722 7584
rect 1146 7104 1462 7105
rect 1146 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1462 7104
rect 1146 7039 1462 7040
rect 2466 7104 2782 7105
rect 2466 7040 2472 7104
rect 2536 7040 2552 7104
rect 2616 7040 2632 7104
rect 2696 7040 2712 7104
rect 2776 7040 2782 7104
rect 2466 7039 2782 7040
rect 3786 7104 4102 7105
rect 3786 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4102 7104
rect 3786 7039 4102 7040
rect 5106 7104 5422 7105
rect 5106 7040 5112 7104
rect 5176 7040 5192 7104
rect 5256 7040 5272 7104
rect 5336 7040 5352 7104
rect 5416 7040 5422 7104
rect 5106 7039 5422 7040
rect 6426 7104 6742 7105
rect 6426 7040 6432 7104
rect 6496 7040 6512 7104
rect 6576 7040 6592 7104
rect 6656 7040 6672 7104
rect 6736 7040 6742 7104
rect 6426 7039 6742 7040
rect 7746 7104 8062 7105
rect 7746 7040 7752 7104
rect 7816 7040 7832 7104
rect 7896 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8062 7104
rect 7746 7039 8062 7040
rect 1806 6560 2122 6561
rect 1806 6496 1812 6560
rect 1876 6496 1892 6560
rect 1956 6496 1972 6560
rect 2036 6496 2052 6560
rect 2116 6496 2122 6560
rect 1806 6495 2122 6496
rect 3126 6560 3442 6561
rect 3126 6496 3132 6560
rect 3196 6496 3212 6560
rect 3276 6496 3292 6560
rect 3356 6496 3372 6560
rect 3436 6496 3442 6560
rect 3126 6495 3442 6496
rect 4446 6560 4762 6561
rect 4446 6496 4452 6560
rect 4516 6496 4532 6560
rect 4596 6496 4612 6560
rect 4676 6496 4692 6560
rect 4756 6496 4762 6560
rect 4446 6495 4762 6496
rect 5766 6560 6082 6561
rect 5766 6496 5772 6560
rect 5836 6496 5852 6560
rect 5916 6496 5932 6560
rect 5996 6496 6012 6560
rect 6076 6496 6082 6560
rect 5766 6495 6082 6496
rect 7086 6560 7402 6561
rect 7086 6496 7092 6560
rect 7156 6496 7172 6560
rect 7236 6496 7252 6560
rect 7316 6496 7332 6560
rect 7396 6496 7402 6560
rect 7086 6495 7402 6496
rect 8406 6560 8722 6561
rect 8406 6496 8412 6560
rect 8476 6496 8492 6560
rect 8556 6496 8572 6560
rect 8636 6496 8652 6560
rect 8716 6496 8722 6560
rect 8406 6495 8722 6496
rect 1146 6016 1462 6017
rect 1146 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1462 6016
rect 1146 5951 1462 5952
rect 2466 6016 2782 6017
rect 2466 5952 2472 6016
rect 2536 5952 2552 6016
rect 2616 5952 2632 6016
rect 2696 5952 2712 6016
rect 2776 5952 2782 6016
rect 2466 5951 2782 5952
rect 3786 6016 4102 6017
rect 3786 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4102 6016
rect 3786 5951 4102 5952
rect 5106 6016 5422 6017
rect 5106 5952 5112 6016
rect 5176 5952 5192 6016
rect 5256 5952 5272 6016
rect 5336 5952 5352 6016
rect 5416 5952 5422 6016
rect 5106 5951 5422 5952
rect 6426 6016 6742 6017
rect 6426 5952 6432 6016
rect 6496 5952 6512 6016
rect 6576 5952 6592 6016
rect 6656 5952 6672 6016
rect 6736 5952 6742 6016
rect 6426 5951 6742 5952
rect 7746 6016 8062 6017
rect 7746 5952 7752 6016
rect 7816 5952 7832 6016
rect 7896 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8062 6016
rect 7746 5951 8062 5952
rect 1806 5472 2122 5473
rect 1806 5408 1812 5472
rect 1876 5408 1892 5472
rect 1956 5408 1972 5472
rect 2036 5408 2052 5472
rect 2116 5408 2122 5472
rect 1806 5407 2122 5408
rect 3126 5472 3442 5473
rect 3126 5408 3132 5472
rect 3196 5408 3212 5472
rect 3276 5408 3292 5472
rect 3356 5408 3372 5472
rect 3436 5408 3442 5472
rect 3126 5407 3442 5408
rect 4446 5472 4762 5473
rect 4446 5408 4452 5472
rect 4516 5408 4532 5472
rect 4596 5408 4612 5472
rect 4676 5408 4692 5472
rect 4756 5408 4762 5472
rect 4446 5407 4762 5408
rect 5766 5472 6082 5473
rect 5766 5408 5772 5472
rect 5836 5408 5852 5472
rect 5916 5408 5932 5472
rect 5996 5408 6012 5472
rect 6076 5408 6082 5472
rect 5766 5407 6082 5408
rect 7086 5472 7402 5473
rect 7086 5408 7092 5472
rect 7156 5408 7172 5472
rect 7236 5408 7252 5472
rect 7316 5408 7332 5472
rect 7396 5408 7402 5472
rect 7086 5407 7402 5408
rect 8406 5472 8722 5473
rect 8406 5408 8412 5472
rect 8476 5408 8492 5472
rect 8556 5408 8572 5472
rect 8636 5408 8652 5472
rect 8716 5408 8722 5472
rect 8406 5407 8722 5408
rect 1146 4928 1462 4929
rect 1146 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1462 4928
rect 1146 4863 1462 4864
rect 2466 4928 2782 4929
rect 2466 4864 2472 4928
rect 2536 4864 2552 4928
rect 2616 4864 2632 4928
rect 2696 4864 2712 4928
rect 2776 4864 2782 4928
rect 2466 4863 2782 4864
rect 3786 4928 4102 4929
rect 3786 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4102 4928
rect 3786 4863 4102 4864
rect 5106 4928 5422 4929
rect 5106 4864 5112 4928
rect 5176 4864 5192 4928
rect 5256 4864 5272 4928
rect 5336 4864 5352 4928
rect 5416 4864 5422 4928
rect 5106 4863 5422 4864
rect 6426 4928 6742 4929
rect 6426 4864 6432 4928
rect 6496 4864 6512 4928
rect 6576 4864 6592 4928
rect 6656 4864 6672 4928
rect 6736 4864 6742 4928
rect 6426 4863 6742 4864
rect 7746 4928 8062 4929
rect 7746 4864 7752 4928
rect 7816 4864 7832 4928
rect 7896 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8062 4928
rect 7746 4863 8062 4864
rect 1806 4384 2122 4385
rect 1806 4320 1812 4384
rect 1876 4320 1892 4384
rect 1956 4320 1972 4384
rect 2036 4320 2052 4384
rect 2116 4320 2122 4384
rect 1806 4319 2122 4320
rect 3126 4384 3442 4385
rect 3126 4320 3132 4384
rect 3196 4320 3212 4384
rect 3276 4320 3292 4384
rect 3356 4320 3372 4384
rect 3436 4320 3442 4384
rect 3126 4319 3442 4320
rect 4446 4384 4762 4385
rect 4446 4320 4452 4384
rect 4516 4320 4532 4384
rect 4596 4320 4612 4384
rect 4676 4320 4692 4384
rect 4756 4320 4762 4384
rect 4446 4319 4762 4320
rect 5766 4384 6082 4385
rect 5766 4320 5772 4384
rect 5836 4320 5852 4384
rect 5916 4320 5932 4384
rect 5996 4320 6012 4384
rect 6076 4320 6082 4384
rect 5766 4319 6082 4320
rect 7086 4384 7402 4385
rect 7086 4320 7092 4384
rect 7156 4320 7172 4384
rect 7236 4320 7252 4384
rect 7316 4320 7332 4384
rect 7396 4320 7402 4384
rect 7086 4319 7402 4320
rect 8406 4384 8722 4385
rect 8406 4320 8412 4384
rect 8476 4320 8492 4384
rect 8556 4320 8572 4384
rect 8636 4320 8652 4384
rect 8716 4320 8722 4384
rect 8406 4319 8722 4320
rect 4521 4042 4587 4045
rect 5441 4042 5507 4045
rect 4521 4040 5507 4042
rect 4521 3984 4526 4040
rect 4582 3984 5446 4040
rect 5502 3984 5507 4040
rect 4521 3982 5507 3984
rect 4521 3979 4587 3982
rect 5441 3979 5507 3982
rect 1146 3840 1462 3841
rect 1146 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1462 3840
rect 1146 3775 1462 3776
rect 2466 3840 2782 3841
rect 2466 3776 2472 3840
rect 2536 3776 2552 3840
rect 2616 3776 2632 3840
rect 2696 3776 2712 3840
rect 2776 3776 2782 3840
rect 2466 3775 2782 3776
rect 3786 3840 4102 3841
rect 3786 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4102 3840
rect 3786 3775 4102 3776
rect 5106 3840 5422 3841
rect 5106 3776 5112 3840
rect 5176 3776 5192 3840
rect 5256 3776 5272 3840
rect 5336 3776 5352 3840
rect 5416 3776 5422 3840
rect 5106 3775 5422 3776
rect 6426 3840 6742 3841
rect 6426 3776 6432 3840
rect 6496 3776 6512 3840
rect 6576 3776 6592 3840
rect 6656 3776 6672 3840
rect 6736 3776 6742 3840
rect 6426 3775 6742 3776
rect 7746 3840 8062 3841
rect 7746 3776 7752 3840
rect 7816 3776 7832 3840
rect 7896 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8062 3840
rect 7746 3775 8062 3776
rect 1806 3296 2122 3297
rect 1806 3232 1812 3296
rect 1876 3232 1892 3296
rect 1956 3232 1972 3296
rect 2036 3232 2052 3296
rect 2116 3232 2122 3296
rect 1806 3231 2122 3232
rect 3126 3296 3442 3297
rect 3126 3232 3132 3296
rect 3196 3232 3212 3296
rect 3276 3232 3292 3296
rect 3356 3232 3372 3296
rect 3436 3232 3442 3296
rect 3126 3231 3442 3232
rect 4446 3296 4762 3297
rect 4446 3232 4452 3296
rect 4516 3232 4532 3296
rect 4596 3232 4612 3296
rect 4676 3232 4692 3296
rect 4756 3232 4762 3296
rect 4446 3231 4762 3232
rect 5766 3296 6082 3297
rect 5766 3232 5772 3296
rect 5836 3232 5852 3296
rect 5916 3232 5932 3296
rect 5996 3232 6012 3296
rect 6076 3232 6082 3296
rect 5766 3231 6082 3232
rect 7086 3296 7402 3297
rect 7086 3232 7092 3296
rect 7156 3232 7172 3296
rect 7236 3232 7252 3296
rect 7316 3232 7332 3296
rect 7396 3232 7402 3296
rect 7086 3231 7402 3232
rect 8406 3296 8722 3297
rect 8406 3232 8412 3296
rect 8476 3232 8492 3296
rect 8556 3232 8572 3296
rect 8636 3232 8652 3296
rect 8716 3232 8722 3296
rect 8406 3231 8722 3232
rect 1142 2753 1458 2770
rect 2462 2753 2778 2768
rect 3782 2753 4098 2766
rect 5104 2753 5420 2768
rect 6412 2753 6728 2782
rect 7754 2753 8070 2782
rect 1142 2752 1462 2753
rect 1142 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1462 2752
rect 1142 2687 1462 2688
rect 2462 2752 2782 2753
rect 2462 2688 2472 2752
rect 2536 2688 2552 2752
rect 2616 2688 2632 2752
rect 2696 2688 2712 2752
rect 2776 2688 2782 2752
rect 2462 2687 2782 2688
rect 3782 2752 4102 2753
rect 3782 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4102 2752
rect 3782 2687 4102 2688
rect 5104 2752 5422 2753
rect 5104 2688 5112 2752
rect 5176 2688 5192 2752
rect 5256 2688 5272 2752
rect 5336 2688 5352 2752
rect 5416 2688 5422 2752
rect 5104 2687 5422 2688
rect 6412 2752 6742 2753
rect 6412 2688 6432 2752
rect 6496 2688 6512 2752
rect 6576 2688 6592 2752
rect 6656 2688 6672 2752
rect 6736 2688 6742 2752
rect 6412 2687 6742 2688
rect 7746 2752 8070 2753
rect 7746 2688 7752 2752
rect 7816 2688 7832 2752
rect 7896 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8070 2752
rect 7746 2687 8070 2688
rect 1142 2066 1458 2687
rect 1806 2208 2122 2209
rect 1806 2144 1812 2208
rect 1876 2144 1892 2208
rect 1956 2144 1972 2208
rect 2036 2144 2052 2208
rect 2116 2144 2122 2208
rect 1806 2143 2122 2144
rect 2462 2066 2778 2687
rect 3126 2208 3442 2209
rect 3126 2144 3132 2208
rect 3196 2144 3212 2208
rect 3276 2144 3292 2208
rect 3356 2144 3372 2208
rect 3436 2144 3442 2208
rect 3126 2143 3442 2144
rect 3782 2066 4098 2687
rect 4446 2208 4762 2209
rect 4446 2144 4452 2208
rect 4516 2144 4532 2208
rect 4596 2144 4612 2208
rect 4676 2144 4692 2208
rect 4756 2144 4762 2208
rect 4446 2143 4762 2144
rect 5104 2066 5420 2687
rect 5766 2208 6082 2209
rect 5766 2144 5772 2208
rect 5836 2144 5852 2208
rect 5916 2144 5932 2208
rect 5996 2144 6012 2208
rect 6076 2144 6082 2208
rect 5766 2143 6082 2144
rect 6412 2066 6728 2687
rect 7086 2208 7402 2209
rect 7086 2144 7092 2208
rect 7156 2144 7172 2208
rect 7236 2144 7252 2208
rect 7316 2144 7332 2208
rect 7396 2144 7402 2208
rect 7086 2143 7402 2144
rect 7754 2066 8070 2687
rect 8406 2208 8722 2209
rect 8406 2144 8412 2208
rect 8476 2144 8492 2208
rect 8556 2144 8572 2208
rect 8636 2144 8652 2208
rect 8716 2144 8722 2208
rect 8406 2143 8722 2144
rect 1134 2018 8070 2066
rect 1134 1820 1358 2018
rect 7744 1820 8070 2018
rect 1134 1750 8070 1820
<< via3 >>
rect 2136 10006 8522 10204
rect 1812 9820 1876 9824
rect 1812 9764 1816 9820
rect 1816 9764 1872 9820
rect 1872 9764 1876 9820
rect 1812 9760 1876 9764
rect 1892 9820 1956 9824
rect 1892 9764 1896 9820
rect 1896 9764 1952 9820
rect 1952 9764 1956 9820
rect 1892 9760 1956 9764
rect 1972 9820 2036 9824
rect 1972 9764 1976 9820
rect 1976 9764 2032 9820
rect 2032 9764 2036 9820
rect 1972 9760 2036 9764
rect 2052 9820 2116 9824
rect 2052 9764 2056 9820
rect 2056 9764 2112 9820
rect 2112 9764 2116 9820
rect 2052 9760 2116 9764
rect 3132 9820 3196 9824
rect 3132 9764 3136 9820
rect 3136 9764 3192 9820
rect 3192 9764 3196 9820
rect 3132 9760 3196 9764
rect 3212 9820 3276 9824
rect 3212 9764 3216 9820
rect 3216 9764 3272 9820
rect 3272 9764 3276 9820
rect 3212 9760 3276 9764
rect 3292 9820 3356 9824
rect 3292 9764 3296 9820
rect 3296 9764 3352 9820
rect 3352 9764 3356 9820
rect 3292 9760 3356 9764
rect 3372 9820 3436 9824
rect 3372 9764 3376 9820
rect 3376 9764 3432 9820
rect 3432 9764 3436 9820
rect 3372 9760 3436 9764
rect 4452 9820 4516 9824
rect 4452 9764 4456 9820
rect 4456 9764 4512 9820
rect 4512 9764 4516 9820
rect 4452 9760 4516 9764
rect 4532 9820 4596 9824
rect 4532 9764 4536 9820
rect 4536 9764 4592 9820
rect 4592 9764 4596 9820
rect 4532 9760 4596 9764
rect 4612 9820 4676 9824
rect 4612 9764 4616 9820
rect 4616 9764 4672 9820
rect 4672 9764 4676 9820
rect 4612 9760 4676 9764
rect 4692 9820 4756 9824
rect 4692 9764 4696 9820
rect 4696 9764 4752 9820
rect 4752 9764 4756 9820
rect 4692 9760 4756 9764
rect 5772 9820 5836 9824
rect 5772 9764 5776 9820
rect 5776 9764 5832 9820
rect 5832 9764 5836 9820
rect 5772 9760 5836 9764
rect 5852 9820 5916 9824
rect 5852 9764 5856 9820
rect 5856 9764 5912 9820
rect 5912 9764 5916 9820
rect 5852 9760 5916 9764
rect 5932 9820 5996 9824
rect 5932 9764 5936 9820
rect 5936 9764 5992 9820
rect 5992 9764 5996 9820
rect 5932 9760 5996 9764
rect 6012 9820 6076 9824
rect 6012 9764 6016 9820
rect 6016 9764 6072 9820
rect 6072 9764 6076 9820
rect 6012 9760 6076 9764
rect 7092 9820 7156 9824
rect 7092 9764 7096 9820
rect 7096 9764 7152 9820
rect 7152 9764 7156 9820
rect 7092 9760 7156 9764
rect 7172 9820 7236 9824
rect 7172 9764 7176 9820
rect 7176 9764 7232 9820
rect 7232 9764 7236 9820
rect 7172 9760 7236 9764
rect 7252 9820 7316 9824
rect 7252 9764 7256 9820
rect 7256 9764 7312 9820
rect 7312 9764 7316 9820
rect 7252 9760 7316 9764
rect 7332 9820 7396 9824
rect 7332 9764 7336 9820
rect 7336 9764 7392 9820
rect 7392 9764 7396 9820
rect 7332 9760 7396 9764
rect 8412 9820 8476 9824
rect 8412 9764 8416 9820
rect 8416 9764 8472 9820
rect 8472 9764 8476 9820
rect 8412 9760 8476 9764
rect 8492 9820 8556 9824
rect 8492 9764 8496 9820
rect 8496 9764 8552 9820
rect 8552 9764 8556 9820
rect 8492 9760 8556 9764
rect 8572 9820 8636 9824
rect 8572 9764 8576 9820
rect 8576 9764 8632 9820
rect 8632 9764 8636 9820
rect 8572 9760 8636 9764
rect 8652 9820 8716 9824
rect 8652 9764 8656 9820
rect 8656 9764 8712 9820
rect 8712 9764 8716 9820
rect 8652 9760 8716 9764
rect 1152 9276 1216 9280
rect 1152 9220 1156 9276
rect 1156 9220 1212 9276
rect 1212 9220 1216 9276
rect 1152 9216 1216 9220
rect 1232 9276 1296 9280
rect 1232 9220 1236 9276
rect 1236 9220 1292 9276
rect 1292 9220 1296 9276
rect 1232 9216 1296 9220
rect 1312 9276 1376 9280
rect 1312 9220 1316 9276
rect 1316 9220 1372 9276
rect 1372 9220 1376 9276
rect 1312 9216 1376 9220
rect 1392 9276 1456 9280
rect 1392 9220 1396 9276
rect 1396 9220 1452 9276
rect 1452 9220 1456 9276
rect 1392 9216 1456 9220
rect 2472 9276 2536 9280
rect 2472 9220 2476 9276
rect 2476 9220 2532 9276
rect 2532 9220 2536 9276
rect 2472 9216 2536 9220
rect 2552 9276 2616 9280
rect 2552 9220 2556 9276
rect 2556 9220 2612 9276
rect 2612 9220 2616 9276
rect 2552 9216 2616 9220
rect 2632 9276 2696 9280
rect 2632 9220 2636 9276
rect 2636 9220 2692 9276
rect 2692 9220 2696 9276
rect 2632 9216 2696 9220
rect 2712 9276 2776 9280
rect 2712 9220 2716 9276
rect 2716 9220 2772 9276
rect 2772 9220 2776 9276
rect 2712 9216 2776 9220
rect 3792 9276 3856 9280
rect 3792 9220 3796 9276
rect 3796 9220 3852 9276
rect 3852 9220 3856 9276
rect 3792 9216 3856 9220
rect 3872 9276 3936 9280
rect 3872 9220 3876 9276
rect 3876 9220 3932 9276
rect 3932 9220 3936 9276
rect 3872 9216 3936 9220
rect 3952 9276 4016 9280
rect 3952 9220 3956 9276
rect 3956 9220 4012 9276
rect 4012 9220 4016 9276
rect 3952 9216 4016 9220
rect 4032 9276 4096 9280
rect 4032 9220 4036 9276
rect 4036 9220 4092 9276
rect 4092 9220 4096 9276
rect 4032 9216 4096 9220
rect 5112 9276 5176 9280
rect 5112 9220 5116 9276
rect 5116 9220 5172 9276
rect 5172 9220 5176 9276
rect 5112 9216 5176 9220
rect 5192 9276 5256 9280
rect 5192 9220 5196 9276
rect 5196 9220 5252 9276
rect 5252 9220 5256 9276
rect 5192 9216 5256 9220
rect 5272 9276 5336 9280
rect 5272 9220 5276 9276
rect 5276 9220 5332 9276
rect 5332 9220 5336 9276
rect 5272 9216 5336 9220
rect 5352 9276 5416 9280
rect 5352 9220 5356 9276
rect 5356 9220 5412 9276
rect 5412 9220 5416 9276
rect 5352 9216 5416 9220
rect 6432 9276 6496 9280
rect 6432 9220 6436 9276
rect 6436 9220 6492 9276
rect 6492 9220 6496 9276
rect 6432 9216 6496 9220
rect 6512 9276 6576 9280
rect 6512 9220 6516 9276
rect 6516 9220 6572 9276
rect 6572 9220 6576 9276
rect 6512 9216 6576 9220
rect 6592 9276 6656 9280
rect 6592 9220 6596 9276
rect 6596 9220 6652 9276
rect 6652 9220 6656 9276
rect 6592 9216 6656 9220
rect 6672 9276 6736 9280
rect 6672 9220 6676 9276
rect 6676 9220 6732 9276
rect 6732 9220 6736 9276
rect 6672 9216 6736 9220
rect 7752 9276 7816 9280
rect 7752 9220 7756 9276
rect 7756 9220 7812 9276
rect 7812 9220 7816 9276
rect 7752 9216 7816 9220
rect 7832 9276 7896 9280
rect 7832 9220 7836 9276
rect 7836 9220 7892 9276
rect 7892 9220 7896 9276
rect 7832 9216 7896 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 1812 8732 1876 8736
rect 1812 8676 1816 8732
rect 1816 8676 1872 8732
rect 1872 8676 1876 8732
rect 1812 8672 1876 8676
rect 1892 8732 1956 8736
rect 1892 8676 1896 8732
rect 1896 8676 1952 8732
rect 1952 8676 1956 8732
rect 1892 8672 1956 8676
rect 1972 8732 2036 8736
rect 1972 8676 1976 8732
rect 1976 8676 2032 8732
rect 2032 8676 2036 8732
rect 1972 8672 2036 8676
rect 2052 8732 2116 8736
rect 2052 8676 2056 8732
rect 2056 8676 2112 8732
rect 2112 8676 2116 8732
rect 2052 8672 2116 8676
rect 3132 8732 3196 8736
rect 3132 8676 3136 8732
rect 3136 8676 3192 8732
rect 3192 8676 3196 8732
rect 3132 8672 3196 8676
rect 3212 8732 3276 8736
rect 3212 8676 3216 8732
rect 3216 8676 3272 8732
rect 3272 8676 3276 8732
rect 3212 8672 3276 8676
rect 3292 8732 3356 8736
rect 3292 8676 3296 8732
rect 3296 8676 3352 8732
rect 3352 8676 3356 8732
rect 3292 8672 3356 8676
rect 3372 8732 3436 8736
rect 3372 8676 3376 8732
rect 3376 8676 3432 8732
rect 3432 8676 3436 8732
rect 3372 8672 3436 8676
rect 4452 8732 4516 8736
rect 4452 8676 4456 8732
rect 4456 8676 4512 8732
rect 4512 8676 4516 8732
rect 4452 8672 4516 8676
rect 4532 8732 4596 8736
rect 4532 8676 4536 8732
rect 4536 8676 4592 8732
rect 4592 8676 4596 8732
rect 4532 8672 4596 8676
rect 4612 8732 4676 8736
rect 4612 8676 4616 8732
rect 4616 8676 4672 8732
rect 4672 8676 4676 8732
rect 4612 8672 4676 8676
rect 4692 8732 4756 8736
rect 4692 8676 4696 8732
rect 4696 8676 4752 8732
rect 4752 8676 4756 8732
rect 4692 8672 4756 8676
rect 5772 8732 5836 8736
rect 5772 8676 5776 8732
rect 5776 8676 5832 8732
rect 5832 8676 5836 8732
rect 5772 8672 5836 8676
rect 5852 8732 5916 8736
rect 5852 8676 5856 8732
rect 5856 8676 5912 8732
rect 5912 8676 5916 8732
rect 5852 8672 5916 8676
rect 5932 8732 5996 8736
rect 5932 8676 5936 8732
rect 5936 8676 5992 8732
rect 5992 8676 5996 8732
rect 5932 8672 5996 8676
rect 6012 8732 6076 8736
rect 6012 8676 6016 8732
rect 6016 8676 6072 8732
rect 6072 8676 6076 8732
rect 6012 8672 6076 8676
rect 7092 8732 7156 8736
rect 7092 8676 7096 8732
rect 7096 8676 7152 8732
rect 7152 8676 7156 8732
rect 7092 8672 7156 8676
rect 7172 8732 7236 8736
rect 7172 8676 7176 8732
rect 7176 8676 7232 8732
rect 7232 8676 7236 8732
rect 7172 8672 7236 8676
rect 7252 8732 7316 8736
rect 7252 8676 7256 8732
rect 7256 8676 7312 8732
rect 7312 8676 7316 8732
rect 7252 8672 7316 8676
rect 7332 8732 7396 8736
rect 7332 8676 7336 8732
rect 7336 8676 7392 8732
rect 7392 8676 7396 8732
rect 7332 8672 7396 8676
rect 8412 8732 8476 8736
rect 8412 8676 8416 8732
rect 8416 8676 8472 8732
rect 8472 8676 8476 8732
rect 8412 8672 8476 8676
rect 8492 8732 8556 8736
rect 8492 8676 8496 8732
rect 8496 8676 8552 8732
rect 8552 8676 8556 8732
rect 8492 8672 8556 8676
rect 8572 8732 8636 8736
rect 8572 8676 8576 8732
rect 8576 8676 8632 8732
rect 8632 8676 8636 8732
rect 8572 8672 8636 8676
rect 8652 8732 8716 8736
rect 8652 8676 8656 8732
rect 8656 8676 8712 8732
rect 8712 8676 8716 8732
rect 8652 8672 8716 8676
rect 1152 8188 1216 8192
rect 1152 8132 1156 8188
rect 1156 8132 1212 8188
rect 1212 8132 1216 8188
rect 1152 8128 1216 8132
rect 1232 8188 1296 8192
rect 1232 8132 1236 8188
rect 1236 8132 1292 8188
rect 1292 8132 1296 8188
rect 1232 8128 1296 8132
rect 1312 8188 1376 8192
rect 1312 8132 1316 8188
rect 1316 8132 1372 8188
rect 1372 8132 1376 8188
rect 1312 8128 1376 8132
rect 1392 8188 1456 8192
rect 1392 8132 1396 8188
rect 1396 8132 1452 8188
rect 1452 8132 1456 8188
rect 1392 8128 1456 8132
rect 2472 8188 2536 8192
rect 2472 8132 2476 8188
rect 2476 8132 2532 8188
rect 2532 8132 2536 8188
rect 2472 8128 2536 8132
rect 2552 8188 2616 8192
rect 2552 8132 2556 8188
rect 2556 8132 2612 8188
rect 2612 8132 2616 8188
rect 2552 8128 2616 8132
rect 2632 8188 2696 8192
rect 2632 8132 2636 8188
rect 2636 8132 2692 8188
rect 2692 8132 2696 8188
rect 2632 8128 2696 8132
rect 2712 8188 2776 8192
rect 2712 8132 2716 8188
rect 2716 8132 2772 8188
rect 2772 8132 2776 8188
rect 2712 8128 2776 8132
rect 3792 8188 3856 8192
rect 3792 8132 3796 8188
rect 3796 8132 3852 8188
rect 3852 8132 3856 8188
rect 3792 8128 3856 8132
rect 3872 8188 3936 8192
rect 3872 8132 3876 8188
rect 3876 8132 3932 8188
rect 3932 8132 3936 8188
rect 3872 8128 3936 8132
rect 3952 8188 4016 8192
rect 3952 8132 3956 8188
rect 3956 8132 4012 8188
rect 4012 8132 4016 8188
rect 3952 8128 4016 8132
rect 4032 8188 4096 8192
rect 4032 8132 4036 8188
rect 4036 8132 4092 8188
rect 4092 8132 4096 8188
rect 4032 8128 4096 8132
rect 5112 8188 5176 8192
rect 5112 8132 5116 8188
rect 5116 8132 5172 8188
rect 5172 8132 5176 8188
rect 5112 8128 5176 8132
rect 5192 8188 5256 8192
rect 5192 8132 5196 8188
rect 5196 8132 5252 8188
rect 5252 8132 5256 8188
rect 5192 8128 5256 8132
rect 5272 8188 5336 8192
rect 5272 8132 5276 8188
rect 5276 8132 5332 8188
rect 5332 8132 5336 8188
rect 5272 8128 5336 8132
rect 5352 8188 5416 8192
rect 5352 8132 5356 8188
rect 5356 8132 5412 8188
rect 5412 8132 5416 8188
rect 5352 8128 5416 8132
rect 6432 8188 6496 8192
rect 6432 8132 6436 8188
rect 6436 8132 6492 8188
rect 6492 8132 6496 8188
rect 6432 8128 6496 8132
rect 6512 8188 6576 8192
rect 6512 8132 6516 8188
rect 6516 8132 6572 8188
rect 6572 8132 6576 8188
rect 6512 8128 6576 8132
rect 6592 8188 6656 8192
rect 6592 8132 6596 8188
rect 6596 8132 6652 8188
rect 6652 8132 6656 8188
rect 6592 8128 6656 8132
rect 6672 8188 6736 8192
rect 6672 8132 6676 8188
rect 6676 8132 6732 8188
rect 6732 8132 6736 8188
rect 6672 8128 6736 8132
rect 7752 8188 7816 8192
rect 7752 8132 7756 8188
rect 7756 8132 7812 8188
rect 7812 8132 7816 8188
rect 7752 8128 7816 8132
rect 7832 8188 7896 8192
rect 7832 8132 7836 8188
rect 7836 8132 7892 8188
rect 7892 8132 7896 8188
rect 7832 8128 7896 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 1812 7644 1876 7648
rect 1812 7588 1816 7644
rect 1816 7588 1872 7644
rect 1872 7588 1876 7644
rect 1812 7584 1876 7588
rect 1892 7644 1956 7648
rect 1892 7588 1896 7644
rect 1896 7588 1952 7644
rect 1952 7588 1956 7644
rect 1892 7584 1956 7588
rect 1972 7644 2036 7648
rect 1972 7588 1976 7644
rect 1976 7588 2032 7644
rect 2032 7588 2036 7644
rect 1972 7584 2036 7588
rect 2052 7644 2116 7648
rect 2052 7588 2056 7644
rect 2056 7588 2112 7644
rect 2112 7588 2116 7644
rect 2052 7584 2116 7588
rect 3132 7644 3196 7648
rect 3132 7588 3136 7644
rect 3136 7588 3192 7644
rect 3192 7588 3196 7644
rect 3132 7584 3196 7588
rect 3212 7644 3276 7648
rect 3212 7588 3216 7644
rect 3216 7588 3272 7644
rect 3272 7588 3276 7644
rect 3212 7584 3276 7588
rect 3292 7644 3356 7648
rect 3292 7588 3296 7644
rect 3296 7588 3352 7644
rect 3352 7588 3356 7644
rect 3292 7584 3356 7588
rect 3372 7644 3436 7648
rect 3372 7588 3376 7644
rect 3376 7588 3432 7644
rect 3432 7588 3436 7644
rect 3372 7584 3436 7588
rect 4452 7644 4516 7648
rect 4452 7588 4456 7644
rect 4456 7588 4512 7644
rect 4512 7588 4516 7644
rect 4452 7584 4516 7588
rect 4532 7644 4596 7648
rect 4532 7588 4536 7644
rect 4536 7588 4592 7644
rect 4592 7588 4596 7644
rect 4532 7584 4596 7588
rect 4612 7644 4676 7648
rect 4612 7588 4616 7644
rect 4616 7588 4672 7644
rect 4672 7588 4676 7644
rect 4612 7584 4676 7588
rect 4692 7644 4756 7648
rect 4692 7588 4696 7644
rect 4696 7588 4752 7644
rect 4752 7588 4756 7644
rect 4692 7584 4756 7588
rect 5772 7644 5836 7648
rect 5772 7588 5776 7644
rect 5776 7588 5832 7644
rect 5832 7588 5836 7644
rect 5772 7584 5836 7588
rect 5852 7644 5916 7648
rect 5852 7588 5856 7644
rect 5856 7588 5912 7644
rect 5912 7588 5916 7644
rect 5852 7584 5916 7588
rect 5932 7644 5996 7648
rect 5932 7588 5936 7644
rect 5936 7588 5992 7644
rect 5992 7588 5996 7644
rect 5932 7584 5996 7588
rect 6012 7644 6076 7648
rect 6012 7588 6016 7644
rect 6016 7588 6072 7644
rect 6072 7588 6076 7644
rect 6012 7584 6076 7588
rect 7092 7644 7156 7648
rect 7092 7588 7096 7644
rect 7096 7588 7152 7644
rect 7152 7588 7156 7644
rect 7092 7584 7156 7588
rect 7172 7644 7236 7648
rect 7172 7588 7176 7644
rect 7176 7588 7232 7644
rect 7232 7588 7236 7644
rect 7172 7584 7236 7588
rect 7252 7644 7316 7648
rect 7252 7588 7256 7644
rect 7256 7588 7312 7644
rect 7312 7588 7316 7644
rect 7252 7584 7316 7588
rect 7332 7644 7396 7648
rect 7332 7588 7336 7644
rect 7336 7588 7392 7644
rect 7392 7588 7396 7644
rect 7332 7584 7396 7588
rect 8412 7644 8476 7648
rect 8412 7588 8416 7644
rect 8416 7588 8472 7644
rect 8472 7588 8476 7644
rect 8412 7584 8476 7588
rect 8492 7644 8556 7648
rect 8492 7588 8496 7644
rect 8496 7588 8552 7644
rect 8552 7588 8556 7644
rect 8492 7584 8556 7588
rect 8572 7644 8636 7648
rect 8572 7588 8576 7644
rect 8576 7588 8632 7644
rect 8632 7588 8636 7644
rect 8572 7584 8636 7588
rect 8652 7644 8716 7648
rect 8652 7588 8656 7644
rect 8656 7588 8712 7644
rect 8712 7588 8716 7644
rect 8652 7584 8716 7588
rect 1152 7100 1216 7104
rect 1152 7044 1156 7100
rect 1156 7044 1212 7100
rect 1212 7044 1216 7100
rect 1152 7040 1216 7044
rect 1232 7100 1296 7104
rect 1232 7044 1236 7100
rect 1236 7044 1292 7100
rect 1292 7044 1296 7100
rect 1232 7040 1296 7044
rect 1312 7100 1376 7104
rect 1312 7044 1316 7100
rect 1316 7044 1372 7100
rect 1372 7044 1376 7100
rect 1312 7040 1376 7044
rect 1392 7100 1456 7104
rect 1392 7044 1396 7100
rect 1396 7044 1452 7100
rect 1452 7044 1456 7100
rect 1392 7040 1456 7044
rect 2472 7100 2536 7104
rect 2472 7044 2476 7100
rect 2476 7044 2532 7100
rect 2532 7044 2536 7100
rect 2472 7040 2536 7044
rect 2552 7100 2616 7104
rect 2552 7044 2556 7100
rect 2556 7044 2612 7100
rect 2612 7044 2616 7100
rect 2552 7040 2616 7044
rect 2632 7100 2696 7104
rect 2632 7044 2636 7100
rect 2636 7044 2692 7100
rect 2692 7044 2696 7100
rect 2632 7040 2696 7044
rect 2712 7100 2776 7104
rect 2712 7044 2716 7100
rect 2716 7044 2772 7100
rect 2772 7044 2776 7100
rect 2712 7040 2776 7044
rect 3792 7100 3856 7104
rect 3792 7044 3796 7100
rect 3796 7044 3852 7100
rect 3852 7044 3856 7100
rect 3792 7040 3856 7044
rect 3872 7100 3936 7104
rect 3872 7044 3876 7100
rect 3876 7044 3932 7100
rect 3932 7044 3936 7100
rect 3872 7040 3936 7044
rect 3952 7100 4016 7104
rect 3952 7044 3956 7100
rect 3956 7044 4012 7100
rect 4012 7044 4016 7100
rect 3952 7040 4016 7044
rect 4032 7100 4096 7104
rect 4032 7044 4036 7100
rect 4036 7044 4092 7100
rect 4092 7044 4096 7100
rect 4032 7040 4096 7044
rect 5112 7100 5176 7104
rect 5112 7044 5116 7100
rect 5116 7044 5172 7100
rect 5172 7044 5176 7100
rect 5112 7040 5176 7044
rect 5192 7100 5256 7104
rect 5192 7044 5196 7100
rect 5196 7044 5252 7100
rect 5252 7044 5256 7100
rect 5192 7040 5256 7044
rect 5272 7100 5336 7104
rect 5272 7044 5276 7100
rect 5276 7044 5332 7100
rect 5332 7044 5336 7100
rect 5272 7040 5336 7044
rect 5352 7100 5416 7104
rect 5352 7044 5356 7100
rect 5356 7044 5412 7100
rect 5412 7044 5416 7100
rect 5352 7040 5416 7044
rect 6432 7100 6496 7104
rect 6432 7044 6436 7100
rect 6436 7044 6492 7100
rect 6492 7044 6496 7100
rect 6432 7040 6496 7044
rect 6512 7100 6576 7104
rect 6512 7044 6516 7100
rect 6516 7044 6572 7100
rect 6572 7044 6576 7100
rect 6512 7040 6576 7044
rect 6592 7100 6656 7104
rect 6592 7044 6596 7100
rect 6596 7044 6652 7100
rect 6652 7044 6656 7100
rect 6592 7040 6656 7044
rect 6672 7100 6736 7104
rect 6672 7044 6676 7100
rect 6676 7044 6732 7100
rect 6732 7044 6736 7100
rect 6672 7040 6736 7044
rect 7752 7100 7816 7104
rect 7752 7044 7756 7100
rect 7756 7044 7812 7100
rect 7812 7044 7816 7100
rect 7752 7040 7816 7044
rect 7832 7100 7896 7104
rect 7832 7044 7836 7100
rect 7836 7044 7892 7100
rect 7892 7044 7896 7100
rect 7832 7040 7896 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 1812 6556 1876 6560
rect 1812 6500 1816 6556
rect 1816 6500 1872 6556
rect 1872 6500 1876 6556
rect 1812 6496 1876 6500
rect 1892 6556 1956 6560
rect 1892 6500 1896 6556
rect 1896 6500 1952 6556
rect 1952 6500 1956 6556
rect 1892 6496 1956 6500
rect 1972 6556 2036 6560
rect 1972 6500 1976 6556
rect 1976 6500 2032 6556
rect 2032 6500 2036 6556
rect 1972 6496 2036 6500
rect 2052 6556 2116 6560
rect 2052 6500 2056 6556
rect 2056 6500 2112 6556
rect 2112 6500 2116 6556
rect 2052 6496 2116 6500
rect 3132 6556 3196 6560
rect 3132 6500 3136 6556
rect 3136 6500 3192 6556
rect 3192 6500 3196 6556
rect 3132 6496 3196 6500
rect 3212 6556 3276 6560
rect 3212 6500 3216 6556
rect 3216 6500 3272 6556
rect 3272 6500 3276 6556
rect 3212 6496 3276 6500
rect 3292 6556 3356 6560
rect 3292 6500 3296 6556
rect 3296 6500 3352 6556
rect 3352 6500 3356 6556
rect 3292 6496 3356 6500
rect 3372 6556 3436 6560
rect 3372 6500 3376 6556
rect 3376 6500 3432 6556
rect 3432 6500 3436 6556
rect 3372 6496 3436 6500
rect 4452 6556 4516 6560
rect 4452 6500 4456 6556
rect 4456 6500 4512 6556
rect 4512 6500 4516 6556
rect 4452 6496 4516 6500
rect 4532 6556 4596 6560
rect 4532 6500 4536 6556
rect 4536 6500 4592 6556
rect 4592 6500 4596 6556
rect 4532 6496 4596 6500
rect 4612 6556 4676 6560
rect 4612 6500 4616 6556
rect 4616 6500 4672 6556
rect 4672 6500 4676 6556
rect 4612 6496 4676 6500
rect 4692 6556 4756 6560
rect 4692 6500 4696 6556
rect 4696 6500 4752 6556
rect 4752 6500 4756 6556
rect 4692 6496 4756 6500
rect 5772 6556 5836 6560
rect 5772 6500 5776 6556
rect 5776 6500 5832 6556
rect 5832 6500 5836 6556
rect 5772 6496 5836 6500
rect 5852 6556 5916 6560
rect 5852 6500 5856 6556
rect 5856 6500 5912 6556
rect 5912 6500 5916 6556
rect 5852 6496 5916 6500
rect 5932 6556 5996 6560
rect 5932 6500 5936 6556
rect 5936 6500 5992 6556
rect 5992 6500 5996 6556
rect 5932 6496 5996 6500
rect 6012 6556 6076 6560
rect 6012 6500 6016 6556
rect 6016 6500 6072 6556
rect 6072 6500 6076 6556
rect 6012 6496 6076 6500
rect 7092 6556 7156 6560
rect 7092 6500 7096 6556
rect 7096 6500 7152 6556
rect 7152 6500 7156 6556
rect 7092 6496 7156 6500
rect 7172 6556 7236 6560
rect 7172 6500 7176 6556
rect 7176 6500 7232 6556
rect 7232 6500 7236 6556
rect 7172 6496 7236 6500
rect 7252 6556 7316 6560
rect 7252 6500 7256 6556
rect 7256 6500 7312 6556
rect 7312 6500 7316 6556
rect 7252 6496 7316 6500
rect 7332 6556 7396 6560
rect 7332 6500 7336 6556
rect 7336 6500 7392 6556
rect 7392 6500 7396 6556
rect 7332 6496 7396 6500
rect 8412 6556 8476 6560
rect 8412 6500 8416 6556
rect 8416 6500 8472 6556
rect 8472 6500 8476 6556
rect 8412 6496 8476 6500
rect 8492 6556 8556 6560
rect 8492 6500 8496 6556
rect 8496 6500 8552 6556
rect 8552 6500 8556 6556
rect 8492 6496 8556 6500
rect 8572 6556 8636 6560
rect 8572 6500 8576 6556
rect 8576 6500 8632 6556
rect 8632 6500 8636 6556
rect 8572 6496 8636 6500
rect 8652 6556 8716 6560
rect 8652 6500 8656 6556
rect 8656 6500 8712 6556
rect 8712 6500 8716 6556
rect 8652 6496 8716 6500
rect 1152 6012 1216 6016
rect 1152 5956 1156 6012
rect 1156 5956 1212 6012
rect 1212 5956 1216 6012
rect 1152 5952 1216 5956
rect 1232 6012 1296 6016
rect 1232 5956 1236 6012
rect 1236 5956 1292 6012
rect 1292 5956 1296 6012
rect 1232 5952 1296 5956
rect 1312 6012 1376 6016
rect 1312 5956 1316 6012
rect 1316 5956 1372 6012
rect 1372 5956 1376 6012
rect 1312 5952 1376 5956
rect 1392 6012 1456 6016
rect 1392 5956 1396 6012
rect 1396 5956 1452 6012
rect 1452 5956 1456 6012
rect 1392 5952 1456 5956
rect 2472 6012 2536 6016
rect 2472 5956 2476 6012
rect 2476 5956 2532 6012
rect 2532 5956 2536 6012
rect 2472 5952 2536 5956
rect 2552 6012 2616 6016
rect 2552 5956 2556 6012
rect 2556 5956 2612 6012
rect 2612 5956 2616 6012
rect 2552 5952 2616 5956
rect 2632 6012 2696 6016
rect 2632 5956 2636 6012
rect 2636 5956 2692 6012
rect 2692 5956 2696 6012
rect 2632 5952 2696 5956
rect 2712 6012 2776 6016
rect 2712 5956 2716 6012
rect 2716 5956 2772 6012
rect 2772 5956 2776 6012
rect 2712 5952 2776 5956
rect 3792 6012 3856 6016
rect 3792 5956 3796 6012
rect 3796 5956 3852 6012
rect 3852 5956 3856 6012
rect 3792 5952 3856 5956
rect 3872 6012 3936 6016
rect 3872 5956 3876 6012
rect 3876 5956 3932 6012
rect 3932 5956 3936 6012
rect 3872 5952 3936 5956
rect 3952 6012 4016 6016
rect 3952 5956 3956 6012
rect 3956 5956 4012 6012
rect 4012 5956 4016 6012
rect 3952 5952 4016 5956
rect 4032 6012 4096 6016
rect 4032 5956 4036 6012
rect 4036 5956 4092 6012
rect 4092 5956 4096 6012
rect 4032 5952 4096 5956
rect 5112 6012 5176 6016
rect 5112 5956 5116 6012
rect 5116 5956 5172 6012
rect 5172 5956 5176 6012
rect 5112 5952 5176 5956
rect 5192 6012 5256 6016
rect 5192 5956 5196 6012
rect 5196 5956 5252 6012
rect 5252 5956 5256 6012
rect 5192 5952 5256 5956
rect 5272 6012 5336 6016
rect 5272 5956 5276 6012
rect 5276 5956 5332 6012
rect 5332 5956 5336 6012
rect 5272 5952 5336 5956
rect 5352 6012 5416 6016
rect 5352 5956 5356 6012
rect 5356 5956 5412 6012
rect 5412 5956 5416 6012
rect 5352 5952 5416 5956
rect 6432 6012 6496 6016
rect 6432 5956 6436 6012
rect 6436 5956 6492 6012
rect 6492 5956 6496 6012
rect 6432 5952 6496 5956
rect 6512 6012 6576 6016
rect 6512 5956 6516 6012
rect 6516 5956 6572 6012
rect 6572 5956 6576 6012
rect 6512 5952 6576 5956
rect 6592 6012 6656 6016
rect 6592 5956 6596 6012
rect 6596 5956 6652 6012
rect 6652 5956 6656 6012
rect 6592 5952 6656 5956
rect 6672 6012 6736 6016
rect 6672 5956 6676 6012
rect 6676 5956 6732 6012
rect 6732 5956 6736 6012
rect 6672 5952 6736 5956
rect 7752 6012 7816 6016
rect 7752 5956 7756 6012
rect 7756 5956 7812 6012
rect 7812 5956 7816 6012
rect 7752 5952 7816 5956
rect 7832 6012 7896 6016
rect 7832 5956 7836 6012
rect 7836 5956 7892 6012
rect 7892 5956 7896 6012
rect 7832 5952 7896 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 1812 5468 1876 5472
rect 1812 5412 1816 5468
rect 1816 5412 1872 5468
rect 1872 5412 1876 5468
rect 1812 5408 1876 5412
rect 1892 5468 1956 5472
rect 1892 5412 1896 5468
rect 1896 5412 1952 5468
rect 1952 5412 1956 5468
rect 1892 5408 1956 5412
rect 1972 5468 2036 5472
rect 1972 5412 1976 5468
rect 1976 5412 2032 5468
rect 2032 5412 2036 5468
rect 1972 5408 2036 5412
rect 2052 5468 2116 5472
rect 2052 5412 2056 5468
rect 2056 5412 2112 5468
rect 2112 5412 2116 5468
rect 2052 5408 2116 5412
rect 3132 5468 3196 5472
rect 3132 5412 3136 5468
rect 3136 5412 3192 5468
rect 3192 5412 3196 5468
rect 3132 5408 3196 5412
rect 3212 5468 3276 5472
rect 3212 5412 3216 5468
rect 3216 5412 3272 5468
rect 3272 5412 3276 5468
rect 3212 5408 3276 5412
rect 3292 5468 3356 5472
rect 3292 5412 3296 5468
rect 3296 5412 3352 5468
rect 3352 5412 3356 5468
rect 3292 5408 3356 5412
rect 3372 5468 3436 5472
rect 3372 5412 3376 5468
rect 3376 5412 3432 5468
rect 3432 5412 3436 5468
rect 3372 5408 3436 5412
rect 4452 5468 4516 5472
rect 4452 5412 4456 5468
rect 4456 5412 4512 5468
rect 4512 5412 4516 5468
rect 4452 5408 4516 5412
rect 4532 5468 4596 5472
rect 4532 5412 4536 5468
rect 4536 5412 4592 5468
rect 4592 5412 4596 5468
rect 4532 5408 4596 5412
rect 4612 5468 4676 5472
rect 4612 5412 4616 5468
rect 4616 5412 4672 5468
rect 4672 5412 4676 5468
rect 4612 5408 4676 5412
rect 4692 5468 4756 5472
rect 4692 5412 4696 5468
rect 4696 5412 4752 5468
rect 4752 5412 4756 5468
rect 4692 5408 4756 5412
rect 5772 5468 5836 5472
rect 5772 5412 5776 5468
rect 5776 5412 5832 5468
rect 5832 5412 5836 5468
rect 5772 5408 5836 5412
rect 5852 5468 5916 5472
rect 5852 5412 5856 5468
rect 5856 5412 5912 5468
rect 5912 5412 5916 5468
rect 5852 5408 5916 5412
rect 5932 5468 5996 5472
rect 5932 5412 5936 5468
rect 5936 5412 5992 5468
rect 5992 5412 5996 5468
rect 5932 5408 5996 5412
rect 6012 5468 6076 5472
rect 6012 5412 6016 5468
rect 6016 5412 6072 5468
rect 6072 5412 6076 5468
rect 6012 5408 6076 5412
rect 7092 5468 7156 5472
rect 7092 5412 7096 5468
rect 7096 5412 7152 5468
rect 7152 5412 7156 5468
rect 7092 5408 7156 5412
rect 7172 5468 7236 5472
rect 7172 5412 7176 5468
rect 7176 5412 7232 5468
rect 7232 5412 7236 5468
rect 7172 5408 7236 5412
rect 7252 5468 7316 5472
rect 7252 5412 7256 5468
rect 7256 5412 7312 5468
rect 7312 5412 7316 5468
rect 7252 5408 7316 5412
rect 7332 5468 7396 5472
rect 7332 5412 7336 5468
rect 7336 5412 7392 5468
rect 7392 5412 7396 5468
rect 7332 5408 7396 5412
rect 8412 5468 8476 5472
rect 8412 5412 8416 5468
rect 8416 5412 8472 5468
rect 8472 5412 8476 5468
rect 8412 5408 8476 5412
rect 8492 5468 8556 5472
rect 8492 5412 8496 5468
rect 8496 5412 8552 5468
rect 8552 5412 8556 5468
rect 8492 5408 8556 5412
rect 8572 5468 8636 5472
rect 8572 5412 8576 5468
rect 8576 5412 8632 5468
rect 8632 5412 8636 5468
rect 8572 5408 8636 5412
rect 8652 5468 8716 5472
rect 8652 5412 8656 5468
rect 8656 5412 8712 5468
rect 8712 5412 8716 5468
rect 8652 5408 8716 5412
rect 1152 4924 1216 4928
rect 1152 4868 1156 4924
rect 1156 4868 1212 4924
rect 1212 4868 1216 4924
rect 1152 4864 1216 4868
rect 1232 4924 1296 4928
rect 1232 4868 1236 4924
rect 1236 4868 1292 4924
rect 1292 4868 1296 4924
rect 1232 4864 1296 4868
rect 1312 4924 1376 4928
rect 1312 4868 1316 4924
rect 1316 4868 1372 4924
rect 1372 4868 1376 4924
rect 1312 4864 1376 4868
rect 1392 4924 1456 4928
rect 1392 4868 1396 4924
rect 1396 4868 1452 4924
rect 1452 4868 1456 4924
rect 1392 4864 1456 4868
rect 2472 4924 2536 4928
rect 2472 4868 2476 4924
rect 2476 4868 2532 4924
rect 2532 4868 2536 4924
rect 2472 4864 2536 4868
rect 2552 4924 2616 4928
rect 2552 4868 2556 4924
rect 2556 4868 2612 4924
rect 2612 4868 2616 4924
rect 2552 4864 2616 4868
rect 2632 4924 2696 4928
rect 2632 4868 2636 4924
rect 2636 4868 2692 4924
rect 2692 4868 2696 4924
rect 2632 4864 2696 4868
rect 2712 4924 2776 4928
rect 2712 4868 2716 4924
rect 2716 4868 2772 4924
rect 2772 4868 2776 4924
rect 2712 4864 2776 4868
rect 3792 4924 3856 4928
rect 3792 4868 3796 4924
rect 3796 4868 3852 4924
rect 3852 4868 3856 4924
rect 3792 4864 3856 4868
rect 3872 4924 3936 4928
rect 3872 4868 3876 4924
rect 3876 4868 3932 4924
rect 3932 4868 3936 4924
rect 3872 4864 3936 4868
rect 3952 4924 4016 4928
rect 3952 4868 3956 4924
rect 3956 4868 4012 4924
rect 4012 4868 4016 4924
rect 3952 4864 4016 4868
rect 4032 4924 4096 4928
rect 4032 4868 4036 4924
rect 4036 4868 4092 4924
rect 4092 4868 4096 4924
rect 4032 4864 4096 4868
rect 5112 4924 5176 4928
rect 5112 4868 5116 4924
rect 5116 4868 5172 4924
rect 5172 4868 5176 4924
rect 5112 4864 5176 4868
rect 5192 4924 5256 4928
rect 5192 4868 5196 4924
rect 5196 4868 5252 4924
rect 5252 4868 5256 4924
rect 5192 4864 5256 4868
rect 5272 4924 5336 4928
rect 5272 4868 5276 4924
rect 5276 4868 5332 4924
rect 5332 4868 5336 4924
rect 5272 4864 5336 4868
rect 5352 4924 5416 4928
rect 5352 4868 5356 4924
rect 5356 4868 5412 4924
rect 5412 4868 5416 4924
rect 5352 4864 5416 4868
rect 6432 4924 6496 4928
rect 6432 4868 6436 4924
rect 6436 4868 6492 4924
rect 6492 4868 6496 4924
rect 6432 4864 6496 4868
rect 6512 4924 6576 4928
rect 6512 4868 6516 4924
rect 6516 4868 6572 4924
rect 6572 4868 6576 4924
rect 6512 4864 6576 4868
rect 6592 4924 6656 4928
rect 6592 4868 6596 4924
rect 6596 4868 6652 4924
rect 6652 4868 6656 4924
rect 6592 4864 6656 4868
rect 6672 4924 6736 4928
rect 6672 4868 6676 4924
rect 6676 4868 6732 4924
rect 6732 4868 6736 4924
rect 6672 4864 6736 4868
rect 7752 4924 7816 4928
rect 7752 4868 7756 4924
rect 7756 4868 7812 4924
rect 7812 4868 7816 4924
rect 7752 4864 7816 4868
rect 7832 4924 7896 4928
rect 7832 4868 7836 4924
rect 7836 4868 7892 4924
rect 7892 4868 7896 4924
rect 7832 4864 7896 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 1812 4380 1876 4384
rect 1812 4324 1816 4380
rect 1816 4324 1872 4380
rect 1872 4324 1876 4380
rect 1812 4320 1876 4324
rect 1892 4380 1956 4384
rect 1892 4324 1896 4380
rect 1896 4324 1952 4380
rect 1952 4324 1956 4380
rect 1892 4320 1956 4324
rect 1972 4380 2036 4384
rect 1972 4324 1976 4380
rect 1976 4324 2032 4380
rect 2032 4324 2036 4380
rect 1972 4320 2036 4324
rect 2052 4380 2116 4384
rect 2052 4324 2056 4380
rect 2056 4324 2112 4380
rect 2112 4324 2116 4380
rect 2052 4320 2116 4324
rect 3132 4380 3196 4384
rect 3132 4324 3136 4380
rect 3136 4324 3192 4380
rect 3192 4324 3196 4380
rect 3132 4320 3196 4324
rect 3212 4380 3276 4384
rect 3212 4324 3216 4380
rect 3216 4324 3272 4380
rect 3272 4324 3276 4380
rect 3212 4320 3276 4324
rect 3292 4380 3356 4384
rect 3292 4324 3296 4380
rect 3296 4324 3352 4380
rect 3352 4324 3356 4380
rect 3292 4320 3356 4324
rect 3372 4380 3436 4384
rect 3372 4324 3376 4380
rect 3376 4324 3432 4380
rect 3432 4324 3436 4380
rect 3372 4320 3436 4324
rect 4452 4380 4516 4384
rect 4452 4324 4456 4380
rect 4456 4324 4512 4380
rect 4512 4324 4516 4380
rect 4452 4320 4516 4324
rect 4532 4380 4596 4384
rect 4532 4324 4536 4380
rect 4536 4324 4592 4380
rect 4592 4324 4596 4380
rect 4532 4320 4596 4324
rect 4612 4380 4676 4384
rect 4612 4324 4616 4380
rect 4616 4324 4672 4380
rect 4672 4324 4676 4380
rect 4612 4320 4676 4324
rect 4692 4380 4756 4384
rect 4692 4324 4696 4380
rect 4696 4324 4752 4380
rect 4752 4324 4756 4380
rect 4692 4320 4756 4324
rect 5772 4380 5836 4384
rect 5772 4324 5776 4380
rect 5776 4324 5832 4380
rect 5832 4324 5836 4380
rect 5772 4320 5836 4324
rect 5852 4380 5916 4384
rect 5852 4324 5856 4380
rect 5856 4324 5912 4380
rect 5912 4324 5916 4380
rect 5852 4320 5916 4324
rect 5932 4380 5996 4384
rect 5932 4324 5936 4380
rect 5936 4324 5992 4380
rect 5992 4324 5996 4380
rect 5932 4320 5996 4324
rect 6012 4380 6076 4384
rect 6012 4324 6016 4380
rect 6016 4324 6072 4380
rect 6072 4324 6076 4380
rect 6012 4320 6076 4324
rect 7092 4380 7156 4384
rect 7092 4324 7096 4380
rect 7096 4324 7152 4380
rect 7152 4324 7156 4380
rect 7092 4320 7156 4324
rect 7172 4380 7236 4384
rect 7172 4324 7176 4380
rect 7176 4324 7232 4380
rect 7232 4324 7236 4380
rect 7172 4320 7236 4324
rect 7252 4380 7316 4384
rect 7252 4324 7256 4380
rect 7256 4324 7312 4380
rect 7312 4324 7316 4380
rect 7252 4320 7316 4324
rect 7332 4380 7396 4384
rect 7332 4324 7336 4380
rect 7336 4324 7392 4380
rect 7392 4324 7396 4380
rect 7332 4320 7396 4324
rect 8412 4380 8476 4384
rect 8412 4324 8416 4380
rect 8416 4324 8472 4380
rect 8472 4324 8476 4380
rect 8412 4320 8476 4324
rect 8492 4380 8556 4384
rect 8492 4324 8496 4380
rect 8496 4324 8552 4380
rect 8552 4324 8556 4380
rect 8492 4320 8556 4324
rect 8572 4380 8636 4384
rect 8572 4324 8576 4380
rect 8576 4324 8632 4380
rect 8632 4324 8636 4380
rect 8572 4320 8636 4324
rect 8652 4380 8716 4384
rect 8652 4324 8656 4380
rect 8656 4324 8712 4380
rect 8712 4324 8716 4380
rect 8652 4320 8716 4324
rect 1152 3836 1216 3840
rect 1152 3780 1156 3836
rect 1156 3780 1212 3836
rect 1212 3780 1216 3836
rect 1152 3776 1216 3780
rect 1232 3836 1296 3840
rect 1232 3780 1236 3836
rect 1236 3780 1292 3836
rect 1292 3780 1296 3836
rect 1232 3776 1296 3780
rect 1312 3836 1376 3840
rect 1312 3780 1316 3836
rect 1316 3780 1372 3836
rect 1372 3780 1376 3836
rect 1312 3776 1376 3780
rect 1392 3836 1456 3840
rect 1392 3780 1396 3836
rect 1396 3780 1452 3836
rect 1452 3780 1456 3836
rect 1392 3776 1456 3780
rect 2472 3836 2536 3840
rect 2472 3780 2476 3836
rect 2476 3780 2532 3836
rect 2532 3780 2536 3836
rect 2472 3776 2536 3780
rect 2552 3836 2616 3840
rect 2552 3780 2556 3836
rect 2556 3780 2612 3836
rect 2612 3780 2616 3836
rect 2552 3776 2616 3780
rect 2632 3836 2696 3840
rect 2632 3780 2636 3836
rect 2636 3780 2692 3836
rect 2692 3780 2696 3836
rect 2632 3776 2696 3780
rect 2712 3836 2776 3840
rect 2712 3780 2716 3836
rect 2716 3780 2772 3836
rect 2772 3780 2776 3836
rect 2712 3776 2776 3780
rect 3792 3836 3856 3840
rect 3792 3780 3796 3836
rect 3796 3780 3852 3836
rect 3852 3780 3856 3836
rect 3792 3776 3856 3780
rect 3872 3836 3936 3840
rect 3872 3780 3876 3836
rect 3876 3780 3932 3836
rect 3932 3780 3936 3836
rect 3872 3776 3936 3780
rect 3952 3836 4016 3840
rect 3952 3780 3956 3836
rect 3956 3780 4012 3836
rect 4012 3780 4016 3836
rect 3952 3776 4016 3780
rect 4032 3836 4096 3840
rect 4032 3780 4036 3836
rect 4036 3780 4092 3836
rect 4092 3780 4096 3836
rect 4032 3776 4096 3780
rect 5112 3836 5176 3840
rect 5112 3780 5116 3836
rect 5116 3780 5172 3836
rect 5172 3780 5176 3836
rect 5112 3776 5176 3780
rect 5192 3836 5256 3840
rect 5192 3780 5196 3836
rect 5196 3780 5252 3836
rect 5252 3780 5256 3836
rect 5192 3776 5256 3780
rect 5272 3836 5336 3840
rect 5272 3780 5276 3836
rect 5276 3780 5332 3836
rect 5332 3780 5336 3836
rect 5272 3776 5336 3780
rect 5352 3836 5416 3840
rect 5352 3780 5356 3836
rect 5356 3780 5412 3836
rect 5412 3780 5416 3836
rect 5352 3776 5416 3780
rect 6432 3836 6496 3840
rect 6432 3780 6436 3836
rect 6436 3780 6492 3836
rect 6492 3780 6496 3836
rect 6432 3776 6496 3780
rect 6512 3836 6576 3840
rect 6512 3780 6516 3836
rect 6516 3780 6572 3836
rect 6572 3780 6576 3836
rect 6512 3776 6576 3780
rect 6592 3836 6656 3840
rect 6592 3780 6596 3836
rect 6596 3780 6652 3836
rect 6652 3780 6656 3836
rect 6592 3776 6656 3780
rect 6672 3836 6736 3840
rect 6672 3780 6676 3836
rect 6676 3780 6732 3836
rect 6732 3780 6736 3836
rect 6672 3776 6736 3780
rect 7752 3836 7816 3840
rect 7752 3780 7756 3836
rect 7756 3780 7812 3836
rect 7812 3780 7816 3836
rect 7752 3776 7816 3780
rect 7832 3836 7896 3840
rect 7832 3780 7836 3836
rect 7836 3780 7892 3836
rect 7892 3780 7896 3836
rect 7832 3776 7896 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 1812 3292 1876 3296
rect 1812 3236 1816 3292
rect 1816 3236 1872 3292
rect 1872 3236 1876 3292
rect 1812 3232 1876 3236
rect 1892 3292 1956 3296
rect 1892 3236 1896 3292
rect 1896 3236 1952 3292
rect 1952 3236 1956 3292
rect 1892 3232 1956 3236
rect 1972 3292 2036 3296
rect 1972 3236 1976 3292
rect 1976 3236 2032 3292
rect 2032 3236 2036 3292
rect 1972 3232 2036 3236
rect 2052 3292 2116 3296
rect 2052 3236 2056 3292
rect 2056 3236 2112 3292
rect 2112 3236 2116 3292
rect 2052 3232 2116 3236
rect 3132 3292 3196 3296
rect 3132 3236 3136 3292
rect 3136 3236 3192 3292
rect 3192 3236 3196 3292
rect 3132 3232 3196 3236
rect 3212 3292 3276 3296
rect 3212 3236 3216 3292
rect 3216 3236 3272 3292
rect 3272 3236 3276 3292
rect 3212 3232 3276 3236
rect 3292 3292 3356 3296
rect 3292 3236 3296 3292
rect 3296 3236 3352 3292
rect 3352 3236 3356 3292
rect 3292 3232 3356 3236
rect 3372 3292 3436 3296
rect 3372 3236 3376 3292
rect 3376 3236 3432 3292
rect 3432 3236 3436 3292
rect 3372 3232 3436 3236
rect 4452 3292 4516 3296
rect 4452 3236 4456 3292
rect 4456 3236 4512 3292
rect 4512 3236 4516 3292
rect 4452 3232 4516 3236
rect 4532 3292 4596 3296
rect 4532 3236 4536 3292
rect 4536 3236 4592 3292
rect 4592 3236 4596 3292
rect 4532 3232 4596 3236
rect 4612 3292 4676 3296
rect 4612 3236 4616 3292
rect 4616 3236 4672 3292
rect 4672 3236 4676 3292
rect 4612 3232 4676 3236
rect 4692 3292 4756 3296
rect 4692 3236 4696 3292
rect 4696 3236 4752 3292
rect 4752 3236 4756 3292
rect 4692 3232 4756 3236
rect 5772 3292 5836 3296
rect 5772 3236 5776 3292
rect 5776 3236 5832 3292
rect 5832 3236 5836 3292
rect 5772 3232 5836 3236
rect 5852 3292 5916 3296
rect 5852 3236 5856 3292
rect 5856 3236 5912 3292
rect 5912 3236 5916 3292
rect 5852 3232 5916 3236
rect 5932 3292 5996 3296
rect 5932 3236 5936 3292
rect 5936 3236 5992 3292
rect 5992 3236 5996 3292
rect 5932 3232 5996 3236
rect 6012 3292 6076 3296
rect 6012 3236 6016 3292
rect 6016 3236 6072 3292
rect 6072 3236 6076 3292
rect 6012 3232 6076 3236
rect 7092 3292 7156 3296
rect 7092 3236 7096 3292
rect 7096 3236 7152 3292
rect 7152 3236 7156 3292
rect 7092 3232 7156 3236
rect 7172 3292 7236 3296
rect 7172 3236 7176 3292
rect 7176 3236 7232 3292
rect 7232 3236 7236 3292
rect 7172 3232 7236 3236
rect 7252 3292 7316 3296
rect 7252 3236 7256 3292
rect 7256 3236 7312 3292
rect 7312 3236 7316 3292
rect 7252 3232 7316 3236
rect 7332 3292 7396 3296
rect 7332 3236 7336 3292
rect 7336 3236 7392 3292
rect 7392 3236 7396 3292
rect 7332 3232 7396 3236
rect 8412 3292 8476 3296
rect 8412 3236 8416 3292
rect 8416 3236 8472 3292
rect 8472 3236 8476 3292
rect 8412 3232 8476 3236
rect 8492 3292 8556 3296
rect 8492 3236 8496 3292
rect 8496 3236 8552 3292
rect 8552 3236 8556 3292
rect 8492 3232 8556 3236
rect 8572 3292 8636 3296
rect 8572 3236 8576 3292
rect 8576 3236 8632 3292
rect 8632 3236 8636 3292
rect 8572 3232 8636 3236
rect 8652 3292 8716 3296
rect 8652 3236 8656 3292
rect 8656 3236 8712 3292
rect 8712 3236 8716 3292
rect 8652 3232 8716 3236
rect 1152 2748 1216 2752
rect 1152 2692 1156 2748
rect 1156 2692 1212 2748
rect 1212 2692 1216 2748
rect 1152 2688 1216 2692
rect 1232 2748 1296 2752
rect 1232 2692 1236 2748
rect 1236 2692 1292 2748
rect 1292 2692 1296 2748
rect 1232 2688 1296 2692
rect 1312 2748 1376 2752
rect 1312 2692 1316 2748
rect 1316 2692 1372 2748
rect 1372 2692 1376 2748
rect 1312 2688 1376 2692
rect 1392 2748 1456 2752
rect 1392 2692 1396 2748
rect 1396 2692 1452 2748
rect 1452 2692 1456 2748
rect 1392 2688 1456 2692
rect 2472 2748 2536 2752
rect 2472 2692 2476 2748
rect 2476 2692 2532 2748
rect 2532 2692 2536 2748
rect 2472 2688 2536 2692
rect 2552 2748 2616 2752
rect 2552 2692 2556 2748
rect 2556 2692 2612 2748
rect 2612 2692 2616 2748
rect 2552 2688 2616 2692
rect 2632 2748 2696 2752
rect 2632 2692 2636 2748
rect 2636 2692 2692 2748
rect 2692 2692 2696 2748
rect 2632 2688 2696 2692
rect 2712 2748 2776 2752
rect 2712 2692 2716 2748
rect 2716 2692 2772 2748
rect 2772 2692 2776 2748
rect 2712 2688 2776 2692
rect 3792 2748 3856 2752
rect 3792 2692 3796 2748
rect 3796 2692 3852 2748
rect 3852 2692 3856 2748
rect 3792 2688 3856 2692
rect 3872 2748 3936 2752
rect 3872 2692 3876 2748
rect 3876 2692 3932 2748
rect 3932 2692 3936 2748
rect 3872 2688 3936 2692
rect 3952 2748 4016 2752
rect 3952 2692 3956 2748
rect 3956 2692 4012 2748
rect 4012 2692 4016 2748
rect 3952 2688 4016 2692
rect 4032 2748 4096 2752
rect 4032 2692 4036 2748
rect 4036 2692 4092 2748
rect 4092 2692 4096 2748
rect 4032 2688 4096 2692
rect 5112 2748 5176 2752
rect 5112 2692 5116 2748
rect 5116 2692 5172 2748
rect 5172 2692 5176 2748
rect 5112 2688 5176 2692
rect 5192 2748 5256 2752
rect 5192 2692 5196 2748
rect 5196 2692 5252 2748
rect 5252 2692 5256 2748
rect 5192 2688 5256 2692
rect 5272 2748 5336 2752
rect 5272 2692 5276 2748
rect 5276 2692 5332 2748
rect 5332 2692 5336 2748
rect 5272 2688 5336 2692
rect 5352 2748 5416 2752
rect 5352 2692 5356 2748
rect 5356 2692 5412 2748
rect 5412 2692 5416 2748
rect 5352 2688 5416 2692
rect 6432 2748 6496 2752
rect 6432 2692 6436 2748
rect 6436 2692 6492 2748
rect 6492 2692 6496 2748
rect 6432 2688 6496 2692
rect 6512 2748 6576 2752
rect 6512 2692 6516 2748
rect 6516 2692 6572 2748
rect 6572 2692 6576 2748
rect 6512 2688 6576 2692
rect 6592 2748 6656 2752
rect 6592 2692 6596 2748
rect 6596 2692 6652 2748
rect 6652 2692 6656 2748
rect 6592 2688 6656 2692
rect 6672 2748 6736 2752
rect 6672 2692 6676 2748
rect 6676 2692 6732 2748
rect 6732 2692 6736 2748
rect 6672 2688 6736 2692
rect 7752 2748 7816 2752
rect 7752 2692 7756 2748
rect 7756 2692 7812 2748
rect 7812 2692 7816 2748
rect 7752 2688 7816 2692
rect 7832 2748 7896 2752
rect 7832 2692 7836 2748
rect 7836 2692 7892 2748
rect 7892 2692 7896 2748
rect 7832 2688 7896 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 1812 2204 1876 2208
rect 1812 2148 1816 2204
rect 1816 2148 1872 2204
rect 1872 2148 1876 2204
rect 1812 2144 1876 2148
rect 1892 2204 1956 2208
rect 1892 2148 1896 2204
rect 1896 2148 1952 2204
rect 1952 2148 1956 2204
rect 1892 2144 1956 2148
rect 1972 2204 2036 2208
rect 1972 2148 1976 2204
rect 1976 2148 2032 2204
rect 2032 2148 2036 2204
rect 1972 2144 2036 2148
rect 2052 2204 2116 2208
rect 2052 2148 2056 2204
rect 2056 2148 2112 2204
rect 2112 2148 2116 2204
rect 2052 2144 2116 2148
rect 3132 2204 3196 2208
rect 3132 2148 3136 2204
rect 3136 2148 3192 2204
rect 3192 2148 3196 2204
rect 3132 2144 3196 2148
rect 3212 2204 3276 2208
rect 3212 2148 3216 2204
rect 3216 2148 3272 2204
rect 3272 2148 3276 2204
rect 3212 2144 3276 2148
rect 3292 2204 3356 2208
rect 3292 2148 3296 2204
rect 3296 2148 3352 2204
rect 3352 2148 3356 2204
rect 3292 2144 3356 2148
rect 3372 2204 3436 2208
rect 3372 2148 3376 2204
rect 3376 2148 3432 2204
rect 3432 2148 3436 2204
rect 3372 2144 3436 2148
rect 4452 2204 4516 2208
rect 4452 2148 4456 2204
rect 4456 2148 4512 2204
rect 4512 2148 4516 2204
rect 4452 2144 4516 2148
rect 4532 2204 4596 2208
rect 4532 2148 4536 2204
rect 4536 2148 4592 2204
rect 4592 2148 4596 2204
rect 4532 2144 4596 2148
rect 4612 2204 4676 2208
rect 4612 2148 4616 2204
rect 4616 2148 4672 2204
rect 4672 2148 4676 2204
rect 4612 2144 4676 2148
rect 4692 2204 4756 2208
rect 4692 2148 4696 2204
rect 4696 2148 4752 2204
rect 4752 2148 4756 2204
rect 4692 2144 4756 2148
rect 5772 2204 5836 2208
rect 5772 2148 5776 2204
rect 5776 2148 5832 2204
rect 5832 2148 5836 2204
rect 5772 2144 5836 2148
rect 5852 2204 5916 2208
rect 5852 2148 5856 2204
rect 5856 2148 5912 2204
rect 5912 2148 5916 2204
rect 5852 2144 5916 2148
rect 5932 2204 5996 2208
rect 5932 2148 5936 2204
rect 5936 2148 5992 2204
rect 5992 2148 5996 2204
rect 5932 2144 5996 2148
rect 6012 2204 6076 2208
rect 6012 2148 6016 2204
rect 6016 2148 6072 2204
rect 6072 2148 6076 2204
rect 6012 2144 6076 2148
rect 7092 2204 7156 2208
rect 7092 2148 7096 2204
rect 7096 2148 7152 2204
rect 7152 2148 7156 2204
rect 7092 2144 7156 2148
rect 7172 2204 7236 2208
rect 7172 2148 7176 2204
rect 7176 2148 7232 2204
rect 7232 2148 7236 2204
rect 7172 2144 7236 2148
rect 7252 2204 7316 2208
rect 7252 2148 7256 2204
rect 7256 2148 7312 2204
rect 7312 2148 7316 2204
rect 7252 2144 7316 2148
rect 7332 2204 7396 2208
rect 7332 2148 7336 2204
rect 7336 2148 7392 2204
rect 7392 2148 7396 2204
rect 7332 2144 7396 2148
rect 8412 2204 8476 2208
rect 8412 2148 8416 2204
rect 8416 2148 8472 2204
rect 8472 2148 8476 2204
rect 8412 2144 8476 2148
rect 8492 2204 8556 2208
rect 8492 2148 8496 2204
rect 8496 2148 8552 2204
rect 8552 2148 8556 2204
rect 8492 2144 8556 2148
rect 8572 2204 8636 2208
rect 8572 2148 8576 2204
rect 8576 2148 8632 2204
rect 8632 2148 8636 2204
rect 8572 2144 8636 2148
rect 8652 2204 8716 2208
rect 8652 2148 8656 2204
rect 8656 2148 8712 2204
rect 8712 2148 8716 2204
rect 8652 2144 8716 2148
rect 1358 1820 7744 2018
<< metal4 >>
rect 1800 10204 8722 10260
rect 1800 10006 2136 10204
rect 8522 10006 8722 10204
rect 1800 9944 8722 10006
rect 1800 9840 2084 9944
rect 1144 9280 1464 9840
rect 1800 9824 2124 9840
rect 1144 9216 1152 9280
rect 1216 9216 1232 9280
rect 1296 9216 1312 9280
rect 1376 9216 1392 9280
rect 1456 9216 1464 9280
rect 1144 9094 1464 9216
rect 1144 8858 1186 9094
rect 1422 8858 1464 9094
rect 1144 8192 1464 8858
rect 1144 8128 1152 8192
rect 1216 8128 1232 8192
rect 1296 8128 1312 8192
rect 1376 8128 1392 8192
rect 1456 8128 1464 8192
rect 1144 7774 1464 8128
rect 1144 7538 1186 7774
rect 1422 7538 1464 7774
rect 1144 7104 1464 7538
rect 1144 7040 1152 7104
rect 1216 7040 1232 7104
rect 1296 7040 1312 7104
rect 1376 7040 1392 7104
rect 1456 7040 1464 7104
rect 1144 6454 1464 7040
rect 1144 6218 1186 6454
rect 1422 6218 1464 6454
rect 1144 6016 1464 6218
rect 1144 5952 1152 6016
rect 1216 5952 1232 6016
rect 1296 5952 1312 6016
rect 1376 5952 1392 6016
rect 1456 5952 1464 6016
rect 1144 5134 1464 5952
rect 1144 4928 1186 5134
rect 1422 4928 1464 5134
rect 1144 4864 1152 4928
rect 1216 4864 1232 4898
rect 1296 4864 1312 4898
rect 1376 4864 1392 4898
rect 1456 4864 1464 4928
rect 1144 3840 1464 4864
rect 1144 3776 1152 3840
rect 1216 3814 1232 3840
rect 1296 3814 1312 3840
rect 1376 3814 1392 3840
rect 1456 3776 1464 3840
rect 1144 3578 1186 3776
rect 1422 3578 1464 3776
rect 1144 2752 1464 3578
rect 1144 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1464 2752
rect 1142 2494 1464 2688
rect 1142 2258 1186 2494
rect 1422 2258 1464 2494
rect 1142 2128 1464 2258
rect 1804 9760 1812 9824
rect 1876 9760 1892 9824
rect 1956 9760 1972 9824
rect 2036 9760 2052 9824
rect 2116 9760 2124 9824
rect 1804 9754 2124 9760
rect 1804 9518 1846 9754
rect 2082 9518 2124 9754
rect 1804 8736 2124 9518
rect 1804 8672 1812 8736
rect 1876 8672 1892 8736
rect 1956 8672 1972 8736
rect 2036 8672 2052 8736
rect 2116 8672 2124 8736
rect 1804 8434 2124 8672
rect 1804 8198 1846 8434
rect 2082 8198 2124 8434
rect 1804 7648 2124 8198
rect 1804 7584 1812 7648
rect 1876 7584 1892 7648
rect 1956 7584 1972 7648
rect 2036 7584 2052 7648
rect 2116 7584 2124 7648
rect 1804 7114 2124 7584
rect 1804 6878 1846 7114
rect 2082 6878 2124 7114
rect 1804 6560 2124 6878
rect 1804 6496 1812 6560
rect 1876 6496 1892 6560
rect 1956 6496 1972 6560
rect 2036 6496 2052 6560
rect 2116 6496 2124 6560
rect 1804 5794 2124 6496
rect 1804 5558 1846 5794
rect 2082 5558 2124 5794
rect 1804 5472 2124 5558
rect 1804 5408 1812 5472
rect 1876 5408 1892 5472
rect 1956 5408 1972 5472
rect 2036 5408 2052 5472
rect 2116 5408 2124 5472
rect 1804 4474 2124 5408
rect 1804 4384 1846 4474
rect 2082 4384 2124 4474
rect 1804 4320 1812 4384
rect 2116 4320 2124 4384
rect 1804 4238 1846 4320
rect 2082 4238 2124 4320
rect 1804 3296 2124 4238
rect 1804 3232 1812 3296
rect 1876 3232 1892 3296
rect 1956 3232 1972 3296
rect 2036 3232 2052 3296
rect 2116 3232 2124 3296
rect 1804 3154 2124 3232
rect 1804 2918 1846 3154
rect 2082 2918 2124 3154
rect 1804 2208 2124 2918
rect 2464 9280 2784 9840
rect 3122 9824 3458 9944
rect 5772 9840 6088 9944
rect 7090 9840 7406 9944
rect 8406 9840 8722 9944
rect 2464 9216 2472 9280
rect 2536 9216 2552 9280
rect 2616 9216 2632 9280
rect 2696 9216 2712 9280
rect 2776 9216 2784 9280
rect 2464 9094 2784 9216
rect 2464 8858 2506 9094
rect 2742 8858 2784 9094
rect 2464 8192 2784 8858
rect 2464 8128 2472 8192
rect 2536 8128 2552 8192
rect 2616 8128 2632 8192
rect 2696 8128 2712 8192
rect 2776 8128 2784 8192
rect 2464 7774 2784 8128
rect 2464 7538 2506 7774
rect 2742 7538 2784 7774
rect 2464 7104 2784 7538
rect 2464 7040 2472 7104
rect 2536 7040 2552 7104
rect 2616 7040 2632 7104
rect 2696 7040 2712 7104
rect 2776 7040 2784 7104
rect 2464 6454 2784 7040
rect 2464 6218 2506 6454
rect 2742 6218 2784 6454
rect 2464 6016 2784 6218
rect 2464 5952 2472 6016
rect 2536 5952 2552 6016
rect 2616 5952 2632 6016
rect 2696 5952 2712 6016
rect 2776 5952 2784 6016
rect 2464 5134 2784 5952
rect 2464 4928 2506 5134
rect 2742 4928 2784 5134
rect 2464 4864 2472 4928
rect 2536 4864 2552 4898
rect 2616 4864 2632 4898
rect 2696 4864 2712 4898
rect 2776 4864 2784 4928
rect 2464 3840 2784 4864
rect 2464 3776 2472 3840
rect 2536 3814 2552 3840
rect 2616 3814 2632 3840
rect 2696 3814 2712 3840
rect 2776 3776 2784 3840
rect 2464 3578 2506 3776
rect 2742 3578 2784 3776
rect 2464 2752 2784 3578
rect 2464 2688 2472 2752
rect 2536 2688 2552 2752
rect 2616 2688 2632 2752
rect 2696 2688 2712 2752
rect 2776 2688 2784 2752
rect 1804 2144 1812 2208
rect 1876 2144 1892 2208
rect 1956 2144 1972 2208
rect 2036 2144 2052 2208
rect 2116 2144 2124 2208
rect 1804 2128 2124 2144
rect 2462 2494 2784 2688
rect 2462 2258 2506 2494
rect 2742 2258 2784 2494
rect 2462 2128 2784 2258
rect 3124 9760 3132 9824
rect 3196 9760 3212 9824
rect 3276 9760 3292 9824
rect 3356 9760 3372 9824
rect 3436 9760 3444 9824
rect 3124 9754 3444 9760
rect 3124 9518 3166 9754
rect 3402 9518 3444 9754
rect 3124 8736 3444 9518
rect 3124 8672 3132 8736
rect 3196 8672 3212 8736
rect 3276 8672 3292 8736
rect 3356 8672 3372 8736
rect 3436 8672 3444 8736
rect 3124 8434 3444 8672
rect 3124 8198 3166 8434
rect 3402 8198 3444 8434
rect 3124 7648 3444 8198
rect 3124 7584 3132 7648
rect 3196 7584 3212 7648
rect 3276 7584 3292 7648
rect 3356 7584 3372 7648
rect 3436 7584 3444 7648
rect 3124 7114 3444 7584
rect 3124 6878 3166 7114
rect 3402 6878 3444 7114
rect 3124 6560 3444 6878
rect 3124 6496 3132 6560
rect 3196 6496 3212 6560
rect 3276 6496 3292 6560
rect 3356 6496 3372 6560
rect 3436 6496 3444 6560
rect 3124 5794 3444 6496
rect 3124 5558 3166 5794
rect 3402 5558 3444 5794
rect 3124 5472 3444 5558
rect 3124 5408 3132 5472
rect 3196 5408 3212 5472
rect 3276 5408 3292 5472
rect 3356 5408 3372 5472
rect 3436 5408 3444 5472
rect 3124 4474 3444 5408
rect 3124 4384 3166 4474
rect 3402 4384 3444 4474
rect 3124 4320 3132 4384
rect 3436 4320 3444 4384
rect 3124 4238 3166 4320
rect 3402 4238 3444 4320
rect 3124 3296 3444 4238
rect 3124 3232 3132 3296
rect 3196 3232 3212 3296
rect 3276 3232 3292 3296
rect 3356 3232 3372 3296
rect 3436 3232 3444 3296
rect 3124 3154 3444 3232
rect 3124 2918 3166 3154
rect 3402 2918 3444 3154
rect 3124 2208 3444 2918
rect 3784 9280 4104 9840
rect 3784 9216 3792 9280
rect 3856 9216 3872 9280
rect 3936 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4104 9280
rect 3784 9094 4104 9216
rect 3784 8858 3826 9094
rect 4062 8858 4104 9094
rect 3784 8192 4104 8858
rect 3784 8128 3792 8192
rect 3856 8128 3872 8192
rect 3936 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4104 8192
rect 3784 7774 4104 8128
rect 3784 7538 3826 7774
rect 4062 7538 4104 7774
rect 3784 7104 4104 7538
rect 3784 7040 3792 7104
rect 3856 7040 3872 7104
rect 3936 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4104 7104
rect 3784 6454 4104 7040
rect 3784 6218 3826 6454
rect 4062 6218 4104 6454
rect 3784 6016 4104 6218
rect 3784 5952 3792 6016
rect 3856 5952 3872 6016
rect 3936 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4104 6016
rect 3784 5134 4104 5952
rect 3784 4928 3826 5134
rect 4062 4928 4104 5134
rect 3784 4864 3792 4928
rect 3856 4864 3872 4898
rect 3936 4864 3952 4898
rect 4016 4864 4032 4898
rect 4096 4864 4104 4928
rect 3784 3840 4104 4864
rect 3784 3776 3792 3840
rect 3856 3814 3872 3840
rect 3936 3814 3952 3840
rect 4016 3814 4032 3840
rect 4096 3776 4104 3840
rect 3784 3578 3826 3776
rect 4062 3578 4104 3776
rect 3784 2752 4104 3578
rect 3784 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4104 2752
rect 3124 2144 3132 2208
rect 3196 2144 3212 2208
rect 3276 2144 3292 2208
rect 3356 2144 3372 2208
rect 3436 2144 3444 2208
rect 3124 2128 3444 2144
rect 3782 2494 4104 2688
rect 3782 2258 3826 2494
rect 4062 2258 4104 2494
rect 3782 2128 4104 2258
rect 4444 9824 4764 9840
rect 4444 9760 4452 9824
rect 4516 9760 4532 9824
rect 4596 9760 4612 9824
rect 4676 9760 4692 9824
rect 4756 9760 4764 9824
rect 4444 9754 4764 9760
rect 4444 9518 4486 9754
rect 4722 9518 4764 9754
rect 4444 8736 4764 9518
rect 4444 8672 4452 8736
rect 4516 8672 4532 8736
rect 4596 8672 4612 8736
rect 4676 8672 4692 8736
rect 4756 8672 4764 8736
rect 4444 8434 4764 8672
rect 4444 8198 4486 8434
rect 4722 8198 4764 8434
rect 4444 7648 4764 8198
rect 4444 7584 4452 7648
rect 4516 7584 4532 7648
rect 4596 7584 4612 7648
rect 4676 7584 4692 7648
rect 4756 7584 4764 7648
rect 4444 7114 4764 7584
rect 4444 6878 4486 7114
rect 4722 6878 4764 7114
rect 4444 6560 4764 6878
rect 4444 6496 4452 6560
rect 4516 6496 4532 6560
rect 4596 6496 4612 6560
rect 4676 6496 4692 6560
rect 4756 6496 4764 6560
rect 4444 5794 4764 6496
rect 4444 5558 4486 5794
rect 4722 5558 4764 5794
rect 4444 5472 4764 5558
rect 4444 5408 4452 5472
rect 4516 5408 4532 5472
rect 4596 5408 4612 5472
rect 4676 5408 4692 5472
rect 4756 5408 4764 5472
rect 4444 4474 4764 5408
rect 4444 4384 4486 4474
rect 4722 4384 4764 4474
rect 4444 4320 4452 4384
rect 4756 4320 4764 4384
rect 4444 4238 4486 4320
rect 4722 4238 4764 4320
rect 4444 3296 4764 4238
rect 4444 3232 4452 3296
rect 4516 3232 4532 3296
rect 4596 3232 4612 3296
rect 4676 3232 4692 3296
rect 4756 3232 4764 3296
rect 4444 3154 4764 3232
rect 4444 2918 4486 3154
rect 4722 2918 4764 3154
rect 4444 2208 4764 2918
rect 4444 2144 4452 2208
rect 4516 2144 4532 2208
rect 4596 2144 4612 2208
rect 4676 2144 4692 2208
rect 4756 2144 4764 2208
rect 4444 2128 4764 2144
rect 5104 9280 5424 9840
rect 5104 9216 5112 9280
rect 5176 9216 5192 9280
rect 5256 9216 5272 9280
rect 5336 9216 5352 9280
rect 5416 9216 5424 9280
rect 5104 9094 5424 9216
rect 5104 8858 5146 9094
rect 5382 8858 5424 9094
rect 5104 8192 5424 8858
rect 5104 8128 5112 8192
rect 5176 8128 5192 8192
rect 5256 8128 5272 8192
rect 5336 8128 5352 8192
rect 5416 8128 5424 8192
rect 5104 7774 5424 8128
rect 5104 7538 5146 7774
rect 5382 7538 5424 7774
rect 5104 7104 5424 7538
rect 5104 7040 5112 7104
rect 5176 7040 5192 7104
rect 5256 7040 5272 7104
rect 5336 7040 5352 7104
rect 5416 7040 5424 7104
rect 5104 6454 5424 7040
rect 5104 6218 5146 6454
rect 5382 6218 5424 6454
rect 5104 6016 5424 6218
rect 5104 5952 5112 6016
rect 5176 5952 5192 6016
rect 5256 5952 5272 6016
rect 5336 5952 5352 6016
rect 5416 5952 5424 6016
rect 5104 5134 5424 5952
rect 5104 4928 5146 5134
rect 5382 4928 5424 5134
rect 5104 4864 5112 4928
rect 5176 4864 5192 4898
rect 5256 4864 5272 4898
rect 5336 4864 5352 4898
rect 5416 4864 5424 4928
rect 5104 3840 5424 4864
rect 5104 3776 5112 3840
rect 5176 3814 5192 3840
rect 5256 3814 5272 3840
rect 5336 3814 5352 3840
rect 5416 3776 5424 3840
rect 5104 3578 5146 3776
rect 5382 3578 5424 3776
rect 5104 2752 5424 3578
rect 5104 2688 5112 2752
rect 5176 2688 5192 2752
rect 5256 2688 5272 2752
rect 5336 2688 5352 2752
rect 5416 2688 5424 2752
rect 5104 2494 5424 2688
rect 5104 2258 5146 2494
rect 5382 2258 5424 2494
rect 5104 2128 5424 2258
rect 5764 9824 6088 9840
rect 5764 9760 5772 9824
rect 5836 9760 5852 9824
rect 5916 9760 5932 9824
rect 5996 9760 6012 9824
rect 6076 9760 6084 9824
rect 5764 9754 6084 9760
rect 5764 9518 5806 9754
rect 6042 9518 6084 9754
rect 5764 8736 6084 9518
rect 5764 8672 5772 8736
rect 5836 8672 5852 8736
rect 5916 8672 5932 8736
rect 5996 8672 6012 8736
rect 6076 8672 6084 8736
rect 5764 8434 6084 8672
rect 5764 8198 5806 8434
rect 6042 8198 6084 8434
rect 5764 7648 6084 8198
rect 5764 7584 5772 7648
rect 5836 7584 5852 7648
rect 5916 7584 5932 7648
rect 5996 7584 6012 7648
rect 6076 7584 6084 7648
rect 5764 7114 6084 7584
rect 5764 6878 5806 7114
rect 6042 6878 6084 7114
rect 5764 6560 6084 6878
rect 5764 6496 5772 6560
rect 5836 6496 5852 6560
rect 5916 6496 5932 6560
rect 5996 6496 6012 6560
rect 6076 6496 6084 6560
rect 5764 5794 6084 6496
rect 5764 5558 5806 5794
rect 6042 5558 6084 5794
rect 5764 5472 6084 5558
rect 5764 5408 5772 5472
rect 5836 5408 5852 5472
rect 5916 5408 5932 5472
rect 5996 5408 6012 5472
rect 6076 5408 6084 5472
rect 5764 4474 6084 5408
rect 5764 4384 5806 4474
rect 6042 4384 6084 4474
rect 5764 4320 5772 4384
rect 6076 4320 6084 4384
rect 5764 4238 5806 4320
rect 6042 4238 6084 4320
rect 5764 3296 6084 4238
rect 5764 3232 5772 3296
rect 5836 3232 5852 3296
rect 5916 3232 5932 3296
rect 5996 3232 6012 3296
rect 6076 3232 6084 3296
rect 5764 3154 6084 3232
rect 5764 2918 5806 3154
rect 6042 2918 6084 3154
rect 5764 2208 6084 2918
rect 6424 9280 6744 9840
rect 6424 9216 6432 9280
rect 6496 9216 6512 9280
rect 6576 9216 6592 9280
rect 6656 9216 6672 9280
rect 6736 9216 6744 9280
rect 6424 9094 6744 9216
rect 6424 8858 6466 9094
rect 6702 8858 6744 9094
rect 6424 8192 6744 8858
rect 6424 8128 6432 8192
rect 6496 8128 6512 8192
rect 6576 8128 6592 8192
rect 6656 8128 6672 8192
rect 6736 8128 6744 8192
rect 6424 7774 6744 8128
rect 6424 7538 6466 7774
rect 6702 7538 6744 7774
rect 6424 7104 6744 7538
rect 6424 7040 6432 7104
rect 6496 7040 6512 7104
rect 6576 7040 6592 7104
rect 6656 7040 6672 7104
rect 6736 7040 6744 7104
rect 6424 6454 6744 7040
rect 6424 6218 6466 6454
rect 6702 6218 6744 6454
rect 6424 6016 6744 6218
rect 6424 5952 6432 6016
rect 6496 5952 6512 6016
rect 6576 5952 6592 6016
rect 6656 5952 6672 6016
rect 6736 5952 6744 6016
rect 6424 5134 6744 5952
rect 6424 4928 6466 5134
rect 6702 4928 6744 5134
rect 6424 4864 6432 4928
rect 6496 4864 6512 4898
rect 6576 4864 6592 4898
rect 6656 4864 6672 4898
rect 6736 4864 6744 4928
rect 6424 3840 6744 4864
rect 6424 3776 6432 3840
rect 6496 3814 6512 3840
rect 6576 3814 6592 3840
rect 6656 3814 6672 3840
rect 6736 3776 6744 3840
rect 6424 3578 6466 3776
rect 6702 3578 6744 3776
rect 6424 2752 6744 3578
rect 6424 2688 6432 2752
rect 6496 2688 6512 2752
rect 6576 2688 6592 2752
rect 6656 2688 6672 2752
rect 6736 2688 6744 2752
rect 5764 2144 5772 2208
rect 5836 2144 5852 2208
rect 5916 2144 5932 2208
rect 5996 2144 6012 2208
rect 6076 2144 6084 2208
rect 5764 2128 6084 2144
rect 6412 2494 6744 2688
rect 6412 2258 6466 2494
rect 6702 2258 6744 2494
rect 6412 2128 6744 2258
rect 7084 9824 7406 9840
rect 7084 9760 7092 9824
rect 7156 9760 7172 9824
rect 7236 9760 7252 9824
rect 7316 9760 7332 9824
rect 7396 9760 7404 9824
rect 7084 9754 7404 9760
rect 7084 9518 7126 9754
rect 7362 9518 7404 9754
rect 7084 8736 7404 9518
rect 7084 8672 7092 8736
rect 7156 8672 7172 8736
rect 7236 8672 7252 8736
rect 7316 8672 7332 8736
rect 7396 8672 7404 8736
rect 7084 8434 7404 8672
rect 7084 8198 7126 8434
rect 7362 8198 7404 8434
rect 7084 7648 7404 8198
rect 7084 7584 7092 7648
rect 7156 7584 7172 7648
rect 7236 7584 7252 7648
rect 7316 7584 7332 7648
rect 7396 7584 7404 7648
rect 7084 7114 7404 7584
rect 7084 6878 7126 7114
rect 7362 6878 7404 7114
rect 7084 6560 7404 6878
rect 7084 6496 7092 6560
rect 7156 6496 7172 6560
rect 7236 6496 7252 6560
rect 7316 6496 7332 6560
rect 7396 6496 7404 6560
rect 7084 5794 7404 6496
rect 7084 5558 7126 5794
rect 7362 5558 7404 5794
rect 7084 5472 7404 5558
rect 7084 5408 7092 5472
rect 7156 5408 7172 5472
rect 7236 5408 7252 5472
rect 7316 5408 7332 5472
rect 7396 5408 7404 5472
rect 7084 4474 7404 5408
rect 7084 4384 7126 4474
rect 7362 4384 7404 4474
rect 7084 4320 7092 4384
rect 7396 4320 7404 4384
rect 7084 4238 7126 4320
rect 7362 4238 7404 4320
rect 7084 3296 7404 4238
rect 7084 3232 7092 3296
rect 7156 3232 7172 3296
rect 7236 3232 7252 3296
rect 7316 3232 7332 3296
rect 7396 3232 7404 3296
rect 7084 3154 7404 3232
rect 7084 2918 7126 3154
rect 7362 2918 7404 3154
rect 7084 2208 7404 2918
rect 7084 2144 7092 2208
rect 7156 2144 7172 2208
rect 7236 2144 7252 2208
rect 7316 2144 7332 2208
rect 7396 2144 7404 2208
rect 7084 2128 7404 2144
rect 7744 9280 8064 9840
rect 7744 9216 7752 9280
rect 7816 9216 7832 9280
rect 7896 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8064 9280
rect 7744 9094 8064 9216
rect 7744 8858 7786 9094
rect 8022 8858 8064 9094
rect 7744 8192 8064 8858
rect 7744 8128 7752 8192
rect 7816 8128 7832 8192
rect 7896 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8064 8192
rect 7744 7774 8064 8128
rect 7744 7538 7786 7774
rect 8022 7538 8064 7774
rect 7744 7104 8064 7538
rect 7744 7040 7752 7104
rect 7816 7040 7832 7104
rect 7896 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8064 7104
rect 7744 6454 8064 7040
rect 7744 6218 7786 6454
rect 8022 6218 8064 6454
rect 7744 6016 8064 6218
rect 7744 5952 7752 6016
rect 7816 5952 7832 6016
rect 7896 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8064 6016
rect 7744 5134 8064 5952
rect 7744 4928 7786 5134
rect 8022 4928 8064 5134
rect 7744 4864 7752 4928
rect 7816 4864 7832 4898
rect 7896 4864 7912 4898
rect 7976 4864 7992 4898
rect 8056 4864 8064 4928
rect 7744 3840 8064 4864
rect 7744 3776 7752 3840
rect 7816 3814 7832 3840
rect 7896 3814 7912 3840
rect 7976 3814 7992 3840
rect 8056 3776 8064 3840
rect 7744 3578 7786 3776
rect 8022 3578 8064 3776
rect 7744 2752 8064 3578
rect 7744 2688 7752 2752
rect 7816 2688 7832 2752
rect 7896 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8064 2752
rect 8404 9824 8724 9840
rect 8404 9760 8412 9824
rect 8476 9760 8492 9824
rect 8556 9760 8572 9824
rect 8636 9760 8652 9824
rect 8716 9760 8724 9824
rect 8404 9754 8724 9760
rect 8404 9518 8446 9754
rect 8682 9518 8724 9754
rect 8404 8736 8724 9518
rect 8404 8672 8412 8736
rect 8476 8672 8492 8736
rect 8556 8672 8572 8736
rect 8636 8672 8652 8736
rect 8716 8672 8724 8736
rect 8404 8434 8724 8672
rect 8404 8198 8446 8434
rect 8682 8198 8724 8434
rect 8404 7648 8724 8198
rect 8404 7584 8412 7648
rect 8476 7584 8492 7648
rect 8556 7584 8572 7648
rect 8636 7584 8652 7648
rect 8716 7584 8724 7648
rect 8404 7114 8724 7584
rect 8404 6878 8446 7114
rect 8682 6878 8724 7114
rect 8404 6560 8724 6878
rect 8404 6496 8412 6560
rect 8476 6496 8492 6560
rect 8556 6496 8572 6560
rect 8636 6496 8652 6560
rect 8716 6496 8724 6560
rect 8404 5794 8724 6496
rect 8404 5558 8446 5794
rect 8682 5558 8724 5794
rect 8404 5472 8724 5558
rect 8404 5408 8412 5472
rect 8476 5408 8492 5472
rect 8556 5408 8572 5472
rect 8636 5408 8652 5472
rect 8716 5408 8724 5472
rect 8404 4474 8724 5408
rect 8404 4384 8446 4474
rect 8682 4384 8724 4474
rect 8404 4320 8412 4384
rect 8716 4320 8724 4384
rect 8404 4238 8446 4320
rect 8682 4238 8724 4320
rect 8404 3296 8724 4238
rect 8404 3232 8412 3296
rect 8476 3232 8492 3296
rect 8556 3232 8572 3296
rect 8636 3232 8652 3296
rect 8716 3232 8724 3296
rect 8404 3154 8724 3232
rect 8404 2918 8446 3154
rect 8682 2918 8724 3154
rect 7744 2494 8070 2688
rect 7744 2258 7786 2494
rect 8022 2258 8070 2494
rect 7744 2128 8070 2258
rect 8404 2208 8724 2918
rect 8404 2144 8412 2208
rect 8476 2144 8492 2208
rect 8556 2144 8572 2208
rect 8636 2144 8652 2208
rect 8716 2144 8724 2208
rect 8404 2128 8724 2144
rect 1142 2066 1458 2128
rect 2462 2066 2778 2128
rect 3782 2066 4098 2128
rect 5104 2066 5420 2128
rect 6412 2066 6728 2128
rect 7754 2066 8070 2128
rect 1134 2018 8070 2066
rect 1134 1820 1358 2018
rect 7744 1820 8070 2018
rect 1134 1750 8070 1820
<< via4 >>
rect 1186 8858 1422 9094
rect 1186 7538 1422 7774
rect 1186 6218 1422 6454
rect 1186 4928 1422 5134
rect 1186 4898 1216 4928
rect 1216 4898 1232 4928
rect 1232 4898 1296 4928
rect 1296 4898 1312 4928
rect 1312 4898 1376 4928
rect 1376 4898 1392 4928
rect 1392 4898 1422 4928
rect 1186 3776 1216 3814
rect 1216 3776 1232 3814
rect 1232 3776 1296 3814
rect 1296 3776 1312 3814
rect 1312 3776 1376 3814
rect 1376 3776 1392 3814
rect 1392 3776 1422 3814
rect 1186 3578 1422 3776
rect 1186 2258 1422 2494
rect 1846 9518 2082 9754
rect 1846 8198 2082 8434
rect 1846 6878 2082 7114
rect 1846 5558 2082 5794
rect 1846 4384 2082 4474
rect 1846 4320 1876 4384
rect 1876 4320 1892 4384
rect 1892 4320 1956 4384
rect 1956 4320 1972 4384
rect 1972 4320 2036 4384
rect 2036 4320 2052 4384
rect 2052 4320 2082 4384
rect 1846 4238 2082 4320
rect 1846 2918 2082 3154
rect 2506 8858 2742 9094
rect 2506 7538 2742 7774
rect 2506 6218 2742 6454
rect 2506 4928 2742 5134
rect 2506 4898 2536 4928
rect 2536 4898 2552 4928
rect 2552 4898 2616 4928
rect 2616 4898 2632 4928
rect 2632 4898 2696 4928
rect 2696 4898 2712 4928
rect 2712 4898 2742 4928
rect 2506 3776 2536 3814
rect 2536 3776 2552 3814
rect 2552 3776 2616 3814
rect 2616 3776 2632 3814
rect 2632 3776 2696 3814
rect 2696 3776 2712 3814
rect 2712 3776 2742 3814
rect 2506 3578 2742 3776
rect 2506 2258 2742 2494
rect 3166 9518 3402 9754
rect 3166 8198 3402 8434
rect 3166 6878 3402 7114
rect 3166 5558 3402 5794
rect 3166 4384 3402 4474
rect 3166 4320 3196 4384
rect 3196 4320 3212 4384
rect 3212 4320 3276 4384
rect 3276 4320 3292 4384
rect 3292 4320 3356 4384
rect 3356 4320 3372 4384
rect 3372 4320 3402 4384
rect 3166 4238 3402 4320
rect 3166 2918 3402 3154
rect 3826 8858 4062 9094
rect 3826 7538 4062 7774
rect 3826 6218 4062 6454
rect 3826 4928 4062 5134
rect 3826 4898 3856 4928
rect 3856 4898 3872 4928
rect 3872 4898 3936 4928
rect 3936 4898 3952 4928
rect 3952 4898 4016 4928
rect 4016 4898 4032 4928
rect 4032 4898 4062 4928
rect 3826 3776 3856 3814
rect 3856 3776 3872 3814
rect 3872 3776 3936 3814
rect 3936 3776 3952 3814
rect 3952 3776 4016 3814
rect 4016 3776 4032 3814
rect 4032 3776 4062 3814
rect 3826 3578 4062 3776
rect 3826 2258 4062 2494
rect 4486 9518 4722 9754
rect 4486 8198 4722 8434
rect 4486 6878 4722 7114
rect 4486 5558 4722 5794
rect 4486 4384 4722 4474
rect 4486 4320 4516 4384
rect 4516 4320 4532 4384
rect 4532 4320 4596 4384
rect 4596 4320 4612 4384
rect 4612 4320 4676 4384
rect 4676 4320 4692 4384
rect 4692 4320 4722 4384
rect 4486 4238 4722 4320
rect 4486 2918 4722 3154
rect 5146 8858 5382 9094
rect 5146 7538 5382 7774
rect 5146 6218 5382 6454
rect 5146 4928 5382 5134
rect 5146 4898 5176 4928
rect 5176 4898 5192 4928
rect 5192 4898 5256 4928
rect 5256 4898 5272 4928
rect 5272 4898 5336 4928
rect 5336 4898 5352 4928
rect 5352 4898 5382 4928
rect 5146 3776 5176 3814
rect 5176 3776 5192 3814
rect 5192 3776 5256 3814
rect 5256 3776 5272 3814
rect 5272 3776 5336 3814
rect 5336 3776 5352 3814
rect 5352 3776 5382 3814
rect 5146 3578 5382 3776
rect 5146 2258 5382 2494
rect 5806 9518 6042 9754
rect 5806 8198 6042 8434
rect 5806 6878 6042 7114
rect 5806 5558 6042 5794
rect 5806 4384 6042 4474
rect 5806 4320 5836 4384
rect 5836 4320 5852 4384
rect 5852 4320 5916 4384
rect 5916 4320 5932 4384
rect 5932 4320 5996 4384
rect 5996 4320 6012 4384
rect 6012 4320 6042 4384
rect 5806 4238 6042 4320
rect 5806 2918 6042 3154
rect 6466 8858 6702 9094
rect 6466 7538 6702 7774
rect 6466 6218 6702 6454
rect 6466 4928 6702 5134
rect 6466 4898 6496 4928
rect 6496 4898 6512 4928
rect 6512 4898 6576 4928
rect 6576 4898 6592 4928
rect 6592 4898 6656 4928
rect 6656 4898 6672 4928
rect 6672 4898 6702 4928
rect 6466 3776 6496 3814
rect 6496 3776 6512 3814
rect 6512 3776 6576 3814
rect 6576 3776 6592 3814
rect 6592 3776 6656 3814
rect 6656 3776 6672 3814
rect 6672 3776 6702 3814
rect 6466 3578 6702 3776
rect 6466 2258 6702 2494
rect 7126 9518 7362 9754
rect 7126 8198 7362 8434
rect 7126 6878 7362 7114
rect 7126 5558 7362 5794
rect 7126 4384 7362 4474
rect 7126 4320 7156 4384
rect 7156 4320 7172 4384
rect 7172 4320 7236 4384
rect 7236 4320 7252 4384
rect 7252 4320 7316 4384
rect 7316 4320 7332 4384
rect 7332 4320 7362 4384
rect 7126 4238 7362 4320
rect 7126 2918 7362 3154
rect 7786 8858 8022 9094
rect 7786 7538 8022 7774
rect 7786 6218 8022 6454
rect 7786 4928 8022 5134
rect 7786 4898 7816 4928
rect 7816 4898 7832 4928
rect 7832 4898 7896 4928
rect 7896 4898 7912 4928
rect 7912 4898 7976 4928
rect 7976 4898 7992 4928
rect 7992 4898 8022 4928
rect 7786 3776 7816 3814
rect 7816 3776 7832 3814
rect 7832 3776 7896 3814
rect 7896 3776 7912 3814
rect 7912 3776 7976 3814
rect 7976 3776 7992 3814
rect 7992 3776 8022 3814
rect 7786 3578 8022 3776
rect 8446 9518 8682 9754
rect 8446 8198 8682 8434
rect 8446 6878 8682 7114
rect 8446 5558 8682 5794
rect 8446 4384 8682 4474
rect 8446 4320 8476 4384
rect 8476 4320 8492 4384
rect 8492 4320 8556 4384
rect 8556 4320 8572 4384
rect 8572 4320 8636 4384
rect 8636 4320 8652 4384
rect 8652 4320 8682 4384
rect 8446 4238 8682 4320
rect 8446 2918 8682 3154
rect 7786 2258 8022 2494
<< metal5 >>
rect 1056 9754 8788 9796
rect 1056 9518 1846 9754
rect 2082 9518 3166 9754
rect 3402 9518 4486 9754
rect 4722 9518 5806 9754
rect 6042 9518 7126 9754
rect 7362 9518 8446 9754
rect 8682 9518 8788 9754
rect 1056 9476 8788 9518
rect 1056 9094 8788 9136
rect 1056 8858 1186 9094
rect 1422 8858 2506 9094
rect 2742 8858 3826 9094
rect 4062 8858 5146 9094
rect 5382 8858 6466 9094
rect 6702 8858 7786 9094
rect 8022 8858 8788 9094
rect 1056 8816 8788 8858
rect 1056 8434 8788 8476
rect 1056 8198 1846 8434
rect 2082 8198 3166 8434
rect 3402 8198 4486 8434
rect 4722 8198 5806 8434
rect 6042 8198 7126 8434
rect 7362 8198 8446 8434
rect 8682 8198 8788 8434
rect 1056 8156 8788 8198
rect 1056 7774 8788 7816
rect 1056 7538 1186 7774
rect 1422 7538 2506 7774
rect 2742 7538 3826 7774
rect 4062 7538 5146 7774
rect 5382 7538 6466 7774
rect 6702 7538 7786 7774
rect 8022 7538 8788 7774
rect 1056 7496 8788 7538
rect 1056 7114 8788 7156
rect 1056 6878 1846 7114
rect 2082 6878 3166 7114
rect 3402 6878 4486 7114
rect 4722 6878 5806 7114
rect 6042 6878 7126 7114
rect 7362 6878 8446 7114
rect 8682 6878 8788 7114
rect 1056 6836 8788 6878
rect 1056 6454 8788 6496
rect 1056 6218 1186 6454
rect 1422 6218 2506 6454
rect 2742 6218 3826 6454
rect 4062 6218 5146 6454
rect 5382 6218 6466 6454
rect 6702 6218 7786 6454
rect 8022 6218 8788 6454
rect 1056 6176 8788 6218
rect 1056 5794 8788 5836
rect 1056 5558 1846 5794
rect 2082 5558 3166 5794
rect 3402 5558 4486 5794
rect 4722 5558 5806 5794
rect 6042 5558 7126 5794
rect 7362 5558 8446 5794
rect 8682 5558 8788 5794
rect 1056 5516 8788 5558
rect 1056 5134 8788 5176
rect 1056 4898 1186 5134
rect 1422 4898 2506 5134
rect 2742 4898 3826 5134
rect 4062 4898 5146 5134
rect 5382 4898 6466 5134
rect 6702 4898 7786 5134
rect 8022 4898 8788 5134
rect 1056 4856 8788 4898
rect 1056 4474 8788 4516
rect 1056 4238 1846 4474
rect 2082 4238 3166 4474
rect 3402 4238 4486 4474
rect 4722 4238 5806 4474
rect 6042 4238 7126 4474
rect 7362 4238 8446 4474
rect 8682 4238 8788 4474
rect 1056 4196 8788 4238
rect 1056 3814 8788 3856
rect 1056 3578 1186 3814
rect 1422 3578 2506 3814
rect 2742 3578 3826 3814
rect 4062 3578 5146 3814
rect 5382 3578 6466 3814
rect 6702 3578 7786 3814
rect 8022 3578 8788 3814
rect 1056 3536 8788 3578
rect 1056 3154 8788 3196
rect 1056 2918 1846 3154
rect 2082 2918 3166 3154
rect 3402 2918 4486 3154
rect 4722 2918 5806 3154
rect 6042 2918 7126 3154
rect 7362 2918 8446 3154
rect 8682 2918 8788 3154
rect 1056 2876 8788 2918
rect 1056 2494 8788 2536
rect 1056 2258 1186 2494
rect 1422 2258 2506 2494
rect 2742 2258 3826 2494
rect 4062 2258 5146 2494
rect 5382 2258 6466 2494
rect 6702 2258 7786 2494
rect 8022 2258 8788 2494
rect 1056 2216 8788 2258
use sky130_fd_sc_hd__xor2_1  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1840 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2208 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _29_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _31_
timestamp 1704896540
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3588 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _33_
timestamp 1704896540
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _34_
timestamp 1704896540
transform 1 0 3772 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _35_
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2392 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _37_
timestamp 1704896540
transform -1 0 3772 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4140 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _42_
timestamp 1704896540
transform -1 0 5152 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _43_
timestamp 1704896540
transform 1 0 4232 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _44_
timestamp 1704896540
transform -1 0 4968 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _45_
timestamp 1704896540
transform -1 0 6164 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _46_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _47_
timestamp 1704896540
transform -1 0 6992 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _48_
timestamp 1704896540
transform -1 0 7636 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _49_
timestamp 1704896540
transform 1 0 6992 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1704896540
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _51_
timestamp 1704896540
transform -1 0 8280 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _52_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3312 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _53_
timestamp 1704896540
transform -1 0 3312 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _54_
timestamp 1704896540
transform 1 0 1656 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _55_
timestamp 1704896540
transform 1 0 1932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _56_
timestamp 1704896540
transform 1 0 2208 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _57_
timestamp 1704896540
transform -1 0 5796 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _58_
timestamp 1704896540
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _59_
timestamp 1704896540
transform 1 0 5152 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _60_
timestamp 1704896540
transform 1 0 6624 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _61_
timestamp 1704896540
transform 1 0 6624 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6072 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 3588 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 5704 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_16
timestamp 1704896540
transform 1 0 2576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_36
timestamp 1704896540
transform 1 0 4416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_40
timestamp 1704896540
transform 1 0 4784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_46
timestamp 1704896540
transform 1 0 5336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50
timestamp 1704896540
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_60
timestamp 1704896540
transform 1 0 6624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_66
timestamp 1704896540
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_70
timestamp 1704896540
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_46
timestamp 1704896540
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_78
timestamp 1704896540
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25
timestamp 1704896540
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_76
timestamp 1704896540
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_29
timestamp 1704896540
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_76
timestamp 1704896540
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_33
timestamp 1704896540
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_70
timestamp 1704896540
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_78
timestamp 1704896540
transform 1 0 8280 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_73
timestamp 1704896540
transform 1 0 7820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_79
timestamp 1704896540
transform 1 0 8372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_33
timestamp 1704896540
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_54
timestamp 1704896540
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_66
timestamp 1704896540
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_78
timestamp 1704896540
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_77
timestamp 1704896540
transform 1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_11
timestamp 1704896540
transform 1 0 2116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_24
timestamp 1704896540
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_77
timestamp 1704896540
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_24
timestamp 1704896540
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_36
timestamp 1704896540
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 1704896540
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_69
timestamp 1704896540
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_77
timestamp 1704896540
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 1704896540
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_24
timestamp 1704896540
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_77
timestamp 1704896540
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_7
timestamp 1704896540
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_77
timestamp 1704896540
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_77
timestamp 1704896540
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_18
timestamp 1704896540
transform 1 0 2760 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 1704896540
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_29
timestamp 1704896540
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1704896540
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1704896540
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_69
timestamp 1704896540
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_77
timestamp 1704896540
transform 1 0 8188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output2
timestamp 1704896540
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output3
timestamp 1704896540
transform -1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output4
timestamp 1704896540
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1704896540
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output6
timestamp 1704896540
transform -1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1704896540
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1704896540
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1704896540
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output10
timestamp 1704896540
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output11
timestamp 1704896540
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_14
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_15
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_16
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 8740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_17
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_18
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 8740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_19
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_20
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 8740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_21
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_22
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 8740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_23
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 8740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_24
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 8740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_25
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_26
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 8740 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_27
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_32
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_33
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_34
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_35
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_36
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_37
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_38
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_39
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_40
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_41
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_42
timestamp 1704896540
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_43
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
<< labels >>
rlabel metal1 s 4922 9792 4922 9792 4 VGND
rlabel metal1 s 4922 9248 4922 9248 4 VPWR
rlabel metal2 s 2898 8058 2898 8058 4 _00_
rlabel metal1 s 3036 6970 3036 6970 4 _01_
rlabel metal1 s 1876 4114 1876 4114 4 _02_
rlabel metal2 s 2438 3298 2438 3298 4 _03_
rlabel metal1 s 3128 4046 3128 4046 4 _04_
rlabel metal1 s 5673 5270 5673 5270 4 _05_
rlabel metal1 s 4998 4182 4998 4182 4 _06_
rlabel metal1 s 5561 3434 5561 3434 4 _07_
rlabel metal1 s 7263 4182 7263 4182 4 _08_
rlabel metal2 s 7682 3196 7682 3196 4 _09_
rlabel metal1 s 2622 6664 2622 6664 4 _10_
rlabel metal1 s 1978 4556 1978 4556 4 _11_
rlabel metal2 s 3082 7140 3082 7140 4 _12_
rlabel metal2 s 1426 4284 1426 4284 4 _13_
rlabel metal2 s 1610 3604 1610 3604 4 _14_
rlabel metal1 s 6762 3162 6762 3162 4 _15_
rlabel metal1 s 2691 3026 2691 3026 4 _16_
rlabel metal2 s 4462 4794 4462 4794 4 _17_
rlabel metal2 s 4186 4556 4186 4556 4 _18_
rlabel metal1 s 5152 5202 5152 5202 4 _19_
rlabel metal1 s 4501 3468 4501 3468 4 _20_
rlabel metal1 s 4784 4590 4784 4590 4 _21_
rlabel metal2 s 5566 3808 5566 3808 4 _22_
rlabel metal1 s 6716 2822 6716 2822 4 _23_
rlabel metal1 s 7544 3162 7544 3162 4 _24_
rlabel metal1 s 7636 5202 7636 5202 4 _25_
rlabel metal1 s 6440 5678 6440 5678 4 clk
rlabel metal1 s 5106 5542 5106 5542 4 clknet_0_clk
rlabel metal2 s 2254 5270 2254 5270 4 clknet_1_0__leaf_clk
rlabel metal2 s 6670 4284 6670 4284 4 clknet_1_1__leaf_clk
rlabel metal1 s 2576 9554 2576 9554 4 enable
rlabel metal1 s 2308 6630 2308 6630 4 net1
rlabel metal1 s 8372 2414 8372 2414 4 net10
rlabel metal1 s 8050 2414 8050 2414 4 net11
rlabel metal1 s 1886 6698 1886 6698 4 net2
rlabel metal1 s 1840 2414 1840 2414 4 net3
rlabel metal1 s 2944 2414 2944 2414 4 net4
rlabel metal1 s 3864 2414 3864 2414 4 net5
rlabel metal1 s 6118 2856 6118 2856 4 net6
rlabel metal1 s 5474 5338 5474 5338 4 net7
rlabel metal1 s 6210 2414 6210 2414 4 net8
rlabel metal1 s 7544 2414 7544 2414 4 net9
flabel metal5 s 1056 9476 8788 9796 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8156 8788 8476 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6836 8788 7156 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 5516 8788 5836 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4196 8788 4516 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 2876 8788 3196 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 8404 2128 8724 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7084 2128 7404 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5764 2128 6084 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4444 2128 4764 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3124 2128 3444 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1804 2128 2124 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8816 8788 9136 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 7496 8788 7816 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 6176 8788 6496 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4856 8788 5176 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3536 8788 3856 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 2216 8788 2536 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 7744 2128 8064 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 6424 2128 6744 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5104 2128 5424 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3784 2128 4104 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2464 2128 2784 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1144 2128 1464 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 2410 10086 2466 10886 0 FreeSans 280 90 0 0 enable
port 4 nsew
flabel metal2 s 6918 9990 6974 10790 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 9034 982 9090 1782 0 FreeSans 280 90 0 0 counter[9]
port 14 nsew
flabel metal2 s 8114 982 8170 1782 0 FreeSans 280 90 0 0 counter[8]
port 13 nsew
flabel metal2 s 7194 982 7250 1782 0 FreeSans 280 90 0 0 counter[7]
port 12 nsew
flabel metal2 s 6274 982 6330 1782 0 FreeSans 280 90 0 0 counter[6]
port 11 nsew
flabel metal2 s 5354 982 5410 1782 0 FreeSans 280 90 0 0 counter[5]
port 10 nsew
flabel metal2 s 4434 982 4490 1782 0 FreeSans 280 90 0 0 counter[4]
port 9 nsew
flabel metal2 s 3514 982 3570 1782 0 FreeSans 280 90 0 0 counter[3]
port 8 nsew
flabel metal2 s 2594 982 2650 1782 0 FreeSans 280 90 0 0 counter[2]
port 7 nsew
flabel metal2 s 1674 982 1730 1782 0 FreeSans 280 90 0 0 counter[1]
port 6 nsew
flabel metal2 s 754 982 810 1782 0 FreeSans 280 90 0 0 counter[0]
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 9882 12026
string GDS_END 320138
<< end >>
