* NGSPICE file created from sky130_fd_sc_hd__inv_2_parax.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y.t2 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND.t1 A.t1 Y.t0 VNB.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y.t3 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR.t0 A.t3 Y.t1 VPB.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R0 A.n0 A.t3 212.081
R1 A.n1 A.t0 212.081
R2 A A.n1 189.073
R3 A.n0 A.t1 139.78
R4 A.n1 A.t2 139.78
R5 A.n1 A.n0 61.346
R6 VPWR.n0 VPWR.t0 262.851
R7 VPWR.n0 VPWR.t1 259.721
R8 VPWR VPWR.n0 0.491471
R9 Y.n2 Y.n1 208.965
R10 Y Y.n0 96.8352
R11 Y.n1 Y.t1 26.5955
R12 Y.n1 Y.t2 26.5955
R13 Y.n0 Y.t0 24.9236
R14 Y.n0 Y.t3 24.9236
R15 Y.n3 Y 11.2645
R16 Y Y.n3 6.1445
R17 Y.n3 Y 4.65505
R18 Y Y.n2 2.0485
R19 Y.n2 Y 1.55202
R20 VPB.t1 VPB.t0 248.599
R21 VPB VPB.t1 198.287
R22 VGND.n0 VGND.t1 169.418
R23 VGND.n0 VGND.t0 166.787
R24 VGND VGND.n0 0.491471
R25 VNB.t0 VNB.t1 1196.12
R26 VNB VNB.t0 954.045
C0 VGND Y 0.154601f
C1 VPB Y 0.006097f
C2 A VPWR 0.06305f
C3 VGND VPB 0.006491f
C4 VPWR Y 0.209105f
C5 A Y 0.089386f
C6 VPWR VGND 0.042274f
C7 A VGND 0.063754f
C8 VPWR VPB 0.052063f
C9 A VPB 0.074183f
C10 VGND VNB 0.266187f
C11 Y VNB 0.03316f
C12 VPWR VNB 0.246044f
C13 A VNB 0.262807f
C14 VPB VNB 0.338976f
.ends

