magic
tech sky130A
magscale 1 2
timestamp 1728255086
<< viali >>
rect 11962 -236 12230 -190
rect 13048 -232 13316 -186
rect 14108 -236 14376 -190
rect 15156 -230 15424 -184
<< metal1 >>
rect 11442 4474 11642 4674
rect 11670 4610 11870 4674
rect 11670 4520 11702 4610
rect 11814 4520 11870 4610
rect 11670 4474 11870 4520
rect 11908 4478 12108 4678
rect 12224 4606 12424 4674
rect 12224 4516 12248 4606
rect 12388 4516 12424 4606
rect 11488 4222 11610 4474
rect 11910 4382 11996 4478
rect 12224 4474 12424 4516
rect 12498 4472 12698 4672
rect 12730 4616 12930 4674
rect 12730 4518 12774 4616
rect 12868 4518 12930 4616
rect 12730 4474 12930 4518
rect 12964 4476 13164 4676
rect 11824 4314 11996 4382
rect 11910 4246 11996 4314
rect 12562 4220 12694 4472
rect 12964 4388 13042 4476
rect 13542 4468 13742 4668
rect 13776 4614 13976 4670
rect 13776 4516 13836 4614
rect 13940 4516 13976 4614
rect 13776 4470 13976 4516
rect 14010 4470 14210 4670
rect 14572 4482 14772 4682
rect 14800 4642 15000 4682
rect 14800 4532 14884 4642
rect 14978 4532 15000 4642
rect 14800 4482 15000 4532
rect 15044 4482 15244 4682
rect 12900 4310 13042 4388
rect 12964 4246 13042 4310
rect 13594 4214 13740 4468
rect 14036 4380 14124 4470
rect 13956 4254 14124 4380
rect 14036 4238 14124 4254
rect 14620 4194 14772 4482
rect 15046 4246 15170 4482
rect 11456 4004 11466 4094
rect 11560 4004 11570 4094
rect 11684 3980 11694 4070
rect 11806 3980 11816 4070
rect 12532 4000 12542 4090
rect 12636 4000 12646 4090
rect 12762 4000 12772 4098
rect 12866 4000 12876 4098
rect 13604 3994 13614 4084
rect 13708 3994 13718 4084
rect 13826 3992 13836 4090
rect 13940 3992 13950 4090
rect 14676 4000 14686 4090
rect 14780 4000 14790 4090
rect 14864 3952 14874 4118
rect 15012 3952 15022 4118
rect 11414 -262 11614 -62
rect 11678 -156 11688 -48
rect 11658 -192 11688 -156
rect 11844 -156 11854 -48
rect 11844 -192 11858 -156
rect 11658 -356 11858 -192
rect 11918 -242 11928 -178
rect 12266 -242 12276 -178
rect 12482 -258 12682 -58
rect 12744 -184 12754 -40
rect 12910 -184 12920 -40
rect 12996 -238 13006 -174
rect 13344 -238 13354 -174
rect 13552 -294 13752 -94
rect 13812 -190 13822 -46
rect 13978 -190 13988 -46
rect 14066 -246 14076 -182
rect 14414 -246 14424 -182
rect 14610 -296 14810 -130
rect 14862 -192 14872 -48
rect 15028 -192 15038 -48
rect 15102 -238 15112 -174
rect 15450 -238 15460 -174
<< via1 >>
rect 11702 4520 11814 4610
rect 12248 4516 12388 4606
rect 12774 4518 12868 4616
rect 13836 4516 13940 4614
rect 14884 4532 14978 4642
rect 11466 4004 11560 4094
rect 11694 3980 11806 4070
rect 12542 4000 12636 4090
rect 12772 4000 12866 4098
rect 13614 3994 13708 4084
rect 13836 3992 13940 4090
rect 14686 4000 14780 4090
rect 14874 3952 15012 4118
rect 11688 -192 11844 -48
rect 11928 -190 12266 -178
rect 11928 -236 11962 -190
rect 11962 -236 12230 -190
rect 12230 -236 12266 -190
rect 11928 -242 12266 -236
rect 12754 -184 12910 -40
rect 13006 -186 13344 -174
rect 13006 -232 13048 -186
rect 13048 -232 13316 -186
rect 13316 -232 13344 -186
rect 13006 -238 13344 -232
rect 13822 -190 13978 -46
rect 14076 -190 14414 -182
rect 14076 -236 14108 -190
rect 14108 -236 14376 -190
rect 14376 -236 14414 -190
rect 14076 -246 14414 -236
rect 14872 -192 15028 -48
rect 15112 -184 15450 -174
rect 15112 -230 15156 -184
rect 15156 -230 15424 -184
rect 15424 -230 15450 -184
rect 15112 -238 15450 -230
<< metal2 >>
rect 14884 4642 14978 4652
rect 11702 4610 11814 4620
rect 12774 4616 12868 4626
rect 11702 4510 11814 4520
rect 12248 4606 12388 4616
rect 12248 4506 12388 4516
rect 12774 4508 12868 4518
rect 13836 4614 13940 4624
rect 14884 4522 14978 4532
rect 13836 4506 13940 4516
rect 14874 4118 15012 4128
rect 11466 4094 11560 4104
rect 12542 4090 12636 4100
rect 11466 3994 11560 4004
rect 11694 4070 11806 4080
rect 12542 3990 12636 4000
rect 12772 4098 12866 4108
rect 12772 3990 12866 4000
rect 13614 4084 13708 4094
rect 13614 3984 13708 3994
rect 13836 4090 13940 4100
rect 13836 3982 13940 3992
rect 14686 4090 14780 4100
rect 14686 3990 14780 4000
rect 11694 3970 11806 3980
rect 14874 3942 15012 3952
rect 11658 -8 15056 -2
rect 11658 -40 15058 -8
rect 11658 -48 12754 -40
rect 11658 -158 11688 -48
rect 11844 -158 12754 -48
rect 11688 -202 11844 -192
rect 11904 -178 12292 -158
rect 11904 -242 11928 -178
rect 12266 -242 12292 -178
rect 12910 -46 15058 -40
rect 12910 -158 13822 -46
rect 12754 -194 12910 -184
rect 12972 -174 13360 -158
rect 11904 -246 12292 -242
rect 12972 -238 13006 -174
rect 13344 -238 13360 -174
rect 13978 -48 15058 -46
rect 13978 -158 14872 -48
rect 13822 -200 13978 -190
rect 14046 -182 14434 -158
rect 12972 -246 13360 -238
rect 14046 -246 14076 -182
rect 14414 -246 14434 -182
rect 15028 -156 15058 -48
rect 15028 -174 15490 -156
rect 15028 -192 15112 -174
rect 14872 -202 15112 -192
rect 15026 -238 15112 -202
rect 15450 -238 15490 -174
rect 15026 -246 15490 -238
rect 11928 -252 12266 -246
rect 13006 -248 13344 -246
rect 14046 -250 14434 -246
rect 15112 -248 15450 -246
rect 14076 -256 14414 -250
<< via2 >>
rect 11702 4520 11814 4610
rect 12248 4516 12388 4606
rect 12774 4518 12868 4616
rect 13836 4516 13940 4614
rect 14884 4532 14978 4642
rect 11466 4004 11560 4094
rect 11694 3980 11806 4070
rect 12542 4000 12636 4090
rect 12772 4000 12866 4098
rect 13614 3994 13708 4084
rect 13836 3992 13940 4090
rect 14686 4000 14780 4090
rect 14876 3984 14980 4104
<< metal3 >>
rect 14874 4644 14988 4647
rect 14870 4642 14990 4644
rect 12764 4616 12878 4621
rect 13834 4619 13942 4622
rect 11692 4610 11824 4615
rect 11692 4520 11702 4610
rect 11814 4520 11824 4610
rect 11692 4515 11824 4520
rect 12238 4606 12398 4611
rect 12238 4516 12248 4606
rect 12388 4532 12398 4606
rect 12388 4516 12414 4532
rect 11456 4094 11570 4099
rect 11456 4004 11466 4094
rect 11560 4004 11570 4094
rect 11700 4075 11790 4515
rect 12238 4511 12414 4516
rect 12764 4518 12774 4616
rect 12868 4518 12878 4616
rect 12764 4513 12878 4518
rect 13826 4614 13950 4619
rect 13826 4516 13836 4614
rect 13940 4516 13950 4614
rect 11456 3999 11570 4004
rect 11684 4070 11816 4075
rect 11464 3898 11562 3999
rect 11684 3980 11694 4070
rect 11806 3980 11816 4070
rect 11684 3975 11816 3980
rect 11700 3958 11790 3975
rect 12244 3898 12414 4511
rect 12772 4103 12872 4513
rect 13826 4511 13950 4516
rect 14870 4532 14884 4642
rect 14978 4532 14990 4642
rect 12762 4098 12876 4103
rect 12532 4090 12646 4095
rect 12532 4000 12542 4090
rect 12636 4000 12646 4090
rect 12532 3995 12646 4000
rect 12762 4000 12772 4098
rect 12866 4000 12876 4098
rect 13834 4095 13942 4511
rect 14870 4109 14990 4532
rect 14866 4104 14990 4109
rect 13826 4090 13950 4095
rect 13612 4089 13710 4090
rect 12762 3995 12876 4000
rect 13604 4084 13718 4089
rect 12540 3898 12638 3995
rect 12772 3970 12872 3995
rect 13604 3994 13614 4084
rect 13708 3994 13718 4084
rect 13604 3989 13718 3994
rect 13826 3992 13836 4090
rect 13940 3992 13950 4090
rect 14676 4090 14790 4095
rect 14676 4000 14686 4090
rect 14780 4000 14790 4090
rect 14676 3995 14790 4000
rect 13612 3898 13710 3989
rect 13826 3987 13950 3992
rect 13834 3974 13942 3987
rect 14682 3898 14780 3995
rect 14866 3984 14876 4104
rect 14980 3984 14990 4104
rect 14866 3979 14990 3984
rect 14870 3954 14990 3979
rect 11428 3790 14794 3898
use passgate  x1
timestamp 1725640011
transform 0 1 12256 -1 0 7822
box 3356 -890 8072 137
use passgate  x2
timestamp 1725640011
transform 0 1 13326 -1 0 7824
box 3356 -890 8072 137
use passgate  x3
timestamp 1725640011
transform 0 1 14396 -1 0 7818
box 3356 -890 8072 137
use passgate  x4
timestamp 1725640011
transform 0 1 15452 -1 0 7826
box 3356 -890 8072 137
<< labels >>
flabel metal1 11442 4474 11642 4674 0 FreeSans 256 0 0 0 A1
port 0 nsew
flabel metal1 11670 4474 11870 4674 0 FreeSans 256 0 0 0 GN1
port 1 nsew
flabel metal1 11908 4478 12108 4678 0 FreeSans 256 0 0 0 GP1
port 2 nsew
flabel metal1 11414 -262 11614 -62 0 FreeSans 256 0 0 0 Z1
port 3 nsew
flabel metal1 12498 4472 12698 4672 0 FreeSans 256 0 0 0 A2
port 4 nsew
flabel metal1 12730 4474 12930 4674 0 FreeSans 256 0 0 0 GN2
port 5 nsew
flabel metal1 12964 4476 13164 4676 0 FreeSans 256 0 0 0 GP2
port 6 nsew
flabel metal1 12482 -258 12682 -58 0 FreeSans 256 0 0 0 Z2
port 7 nsew
flabel metal1 13542 4468 13742 4668 0 FreeSans 256 0 0 0 A3
port 8 nsew
flabel metal1 13776 4470 13976 4670 0 FreeSans 256 0 0 0 GN3
port 9 nsew
flabel metal1 14010 4470 14210 4670 0 FreeSans 256 0 0 0 GP3
port 10 nsew
flabel metal1 13552 -294 13752 -94 0 FreeSans 256 0 0 0 Z3
port 11 nsew
flabel metal1 14586 4502 14752 4664 0 FreeSans 640 0 0 0 A4
port 12 nsew
flabel metal1 14800 4482 15000 4682 0 FreeSans 256 0 0 0 GN4
port 13 nsew
flabel metal1 15044 4482 15244 4682 0 FreeSans 256 0 0 0 GP4
port 14 nsew
flabel metal1 14610 -296 14810 -130 0 FreeSans 640 0 0 0 Z4
port 15 nsew
flabel metal1 11658 -356 11858 -156 0 FreeSans 256 0 0 0 VDD
port 16 nsew
flabel metal1 12224 4474 12424 4674 0 FreeSans 256 0 0 0 VSS
port 17 nsew
<< end >>
