* NGSPICE file created from mux4onehot_b_parax.ext - technology: sky130A

.subckt mux4onehot_b_parax select1 select2 A1 A3 Z1 A2 A4 select0 Z4 Z3 VPWR Z2 VGND
+ nselect2
X0 A2.t1 x2.GP2.t4 Z2.t0 VPWR.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X1 VPWR.t5 a_5275_n4059# a_5275_n4235# VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X2 A1.t2 x2.GP1.t4 Z1.t2 VPWR.t53 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X3 VGND.t56 select0.t0 a_5275_n3507# VGND.t55 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X4 a_5275_n3683# a_5275_n3507# a_5301_n3555# VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X5 A4.t3 x2.GP4.t4 Z4.t2 VPWR.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X6 VGND.t17 select1.t0 x1.nSEL1 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X7 VGND.t32 x2.GN2 x2.GP2.t3 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X8 x1.nSEL0 select0.t1 VGND.t54 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X9 VGND.t27 a_5275_n4651# x2.GN1.t1 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X10 VPWR.t52 select0.t2 x1.nSEL0 VPWR.t51 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X11 x2.GP1.t0 x2.GN1.t2 VGND.t37 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X12 VGND.t43 x2.GN1.t3 x2.GP1.t1 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X13 x2.GP4.t0 x2.GN4.t2 VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X14 VPWR.t63 x2.GN4.t3 x2.GP4.t3 VPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X15 a_5275_n4059# select1.t1 VPWR.t18 VPWR.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X16 VGND.t11 VPWR.t71 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X17 a_5301_n4107# select0.t3 VGND.t52 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X18 VGND.t61 a_5275_n4235# x2.GN2 VGND.t60 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X19 a_5275_n4651# x1.nSEL1 VPWR.t14 VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X20 VGND.t8 VPWR.t72 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X21 a_5275_n3507# select0.t4 VPWR.t16 VPWR.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X22 a_5275_n4235# select0.t5 VPWR.t44 VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X23 VPWR.t42 x1.nSEL0 a_5275_n4651# VPWR.t41 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X24 VPWR.t50 a_5275_n3507# a_5275_n3683# VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X25 VPWR.t48 a_5275_n3683# x2.GN3 VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X26 VGND.t39 a_5275_n2995# x2.GN4.t1 VGND.t38 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X27 nselect2.t1 select2.t0 VPWR.t40 VPWR.t39 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X28 A3.t3 x2.GP3 Z3.t2 VPWR.t70 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X29 VGND.t50 select0.t6 x1.nSEL0 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X30 Z3.t0 x2.GN3 A3.t1 VGND.t25 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X31 Z3.t1 x2.GN3 A3.t0 VGND.t25 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X32 VPWR.t65 select2.t1 nselect2.t0 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X33 x2.GP4.t1 x2.GN4.t4 VGND.t45 VGND.t44 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X34 x2.GP3 x2.GN3 VPWR.t30 VPWR.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X35 x1.nSEL1 select1.t2 VPWR.t67 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X36 x2.GP2.t0 x2.GN2 VPWR.t36 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X37 VPWR.t12 VGND.t68 VPWR.t11 VPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X38 VGND.t65 x2.GN4.t5 x2.GP4.t2 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X39 VGND.t5 VPWR.t73 VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X40 a_5329_n4513# x1.nSEL1 VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X41 VPWR.t2 VGND.t69 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X42 a_5275_n4651# x1.nSEL0 a_5329_n4513# VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X43 A4.t2 x2.GP4.t5 Z4.t3 VPWR.t3 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X44 a_5275_n2995# select0.t7 VPWR.t21 VPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X45 VPWR.t28 x2.GN3 x2.GP3 VPWR.t27 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X46 VPWR.t32 a_5275_n4651# x2.GN1.t0 VPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X47 Z4.t1 x2.GN4.t6 A4.t1 VGND.t12 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X48 VGND.t2 VPWR.t74 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X49 Z4.t0 x2.GN4.t7 A4.t0 VGND.t12 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X50 VPWR.t7 select1.t3 a_5275_n2995# VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X51 a_5275_n3683# select1.t4 VPWR.t56 VPWR.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X52 nselect2.t3 select2.t2 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X53 a_5275_n4235# a_5275_n4059# a_5301_n4107# VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X54 VGND.t35 select2.t3 nselect2.t2 VGND.t34 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X55 x2.GP3 x2.GN3 VGND.t24 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X56 VPWR.t59 VGND.t70 VPWR.t58 VPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X57 A2.t0 x2.GP2.t5 Z2.t1 VPWR.t19 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X58 VPWR.t61 select1.t5 x1.nSEL1 VPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X59 x1.nSEL1 select1.t6 VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X60 x2.GP2.t2 x2.GN2 VGND.t30 VGND.t29 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X61 VPWR.t55 a_5275_n4235# x2.GN2 VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X62 Z2.t2 x2.GN2 A2.t3 VGND.t28 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X63 a_5329_n2857# select0.t8 VGND.t48 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X64 A1.t1 x2.GP1.t5 Z1.t1 VPWR.t53 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X65 Z2.t3 x2.GN2 A2.t2 VGND.t28 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X66 VPWR.t38 a_5275_n2995# x2.GN4.t0 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X67 VPWR.t24 VGND.t71 VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X68 VGND.t22 x2.GN3 x2.GP3 VGND.t21 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X69 VPWR.t34 x2.GN2 x2.GP2.t1 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X70 x1.nSEL0 select0.t9 VPWR.t26 VPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X71 Z1.t3 x2.GN1.t4 A1.t3 VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X72 x2.GP1.t2 x2.GN1.t5 VPWR.t46 VPWR.t45 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X73 Z1.t0 x2.GN1.t6 A1.t0 VGND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X74 a_5275_n2995# select1.t7 a_5329_n2857# VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X75 a_5301_n3555# select1.t8 VGND.t41 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X76 VGND.t58 a_5275_n3683# x2.GN3 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X77 VGND.t63 select1.t9 a_5275_n4059# VGND.t62 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X78 VPWR.t69 x2.GN1.t7 x2.GP1.t3 VPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X79 A3.t2 x2.GP3 Z3.t3 VPWR.t70 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
R0 x2.GP2.n4 x2.GP2.t4 450.938
R1 x2.GP2.n4 x2.GP2.t5 445.666
R2 x2.GP2.n5 x2.GP2.n3 195.958
R3 x2.GP2.n1 x2.GP2.n0 101.49
R4 x2.GP2.n3 x2.GP2.t1 26.5955
R5 x2.GP2.n3 x2.GP2.t0 26.5955
R6 x2.GP2.n0 x2.GP2.t3 24.9236
R7 x2.GP2.n0 x2.GP2.t2 24.9236
R8 x1.gpo1 x2.x2.GP 13.129
R9 x2.GP2.n5 x1.gpo1 11.995
R10 x2.GP2.n2 x1.x12.Y 10.7525
R11 x1.x12.Y x2.GP2.n5 7.96524
R12 x2.GP2.n2 x1.x12.Y 6.6565
R13 x1.x12.Y x2.GP2.n2 5.04292
R14 x2.x2.GP x2.GP2.n4 2.94361
R15 x1.x12.Y x2.GP2.n1 2.5605
R16 x2.GP2.n1 x1.x12.Y 1.93989
R17 Z2.n1 Z2.t1 23.6581
R18 Z2.n3 Z2.t0 23.3739
R19 Z2.n1 Z2.t2 10.7528
R20 Z2.n0 Z2.t3 10.6417
R21 Z2.n2 Z2.n1 1.30064
R22 Z2.n5 Z2.n4 0.936641
R23 Z2.n3 Z2.n2 0.726502
R24 Z2.n2 Z2.n0 0.512491
R25 Z2.n4 Z2.n0 0.359663
R26 Z2.n4 Z2.n3 0.216071
R27 Z2.n5 Z2 0.0776605
R28 Z2 Z2.n5 0.0561931
R29 A2.n1 A2.t1 26.3998
R30 A2.n1 A2.t0 23.5483
R31 A2.n0 A2.t2 12.7127
R32 A2.n0 A2.t3 10.8578
R33 A2.n2 A2.n1 3.12177
R34 A2.n2 A2.n0 1.81453
R35 A2.n3 A2.n2 1.1255
R36 A2.n3 A2 0.219402
R37 A2 A2.n3 0.0655
R38 VPWR.n57 VPWR.n55 8629.41
R39 VPWR.n60 VPWR.n54 8629.41
R40 VPWR.n40 VPWR.n39 8629.41
R41 VPWR.n42 VPWR.n37 8629.41
R42 VPWR.n23 VPWR.n22 8629.41
R43 VPWR.n25 VPWR.n20 8629.41
R44 VPWR.n6 VPWR.n4 8629.41
R45 VPWR.n9 VPWR.n3 8629.41
R46 VPWR.n56 VPWR.n53 920.471
R47 VPWR.n43 VPWR.n36 920.471
R48 VPWR.n26 VPWR.n19 920.471
R49 VPWR.n5 VPWR.n2 920.471
R50 VPWR.n62 VPWR.n53 914.447
R51 VPWR.n45 VPWR.n43 914.447
R52 VPWR.n28 VPWR.n26 914.447
R53 VPWR.n11 VPWR.n2 914.447
R54 VPWR.t58 VPWR.n127 804.731
R55 VPWR.n129 VPWR.t58 751.692
R56 VPWR.n101 VPWR.t7 671.408
R57 VPWR.n90 VPWR.t42 671.408
R58 VPWR VPWR.t57 630.375
R59 VPWR.n160 VPWR.n159 602.456
R60 VPWR.n182 VPWR.n70 602.456
R61 VPWR.n74 VPWR.n73 585
R62 VPWR.n76 VPWR.n75 585
R63 VPWR.n56 VPWR.n51 480.764
R64 VPWR.n36 VPWR.n34 480.764
R65 VPWR.n19 VPWR.n17 480.764
R66 VPWR.n5 VPWR.n1 480.764
R67 VPWR VPWR.t22 458.724
R68 VPWR.t57 VPWR 458.724
R69 VPWR.n122 VPWR.t64 420.25
R70 VPWR.n118 VPWR.t23 388.656
R71 VPWR.n153 VPWR.t24 388.656
R72 VPWR.n131 VPWR.t59 388.656
R73 VPWR.n104 VPWR.t1 388.656
R74 VPWR.n113 VPWR.t2 388.656
R75 VPWR.n78 VPWR.t11 388.656
R76 VPWR.n83 VPWR.t12 388.656
R77 VPWR.n64 VPWR.n51 379.2
R78 VPWR.n47 VPWR.n34 379.2
R79 VPWR.n30 VPWR.n17 379.2
R80 VPWR.n13 VPWR.n1 379.2
R81 VPWR VPWR.t60 369.938
R82 VPWR VPWR.t51 369.938
R83 VPWR.n107 VPWR.n100 322.329
R84 VPWR.n85 VPWR.n81 322.329
R85 VPWR.n164 VPWR.n162 259.697
R86 VPWR.n140 VPWR.t52 255.905
R87 VPWR.n145 VPWR.t61 255.905
R88 VPWR.n121 VPWR.t65 255.905
R89 VPWR.n161 VPWR.t28 255.905
R90 VPWR.n111 VPWR.t63 254.475
R91 VPWR.n136 VPWR.t26 252.95
R92 VPWR.n141 VPWR.t67 252.95
R93 VPWR.n146 VPWR.t40 252.95
R94 VPWR.n181 VPWR.t36 252.95
R95 VPWR.n160 VPWR.t9 251.516
R96 VPWR.n71 VPWR.t69 250.724
R97 VPWR.n69 VPWR.t34 250.724
R98 VPWR.t64 VPWR.t39 248.599
R99 VPWR.t60 VPWR.t66 248.599
R100 VPWR.t51 VPWR.t25 248.599
R101 VPWR.n176 VPWR.t46 248.219
R102 VPWR.n163 VPWR.t30 248.219
R103 VPWR.n122 VPWR 221.964
R104 VPWR.n129 VPWR.t73 215.827
R105 VPWR.n111 VPWR.n110 213.119
R106 VPWR.n151 VPWR.n122 213.119
R107 VPWR.n119 VPWR.t74 210.964
R108 VPWR.n105 VPWR.t72 210.964
R109 VPWR.n80 VPWR.t71 210.964
R110 VPWR.n171 VPWR.n170 209.368
R111 VPWR.t39 VPWR 198.287
R112 VPWR.t66 VPWR 198.287
R113 VPWR.t25 VPWR 198.287
R114 VPWR.n173 VPWR.n172 183.673
R115 VPWR VPWR.t37 182.952
R116 VPWR VPWR.n171 182.952
R117 VPWR.t31 VPWR 182.952
R118 VPWR.n75 VPWR.n74 159.476
R119 VPWR.n162 VPWR.t56 157.014
R120 VPWR.t68 VPWR.t43 154.417
R121 VPWR.t49 VPWR.t27 147.703
R122 VPWR.t20 VPWR.t6 140.989
R123 VPWR.t27 VPWR.t29 140.989
R124 VPWR.t35 VPWR.t33 140.989
R125 VPWR.t45 VPWR.t68 140.989
R126 VPWR.t41 VPWR.t13 140.989
R127 VPWR.n162 VPWR.t48 137.079
R128 VPWR.n110 VPWR 125.883
R129 VPWR.n172 VPWR 125.883
R130 VPWR.n100 VPWR.t21 116.341
R131 VPWR.n81 VPWR.t14 116.341
R132 VPWR.t6 VPWR 112.457
R133 VPWR.t29 VPWR 112.457
R134 VPWR VPWR.t41 112.457
R135 VPWR VPWR.t54 109.1
R136 VPWR.t0 VPWR.t20 104.064
R137 VPWR.t13 VPWR.t10 104.064
R138 VPWR.t15 VPWR 102.385
R139 VPWR.t62 VPWR 99.0288
R140 VPWR.n159 VPWR.t50 96.1553
R141 VPWR.n70 VPWR.t5 96.1553
R142 VPWR VPWR.t4 92.315
R143 VPWR.n74 VPWR.t44 86.7743
R144 VPWR.n110 VPWR.t62 83.9228
R145 VPWR.n171 VPWR.t47 80.5659
R146 VPWR.t37 VPWR.t0 77.209
R147 VPWR.t10 VPWR.t31 77.209
R148 VPWR.n75 VPWR.t55 66.8398
R149 VPWR.n63 VPWR.n62 66.6358
R150 VPWR.n46 VPWR.n45 66.6358
R151 VPWR.n29 VPWR.n28 66.6358
R152 VPWR.n12 VPWR.n11 66.6358
R153 VPWR.n159 VPWR.t16 63.3219
R154 VPWR.n70 VPWR.t18 63.3219
R155 VPWR VPWR.t49 62.103
R156 VPWR.n57 VPWR.n56 61.6672
R157 VPWR.n61 VPWR.n60 61.6672
R158 VPWR.n40 VPWR.n36 61.6672
R159 VPWR.n37 VPWR.n35 61.6672
R160 VPWR.n23 VPWR.n19 61.6672
R161 VPWR.n20 VPWR.n18 61.6672
R162 VPWR.n6 VPWR.n5 61.6672
R163 VPWR.n10 VPWR.n9 61.6672
R164 VPWR.n58 VPWR.n57 60.9564
R165 VPWR.n60 VPWR.n59 60.9564
R166 VPWR.n41 VPWR.n40 60.9564
R167 VPWR.n38 VPWR.n37 60.9564
R168 VPWR.n24 VPWR.n23 60.9564
R169 VPWR.n21 VPWR.n20 60.9564
R170 VPWR.n7 VPWR.n6 60.9564
R171 VPWR.n9 VPWR.n8 60.9564
R172 VPWR.n46 VPWR.n35 60.6123
R173 VPWR.n29 VPWR.n18 60.6123
R174 VPWR.n63 VPWR.n52 59.4829
R175 VPWR.n12 VPWR.n0 58.7299
R176 VPWR.t43 VPWR 55.3892
R177 VPWR.t17 VPWR 52.0323
R178 VPWR VPWR.t47 45.3185
R179 VPWR VPWR.t8 41.9616
R180 VPWR.n58 VPWR.n54 38.5759
R181 VPWR.n59 VPWR.n55 38.5759
R182 VPWR.n42 VPWR.n41 38.5759
R183 VPWR.n39 VPWR.n38 38.5759
R184 VPWR.n25 VPWR.n24 38.5759
R185 VPWR.n22 VPWR.n21 38.5759
R186 VPWR.n7 VPWR.n3 38.5759
R187 VPWR.n8 VPWR.n4 38.5759
R188 VPWR.n170 VPWR.n92 34.6358
R189 VPWR.n170 VPWR.n93 34.6358
R190 VPWR.n175 VPWR.n174 34.6358
R191 VPWR.n172 VPWR 28.5341
R192 VPWR.n100 VPWR.t38 28.4453
R193 VPWR.n81 VPWR.t32 28.4453
R194 VPWR.n177 VPWR.n176 28.3534
R195 VPWR.n174 VPWR.n173 25.6953
R196 VPWR.n140 VPWR.n125 25.224
R197 VPWR.n136 VPWR.n125 25.224
R198 VPWR.n145 VPWR.n124 25.224
R199 VPWR.n141 VPWR.n124 25.224
R200 VPWR.n147 VPWR.n121 25.224
R201 VPWR.n147 VPWR.n146 25.224
R202 VPWR.n165 VPWR.n161 25.224
R203 VPWR.n111 VPWR.n95 23.7181
R204 VPWR VPWR.n101 23.252
R205 VPWR.n160 VPWR.n95 21.4593
R206 VPWR.n141 VPWR.n140 20.3299
R207 VPWR.n146 VPWR.n145 20.3299
R208 VPWR.t4 VPWR.t35 20.1418
R209 VPWR.n182 VPWR.n69 19.9534
R210 VPWR.n181 VPWR.n180 19.8181
R211 VPWR.n151 VPWR.n121 17.3181
R212 VPWR.n164 VPWR.n163 17.3181
R213 VPWR.n161 VPWR.n160 16.5652
R214 VPWR.n165 VPWR.n164 16.5652
R215 VPWR.n136 VPWR.n135 15.8123
R216 VPWR.n152 VPWR.n151 14.2735
R217 VPWR.n112 VPWR.n111 14.2735
R218 VPWR.n174 VPWR.n90 13.9299
R219 VPWR.n67 VPWR.n66 13.6791
R220 VPWR.n182 VPWR.n181 13.5534
R221 VPWR.n117 VPWR.n116 11.4366
R222 VPWR.n65 VPWR.n64 11.3235
R223 VPWR.n48 VPWR.n47 11.3235
R224 VPWR.n31 VPWR.n30 11.3235
R225 VPWR.n14 VPWR.n13 11.3235
R226 VPWR.n173 VPWR.n91 11.2937
R227 VPWR.n157 VPWR.n156 11.2737
R228 VPWR.t8 VPWR.t15 10.0712
R229 VPWR.n131 VPWR.n128 9.60526
R230 VPWR.n118 VPWR.n117 9.60526
R231 VPWR.n83 VPWR.n82 9.60526
R232 VPWR.n120 VPWR.n96 9.3005
R233 VPWR.n155 VPWR.n154 9.3005
R234 VPWR.n152 VPWR.n97 9.3005
R235 VPWR.n151 VPWR.n150 9.3005
R236 VPWR.n146 VPWR.n123 9.3005
R237 VPWR.n142 VPWR.n141 9.3005
R238 VPWR.n137 VPWR.n136 9.3005
R239 VPWR.n133 VPWR.n132 9.3005
R240 VPWR.n138 VPWR.n125 9.3005
R241 VPWR.n140 VPWR.n139 9.3005
R242 VPWR.n143 VPWR.n124 9.3005
R243 VPWR.n145 VPWR.n144 9.3005
R244 VPWR.n148 VPWR.n147 9.3005
R245 VPWR.n149 VPWR.n121 9.3005
R246 VPWR.n178 VPWR.n177 9.3005
R247 VPWR.n183 VPWR.n182 9.3005
R248 VPWR.n167 VPWR.n92 9.3005
R249 VPWR.n160 VPWR.n158 9.3005
R250 VPWR.n111 VPWR.n109 9.3005
R251 VPWR.n103 VPWR.n102 9.3005
R252 VPWR.n106 VPWR.n98 9.3005
R253 VPWR.n115 VPWR.n114 9.3005
R254 VPWR.n112 VPWR.n99 9.3005
R255 VPWR.n108 VPWR.n95 9.3005
R256 VPWR.n161 VPWR.n94 9.3005
R257 VPWR.n166 VPWR.n165 9.3005
R258 VPWR.n170 VPWR.n169 9.3005
R259 VPWR.n168 VPWR.n93 9.3005
R260 VPWR.n181 VPWR.n68 9.3005
R261 VPWR.n180 VPWR.n179 9.3005
R262 VPWR.n175 VPWR.n72 9.3005
R263 VPWR.n174 VPWR.n77 9.3005
R264 VPWR.n89 VPWR.n88 9.3005
R265 VPWR.n87 VPWR.n86 9.3005
R266 VPWR.n84 VPWR.n79 9.3005
R267 VPWR.n15 VPWR.n0 8.23557
R268 VPWR.n76 VPWR.n73 6.8005
R269 VPWR.n135 VPWR.n127 6.48583
R270 VPWR.n62 VPWR.n61 6.02403
R271 VPWR.n11 VPWR.n10 6.02403
R272 VPWR.n130 VPWR.n129 5.8885
R273 VPWR.n44 VPWR.n35 4.89462
R274 VPWR.n28 VPWR.n27 4.89462
R275 VPWR.n154 VPWR.n120 4.67352
R276 VPWR.n135 VPWR.n134 4.62124
R277 VPWR.n132 VPWR.n131 4.36875
R278 VPWR.n154 VPWR.n153 4.36875
R279 VPWR.n114 VPWR.n113 4.36875
R280 VPWR.n84 VPWR.n83 4.36875
R281 VPWR.t33 VPWR.t17 3.35739
R282 VPWR.t54 VPWR.t45 3.35739
R283 VPWR.n44 VPWR.n33 3.23917
R284 VPWR.n27 VPWR.n16 3.23136
R285 VPWR.n52 VPWR.n50 3.22655
R286 VPWR.n132 VPWR.n130 3.2005
R287 VPWR.n54 VPWR.n53 2.84665
R288 VPWR.n55 VPWR.n51 2.84665
R289 VPWR.n43 VPWR.n42 2.84665
R290 VPWR.n39 VPWR.n34 2.84665
R291 VPWR.n26 VPWR.n25 2.84665
R292 VPWR.n22 VPWR.n17 2.84665
R293 VPWR.n3 VPWR.n2 2.84665
R294 VPWR.n4 VPWR.n1 2.84665
R295 VPWR.n130 VPWR.n127 2.8165
R296 VPWR.n107 VPWR.n106 2.54018
R297 VPWR.n86 VPWR.n85 2.54018
R298 VPWR.n120 VPWR.n119 2.33701
R299 VPWR.n106 VPWR.n105 2.33701
R300 VPWR.n86 VPWR.n80 2.33701
R301 VPWR.n64 VPWR.n63 2.28169
R302 VPWR.n47 VPWR.n46 2.28169
R303 VPWR.n30 VPWR.n29 2.28169
R304 VPWR.n13 VPWR.n12 2.28169
R305 VPWR.n114 VPWR.n107 2.13383
R306 VPWR.n85 VPWR.n84 2.13383
R307 VPWR.n119 VPWR.n118 2.03225
R308 VPWR.n105 VPWR.n104 2.03225
R309 VPWR.n80 VPWR.n78 2.03225
R310 VPWR.n10 VPWR.n0 1.88285
R311 VPWR.n185 VPWR.n184 1.753
R312 VPWR.n93 VPWR.n69 1.50638
R313 VPWR.n177 VPWR.n76 1.4005
R314 VPWR.n103 VPWR.n101 1.37193
R315 VPWR.n90 VPWR.n89 1.37193
R316 VPWR.n49 VPWR.n48 1.143
R317 VPWR.n32 VPWR.n31 1.143
R318 VPWR.n66 VPWR.n65 1.13925
R319 VPWR.n15 VPWR.n14 1.13675
R320 VPWR.n61 VPWR.n52 1.12991
R321 VPWR.n45 VPWR.n44 1.12991
R322 VPWR.n27 VPWR.n18 1.12991
R323 VPWR.n126 VPWR 1.06099
R324 VPWR.n33 VPWR.n32 0.862816
R325 VPWR.n16 VPWR.n15 0.770881
R326 VPWR.n163 VPWR.n92 0.753441
R327 VPWR.n176 VPWR.n175 0.753441
R328 VPWR.n50 VPWR.n49 0.729231
R329 VPWR.n73 VPWR.n71 0.6005
R330 VPWR.n185 VPWR.n67 0.511794
R331 VPWR VPWR.n185 0.460219
R332 VPWR.n66 VPWR.n50 0.405788
R333 VPWR.n180 VPWR.n71 0.4005
R334 VPWR.n32 VPWR.n16 0.392323
R335 VPWR.n49 VPWR.n33 0.360318
R336 VPWR.n153 VPWR.n152 0.305262
R337 VPWR.n104 VPWR.n103 0.305262
R338 VPWR.n113 VPWR.n112 0.305262
R339 VPWR.n89 VPWR.n78 0.305262
R340 VPWR.t53 VPWR.n58 0.27666
R341 VPWR.n59 VPWR.t53 0.27666
R342 VPWR.n41 VPWR.t19 0.27666
R343 VPWR.n38 VPWR.t19 0.27666
R344 VPWR.n24 VPWR.t70 0.27666
R345 VPWR.n21 VPWR.t70 0.27666
R346 VPWR.t3 VPWR.n7 0.27666
R347 VPWR.n8 VPWR.t3 0.27666
R348 VPWR.n134 VPWR.n133 0.180304
R349 VPWR.n134 VPWR 0.120408
R350 VPWR.n117 VPWR.n96 0.120292
R351 VPWR.n155 VPWR.n97 0.120292
R352 VPWR.n149 VPWR.n148 0.120292
R353 VPWR.n148 VPWR.n123 0.120292
R354 VPWR.n144 VPWR.n143 0.120292
R355 VPWR.n143 VPWR.n142 0.120292
R356 VPWR.n139 VPWR.n138 0.120292
R357 VPWR.n138 VPWR.n137 0.120292
R358 VPWR.n133 VPWR.n128 0.120292
R359 VPWR.n102 VPWR.n98 0.120292
R360 VPWR.n115 VPWR.n99 0.120292
R361 VPWR.n166 VPWR.n94 0.120292
R362 VPWR.n167 VPWR.n166 0.120292
R363 VPWR.n183 VPWR.n68 0.120292
R364 VPWR.n179 VPWR.n178 0.120292
R365 VPWR.n178 VPWR.n72 0.120292
R366 VPWR.n88 VPWR.n87 0.120292
R367 VPWR.n87 VPWR.n79 0.120292
R368 VPWR.n82 VPWR.n79 0.120292
R369 VPWR.n156 VPWR.n96 0.11899
R370 VPWR.n102 VPWR 0.0981562
R371 VPWR.n157 VPWR 0.0955521
R372 VPWR.n116 VPWR.n98 0.0916458
R373 VPWR.n65 VPWR 0.06425
R374 VPWR.n48 VPWR 0.06425
R375 VPWR.n31 VPWR 0.06425
R376 VPWR.n14 VPWR 0.06425
R377 VPWR.n150 VPWR 0.0603958
R378 VPWR VPWR.n149 0.0603958
R379 VPWR.n144 VPWR 0.0603958
R380 VPWR.n139 VPWR 0.0603958
R381 VPWR.n109 VPWR 0.0603958
R382 VPWR VPWR.n108 0.0603958
R383 VPWR VPWR.n94 0.0603958
R384 VPWR.n169 VPWR 0.0603958
R385 VPWR VPWR.n168 0.0603958
R386 VPWR.n179 VPWR 0.0603958
R387 VPWR.n88 VPWR 0.0603958
R388 VPWR.n91 VPWR 0.0590938
R389 VPWR.n184 VPWR 0.0525833
R390 VPWR.n184 VPWR.n183 0.0460729
R391 VPWR.n109 VPWR 0.0382604
R392 VPWR VPWR.n126 0.0369583
R393 VPWR.n150 VPWR 0.03175
R394 VPWR.n169 VPWR 0.03175
R395 VPWR.n116 VPWR.n115 0.0291458
R396 VPWR.n67 VPWR 0.0236148
R397 VPWR VPWR.n97 0.0226354
R398 VPWR VPWR.n123 0.0226354
R399 VPWR.n142 VPWR 0.0226354
R400 VPWR.n137 VPWR 0.0226354
R401 VPWR.n128 VPWR 0.0226354
R402 VPWR VPWR.n99 0.0226354
R403 VPWR.n108 VPWR 0.0226354
R404 VPWR.n158 VPWR 0.0226354
R405 VPWR VPWR.n167 0.0226354
R406 VPWR.n168 VPWR 0.0226354
R407 VPWR VPWR.n68 0.0226354
R408 VPWR VPWR.n72 0.0226354
R409 VPWR VPWR.n77 0.0226354
R410 VPWR.n82 VPWR 0.0226354
R411 VPWR.n158 VPWR.n157 0.00310417
R412 VPWR.n156 VPWR.n155 0.00180208
R413 VPWR.n126 VPWR 0.00180208
R414 VPWR.n91 VPWR.n77 0.00180208
R415 x2.GP1.n4 x2.GP1.t4 450.938
R416 x2.GP1.n4 x2.GP1.t5 445.666
R417 x2.GP1.n5 x2.GP1.n3 195.832
R418 x2.GP1.n1 x2.GP1.n0 101.49
R419 x2.GP1.n3 x2.GP1.t3 26.5955
R420 x2.GP1.n3 x2.GP1.t2 26.5955
R421 x2.GP1.n0 x2.GP1.t1 24.9236
R422 x2.GP1.n0 x2.GP1.t0 24.9236
R423 x2.GP1.n5 x1.gpo0 11.8923
R424 x1.gpo0 x2.x1.GP 11.5413
R425 x2.GP1.n2 x1.x11.Y 10.7525
R426 x1.x11.Y x2.GP1.n5 8.09215
R427 x2.GP1.n2 x1.x11.Y 6.6565
R428 x1.x11.Y x2.GP1.n2 5.04292
R429 x2.x1.GP x2.GP1.n4 2.90754
R430 x1.x11.Y x2.GP1.n1 2.5605
R431 x2.GP1.n1 x1.x11.Y 1.93989
R432 Z1.n1 Z1.t1 23.6581
R433 Z1.n3 Z1.t2 23.3739
R434 Z1.n1 Z1.t3 10.7528
R435 Z1.n0 Z1.t0 10.6417
R436 Z1.n2 Z1.n1 1.30064
R437 Z1 Z1.n4 0.983856
R438 Z1.n3 Z1.n2 0.726502
R439 Z1.n2 Z1.n0 0.512491
R440 Z1.n4 Z1.n0 0.359663
R441 Z1.n4 Z1.n3 0.216071
R442 A1.n1 A1.t2 26.3998
R443 A1.n1 A1.t1 23.5483
R444 A1.n0 A1.t0 12.7127
R445 A1.n0 A1.t3 10.8578
R446 A1.n2 A1.n1 3.12177
R447 A1.n2 A1.n0 1.81453
R448 A1.n3 A1.n2 1.1255
R449 A1.n3 A1 0.21174
R450 A1 A1.n3 0.0655
R451 select0.n5 select0.t4 327.99
R452 select0.n9 select0.t3 293.969
R453 select0.n3 select0.t7 261.887
R454 select0.n1 select0.t9 212.081
R455 select0.n0 select0.t2 212.081
R456 select0.n5 select0.t0 199.457
R457 select0.n2 select0.n1 183.185
R458 select0.n3 select0.t8 155.847
R459 select0 select0.n9 154.065
R460 select0.n6 select0.n5 152
R461 select0.n4 select0.n3 152
R462 select0.n1 select0.t1 139.78
R463 select0.n0 select0.t6 139.78
R464 select0.n9 select0.t5 138.338
R465 select0.n1 select0.n0 61.346
R466 select0.n10 select0 13.4199
R467 select0.n8 select0.n4 11.9062
R468 select0.n11 select0.n8 11.7395
R469 select0.n12 select0.n11 11.5949
R470 select0.n12 select0.n2 9.68118
R471 select0.n7 select0 9.17383
R472 select0.n2 select0 5.8885
R473 select0.n10 select0 5.57469
R474 select0.n8 select0.n7 4.6505
R475 select0.n11 select0.n10 4.6505
R476 select0.n7 select0.n6 2.98717
R477 select0.n6 select0 2.34717
R478 select0.n4 select0 2.07109
R479 select0 select0.n12 0.559212
R480 VGND.n182 VGND.n181 545142
R481 VGND.n42 VGND.n41 20148.7
R482 VGND.n55 VGND.n10 19433.3
R483 VGND.n49 VGND.n48 19054.3
R484 VGND VGND.n180 11981.2
R485 VGND.n50 VGND.n11 11744.7
R486 VGND.n54 VGND.n11 11744.7
R487 VGND.n50 VGND.n12 11744.7
R488 VGND.n54 VGND.n12 11744.7
R489 VGND.n36 VGND.n22 11744.7
R490 VGND.n40 VGND.n22 11744.7
R491 VGND.n36 VGND.n23 11744.7
R492 VGND.n40 VGND.n23 11744.7
R493 VGND.n43 VGND.n16 11744.7
R494 VGND.n47 VGND.n16 11744.7
R495 VGND.n43 VGND.n17 11744.7
R496 VGND.n47 VGND.n17 11744.7
R497 VGND.n184 VGND.n4 11744.7
R498 VGND.n184 VGND.n5 11744.7
R499 VGND.n9 VGND.n5 11744.7
R500 VGND.n9 VGND.n4 11744.7
R501 VGND.n56 VGND.n7 5416.06
R502 VGND.n21 VGND.n7 5357.62
R503 VGND.n180 VGND.n56 3878.48
R504 VGND.n183 VGND.n182 2174.55
R505 VGND VGND.t55 1289.66
R506 VGND.n179 VGND.n178 1198.25
R507 VGND.n137 VGND.n135 1198.25
R508 VGND.n146 VGND.n6 1194.5
R509 VGND.n165 VGND.n164 1171.32
R510 VGND VGND.n6 918.774
R511 VGND.t26 VGND 918.774
R512 VGND.t40 VGND.t57 826.054
R513 VGND.t51 VGND.t60 826.054
R514 VGND.t62 VGND.t16 792.337
R515 VGND.n45 VGND.n44 767.294
R516 VGND.n8 VGND.n3 767.294
R517 VGND.n52 VGND.n51 763.106
R518 VGND.n38 VGND.n37 763.106
R519 VGND.n51 VGND.n15 732.236
R520 VGND.n37 VGND.n34 732.236
R521 VGND.n44 VGND.n20 732.236
R522 VGND.n8 VGND.n1 732.236
R523 VGND.n181 VGND.n6 708.047
R524 VGND.t34 VGND.t19 708.047
R525 VGND.t16 VGND.t66 708.047
R526 VGND.t49 VGND.t53 708.047
R527 VGND.t46 VGND.t14 708.047
R528 VGND.n164 VGND.t9 681.482
R529 VGND.t19 VGND 564.751
R530 VGND.t53 VGND 564.751
R531 VGND VGND.t46 564.751
R532 VGND.n182 VGND 564.751
R533 VGND.t38 VGND.t47 554.492
R534 VGND.t14 VGND.t3 522.606
R535 VGND.n181 VGND.t38 513.419
R536 VGND.t13 VGND 480.461
R537 VGND.t6 VGND 459.26
R538 VGND.t9 VGND 459.26
R539 VGND.t47 VGND.t33 431.272
R540 VGND.t3 VGND.t26 387.74
R541 VGND VGND.t64 370.37
R542 VGND VGND.t21 370.37
R543 VGND.t42 VGND 370.37
R544 VGND.t33 VGND 343.991
R545 VGND.n135 VGND.t59 337.166
R546 VGND.n179 VGND.n57 334.815
R547 VGND.n46 VGND.n45 325.502
R548 VGND.n185 VGND.n3 325.502
R549 VGND.n135 VGND.t40 320.307
R550 VGND.n53 VGND.n52 304.204
R551 VGND.n39 VGND.n38 304.204
R552 VGND.t59 VGND 295.019
R553 VGND.n180 VGND.t6 278.519
R554 VGND VGND.t62 261.303
R555 VGND.t64 VGND.t44 248.889
R556 VGND.t21 VGND.t23 248.889
R557 VGND.t29 VGND.t31 248.889
R558 VGND.t36 VGND.t42 248.889
R559 VGND.t0 VGND 244.445
R560 VGND.n53 VGND.n13 242.448
R561 VGND.n39 VGND.n24 242.448
R562 VGND.n46 VGND.n18 242.448
R563 VGND.n186 VGND.n185 242.448
R564 VGND.n10 VGND.t18 241.579
R565 VGND.n153 VGND.t63 240.575
R566 VGND.n133 VGND.t56 237.327
R567 VGND VGND.n179 222.222
R568 VGND.n164 VGND 222.222
R569 VGND.n112 VGND.t68 218.308
R570 VGND.n88 VGND.t69 218.308
R571 VGND.n70 VGND.t70 218.308
R572 VGND.n140 VGND.t71 218.308
R573 VGND.n109 VGND.t10 214.456
R574 VGND.n111 VGND.t11 214.456
R575 VGND.n122 VGND.t7 214.456
R576 VGND.n89 VGND.t8 214.456
R577 VGND.n65 VGND.t4 214.456
R578 VGND.n69 VGND.t5 214.456
R579 VGND.n145 VGND.t1 214.456
R580 VGND.n139 VGND.t2 214.456
R581 VGND.n127 VGND.n126 204.457
R582 VGND.n78 VGND.n77 200.231
R583 VGND.n83 VGND.n82 200.231
R584 VGND.n72 VGND.n67 200.105
R585 VGND.t44 VGND 198.519
R586 VGND.t23 VGND 198.519
R587 VGND VGND.t29 198.519
R588 VGND VGND.t36 198.519
R589 VGND.n45 VGND.n17 195
R590 VGND.t25 VGND.n17 195
R591 VGND.n19 VGND.n16 195
R592 VGND.t25 VGND.n16 195
R593 VGND.n38 VGND.n23 195
R594 VGND.t12 VGND.n23 195
R595 VGND.n33 VGND.n22 195
R596 VGND.t12 VGND.n22 195
R597 VGND.n52 VGND.n12 195
R598 VGND.n12 VGND.t28 195
R599 VGND.n14 VGND.n11 195
R600 VGND.n11 VGND.t28 195
R601 VGND.n4 VGND.n2 195
R602 VGND.n57 VGND.n4 195
R603 VGND.n5 VGND.n3 195
R604 VGND.t18 VGND.n5 195
R605 VGND VGND.t51 177.012
R606 VGND.n36 VGND.n35 174.921
R607 VGND.n42 VGND.t25 163.988
R608 VGND.n49 VGND.t28 163.85
R609 VGND.n100 VGND.t65 162.471
R610 VGND.n95 VGND.t22 162.471
R611 VGND.n177 VGND.t32 162.471
R612 VGND.n172 VGND.t43 162.471
R613 VGND.n154 VGND.t17 162.471
R614 VGND.n78 VGND.t50 160.046
R615 VGND.n83 VGND.t35 160.046
R616 VGND.n91 VGND.t45 160.017
R617 VGND.n58 VGND.t24 160.017
R618 VGND.n61 VGND.t30 160.017
R619 VGND.n170 VGND.t37 160.017
R620 VGND.n161 VGND.t54 160.017
R621 VGND.n156 VGND.t67 160.017
R622 VGND.n153 VGND.t20 158.534
R623 VGND.n184 VGND.n183 152.552
R624 VGND VGND.t18 121.481
R625 VGND.n41 VGND.n21 105.025
R626 VGND.n48 VGND.n7 98.5767
R627 VGND.n56 VGND.n55 98.4942
R628 VGND.t31 VGND.n57 85.9264
R629 VGND.t66 VGND.t13 84.2917
R630 VGND.n67 VGND.t15 72.8576
R631 VGND.n126 VGND.t48 72.8576
R632 VGND.t25 VGND.n7 65.4109
R633 VGND.n56 VGND.t28 65.3562
R634 VGND.n35 VGND.n21 58.925
R635 VGND.n77 VGND.t52 58.5719
R636 VGND.n82 VGND.t41 58.5719
R637 VGND.t57 VGND.t34 50.5752
R638 VGND.t60 VGND.t49 50.5752
R639 VGND.n125 VGND 43.9579
R640 VGND.n128 VGND.n125 34.6358
R641 VGND.n132 VGND.n85 34.6358
R642 VGND.n15 VGND.n14 30.8711
R643 VGND.n34 VGND.n33 30.8711
R644 VGND.n20 VGND.n19 30.8711
R645 VGND.n2 VGND.n1 30.8711
R646 VGND.n165 VGND.n63 26.9246
R647 VGND.n146 VGND.n132 25.6926
R648 VGND.n77 VGND.t61 25.4291
R649 VGND.n82 VGND.t58 25.4291
R650 VGND.n100 VGND.n99 25.224
R651 VGND.n99 VGND.n91 25.224
R652 VGND.n95 VGND.n94 25.224
R653 VGND.n94 VGND.n58 25.224
R654 VGND.n177 VGND.n176 25.224
R655 VGND.n176 VGND.n61 25.224
R656 VGND.n172 VGND.n171 25.224
R657 VGND.n171 VGND.n170 25.224
R658 VGND.n161 VGND.n160 25.224
R659 VGND.n155 VGND.n154 25.224
R660 VGND.n156 VGND.n155 25.224
R661 VGND.n183 VGND.t18 24.1956
R662 VGND.n153 VGND.n152 24.0946
R663 VGND.n67 VGND.t27 22.3257
R664 VGND.n126 VGND.t39 22.3257
R665 VGND.n160 VGND.n78 21.4593
R666 VGND.n152 VGND.n83 21.4593
R667 VGND.n95 VGND.n91 20.3299
R668 VGND.n172 VGND.n61 20.3299
R669 VGND.n101 VGND.n100 19.2926
R670 VGND.n161 VGND.n76 17.7867
R671 VGND.n178 VGND.n177 17.3181
R672 VGND.t55 VGND.t0 16.8587
R673 VGND.n178 VGND.n58 15.8123
R674 VGND.n170 VGND.n63 15.8123
R675 VGND.n108 VGND.n63 14.775
R676 VGND.n138 VGND.n137 14.775
R677 VGND.n154 VGND.n153 13.5534
R678 VGND.n124 VGND.n123 11.2844
R679 VGND.n47 VGND.n46 11.0382
R680 VGND.n48 VGND.n47 11.0382
R681 VGND.n44 VGND.n43 11.0382
R682 VGND.n43 VGND.n42 11.0382
R683 VGND.n40 VGND.n39 11.0382
R684 VGND.n41 VGND.n40 11.0382
R685 VGND.n37 VGND.n36 11.0382
R686 VGND.n54 VGND.n53 11.0382
R687 VGND.n55 VGND.n54 11.0382
R688 VGND.n51 VGND.n50 11.0382
R689 VGND.n50 VGND.n49 11.0382
R690 VGND.n9 VGND.n8 11.0382
R691 VGND.n10 VGND.n9 11.0382
R692 VGND.n185 VGND.n184 11.0382
R693 VGND.n14 VGND.n13 10.9181
R694 VGND.n33 VGND.n24 10.9181
R695 VGND.n19 VGND.n18 10.9181
R696 VGND.n186 VGND.n2 10.9181
R697 VGND.n27 VGND.n15 10.4476
R698 VGND.n34 VGND.n32 10.4476
R699 VGND.n25 VGND.n20 10.4476
R700 VGND.n187 VGND.n1 10.4476
R701 VGND.n156 VGND.n78 10.1652
R702 VGND.n111 VGND.n106 9.70901
R703 VGND.n123 VGND.n122 9.70901
R704 VGND.n69 VGND.n68 9.70901
R705 VGND.n127 VGND.n85 9.41227
R706 VGND.n166 VGND.n165 9.3005
R707 VGND.n170 VGND.n169 9.3005
R708 VGND.n174 VGND.n61 9.3005
R709 VGND.n178 VGND.n59 9.3005
R710 VGND.n92 VGND.n58 9.3005
R711 VGND.n97 VGND.n91 9.3005
R712 VGND.n102 VGND.n101 9.3005
R713 VGND.n120 VGND.n119 9.3005
R714 VGND.n121 VGND.n87 9.3005
R715 VGND.n100 VGND.n90 9.3005
R716 VGND.n99 VGND.n98 9.3005
R717 VGND.n96 VGND.n95 9.3005
R718 VGND.n94 VGND.n93 9.3005
R719 VGND.n177 VGND.n60 9.3005
R720 VGND.n176 VGND.n175 9.3005
R721 VGND.n173 VGND.n172 9.3005
R722 VGND.n171 VGND.n62 9.3005
R723 VGND.n114 VGND.n113 9.3005
R724 VGND.n110 VGND.n105 9.3005
R725 VGND.n108 VGND.n107 9.3005
R726 VGND.n168 VGND.n63 9.3005
R727 VGND.n147 VGND.n146 9.3005
R728 VGND.n144 VGND.n143 9.3005
R729 VGND.n84 VGND.n83 9.3005
R730 VGND.n153 VGND.n81 9.3005
R731 VGND.n158 VGND.n78 9.3005
R732 VGND.n71 VGND.n66 9.3005
R733 VGND.n74 VGND.n73 9.3005
R734 VGND.n76 VGND.n75 9.3005
R735 VGND.n162 VGND.n161 9.3005
R736 VGND.n160 VGND.n159 9.3005
R737 VGND.n157 VGND.n156 9.3005
R738 VGND.n155 VGND.n79 9.3005
R739 VGND.n154 VGND.n80 9.3005
R740 VGND.n152 VGND.n151 9.3005
R741 VGND.n138 VGND.n134 9.3005
R742 VGND.n142 VGND.n141 9.3005
R743 VGND.n132 VGND.n131 9.3005
R744 VGND.n130 VGND.n85 9.3005
R745 VGND.n129 VGND.n128 9.3005
R746 VGND.n125 VGND.n86 9.3005
R747 VGND.n137 VGND.n136 9.3005
R748 VGND.n31 VGND.n30 8.45078
R749 VGND.n188 VGND.n0 8.30267
R750 VGND.n29 VGND.n28 7.97888
R751 VGND.n30 VGND.n26 7.97601
R752 VGND.n28 VGND.n27 7.16724
R753 VGND.n32 VGND.n31 7.16724
R754 VGND.n26 VGND.n25 7.16724
R755 VGND.n188 VGND.n187 7.16724
R756 VGND.n137 VGND.n83 7.15344
R757 VGND.n167 VGND.n163 6.50373
R758 VGND.n128 VGND.n127 6.4005
R759 VGND.n113 VGND.n110 6.26433
R760 VGND.n121 VGND.n120 6.26433
R761 VGND.n110 VGND.n109 5.85582
R762 VGND.n122 VGND.n121 5.85582
R763 VGND.n73 VGND.n65 5.85582
R764 VGND.n145 VGND.n144 5.85582
R765 VGND.n141 VGND.n133 5.85582
R766 VGND.n168 VGND.n167 4.788
R767 VGND.n27 VGND.n13 4.73093
R768 VGND.n32 VGND.n24 4.73093
R769 VGND.n25 VGND.n18 4.73093
R770 VGND.n187 VGND.n186 4.73093
R771 VGND.n167 VGND.n166 4.50726
R772 VGND.n103 VGND 4.01425
R773 VGND.n72 VGND.n71 3.40476
R774 VGND.n113 VGND.n112 3.13241
R775 VGND.n120 VGND.n88 3.13241
R776 VGND.n71 VGND.n70 3.13241
R777 VGND.n141 VGND.n140 3.13241
R778 VGND.n149 VGND.n148 2.88636
R779 VGND.n73 VGND.n72 2.86007
R780 VGND.n112 VGND.n111 2.7239
R781 VGND.n89 VGND.n88 2.7239
R782 VGND.n70 VGND.n69 2.7239
R783 VGND.n140 VGND.n139 2.7239
R784 VGND.n118 VGND.n117 1.753
R785 VGND.n116 VGND.n115 1.753
R786 VGND.n150 VGND.n149 1.21169
R787 VGND.n117 VGND.n116 0.761313
R788 VGND.n117 VGND.n104 0.591917
R789 VGND.n149 VGND 0.531208
R790 VGND.n104 VGND.n103 0.506165
R791 VGND.n30 VGND.n29 0.467019
R792 VGND.n109 VGND.n108 0.409011
R793 VGND.n101 VGND.n89 0.409011
R794 VGND.n76 VGND.n65 0.409011
R795 VGND.n146 VGND.n145 0.409011
R796 VGND.n144 VGND.n133 0.409011
R797 VGND.n139 VGND.n138 0.409011
R798 VGND.n103 VGND.n0 0.198729
R799 VGND.n166 VGND.n64 0.1255
R800 VGND.n123 VGND.n87 0.120292
R801 VGND.n119 VGND.n87 0.120292
R802 VGND.n98 VGND.n90 0.120292
R803 VGND.n98 VGND.n97 0.120292
R804 VGND.n96 VGND.n93 0.120292
R805 VGND.n93 VGND.n92 0.120292
R806 VGND.n175 VGND.n60 0.120292
R807 VGND.n175 VGND.n174 0.120292
R808 VGND.n173 VGND.n62 0.120292
R809 VGND.n169 VGND.n62 0.120292
R810 VGND.n107 VGND.n105 0.120292
R811 VGND.n114 VGND.n106 0.120292
R812 VGND.n129 VGND.n86 0.120292
R813 VGND.n130 VGND.n129 0.120292
R814 VGND.n131 VGND.n130 0.120292
R815 VGND.n142 VGND.n134 0.120292
R816 VGND.n80 VGND.n79 0.120292
R817 VGND.n157 VGND.n79 0.120292
R818 VGND.n159 VGND.n158 0.120292
R819 VGND.n75 VGND.n74 0.120292
R820 VGND.n74 VGND.n66 0.120292
R821 VGND.n68 VGND.n66 0.120292
R822 VGND VGND.n142 0.0981562
R823 VGND VGND.n124 0.09425
R824 VGND.n116 VGND 0.0881354
R825 VGND.n29 VGND.n0 0.0766574
R826 VGND.n115 VGND.n114 0.0721146
R827 VGND.n151 VGND.n150 0.0708125
R828 VGND.n28 VGND 0.064875
R829 VGND.n26 VGND 0.064875
R830 VGND VGND.n188 0.064875
R831 VGND.n31 VGND 0.063625
R832 VGND.n119 VGND.n118 0.0616979
R833 VGND.n90 VGND 0.0603958
R834 VGND VGND.n96 0.0603958
R835 VGND VGND.n59 0.0603958
R836 VGND.n60 VGND 0.0603958
R837 VGND VGND.n173 0.0603958
R838 VGND VGND.n168 0.0603958
R839 VGND.n107 VGND 0.0603958
R840 VGND.n131 VGND 0.0603958
R841 VGND.n143 VGND 0.0603958
R842 VGND.n136 VGND 0.0603958
R843 VGND VGND.n84 0.0603958
R844 VGND.n151 VGND 0.0603958
R845 VGND VGND.n81 0.0603958
R846 VGND VGND.n80 0.0603958
R847 VGND.n158 VGND 0.0603958
R848 VGND.n159 VGND 0.0603958
R849 VGND.n75 VGND 0.0603958
R850 VGND.n118 VGND.n102 0.0590938
R851 VGND.n163 VGND 0.0590938
R852 VGND.n150 VGND.n84 0.0499792
R853 VGND.n115 VGND.n105 0.0486771
R854 VGND.n148 VGND 0.0460729
R855 VGND.n147 VGND 0.0343542
R856 VGND VGND.n59 0.0330521
R857 VGND.n136 VGND 0.0330521
R858 VGND VGND.n64 0.03175
R859 VGND.n104 VGND 0.0292529
R860 VGND.n35 VGND.t12 0.028591
R861 VGND.n102 VGND 0.0226354
R862 VGND.n97 VGND 0.0226354
R863 VGND.n92 VGND 0.0226354
R864 VGND.n174 VGND 0.0226354
R865 VGND.n169 VGND 0.0226354
R866 VGND.n106 VGND 0.0226354
R867 VGND.n143 VGND 0.0226354
R868 VGND VGND.n134 0.0226354
R869 VGND.n81 VGND 0.0226354
R870 VGND VGND.n157 0.0226354
R871 VGND.n162 VGND 0.0226354
R872 VGND.n68 VGND 0.0226354
R873 VGND.n148 VGND.n147 0.0148229
R874 VGND.n124 VGND.n86 0.00440625
R875 VGND.n168 VGND.n64 0.00180208
R876 VGND.n163 VGND.n162 0.00180208
R877 x2.GP4.n2 x2.GP4.t4 450.938
R878 x2.GP4.n2 x2.GP4.t5 445.666
R879 x1.x14.Y x2.GP4.n4 203.923
R880 x2.GP4.n0 x2.GP4.n1 101.49
R881 x2.GP4.n4 x2.GP4.t3 26.5955
R882 x2.GP4.n4 x2.GP4.t0 26.5955
R883 x2.GP4.n1 x2.GP4.t2 24.9236
R884 x2.GP4.n1 x2.GP4.t1 24.9236
R885 x1.gpo3 x2.x4.GP 16.5752
R886 x2.GP4.n3 x1.x14.Y 10.7525
R887 x2.GP4.n0 x1.gpo3 7.7042
R888 x2.GP4.n3 x1.x14.Y 6.6565
R889 x1.x14.Y x2.GP4.n3 5.04292
R890 x2.x4.GP x2.GP4.n2 2.95993
R891 x1.x14.Y x2.GP4.n0 2.5605
R892 x2.GP4.n0 x1.x14.Y 1.93989
R893 Z4.n1 Z4.t3 23.6581
R894 Z4.n3 Z4.t2 23.3739
R895 Z4.n1 Z4.t0 10.7528
R896 Z4.n0 Z4.t1 10.6417
R897 Z4.n2 Z4.n1 1.30064
R898 Z4 Z4.n4 0.983856
R899 Z4.n3 Z4.n2 0.726502
R900 Z4.n2 Z4.n0 0.512491
R901 Z4.n4 Z4.n0 0.359663
R902 Z4.n4 Z4.n3 0.216071
R903 A4.n1 A4.t3 26.3998
R904 A4.n1 A4.t2 23.5483
R905 A4.n0 A4.t1 12.7127
R906 A4.n0 A4.t0 10.8578
R907 A4.n2 A4.n1 3.12177
R908 A4.n2 A4.n0 1.81453
R909 A4.n3 A4.n2 1.1255
R910 A4 A4.n3 0.203263
R911 A4.n3 A4 0.0655
R912 select1.n10 select1.t1 327.99
R913 select1.n3 select1.t8 293.969
R914 select1.n6 select1.t3 256.07
R915 select1.n1 select1.t2 212.081
R916 select1.n0 select1.t5 212.081
R917 select1.n10 select1.t9 199.457
R918 select1.n2 select1.n1 182.929
R919 select1 select1.n3 154.065
R920 select1.n11 select1.n10 152
R921 select1.n7 select1.n6 152
R922 select1.n6 select1.t7 150.03
R923 select1.n1 select1.t6 139.78
R924 select1.n0 select1.t0 139.78
R925 select1.n3 select1.t4 138.338
R926 select1.n1 select1.n0 61.346
R927 select1.n5 select1 22.1096
R928 select1.n14 select1.n13 14.6836
R929 select1.n13 select1.n12 14.6704
R930 select1.n12 select1 13.8672
R931 select1.n4 select1 13.8328
R932 select1.n11 select1 12.1605
R933 select1.n14 select1.n2 10.6811
R934 select1.n7 select1.n5 10.4374
R935 select1.n9 select1.n8 8.15359
R936 select1.n2 select1 6.1445
R937 select1.n4 select1 5.16179
R938 select1.n9 select1.n4 4.65206
R939 select1.n8 select1 3.93896
R940 select1 select1.n11 2.34717
R941 select1.n5 select1 2.16665
R942 select1.n8 select1.n7 1.57588
R943 select1.n13 select1.n9 0.79438
R944 select1.n12 select1 0.6405
R945 select1 select1.n14 0.248606
R946 x2.GN1.n1 x2.GN1.t6 377.486
R947 x2.GN1.n1 x2.GN1.t4 374.202
R948 x2.GN1.n7 x2.GN1.t0 339.418
R949 x2.GN1.n0 x2.GN1.t1 274.06
R950 x2.GN1.n4 x2.GN1.t5 212.081
R951 x2.GN1.n3 x2.GN1.t7 212.081
R952 x2.GN1.n5 x2.GN1.n4 182.673
R953 x2.GN1.n4 x2.GN1.t2 139.78
R954 x2.GN1.n3 x2.GN1.t3 139.78
R955 x2.GN1.n4 x2.GN1.n3 61.346
R956 x2.GN1 x2.GN1.n5 15.8606
R957 x2.GN1 x2.GN1.n6 13.8044
R958 x2.GN1.n2 x2.GN1 11.5859
R959 x2.GN1 x2.GN1.n0 11.0989
R960 x2.GN1 x2.GN1.n2 10.8756
R961 x2.GN1.n6 x2.GN1 8.1246
R962 x2.GN1.n8 x2.GN1 6.6565
R963 x2.GN1.n5 x2.GN1 6.4005
R964 x2.GN1.n0 x2.GN1 6.1445
R965 x2.GN1.n2 x2.GN1 4.55738
R966 x2.GN1.n8 x2.GN1.n7 4.0914
R967 x2.GN1 x2.GN1.n8 3.61789
R968 x2.GN1.n6 x2.GN1 3.26325
R969 x2.GN1.n0 x2.GN1 2.86947
R970 x2.GN1 x2.GN1.n1 2.04102
R971 x2.GN1.n7 x2.GN1 1.74382
R972 x2.GN4.n1 x2.GN4.t6 377.486
R973 x2.GN4.n1 x2.GN4.t7 374.202
R974 x2.GN4.n7 x2.GN4.t0 339.418
R975 x2.GN4.n0 x2.GN4.t1 274.06
R976 x2.GN4.n4 x2.GN4.t2 212.081
R977 x2.GN4.n3 x2.GN4.t3 212.081
R978 x2.GN4.n5 x2.GN4.n4 184.977
R979 x2.GN4.n4 x2.GN4.t4 139.78
R980 x2.GN4.n3 x2.GN4.t5 139.78
R981 x2.GN4.n4 x2.GN4.n3 61.346
R982 x2.GN4.n6 x2.GN4 18.2601
R983 x2.GN4 x2.GN4.n2 17.2682
R984 x2.GN4 x2.GN4.n5 15.0136
R985 x2.GN4 x2.GN4.n0 11.2645
R986 x2.GN4 x2.GN4.n6 8.9605
R987 x2.GN4.n6 x2.GN4 8.4485
R988 x2.GN4.n2 x2.GN4 8.16743
R989 x2.GN4.n8 x2.GN4 6.6565
R990 x2.GN4.n0 x2.GN4 6.1445
R991 x2.GN4.n2 x2.GN4 4.58237
R992 x2.GN4.n5 x2.GN4 4.0965
R993 x2.GN4.n8 x2.GN4.n7 4.0914
R994 x2.GN4 x2.GN4.n8 3.61789
R995 x2.GN4.n0 x2.GN4 2.86947
R996 x2.GN4 x2.GN4.n1 2.04102
R997 x2.GN4.n7 x2.GN4 1.74382
R998 select2.n1 select2.t0 212.081
R999 select2.n0 select2.t1 212.081
R1000 select2.n2 select2.n1 183.441
R1001 select2.n1 select2.t2 139.78
R1002 select2.n0 select2.t3 139.78
R1003 select2.n1 select2.n0 61.346
R1004 select2 select2.n2 11.4331
R1005 select2.n2 select2 5.6325
R1006 nselect2.n5 nselect2.n4 196.339
R1007 nselect2.n1 nselect2.n0 101.49
R1008 nselect2.n4 nselect2.t0 26.5955
R1009 nselect2.n4 nselect2.t1 26.5955
R1010 nselect2.n0 nselect2.t2 24.9236
R1011 nselect2.n0 nselect2.t3 24.9236
R1012 nselect2.n2 nselect2 13.5685
R1013 nselect2.n3 nselect2 10.7525
R1014 nselect2.n6 nselect2.n2 9.50196
R1015 nselect2.n6 nselect2.n5 7.64514
R1016 nselect2.n5 nselect2 7.58449
R1017 nselect2.n3 nselect2 6.6565
R1018 nselect2 nselect2.n3 5.04292
R1019 nselect2 nselect2.n2 3.8405
R1020 nselect2 nselect2.n1 2.5605
R1021 nselect2.n1 nselect2 1.93989
R1022 nselect2 nselect2.n6 1.81877
R1023 Z3.n1 Z3.t2 23.6581
R1024 Z3.n3 Z3.t3 23.3739
R1025 Z3.n1 Z3.t0 10.7528
R1026 Z3.n0 Z3.t1 10.6417
R1027 Z3.n2 Z3.n1 1.30064
R1028 Z3.n5 Z3.n4 0.924585
R1029 Z3.n3 Z3.n2 0.726502
R1030 Z3.n2 Z3.n0 0.512491
R1031 Z3.n4 Z3.n0 0.359663
R1032 Z3.n4 Z3.n3 0.216071
R1033 Z3.n5 Z3 0.0656042
R1034 Z3 Z3.n5 0.0376287
R1035 A3.n1 A3.t2 26.3998
R1036 A3.n1 A3.t3 23.5483
R1037 A3.n0 A3.t0 12.7127
R1038 A3.n0 A3.t1 10.8578
R1039 A3.n2 A3.n1 3.12177
R1040 A3.n2 A3.n0 1.81453
R1041 A3.n3 A3.n2 1.1255
R1042 A3.n3 A3 0.210543
R1043 A3 A3.n3 0.0655
C0 x2.GN1 a_5275_n4651# 0.12869f
C1 x2.GN4 a_5329_n2857# 0.001562f
C2 x2.GN2 a_5329_n2857# 8.14e-21
C3 x2.GN3 a_5275_n4059# 0.048646f
C4 a_5275_n3683# x2.GP3 0.00144f
C5 a_5275_n4235# select2 8.66e-20
C6 a_5275_n4235# select0 0.246189f
C7 a_5275_n4235# select1 0.03417f
C8 a_5275_n4235# VPWR 0.161854f
C9 a_5275_n3683# x1.nSEL0 1.91e-20
C10 a_5329_n2857# x2.GN3 1.07e-20
C11 x2.GN4 x2.GN1 0.001075f
C12 x2.GN2 x2.GN1 0.065209f
C13 a_5275_n3683# x1.nSEL1 7.84e-19
C14 a_5275_n4235# a_5275_n4651# 0.002207f
C15 a_5301_n4107# VPWR 4.32e-19
C16 a_5275_n3683# a_5275_n4059# 3.02e-19
C17 x1.nSEL0 x1.nSEL1 0.352716f
C18 x2.GN1 x2.GN3 0.00286f
C19 a_5275_n3507# A1 5.02e-20
C20 a_5275_n3507# nselect2 6.01e-20
C21 a_5275_n3507# select0 0.279858f
C22 a_5275_n3507# select1 0.127717f
C23 a_5275_n3507# VPWR 0.262185f
C24 x1.nSEL0 a_5275_n4059# 0.001174f
C25 a_5275_n4235# x2.GN2 0.106186f
C26 x1.nSEL1 a_5275_n4059# 0.041068f
C27 select0 a_5301_n3555# 0.001558f
C28 VPWR a_5301_n3555# 0.001496f
C29 a_5275_n4235# x2.GN3 6.68e-19
C30 nselect2 a_5275_n2995# 9.77e-20
C31 a_5301_n4107# x2.GN2 0.002418f
C32 select0 a_5275_n2995# 0.220366f
C33 a_5275_n3683# x2.GN1 6.43e-20
C34 select1 a_5275_n2995# 0.125445f
C35 VPWR a_5275_n2995# 0.217381f
C36 x2.GN1 x2.GP3 0.002439f
C37 a_5275_n3507# x2.GN4 0.003699f
C38 a_5275_n3507# x2.GN2 5.62e-20
C39 x1.nSEL0 x2.GN1 0.004383f
C40 x2.GN1 x1.nSEL1 0.034891f
C41 a_5301_n4107# x2.GN3 5.17e-20
C42 Z4 A4 4.51497f
C43 Z3 Z4 0.002229f
C44 Z4 A3 0.005563f
C45 A3 A4 2.08862f
C46 x2.GN1 a_5275_n4059# 1.46e-19
C47 Z3 A3 4.51555f
C48 A2 A4 2.39e-19
C49 VPWR Z4 2.81281f
C50 a_5275_n3507# x2.GN3 0.004288f
C51 Z3 Z2 7.65e-19
C52 Z2 A3 1.49e-20
C53 A2 A3 1.81997f
C54 Z3 A2 0.004565f
C55 A2 Z2 4.51569f
C56 x2.GN4 a_5301_n3555# 3.22e-19
C57 A1 Z3 4.74e-21
C58 x2.GN2 a_5301_n3555# 3.11e-20
C59 VPWR A4 1.54289f
C60 A1 Z2 0.004942f
C61 Z3 VPWR 2.85668f
C62 VPWR A3 1.61205f
C63 A1 A2 1.81909f
C64 x2.GN4 a_5275_n2995# 0.134079f
C65 x2.GN2 a_5275_n2995# 7.58e-21
C66 a_5275_n4235# x1.nSEL0 0.03096f
C67 VPWR Z2 2.85288f
C68 A2 VPWR 1.61513f
C69 A1 Z1 4.51491f
C70 m3_10270_n3216# A4 0.091998f
C71 Z1 select0 4.1e-22
C72 m3_9240_n3230# A4 6.07e-21
C73 A1 select0 3.49e-20
C74 select2 nselect2 0.150826f
C75 VPWR Z1 2.90992f
C76 select0 nselect2 1.88e-19
C77 select2 select0 0.368835f
C78 A1 select1 1.45e-21
C79 A1 VPWR 1.98654f
C80 VPWR nselect2 1.06761f
C81 a_5275_n4235# x1.nSEL1 0.073392f
C82 m3_9240_n3230# A3 0.097296f
C83 select1 nselect2 0.001177f
C84 select2 select1 0.139336f
C85 select2 VPWR 0.231538f
C86 select1 select0 1.66811f
C87 VPWR select0 1.09594f
C88 VPWR select1 2.64545f
C89 A2 m3_8196_n3226# 0.1002f
C90 x2.GN3 a_5301_n3555# 0.001073f
C91 a_5275_n4235# a_5275_n4059# 0.185422f
C92 select2 m2_5406_n4650# 4.4e-19
C93 m2_5406_n4650# select0 0.130999f
C94 x2.GN3 a_5275_n2995# 1.07e-20
C95 a_5329_n4513# select0 9.55e-19
C96 m2_5406_n4650# VPWR 0.139545f
C97 m2_5406_n4650# select1 0.183786f
C98 a_5329_n4513# VPWR 9.09e-19
C99 a_5301_n4107# x1.nSEL0 2.51e-19
C100 select0 a_5275_n4651# 0.048888f
C101 m3_10270_n3216# m3_9240_n3230# 0.003741f
C102 a_5275_n3507# a_5275_n3683# 0.185422f
C103 VPWR a_5275_n4651# 0.210313f
C104 select1 a_5275_n4651# 0.02803f
C105 a_5275_n3507# x2.GP3 5.21e-19
C106 a_5301_n4107# x1.nSEL1 9.57e-19
C107 m3_9240_n3230# m3_8196_n3226# 0.003764f
C108 x2.GN4 Z4 0.443708f
C109 a_5275_n3507# x1.nSEL0 1.21e-20
C110 m2_5406_n4650# a_5275_n4651# 0.01297f
C111 x2.GN4 A4 3.83736f
C112 a_5329_n4513# a_5275_n4651# 0.006584f
C113 x2.GN4 Z3 0.00128f
C114 x2.GN4 A3 0.187073f
C115 Z3 x2.GN2 2.12e-20
C116 x2.GN2 A3 0.004147f
C117 a_5275_n3507# x1.nSEL1 1.59e-19
C118 x2.GN4 A2 3.42e-19
C119 x2.GN2 Z2 0.427019f
C120 x2.GN2 A2 3.81441f
C121 x2.GN4 A1 0.001437f
C122 x2.GN2 Z1 7.73e-19
C123 A1 x2.GN2 0.157008f
C124 x2.GN4 nselect2 1.53e-20
C125 x2.GN4 select0 0.218396f
C126 select2 x2.GN2 0.001308f
C127 x2.GN2 select0 0.114345f
C128 a_5275_n3683# a_5301_n3555# 0.004764f
C129 x2.GN4 VPWR 1.23434f
C130 x2.GN4 select1 0.059813f
C131 x2.GN2 select1 0.108649f
C132 x2.GN2 VPWR 0.600374f
C133 x2.GN3 Z4 1.95e-20
C134 x2.GP3 a_5301_n3555# 4.39e-19
C135 x2.GN4 m3_10270_n3216# 0.084813f
C136 x2.GN4 m3_9240_n3230# 7.07e-19
C137 x2.GN2 m3_9240_n3230# 0.016745f
C138 x2.GN3 A4 0.004656f
C139 a_5275_n4235# x2.GN1 0.012466f
C140 Z3 x2.GN3 0.427085f
C141 x2.GN3 A3 3.80482f
C142 x2.GN4 m3_8196_n3226# 7.17e-19
C143 x2.GN2 m3_8196_n3226# 0.099332f
C144 x2.GN3 Z2 0.00126f
C145 A2 x2.GN3 0.164396f
C146 a_5329_n4513# x2.GN2 8.86e-19
C147 x2.GN2 a_5275_n4651# 0.039612f
C148 Z1 x2.GN3 4.42e-20
C149 x1.nSEL1 a_5301_n3555# 4.08e-19
C150 A1 x2.GN3 0.002069f
C151 x2.GN3 nselect2 7.39e-21
C152 select2 x2.GN3 0.001055f
C153 x2.GN3 select0 0.254198f
C154 x2.GN3 select1 0.272312f
C155 VPWR x2.GN3 0.649708f
C156 m3_10270_n3216# x2.GN3 0.016026f
C157 m3_9240_n3230# x2.GN3 0.087318f
C158 a_5301_n4107# x2.GN1 1.22e-20
C159 x2.GN3 m3_8196_n3226# 0.001446f
C160 x2.GP3 Z4 0.071646f
C161 x2.GN4 x2.GN2 8.84e-19
C162 a_5275_n3507# x2.GN1 3.78e-20
C163 x2.GP3 A4 0.161499f
C164 Z3 x2.GP3 0.278332f
C165 x2.GP3 A3 4.01143f
C166 x2.GP3 Z2 1.03e-20
C167 A1 a_5275_n3683# 1.55e-21
C168 A2 x2.GP3 0.001826f
C169 a_5275_n3683# nselect2 1.29e-19
C170 select2 a_5275_n3683# 0.009143f
C171 a_5275_n3683# select0 0.086353f
C172 a_5329_n2857# a_5275_n2995# 0.006584f
C173 a_5275_n3683# VPWR 0.171441f
C174 a_5275_n3683# select1 0.261734f
C175 Z1 x2.GP3 7.56e-20
C176 A1 x2.GP3 0.001277f
C177 x2.GP3 select0 2.82e-19
C178 x2.GP3 select1 0.003386f
C179 VPWR x2.GP3 1.78272f
C180 x2.GN4 x2.GN3 0.07149f
C181 a_5275_n4235# a_5301_n4107# 0.004764f
C182 x2.GN2 x2.GN3 0.067572f
C183 A1 x1.nSEL0 1.93e-21
C184 select2 x1.nSEL0 0.131218f
C185 m3_10270_n3216# x2.GP3 0.006132f
C186 x1.nSEL0 select0 0.324538f
C187 x1.nSEL0 select1 0.137403f
C188 m3_9240_n3230# x2.GP3 0.002824f
C189 x1.nSEL0 VPWR 0.391764f
C190 x1.nSEL1 nselect2 0.047548f
C191 select2 x1.nSEL1 0.164723f
C192 select0 x1.nSEL1 0.168464f
C193 x2.GP3 m3_8196_n3226# 9.67e-19
C194 select1 x1.nSEL1 0.272823f
C195 VPWR x1.nSEL1 0.481997f
C196 m2_5406_n4650# x1.nSEL0 3.43e-19
C197 x1.nSEL0 a_5275_n4651# 0.081627f
C198 select2 a_5275_n4059# 1.67e-19
C199 select0 a_5275_n4059# 0.143958f
C200 select1 a_5275_n4059# 0.254026f
C201 VPWR a_5275_n4059# 0.19314f
C202 m2_5406_n4650# x1.nSEL1 0.00815f
C203 a_5329_n4513# x1.nSEL1 0.00175f
C204 x1.nSEL1 a_5275_n4651# 0.193944f
C205 x2.GN4 a_5275_n3683# 6.84e-19
C206 x2.GN2 a_5275_n3683# 1.63e-19
C207 x2.GN4 x2.GP3 3.44338f
C208 x2.GN2 x2.GP3 0.004319f
C209 a_5329_n2857# select0 1.4e-19
C210 VPWR a_5329_n2857# 8.97e-19
C211 a_5329_n2857# select1 8.84e-19
C212 x2.GN4 x1.nSEL0 2.26e-20
C213 x2.GN2 x1.nSEL0 0.154394f
C214 x2.GN2 x1.nSEL1 0.209956f
C215 a_5275_n3683# x2.GN3 0.104343f
C216 x2.GN1 Z2 4.77e-21
C217 A2 x2.GN1 1.78e-19
C218 x2.GP3 x2.GN3 2.868f
C219 x2.GN1 Z1 0.428262f
C220 A1 x2.GN1 4.61808f
C221 select2 x2.GN1 0.009187f
C222 x2.GN1 select0 0.020307f
C223 x2.GN1 select1 0.312198f
C224 VPWR x2.GN1 1.36505f
C225 x2.GN2 a_5275_n4059# 0.017018f
C226 x1.nSEL0 x2.GN3 4.01e-20
C227 x2.GN3 x1.nSEL1 0.012418f
C228 m2_5406_n4650# x2.GN1 0.06935f
C229 x2.GN1 m3_8196_n3226# 6.03e-20
C230 a_5329_n4513# x2.GN1 0.001144f
C231 Z4 VGND 2.703709f
C232 A4 VGND 3.673923f
C233 Z3 VGND 2.48903f
C234 A3 VGND 3.139328f
C235 Z2 VGND 2.454758f
C236 A2 VGND 3.238628f
C237 Z1 VGND 2.838278f
C238 A1 VGND 3.972252f
C239 nselect2 VGND 0.47102f
C240 select2 VGND 1.16504f
C241 select0 VGND 1.41757f
C242 select1 VGND 1.610708f
C243 VPWR VGND 56.37729f
C244 m3_10270_n3216# VGND 0.090191f $ **FLOATING
C245 m3_9240_n3230# VGND 0.086003f $ **FLOATING
C246 m3_8196_n3226# VGND 0.168273f $ **FLOATING
C247 m2_5406_n4650# VGND 0.065655f $ **FLOATING
C248 a_5329_n4513# VGND 0.006505f
C249 a_5275_n4651# VGND 0.266782f
C250 x1.nSEL0 VGND 0.649982f
C251 x2.GN1 VGND 6.355386f
C252 a_5301_n4107# VGND 0.004461f
C253 a_5275_n4235# VGND 0.220868f
C254 x1.nSEL1 VGND 0.69132f
C255 x2.GN2 VGND 3.93258f
C256 a_5275_n4059# VGND 0.23458f
C257 x2.GP3 VGND 1.67788f
C258 a_5301_n3555# VGND 0.006801f
C259 x2.GN3 VGND 3.65509f
C260 a_5275_n3683# VGND 0.232764f
C261 a_5275_n3507# VGND 0.249604f
C262 x2.GN4 VGND 7.590769f
C263 a_5329_n2857# VGND 0.006439f
C264 a_5275_n2995# VGND 0.306675f
C265 A3.t0 VGND 0.893857f
C266 A3.t1 VGND 0.513146f
C267 A3.n0 VGND 4.9699f
C268 A3.t2 VGND 0.925152f
C269 A3.t3 VGND 0.654459f
C270 A3.n1 VGND 5.08132f
C271 A3.n2 VGND 0.803733f
C272 A3.n3 VGND 0.264783f
C273 Z3.t1 VGND 0.362117f
C274 Z3.n0 VGND 0.540706f
C275 Z3.t0 VGND 0.369386f
C276 Z3.t2 VGND 0.490183f
C277 Z3.n1 VGND 2.47361f
C278 Z3.n2 VGND 0.836966f
C279 Z3.t3 VGND 0.477048f
C280 Z3.n3 VGND 0.593305f
C281 Z3.n4 VGND 0.728891f
C282 Z3.n5 VGND 0.331987f
C283 x2.GN4.t1 VGND 0.06076f
C284 x2.GN4.n0 VGND 0.070042f
C285 x2.GN4.t6 VGND 0.686652f
C286 x2.GN4.t7 VGND 0.670085f
C287 x2.GN4.n1 VGND 3.00641f
C288 x2.GN4.n2 VGND 1.54718f
C289 x2.GN4.t2 VGND 0.038143f
C290 x2.GN4.t4 VGND 0.022477f
C291 x2.GN4.t3 VGND 0.038143f
C292 x2.GN4.t5 VGND 0.022477f
C293 x2.GN4.n3 VGND 0.063998f
C294 x2.GN4.n4 VGND 0.094806f
C295 x2.GN4.n5 VGND 0.042443f
C296 x2.GN4.n6 VGND 0.343794f
C297 x2.GN4.t0 VGND 0.155177f
C298 x2.GN4.n7 VGND 0.027911f
C299 x2.GN4.n8 VGND 0.031268f
C300 x2.GN1.t1 VGND 0.029997f
C301 x2.GN1.n0 VGND 0.034614f
C302 x2.GN1.t6 VGND 0.338995f
C303 x2.GN1.t4 VGND 0.330816f
C304 x2.GN1.n1 VGND 1.48424f
C305 x2.GN1.n2 VGND 0.51776f
C306 x2.GN1.t5 VGND 0.018831f
C307 x2.GN1.t2 VGND 0.011097f
C308 x2.GN1.t7 VGND 0.018831f
C309 x2.GN1.t3 VGND 0.011097f
C310 x2.GN1.n3 VGND 0.031595f
C311 x2.GN1.n4 VGND 0.046667f
C312 x2.GN1.n5 VGND 0.045389f
C313 x2.GN1.n6 VGND 0.098587f
C314 x2.GN1.t0 VGND 0.076609f
C315 x2.GN1.n7 VGND 0.013779f
C316 x2.GN1.n8 VGND 0.015437f
C317 select1.t2 VGND 0.032343f
C318 select1.t6 VGND 0.019059f
C319 select1.t5 VGND 0.032343f
C320 select1.t0 VGND 0.019059f
C321 select1.n0 VGND 0.054267f
C322 select1.n1 VGND 0.080179f
C323 select1.n2 VGND 0.048819f
C324 select1.t4 VGND 0.014966f
C325 select1.t8 VGND 0.031563f
C326 select1.n3 VGND 0.113336f
C327 select1.n4 VGND 0.021975f
C328 select1.n5 VGND 0.018928f
C329 select1.t3 VGND 0.022802f
C330 select1.t7 VGND 0.015669f
C331 select1.n6 VGND 0.06626f
C332 select1.n7 VGND 0.015263f
C333 select1.n8 VGND 0.109332f
C334 select1.n9 VGND 0.396f
C335 select1.t1 VGND 0.02778f
C336 select1.t9 VGND 0.018863f
C337 select1.n10 VGND 0.065634f
C338 select1.n11 VGND 0.01571f
C339 select1.n12 VGND 0.101902f
C340 select1.n13 VGND 0.457083f
C341 select1.n14 VGND 0.597136f
C342 A4.t1 VGND 0.893325f
C343 A4.t0 VGND 0.512841f
C344 A4.n0 VGND 4.96695f
C345 A4.t3 VGND 0.924602f
C346 A4.t2 VGND 0.65407f
C347 A4.n1 VGND 5.0783f
C348 A4.n2 VGND 0.803255f
C349 A4.n3 VGND 0.258761f
C350 Z4.t1 VGND 0.356817f
C351 Z4.n0 VGND 0.532792f
C352 Z4.t0 VGND 0.363979f
C353 Z4.t3 VGND 0.483009f
C354 Z4.n1 VGND 2.43741f
C355 Z4.n2 VGND 0.824716f
C356 Z4.t2 VGND 0.470066f
C357 Z4.n3 VGND 0.584621f
C358 Z4.n4 VGND 0.742893f
C359 x2.GP4.n0 VGND 0.095571f
C360 x2.x4.GP VGND 2.50543f
C361 x1.gpo3 VGND 1.18077f
C362 x2.GP4.t2 VGND 0.012052f
C363 x2.GP4.t1 VGND 0.012052f
C364 x2.GP4.n1 VGND 0.028739f
C365 x1.x14.Y VGND 0.104168f
C366 x2.GP4.t5 VGND 0.609957f
C367 x2.GP4.t4 VGND 0.626965f
C368 x2.GP4.n2 VGND 2.22891f
C369 x2.GP4.n3 VGND 0.017567f
C370 x2.GP4.t3 VGND 0.018542f
C371 x2.GP4.t0 VGND 0.018542f
C372 x2.GP4.n4 VGND 0.040723f
C373 A1.t0 VGND 0.813767f
C374 A1.t3 VGND 0.467169f
C375 A1.n0 VGND 4.5246f
C376 A1.t2 VGND 0.842259f
C377 A1.t1 VGND 0.59582f
C378 A1.n1 VGND 4.62603f
C379 A1.n2 VGND 0.731718f
C380 A1.n3 VGND 0.224671f
C381 Z1.t0 VGND 0.363377f
C382 Z1.n0 VGND 0.542586f
C383 Z1.t3 VGND 0.370671f
C384 Z1.t1 VGND 0.491889f
C385 Z1.n1 VGND 2.48222f
C386 Z1.n2 VGND 0.839878f
C387 Z1.t2 VGND 0.478707f
C388 Z1.n3 VGND 0.595368f
C389 Z1.n4 VGND 0.756551f
C390 x2.x1.GP VGND 1.98566f
C391 x2.GP1.t1 VGND 0.012716f
C392 x2.GP1.t0 VGND 0.012716f
C393 x2.GP1.n0 VGND 0.03032f
C394 x1.x11.Y VGND 0.046385f
C395 x2.GP1.n1 VGND 0.059566f
C396 x2.GP1.n2 VGND 0.018534f
C397 x2.GP1.t3 VGND 0.019563f
C398 x2.GP1.t2 VGND 0.019563f
C399 x2.GP1.n3 VGND 0.040309f
C400 x2.GP1.t5 VGND 0.643518f
C401 x2.GP1.t4 VGND 0.661463f
C402 x2.GP1.n4 VGND 2.33672f
C403 x1.gpo0 VGND 0.626909f
C404 x2.GP1.n5 VGND 0.086057f
C405 VPWR.n0 VGND 0.03081f
C406 VPWR.n1 VGND 0.137121f
C407 VPWR.n2 VGND 0.066225f
C408 VPWR.n3 VGND 0.557756f
C409 VPWR.n4 VGND 0.557756f
C410 VPWR.n5 VGND 0.091797f
C411 VPWR.n6 VGND 0.067234f
C412 VPWR.t3 VGND 0.741619f
C413 VPWR.n9 VGND 0.067234f
C414 VPWR.n10 VGND 2.85e-19
C415 VPWR.n11 VGND 0.040828f
C416 VPWR.n12 VGND 0.007424f
C417 VPWR.n13 VGND 0.080708f
C418 VPWR.n14 VGND 0.043153f
C419 VPWR.n15 VGND 0.08763f
C420 VPWR.n16 VGND 0.101662f
C421 VPWR.n17 VGND 0.137121f
C422 VPWR.n18 VGND 0.002226f
C423 VPWR.n19 VGND 0.091797f
C424 VPWR.n20 VGND 0.067234f
C425 VPWR.t70 VGND 0.741619f
C426 VPWR.n22 VGND 0.557756f
C427 VPWR.n23 VGND 0.067234f
C428 VPWR.n25 VGND 0.557756f
C429 VPWR.n26 VGND 0.066225f
C430 VPWR.n27 VGND 0.00533f
C431 VPWR.n28 VGND 0.040787f
C432 VPWR.n29 VGND 0.007491f
C433 VPWR.n30 VGND 0.080708f
C434 VPWR.n31 VGND 0.042812f
C435 VPWR.n32 VGND 0.069384f
C436 VPWR.n33 VGND 0.099666f
C437 VPWR.n34 VGND 0.137121f
C438 VPWR.n35 VGND 0.002362f
C439 VPWR.n36 VGND 0.091797f
C440 VPWR.n37 VGND 0.067234f
C441 VPWR.t19 VGND 0.741619f
C442 VPWR.n39 VGND 0.557756f
C443 VPWR.n40 VGND 0.067234f
C444 VPWR.n42 VGND 0.557756f
C445 VPWR.n43 VGND 0.066225f
C446 VPWR.n44 VGND 0.005339f
C447 VPWR.n45 VGND 0.040651f
C448 VPWR.n46 VGND 0.007491f
C449 VPWR.n47 VGND 0.080708f
C450 VPWR.n48 VGND 0.042812f
C451 VPWR.n49 VGND 0.067641f
C452 VPWR.n50 VGND 0.103727f
C453 VPWR.n51 VGND 0.137121f
C454 VPWR.n52 VGND 0.007292f
C455 VPWR.n53 VGND 0.066225f
C456 VPWR.n54 VGND 0.557756f
C457 VPWR.n55 VGND 0.557756f
C458 VPWR.n56 VGND 0.091797f
C459 VPWR.n57 VGND 0.067234f
C460 VPWR.t53 VGND 0.741619f
C461 VPWR.n60 VGND 0.067234f
C462 VPWR.n61 VGND 2.58e-19
C463 VPWR.n62 VGND 0.040828f
C464 VPWR.n63 VGND 0.007451f
C465 VPWR.n64 VGND 0.080708f
C466 VPWR.n65 VGND 0.043126f
C467 VPWR.n66 VGND 0.246672f
C468 VPWR.n67 VGND 0.187384f
C469 VPWR.n68 VGND 0.004178f
C470 VPWR.t34 VGND 0.008431f
C471 VPWR.n69 VGND 0.008293f
C472 VPWR.t18 VGND 9.05e-19
C473 VPWR.t5 VGND 0.001375f
C474 VPWR.n70 VGND 0.002375f
C475 VPWR.t36 VGND 0.008593f
C476 VPWR.t69 VGND 0.008431f
C477 VPWR.n71 VGND 0.008031f
C478 VPWR.n72 VGND 0.004178f
C479 VPWR.n73 VGND 0.003782f
C480 VPWR.t44 VGND 0.001241f
C481 VPWR.n74 VGND 0.003521f
C482 VPWR.t55 VGND 0.005101f
C483 VPWR.n75 VGND 0.004695f
C484 VPWR.n76 VGND 0.00419f
C485 VPWR.t46 VGND 0.008433f
C486 VPWR.n77 VGND 6.9e-19
C487 VPWR.t42 VGND 0.003616f
C488 VPWR.t11 VGND 0.005969f
C489 VPWR.n78 VGND 0.005884f
C490 VPWR.n79 VGND 0.007052f
C491 VPWR.t71 VGND 0.024909f
C492 VPWR.n80 VGND 0.02253f
C493 VPWR.t32 VGND 6.76e-19
C494 VPWR.t14 VGND 0.001812f
C495 VPWR.n81 VGND 0.008269f
C496 VPWR.t12 VGND 0.005969f
C497 VPWR.n82 VGND 0.004367f
C498 VPWR.n83 VGND 0.0163f
C499 VPWR.n84 VGND 0.012878f
C500 VPWR.n85 VGND 0.016727f
C501 VPWR.n86 VGND 0.009658f
C502 VPWR.n87 VGND 0.007052f
C503 VPWR.n88 VGND 0.005289f
C504 VPWR.n89 VGND 0.00332f
C505 VPWR.n90 VGND 0.010459f
C506 VPWR.n91 VGND 0.016397f
C507 VPWR.t47 VGND 0.016948f
C508 VPWR.n92 VGND 0.001276f
C509 VPWR.n93 VGND 0.001303f
C510 VPWR.n94 VGND 0.005289f
C511 VPWR.n95 VGND 0.001629f
C512 VPWR.t9 VGND 0.008547f
C513 VPWR.n96 VGND 0.007014f
C514 VPWR.n97 VGND 0.004178f
C515 VPWR.t74 VGND 0.024909f
C516 VPWR.n98 VGND 0.006209f
C517 VPWR.n99 VGND 0.004178f
C518 VPWR.t38 VGND 6.76e-19
C519 VPWR.t21 VGND 0.001812f
C520 VPWR.n100 VGND 0.008269f
C521 VPWR.t72 VGND 0.024909f
C522 VPWR.t7 VGND 0.003616f
C523 VPWR.n101 VGND 0.011165f
C524 VPWR.n102 VGND 0.006401f
C525 VPWR.n103 VGND 0.00332f
C526 VPWR.t1 VGND 0.005969f
C527 VPWR.n104 VGND 0.005884f
C528 VPWR.n105 VGND 0.02253f
C529 VPWR.n106 VGND 0.009658f
C530 VPWR.n107 VGND 0.016727f
C531 VPWR.t2 VGND 0.005969f
C532 VPWR.t63 VGND 0.008548f
C533 VPWR.n108 VGND 0.002415f
C534 VPWR.n109 VGND 0.002875f
C535 VPWR.t6 VGND 0.034122f
C536 VPWR.t20 VGND 0.032992f
C537 VPWR.t0 VGND 0.024405f
C538 VPWR.t37 VGND 0.035026f
C539 VPWR.t29 VGND 0.034122f
C540 VPWR.t27 VGND 0.038867f
C541 VPWR.t49 VGND 0.028246f
C542 VPWR.t15 VGND 0.01514f
C543 VPWR.t8 VGND 0.007005f
C544 VPWR.t62 VGND 0.024631f
C545 VPWR.n110 VGND 0.032141f
C546 VPWR.n111 VGND 0.02229f
C547 VPWR.n112 VGND 0.006552f
C548 VPWR.n113 VGND 0.010512f
C549 VPWR.n114 VGND 0.012878f
C550 VPWR.n115 VGND 0.004369f
C551 VPWR.n116 VGND 0.034804f
C552 VPWR.n117 VGND 0.047342f
C553 VPWR.t23 VGND 0.005969f
C554 VPWR.n118 VGND 0.011672f
C555 VPWR.n119 VGND 0.02253f
C556 VPWR.n120 VGND 0.013884f
C557 VPWR.t24 VGND 0.005969f
C558 VPWR.t65 VGND 0.008589f
C559 VPWR.n121 VGND 0.010036f
C560 VPWR.t22 VGND 0.076766f
C561 VPWR.t57 VGND 0.047161f
C562 VPWR.t25 VGND 0.019351f
C563 VPWR.t51 VGND 0.026784f
C564 VPWR.t66 VGND 0.019351f
C565 VPWR.t60 VGND 0.026784f
C566 VPWR.t39 VGND 0.019351f
C567 VPWR.t64 VGND 0.028963f
C568 VPWR.n122 VGND 0.031705f
C569 VPWR.n123 VGND 0.004178f
C570 VPWR.n124 VGND 0.001819f
C571 VPWR.t61 VGND 0.008589f
C572 VPWR.n125 VGND 0.001819f
C573 VPWR.t52 VGND 0.008589f
C574 VPWR.n126 VGND 0.122759f
C575 VPWR.n127 VGND 0.007185f
C576 VPWR.n128 VGND 0.004367f
C577 VPWR.t73 VGND 0.025299f
C578 VPWR.t58 VGND 0.005969f
C579 VPWR.n129 VGND 0.025046f
C580 VPWR.n130 VGND 0.012447f
C581 VPWR.t59 VGND 0.005969f
C582 VPWR.n131 VGND 0.0163f
C583 VPWR.n132 VGND 0.014991f
C584 VPWR.n133 VGND 0.009406f
C585 VPWR.n134 VGND 0.00734f
C586 VPWR.n135 VGND 0.007158f
C587 VPWR.t26 VGND 0.008593f
C588 VPWR.n136 VGND 0.010814f
C589 VPWR.n137 VGND 0.004178f
C590 VPWR.n138 VGND 0.007052f
C591 VPWR.n139 VGND 0.005289f
C592 VPWR.n140 VGND 0.010144f
C593 VPWR.t67 VGND 0.008593f
C594 VPWR.n141 VGND 0.010977f
C595 VPWR.n142 VGND 0.004178f
C596 VPWR.n143 VGND 0.007052f
C597 VPWR.n144 VGND 0.005289f
C598 VPWR.n145 VGND 0.010144f
C599 VPWR.t40 VGND 0.008593f
C600 VPWR.n146 VGND 0.010977f
C601 VPWR.n147 VGND 0.001819f
C602 VPWR.n148 VGND 0.007052f
C603 VPWR.n149 VGND 0.005289f
C604 VPWR.n150 VGND 0.002683f
C605 VPWR.n151 VGND 0.014656f
C606 VPWR.n152 VGND 0.006552f
C607 VPWR.n153 VGND 0.010512f
C608 VPWR.n154 VGND 0.017908f
C609 VPWR.n155 VGND 0.003564f
C610 VPWR.n156 VGND 0.032389f
C611 VPWR.n157 VGND 0.031406f
C612 VPWR.n158 VGND 7.28e-19
C613 VPWR.t16 VGND 9.05e-19
C614 VPWR.t50 VGND 0.001375f
C615 VPWR.n159 VGND 0.002375f
C616 VPWR.n160 VGND 0.015943f
C617 VPWR.t28 VGND 0.008589f
C618 VPWR.n161 VGND 0.010009f
C619 VPWR.t56 VGND 0.00283f
C620 VPWR.t48 VGND 0.007522f
C621 VPWR.n162 VGND 0.004267f
C622 VPWR.t30 VGND 0.008433f
C623 VPWR.n163 VGND 0.008897f
C624 VPWR.n164 VGND 0.011444f
C625 VPWR.n165 VGND 0.001507f
C626 VPWR.n166 VGND 0.007052f
C627 VPWR.n167 VGND 0.004178f
C628 VPWR.n168 VGND 0.002415f
C629 VPWR.n169 VGND 0.002683f
C630 VPWR.n170 VGND 0.01436f
C631 VPWR.n171 VGND 0.039157f
C632 VPWR.t17 VGND 0.007457f
C633 VPWR.t33 VGND 0.019434f
C634 VPWR.t35 VGND 0.021693f
C635 VPWR.t4 VGND 0.01514f
C636 VPWR.t43 VGND 0.028246f
C637 VPWR.t68 VGND 0.039771f
C638 VPWR.t45 VGND 0.019434f
C639 VPWR.t54 VGND 0.01514f
C640 VPWR.t31 VGND 0.035026f
C641 VPWR.t10 VGND 0.024405f
C642 VPWR.t13 VGND 0.032992f
C643 VPWR.t41 VGND 0.034122f
C644 VPWR.n172 VGND 0.023237f
C645 VPWR.n173 VGND 0.006751f
C646 VPWR.n174 VGND 0.004805f
C647 VPWR.n175 VGND 0.001276f
C648 VPWR.n176 VGND 0.009362f
C649 VPWR.n177 VGND 0.003571f
C650 VPWR.n178 VGND 0.007052f
C651 VPWR.n179 VGND 0.005289f
C652 VPWR.n180 VGND 0.003144f
C653 VPWR.n181 VGND 0.010688f
C654 VPWR.n182 VGND 0.007648f
C655 VPWR.n183 VGND 0.004868f
C656 VPWR.n184 VGND 0.013764f
C657 VPWR.n185 VGND 0.087548f
C658 A2.t2 VGND 0.763965f
C659 A2.t3 VGND 0.438578f
C660 A2.n0 VGND 4.2477f
C661 A2.t1 VGND 0.790712f
C662 A2.t0 VGND 0.559356f
C663 A2.n1 VGND 4.34292f
C664 A2.n2 VGND 0.686937f
C665 A2.n3 VGND 0.222065f
C666 Z2.t3 VGND 0.363425f
C667 Z2.n0 VGND 0.542659f
C668 Z2.t2 VGND 0.37072f
C669 Z2.t1 VGND 0.491954f
C670 Z2.n1 VGND 2.48255f
C671 Z2.n2 VGND 0.83999f
C672 Z2.t0 VGND 0.478771f
C673 Z2.n3 VGND 0.595448f
C674 Z2.n4 VGND 0.733795f
C675 Z2.n5 VGND 0.3243f
C676 x2.x2.GP VGND 2.76866f
C677 x1.gpo1 VGND 0.998586f
C678 x2.GP2.t3 VGND 0.016016f
C679 x2.GP2.t2 VGND 0.016016f
C680 x2.GP2.n0 VGND 0.03819f
C681 x1.x12.Y VGND 0.058128f
C682 x2.GP2.n1 VGND 0.075027f
C683 x2.GP2.n2 VGND 0.023344f
C684 x2.GP2.t1 VGND 0.02464f
C685 x2.GP2.t0 VGND 0.02464f
C686 x2.GP2.n3 VGND 0.050813f
C687 x2.GP2.t5 VGND 0.810542f
C688 x2.GP2.t4 VGND 0.833144f
C689 x2.GP2.n4 VGND 2.95587f
C690 x2.GP2.n5 VGND 0.106388f
.ends

