magic
tech sky130A
magscale 1 2
timestamp 1729128768
<< metal1 >>
rect 19478 1626 19758 2240
rect 19478 1346 20470 1626
rect 14060 858 14352 864
rect 14352 566 16056 858
rect 20190 570 20470 1346
rect 14060 560 14352 566
rect 15554 -116 15560 80
rect 15756 -116 15888 80
rect 20110 -198 20820 82
rect 22793 -155 28415 55
rect 14090 -726 14377 -720
rect 14377 -1013 15921 -726
rect 14090 -1019 14377 -1013
rect 14819 -1431 14825 -1365
rect 14891 -1431 17179 -1365
rect 14565 -1561 14571 -1495
rect 14637 -1561 17179 -1495
rect 17107 -2305 17173 -1609
rect 17107 -2377 17173 -2371
rect 13714 -3814 14338 -3614
rect 20110 -3652 20390 -198
rect 20664 -1288 20984 -1098
rect 20664 -1614 20984 -1608
rect 23069 -1780 23264 -155
rect 13714 -4693 13914 -3814
rect 18879 -3819 20390 -3652
rect 20110 -3822 20390 -3819
rect 20889 -1975 23264 -1780
rect 28205 -1809 28415 -155
rect 13714 -4893 14336 -4693
rect 20889 -4714 21084 -1975
rect 28205 -2025 28415 -2019
rect 18886 -4886 21084 -4714
rect 18886 -4887 20880 -4886
rect 13714 -5763 13914 -4893
rect 13714 -5963 14300 -5763
rect 18908 -5920 21290 -5816
rect 13714 -6821 13914 -5963
rect 13714 -7021 14298 -6821
rect 18931 -6936 20632 -6825
rect 20521 -11709 20632 -6936
rect 21186 -11476 21290 -5920
rect 21186 -11580 24870 -11476
rect 24974 -11580 24980 -11476
rect 20521 -11819 28547 -11709
rect 28657 -11819 28663 -11709
<< via1 >>
rect 20679 2379 20981 2681
rect 14060 566 14352 858
rect 15560 -116 15756 80
rect 14090 -1013 14377 -726
rect 14825 -1431 14891 -1365
rect 14571 -1561 14637 -1495
rect 17107 -2371 17173 -2305
rect 20664 -1608 20984 -1288
rect 28205 -2019 28415 -1809
rect 24870 -11580 24974 -11476
rect 28547 -11819 28657 -11709
<< metal2 >>
rect 20664 2681 20992 2690
rect 13851 2379 14131 2681
rect 14433 2379 14442 2681
rect 20664 2379 20679 2681
rect 20981 2379 20992 2681
rect 13881 858 14123 2379
rect 20664 2362 20992 2379
rect 13856 566 14060 858
rect 14352 566 14358 858
rect 13881 -726 14123 566
rect 13859 -1013 14090 -726
rect 14377 -1013 14383 -726
rect 13881 -3866 14124 -1013
rect 14551 -1495 14657 2117
rect 14797 -1365 14920 2099
rect 14797 -1431 14825 -1365
rect 14891 -1431 14920 -1365
rect 14797 -1459 14920 -1431
rect 15519 80 15797 89
rect 15519 -116 15560 80
rect 15756 -116 15797 80
rect 14551 -1561 14571 -1495
rect 14637 -1561 14657 -1495
rect 14551 -1581 14657 -1561
rect 15519 -1683 15797 -116
rect 20658 -1608 20664 -1288
rect 20984 -1608 20990 -1288
rect 15519 -1869 15565 -1683
rect 15751 -1869 15797 -1683
rect 15519 -1897 15797 -1869
rect 17107 -2305 17173 -2259
rect 17101 -2371 17107 -2305
rect 17173 -2371 17179 -2305
rect 20664 -2414 20984 -1608
rect 22070 -2393 22310 -1188
rect 23750 -2054 23887 2594
rect 28199 -2019 28205 -1809
rect 28415 -2019 28421 -1809
rect 22066 -2623 22075 -2393
rect 22305 -2623 22314 -2393
rect 22070 -2628 22310 -2623
rect 20664 -2743 20984 -2734
rect 13881 -4530 14262 -3866
rect 13881 -4950 14124 -4530
rect 13881 -5614 14266 -4950
rect 13881 -6028 14124 -5614
rect 13881 -6692 14278 -6028
rect 13881 -6964 14124 -6692
rect 13881 -7700 14236 -6964
rect 13881 -7744 14234 -7700
rect 13881 -10542 14124 -7744
rect 13881 -10545 14335 -10542
rect 13881 -10551 14340 -10545
rect 13881 -10784 14102 -10551
rect 14335 -10784 14340 -10551
rect 13881 -10788 14340 -10784
rect 14102 -10793 14335 -10788
rect 24870 -11476 24974 -11014
rect 24870 -11586 24974 -11580
rect 28547 -11709 28657 -11019
rect 28547 -11825 28657 -11819
<< via2 >>
rect 14131 2379 14433 2681
rect 20684 2384 20976 2676
rect 15565 -1869 15751 -1683
rect 20664 -2734 20984 -2414
rect 22075 -2623 22305 -2393
rect 14102 -10784 14335 -10551
<< metal3 >>
rect 14126 2681 14438 2686
rect 14126 2379 14131 2681
rect 14433 2676 20981 2681
rect 14433 2384 20684 2676
rect 20976 2384 20981 2676
rect 14433 2379 20981 2384
rect 14126 2374 14438 2379
rect 15514 -1678 15818 -1672
rect 15514 -1683 19874 -1678
rect 15514 -1869 15565 -1683
rect 15751 -1869 19874 -1683
rect 15514 -1874 19874 -1869
rect 15514 -2108 15818 -1874
rect 19678 -2532 19874 -1874
rect 22070 -2393 22310 -2388
rect 20659 -2414 20989 -2409
rect 20659 -2532 20664 -2414
rect 19678 -2728 20664 -2532
rect 19678 -2794 19874 -2728
rect 20659 -2734 20664 -2728
rect 20984 -2532 20989 -2414
rect 22070 -2532 22075 -2393
rect 20984 -2623 22075 -2532
rect 22305 -2532 22310 -2393
rect 22305 -2623 23452 -2532
rect 20984 -2728 23452 -2623
rect 29766 -2716 30104 -1679
rect 20984 -2734 20989 -2728
rect 20659 -2739 20989 -2734
rect 22070 -2750 22310 -2728
rect 19269 -2964 19874 -2794
rect 19678 -2968 19874 -2964
rect 14097 -10551 22748 -10546
rect 14097 -10784 14102 -10551
rect 14335 -10784 22748 -10551
rect 14097 -10789 22748 -10784
use ring  x1
timestamp 1725617623
transform 1 0 15830 0 1 242
box -220 -1240 4640 640
use driver  x2
timestamp 1725547227
transform 1 0 17793 0 1 -778
box 2790 -640 5210 3480
use mux4onehot_b  x3
timestamp 1728327329
transform 0 1 22092 -1 0 3487
box 4658 -8054 11287 -2405
use simplecounter  x4
timestamp 1729128768
transform 1 0 21380 0 1 -12570
box 750 982 9094 10886
<< labels >>
flabel metal3 15514 -2108 15818 -1672 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal3 29766 -2134 30104 -1679 0 FreeSans 1600 0 0 0 VSS
port 1 nsew
flabel metal3 14344 -10790 14698 -10550 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal3 14576 2386 14972 2676 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal1 19480 1950 19744 2218 0 FreeSans 1600 0 0 0 enable_ring
port 2 nsew
flabel metal2 23742 2414 23880 2590 0 FreeSans 1600 0 0 0 enable_counter
port 5 nsew
flabel metal2 14551 2001 14657 2107 0 FreeSans 1600 0 0 0 select0
port 3 nsew
flabel metal2 14797 1976 14920 2099 0 FreeSans 1600 0 0 0 select1
port 4 nsew
flabel metal1 13714 -5970 13914 -5770 0 FreeSans 1600 0 0 0 mux_out
port 6 nsew
flabel metal1 27990 -158 28270 52 0 FreeSans 1600 0 0 0 drv_out
flabel metal1 21176 -5906 21266 -5822 0 FreeSans 320 0 0 0 counter3
flabel metal1 20508 -6914 20598 -6830 0 FreeSans 320 0 0 0 counter7
flabel metal1 20172 -154 20376 28 0 FreeSans 320 0 0 0 ring_out
<< end >>
