* NGSPICE file created from tt_um_patdeegan_anamux_parax.ext - technology: sky130A

.subckt tt_um_patdeegan_anamux_parax clk ena rst_n ua[4] ua[5] ua[6] ua[7] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ ui_in[5] ua[0] ua[3] ui_in[1] ua[1] ui_in[4] ui_in[2] ui_in[6] ui_in[0] ua[2] ui_in[3]
+ VSS VDPWR
X0 a_21007_3867# ringtest_0.x4.net2.t2 VSS.t926 VSS.t925 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VSS.t899 VDPWR.t1166 VSS.t898 VSS.t897 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2 VSS.t901 VDPWR.t1167 VSS.t900 VSS.t671 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3 a_24527_5340# a_24361_5340# VSS.t165 VSS.t164 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 ua[2].t3 muxtest_0.x2.x2.GP1.t4 ua[3].t4 VDPWR.t314 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X5 ringtest_0.x4.clknet_0_clk.t15 a_23879_6940# VSS.t642 VSS.t641 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_24135_3867# ringtest_0.x4.net6.t2 VDPWR.t160 VDPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7 VSS.t1093 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t15 VSS.t1092 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VDPWR.t1046 ui_in[1].t0 muxtest_0.x1.x1.nSEL1 VDPWR.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 a_22399_8976# a_21852_8720# a_22052_8875# VDPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X10 muxtest_0.x1.x3.GP1.t3 muxtest_0.x1.x3.GN1 VDPWR.t73 VDPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_27491_4566# ringtest_0.x4._23_ ringtest_0.x4._09_ VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X12 VSS.t550 a_27065_5156# a_27233_5058# VSS.t549 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VDPWR.t1135 ringtest_0.x4._05_ a_24883_6800# VDPWR.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X14 VDPWR.t1039 a_16579_11759# ringtest_0.x3.x2.GN3 VDPWR.t1038 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X15 VDPWR.t754 VSS.t1127 VDPWR.t753 VDPWR.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X16 a_25309_5334# a_24527_5340# a_25225_5334# VDPWR.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_12019_24012# muxtest_0.x2.x1.nSEL1 VSS.t548 VSS.t547 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X18 a_26913_4566# ringtest_0.x4._15_ a_26817_4566# VSS.t575 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X19 VSS.t579 ringtest_0.x4._21_ a_24545_5878# VSS.t578 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 muxtest_0.x1.x3.GP4.t3 muxtest_0.x1.x3.GN4 VDPWR.t1011 VDPWR.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR.t77 VDPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 VDPWR.t361 ringtest_0.x4._15_ a_25925_6788# VDPWR.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_24004_6128# ringtest_0.x4._17_ a_23932_6128# VDPWR.t1143 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X24 VSS.t904 VDPWR.t1168 VSS.t903 VSS.t902 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X25 a_23467_4818# ringtest_0.x4._11_.t4 a_23381_4818# VSS.t854 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X26 a_19114_31955# a_19290_32287# a_19242_32347# VSS.t967 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 VSS.t906 VDPWR.t1169 VSS.t905 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X28 ringtest_0.x4.clknet_1_1__leaf_clk.t14 a_25364_5878# VSS.t1091 VSS.t1090 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 VDPWR.t963 a_21375_3867# ringtest_0.x4.counter[1] VDPWR.t962 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X30 VDPWR.t129 ringtest_0.x4.net5 a_22486_4246# VDPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X31 muxtest_0.x1.x1.nSEL0 ui_in[0].t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X32 VDPWR.t849 a_19842_32287# a_19666_31955# VDPWR.t848 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X33 muxtest_0.R3R4.t9 muxtest_0.x2.x2.GN3 ua[2].t11 VSS.t947 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X34 VDPWR.t751 VSS.t1128 VDPWR.t750 VDPWR.t749 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X35 a_12473_23980# ui_in[4].t0 VDPWR.t789 VDPWR.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X36 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP3 muxtest_0.R1R2.t1 VDPWR.t123 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X37 a_16579_11759# a_16755_12091# a_16707_12151# VSS.t929 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X38 VDPWR.t5 a_13501_23906# muxtest_0.x2.x2.GN4 VDPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X39 VDPWR.t219 a_19289_13081.t2 ringtest_0.drv_out.t18 VDPWR.t218 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X40 VSS.t5 a_21465_9294# ringtest_0.x4.net2.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X41 ringtest_0.x4.clknet_0_clk.t31 a_23879_6940# VDPWR.t425 VDPWR.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X42 VDPWR.t249 a_22021_4220# ringtest_0.x4._03_ VDPWR.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
X43 VSS.t304 ringtest_0.x4.net5 a_23467_4584# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X44 muxtest_0.x2.nselect2 VDPWR.t951 VDPWR.t953 VDPWR.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X45 a_16707_12151# ui_in[4].t1 VSS.t114 VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X46 VSS.t909 VDPWR.t1170 VSS.t908 VSS.t907 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X47 VDPWR.t748 VSS.t1129 VDPWR.t747 VDPWR.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X48 ringtest_0.x4._15_ a_23381_4584# VSS.t829 VSS.t828 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X49 a_23899_5334# ringtest_0.x4._15_ VDPWR.t359 VDPWR.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X50 VDPWR.t330 a_27065_5156# a_27233_5058# VDPWR.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X51 muxtest_0.x1.x3.GP3 muxtest_0.x1.x3.GN3 VDPWR.t852 VDPWR.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X52 VSS.t912 VDPWR.t1171 VSS.t911 VSS.t910 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X53 VSS.t993 ringtest_0.x4.net3.t2 ringtest_0.x4._12_ VSS.t992 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X54 VSS.t11 a_25975_3867# ringtest_0.x4.counter[6] VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X55 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk.t32 VDPWR.t1159 VDPWR.t1158 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X56 muxtest_0.x1.x5.A ui_in[2].t0 ua[3].t8 VDPWR.t772 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X57 ua[1].t1 ringtest_0.x3.x2.GP4.t4 ringtest_0.counter7.t1 VDPWR.t1094 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X58 a_22392_5990# a_22224_6244# VDPWR.t921 VDPWR.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X59 ringtest_0.x4.clknet_1_0__leaf_clk.t31 a_21395_6940# VDPWR.t1086 VDPWR.t1085 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X60 VSS.t1017 ringtest_0.x4._22_ a_26913_4566# VSS.t1016 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X61 a_26640_5334# a_26367_5340# a_26555_5334# VDPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X62 ringtest_0.x4.clknet_1_1__leaf_clk.t31 a_25364_5878# VDPWR.t1131 VDPWR.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X63 VDPWR.t746 VSS.t1130 VDPWR.t745 VDPWR.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X64 VSS.t39 VDPWR.t1172 VSS.t38 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X65 a_21785_8054# ringtest_0.x4.net3.t3 VDPWR.t1018 VDPWR.t1017 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X66 ringtest_0.x4._17_ a_25925_6788# VSS.t479 VSS.t478 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X67 VSS.t359 a_19114_31955# muxtest_0.x1.x3.GN2 VSS.t358 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VDPWR.t183 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR.t182 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X69 VDPWR.t950 VDPWR.t948 ringtest_0.x3.nselect2 VDPWR.t949 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X70 VDPWR.t423 a_23879_6940# ringtest_0.x4.clknet_0_clk.t30 VDPWR.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X71 VSS.t856 ringtest_0.x4.net4 ringtest_0.x4._13_ VSS.t855 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 a_24317_4942# ringtest_0.x4.net6.t3 a_24551_4790# VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X73 VSS.t723 ringtest_0.x4.clknet_0_clk.t32 a_25364_5878# VSS.t722 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X74 VSS.t127 a_22111_10993# ringtest_0.x4.net1 VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X75 VSS.t42 VDPWR.t1173 VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X76 VDPWR.t141 a_27815_3867# ringtest_0.x4.counter[8] VDPWR.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X77 ringtest_0.x4._00_ a_21425_9686# a_21675_9686# VDPWR.t857 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X78 VDPWR.t743 VSS.t1131 VDPWR.t742 VDPWR.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X79 VDPWR.t741 VSS.t1132 VDPWR.t740 VDPWR.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X80 VDPWR.t841 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X81 VDPWR.t175 ringtest_0.x4._00_ a_22399_9142# VDPWR.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X82 VSS.t640 a_23879_6940# ringtest_0.x4.clknet_0_clk.t14 VSS.t639 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X83 a_21675_4790# a_21509_4790# VSS.t557 VSS.t556 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X84 VSS.t1055 ui_in[0].t1 a_19842_32287# VSS.t1054 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 VSS.t45 VDPWR.t1174 VSS.t44 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X86 VDPWR.t1084 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t30 VDPWR.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X87 VSS.t136 a_23399_3867# ringtest_0.counter3.t2 VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X88 VDPWR.t286 a_18662_32213# muxtest_0.x1.x3.GN1 VDPWR.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X89 VDPWR.t941 ringtest_0.x4.net2.t3 a_21507_9686# VDPWR.t940 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 VDPWR.t738 VSS.t1133 VDPWR.t737 VDPWR.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X91 a_27659_4246# ringtest_0.x4.net11 VDPWR.t809 VDPWR.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X92 a_22390_4566# ringtest_0.x4.net5 VSS.t302 VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X93 ringtest_0.x3.x1.nSEL1 ui_in[4].t2 VSS.t116 VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X94 ringtest_0.x4.clknet_1_0__leaf_clk.t15 a_21395_6940# VSS.t1051 VSS.t1050 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X95 a_22649_6244# a_21785_5878# a_22392_5990# VDPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X96 muxtest_0.x1.x3.GP2.t3 muxtest_0.x1.x3.GN2 VDPWR.t179 VDPWR.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X97 ua[3].t9 ui_in[2].t1 muxtest_0.x1.x4.A VSS.t662 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X98 muxtest_0.R5R6.t5 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A VSS.t838 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X99 VSS.t965 a_24329_6640# a_24336_6544# VSS.t964 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X100 a_27303_4246# a_27273_4220# ringtest_0.x4._09_ VDPWR.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X101 VDPWR.t735 VSS.t1134 VDPWR.t734 VDPWR.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X102 ringtest_0.x4.clknet_1_0__leaf_clk.t29 a_21395_6940# VDPWR.t1082 VDPWR.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X103 VSS.t924 ringtest_0.x4.net2.t4 a_21425_9686# VSS.t923 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X104 a_19666_31955# a_19842_32287# a_19794_32347# VSS.t830 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X105 muxtest_0.R3R4.t1 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A VSS.t155 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X106 VDPWR.t885 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X107 a_21845_8816# ringtest_0.x4.clknet_1_0__leaf_clk.t32 VDPWR.t1014 VDPWR.t1013 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X108 VSS.t1049 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t14 VSS.t1048 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X109 a_21672_5334# a_21399_5340# a_21587_5334# VDPWR.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X110 ringtest_0.x4.clknet_1_1__leaf_clk.t30 a_25364_5878# VDPWR.t1129 VDPWR.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X111 VDPWR.t732 VSS.t1135 VDPWR.t731 VDPWR.t730 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X112 a_18662_32213# muxtest_0.x1.x1.nSEL0 a_18836_32319# VSS.t648 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X113 a_16203_12091# ui_in[4].t3 VDPWR.t113 VDPWR.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X114 a_19794_32347# ui_in[1].t1 VSS.t752 VSS.t751 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X115 VDPWR.t729 VSS.t1136 VDPWR.t728 VDPWR.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X116 VDPWR.t813 a_22817_6146# a_22733_6244# VDPWR.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X117 VDPWR.t207 a_17231_12017# ringtest_0.x3.x2.GN4 VDPWR.t206 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X118 VDPWR.t421 a_23879_6940# ringtest_0.x4.clknet_0_clk.t29 VDPWR.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X119 VSS.t1089 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t13 VSS.t1088 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X120 ringtest_0.x3.nselect2 VDPWR.t945 VDPWR.t947 VDPWR.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X121 a_25925_6788# ringtest_0.x4.net6.t4 VDPWR.t162 VDPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X122 a_25975_3867# ringtest_0.x4.net8 VDPWR.t802 VDPWR.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X123 ringtest_0.x4.net10 a_27233_5308# VDPWR.t832 VDPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X124 a_11845_23906# muxtest_0.x2.x1.nSEL1 VDPWR.t329 VDPWR.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X125 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VSS.t514 VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X126 VDPWR.t276 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X127 a_21939_8054# ringtest_0.x4.net3.t4 a_21867_8054# VSS.t994 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X128 a_26721_4246# ringtest_0.x4.net10 a_26627_4246# VDPWR.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X129 a_22116_4902# a_21948_5156# VSS.t847 VSS.t846 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X130 VDPWR.t1080 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t28 VDPWR.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X131 a_25149_4220# ringtest_0.x4.net7 VDPWR.t228 VDPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X132 VDPWR.t891 a_21840_5308# a_21767_5334# VDPWR.t890 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X133 VSS.t48 VDPWR.t1175 VSS.t47 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X134 VSS.t51 VDPWR.t1176 VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X135 VDPWR.t173 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X136 VDPWR.t726 VSS.t1137 VDPWR.t725 VDPWR.t724 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X137 a_24627_6200# ringtest_0.x4._21_ VDPWR.t365 VDPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X138 VSS.t658 ringtest_0.x4._16_.t2 a_24986_5878# VSS.t657 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.06615 ps=0.735 w=0.42 l=0.15
X139 VSS.t54 VDPWR.t1177 VSS.t53 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X140 VDPWR.t349 a_22245_8054# ringtest_0.x4._11_.t3 VDPWR.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X141 a_25977_4220# ringtest_0.x4._11_.t5 VDPWR.t1041 VDPWR.t1040 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X142 VSS.t57 VDPWR.t1178 VSS.t56 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X143 a_26367_4790# a_26201_4790# VSS.t321 VSS.t320 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X144 VDPWR.t723 VSS.t1138 VDPWR.t722 VDPWR.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X145 a_25677_5156# a_24895_4790# a_25593_5156# VDPWR.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 VDPWR.t1142 ringtest_0.x4._17_ a_23349_6422# VDPWR.t1141 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 VDPWR.t357 ringtest_0.x4._15_ a_25977_4220# VDPWR.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X148 VDPWR.t721 VSS.t1139 VDPWR.t720 VDPWR.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X149 VDPWR.t187 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2.t3 VDPWR.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X150 VDPWR.t309 a_24070_5852# a_24004_6128# VDPWR.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X151 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP2.t4 muxtest_0.R6R7.t1 VDPWR.t13 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X152 ua[0].t1 muxtest_0.x2.x2.GN2 ua[2].t1 VSS.t357 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X153 VSS.t587 a_25977_4220# ringtest_0.x4._23_ VSS.t586 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X154 VDPWR.t719 VSS.t1140 VDPWR.t718 VDPWR.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X155 VDPWR.t716 VSS.t1141 VDPWR.t715 VDPWR.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X156 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VSS.t351 VSS.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X157 VDPWR.t87 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X158 a_21425_9686# ringtest_0.x4.net1 VSS.t134 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X159 VSS.t721 a_24317_4942# ringtest_0.x4._20_ VSS.t720 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X160 muxtest_0.x1.x1.nSEL1 ui_in[1].t2 VDPWR.t815 VDPWR.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X161 a_21465_8830# a_21561_8830# VSS.t970 VSS.t881 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X162 ringtest_0.x4.clknet_0_clk.t13 a_23879_6940# VSS.t638 VSS.t637 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X163 a_22295_3867# ringtest_0.x4.net4 VDPWR.t875 VDPWR.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X164 muxtest_0.R7R8.t9 muxtest_0.R6R7.t5 VSS.t643 sky130_fd_pr__res_high_po_1p41 l=1.75
X165 VDPWR.t713 VSS.t1142 VDPWR.t712 VDPWR.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X166 a_26808_4902# a_26640_5156# VDPWR.t199 VDPWR.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X167 VSS.t60 VDPWR.t1179 VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X168 ringtest_0.x4.clknet_1_1__leaf_clk.t29 a_25364_5878# VDPWR.t1127 VDPWR.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X169 VSS.t731 a_26808_5308# a_26766_5712# VSS.t730 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X170 a_25351_5712# a_24361_5340# a_25225_5334# VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X171 VSS.t1047 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t13 VSS.t1046 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X172 VSS.t63 VDPWR.t1180 VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X173 muxtest_0.R7R8.t8 muxtest_0.x2.x2.GN4 ua[2].t13 VSS.t961 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X174 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VSS.t776 VSS.t503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X175 VSS.t66 VDPWR.t1181 VSS.t65 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X176 a_21007_3867# ringtest_0.x4.net2.t5 VDPWR.t939 VDPWR.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X177 ringtest_0.x4.net4 a_22265_5308# VDPWR.t215 VDPWR.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X178 VDPWR.t895 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X179 VSS.t391 a_19289_13081.t3 ringtest_0.drv_out.t10 VSS.t390 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X180 a_22373_5156# a_21509_4790# a_22116_4902# VDPWR.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X181 VDPWR.t710 VSS.t1143 VDPWR.t709 VDPWR.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X182 a_26895_3867# ringtest_0.x4.net9 VSS.t522 VSS.t521 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X183 a_27191_4790# a_26201_4790# a_27065_5156# VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X184 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR.t845 VDPWR.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X185 VDPWR.t708 VSS.t1144 VDPWR.t707 VDPWR.t489 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X186 VSS.t69 VDPWR.t1182 VSS.t68 VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X187 a_22116_4902# a_21948_5156# VDPWR.t863 VDPWR.t862 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X188 VSS.t738 ringtest_0.x4.net8 a_23837_5878# VSS.t737 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X189 VDPWR.t1078 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t27 VDPWR.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X190 a_16755_12091# ui_in[3].t0 VDPWR.t131 VDPWR.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X191 VDPWR.t1125 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t28 VDPWR.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X192 VDPWR.t1138 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 VDPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X193 ringtest_0.x4.clknet_1_0__leaf_clk.t12 a_21395_6940# VSS.t1045 VSS.t1044 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X194 VSS.t72 VDPWR.t1183 VSS.t71 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X195 VSS.t161 a_21007_3867# ringtest_0.x4.counter[0] VSS.t160 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X196 a_22181_5334# a_21399_5340# a_22097_5334# VDPWR.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X197 a_20318_32213# ui_in[1].t3 a_20492_32319# VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X198 VSS.t339 ringtest_0.x4._00_ a_22399_9142# VSS.t338 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X199 a_22224_6244# a_21951_5878# a_22139_5878# VDPWR.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X200 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VSS.t535 VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X201 VSS.t532 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1.t1 VSS.t531 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X202 VDPWR.t127 ringtest_0.x4.net5 a_23381_4584# VDPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 a_26555_5334# ringtest_0.x4._08_ VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X204 ua[2].t5 muxtest_0.x2.x2.GP3 muxtest_0.R3R4.t3 VDPWR.t282 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X205 a_16027_11759# ui_in[3].t1 VDPWR.t56 VDPWR.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X206 VDPWR.t205 a_22541_5058# a_22457_5156# VDPWR.t204 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X207 ringtest_0.x4.clknet_1_1__leaf_clk.t12 a_25364_5878# VSS.t1087 VSS.t1086 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X208 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VSS.t866 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X209 ringtest_0.x4._19_ a_23529_6422# VSS.t93 VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X210 a_26569_6422# ringtest_0.x4._23_ VSS.t607 VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X211 a_24895_4790# a_24729_4790# VDPWR.t144 VDPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X212 VDPWR.t313 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 ringtest_0.ring_out.t4 ringtest_0.x3.x2.GN1 ua[1].t9 VSS.t530 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X214 ringtest_0.drv_out.t9 a_19289_13081.t4 VSS.t393 VSS.t392 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X215 a_23899_5334# ringtest_0.x4.net6.t5 VDPWR.t1026 VDPWR.t1025 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X216 VDPWR.t706 VSS.t1145 VDPWR.t705 VDPWR.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X217 a_24045_6654# a_24336_6544# a_24287_6422# VDPWR.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X218 a_24800_5334# a_24527_5340# a_24715_5334# VDPWR.t816 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X219 muxtest_0.R7R8.t1 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A VSS.t154 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X220 muxtest_0.x2.x2.GP3 muxtest_0.x2.x2.GN3 VSS.t946 VSS.t945 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X221 VSS.t75 VDPWR.t1184 VSS.t74 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X222 a_25925_6788# ringtest_0.x4._11_.t6 VDPWR.t1043 VDPWR.t1042 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X223 ringtest_0.x4.net10 a_27233_5308# VSS.t769 VSS.t768 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X224 VSS.t870 a_21840_5308# a_21798_5712# VSS.t869 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X225 VSS.t140 ui_in[3].t2 muxtest_0.x2.x1.nSEL0 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X226 VDPWR.t703 VSS.t1146 VDPWR.t702 VDPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X227 VDPWR.t1054 a_22392_5990# a_22319_6244# VDPWR.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X228 VSS.t78 VDPWR.t1185 VSS.t77 VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X229 VSS.t477 a_15575_12017# ringtest_0.x3.x2.GN1 VSS.t476 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X230 a_22201_9142# a_21981_9142# VSS.t335 VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X231 ringtest_0.counter7.t3 ringtest_0.x3.x2.GN4 ua[1].t6 VSS.t383 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X232 VDPWR.t226 ringtest_0.x4.net7 a_25925_6788# VDPWR.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X233 VDPWR.t8 a_25975_3867# ringtest_0.x4.counter[6] VDPWR.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X234 VSS.t725 ringtest_0.x4.clknet_0_clk.t33 a_25364_5878# VSS.t724 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X235 VDPWR.t701 VSS.t1147 VDPWR.t700 VDPWR.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X236 VSS.t727 ringtest_0.x4.clknet_0_clk.t34 a_21395_6940# VSS.t726 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X237 a_19114_31955# ui_in[0].t2 VDPWR.t1090 VDPWR.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X238 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VSS.t466 VSS.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X239 VDPWR.t698 VSS.t1148 VDPWR.t697 VDPWR.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X240 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR.t893 VDPWR.t892 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X241 VDPWR.t881 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2.t3 VDPWR.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X242 VDPWR.t1016 ringtest_0.x4.clknet_1_0__leaf_clk.t33 a_21509_4790# VDPWR.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X243 VDPWR.t695 VSS.t1149 VDPWR.t694 VDPWR.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X244 a_21803_9508# a_21465_9294# VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X245 a_22052_9116# a_21852_9416# a_22201_9142# VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X246 VSS.t81 VDPWR.t1186 VSS.t80 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X247 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VSS.t504 VSS.t503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X248 ringtest_0.x4._12_ ringtest_0.x4.net2.t6 a_21132_8918# VSS.t922 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X249 a_22052_8875# a_21852_8720# a_22201_8964# VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X250 a_27065_5156# a_26201_4790# a_26808_4902# VDPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X251 ringtest_0.x4.clknet_1_0__leaf_clk.t11 a_21395_6940# VSS.t1043 VSS.t1042 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X252 a_21587_5334# ringtest_0.x4._02_ VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X253 VSS.t1057 ui_in[0].t3 muxtest_0.x1.x1.nSEL0 VSS.t1056 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X254 VSS.t84 VDPWR.t1187 VSS.t83 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X255 VDPWR.t1 a_21465_9294# ringtest_0.x4.net2.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X256 ringtest_0.x4._25_ a_26749_6422# VDPWR.t268 VDPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X257 VDPWR.t52 a_23399_3867# ringtest_0.counter3.t3 VDPWR.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X258 VDPWR.t1123 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t27 VDPWR.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X259 muxtest_0.x2.x2.GP2.t1 muxtest_0.x2.x2.GN2 VSS.t356 VSS.t355 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X260 ringtest_0.x3.x2.GP1.t0 ringtest_0.x3.x2.GN1 VSS.t529 VSS.t528 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X261 VSS.t87 VDPWR.t1188 VSS.t86 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X262 VDPWR.t693 VSS.t1150 VDPWR.t692 VDPWR.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X263 a_26817_4566# ringtest_0.x4._11_.t7 a_26627_4246# VSS.t1012 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X264 a_22649_6244# a_21951_5878# a_22392_5990# VSS.t740 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X265 VDPWR.t850 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 VDPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X266 VDPWR.t691 VSS.t1151 VDPWR.t690 VDPWR.t536 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X267 VSS.t331 a_21845_9116# a_21852_9416# VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X268 a_21591_6128# ringtest_0.x4._11_.t8 ringtest_0.x4._13_ VDPWR.t1044 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X269 VDPWR.t355 ringtest_0.x4._15_ a_23381_4818# VDPWR.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X270 a_21981_9142# a_21845_9116# a_21561_9116# VDPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X271 VDPWR.t689 VSS.t1152 VDPWR.t688 VDPWR.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X272 VSS.t1085 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t11 VSS.t1084 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X273 VSS.t153 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1.t1 VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X274 muxtest_0.R6R7.t3 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A VSS.t347 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X275 VDPWR.t686 VSS.t1153 VDPWR.t685 VDPWR.t684 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X276 ringtest_0.x4.clknet_0_clk.t12 a_23879_6940# VSS.t636 VSS.t635 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X277 VDPWR.t1145 a_27233_5058# a_27149_5156# VDPWR.t829 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X278 VDPWR.t683 VSS.t1154 VDPWR.t682 VDPWR.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X279 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VSS.t177 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X280 VDPWR.t680 VSS.t1155 VDPWR.t679 VDPWR.t678 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X281 ringtest_0.x4.clknet_1_1__leaf_clk.t26 a_25364_5878# VDPWR.t1121 VDPWR.t1120 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X282 a_26839_6788# a_26569_6422# a_26749_6422# VSS.t850 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X283 VSS.t90 VDPWR.t1189 VSS.t89 VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X284 VSS.t1041 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t10 VSS.t1040 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X285 VSS.t673 VDPWR.t1190 VSS.t672 VSS.t671 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X286 ringtest_0.x4.net8 a_25393_5308# VDPWR.t384 VDPWR.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X287 VSS.t991 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP4.t1 VSS.t990 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X288 a_24479_4790# ringtest_0.x4.net8 VSS.t736 VSS.t735 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X289 ringtest_0.x4.net9 a_25761_5058# VSS.t539 VSS.t538 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X290 a_27191_5712# a_26201_5340# a_27065_5334# VSS.t656 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X291 VSS.t605 ringtest_0.x4._23_ a_27273_4220# VSS.t604 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X292 a_25593_5156# a_24895_4790# a_25336_4902# VSS.t650 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X293 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR.t171 VDPWR.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X294 VSS.t746 ringtest_0.x4.net11 a_27489_3702# VSS.t745 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X295 ringtest_0.drv_out.t8 a_19289_13081.t5 VSS.t395 VSS.t394 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X296 ringtest_0.x3.x2.GP3 ringtest_0.x3.x2.GN3 VSS.t1102 VSS.t1101 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X297 VSS.t676 VDPWR.t1191 VSS.t675 VSS.t674 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X298 ringtest_0.counter3.t5 ringtest_0.x3.x2.GN3 ua[1].t14 VSS.t1100 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X299 ringtest_0.x4.clknet_0_clk.t28 a_23879_6940# VDPWR.t419 VDPWR.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X300 a_24699_6200# ringtest_0.x4.net9 a_24627_6200# VDPWR.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0441 ps=0.63 w=0.42 l=0.15
X301 VSS.t679 VDPWR.t1192 VSS.t678 VSS.t677 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X302 VDPWR.t677 VSS.t1156 VDPWR.t676 VDPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X303 VSS.t681 VDPWR.t1193 muxtest_0.x2.nselect2 VSS.t680 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X304 ringtest_0.x4.clknet_1_0__leaf_clk.t9 a_21395_6940# VSS.t1039 VSS.t1038 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X305 a_24264_6788# a_23949_6654# VSS.t593 VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X306 VSS.t146 a_24135_3867# ringtest_0.x4.counter[4] VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X307 VSS.t684 VDPWR.t1194 VSS.t683 VSS.t682 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X308 VDPWR.t784 ringtest_0.x4.clknet_1_1__leaf_clk.t33 a_26201_4790# VDPWR.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X309 a_21465_8830# a_21561_8830# VDPWR.t993 VDPWR.t992 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X310 a_19666_31955# ui_in[1].t4 VDPWR.t105 VDPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X311 VDPWR.t177 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2.t2 VDPWR.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X312 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP2.t5 muxtest_0.R6R7.t0 VDPWR.t67 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X313 ua[0].t8 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A VSS.t989 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X314 ringtest_0.x4.net5 a_22541_5058# VSS.t375 VSS.t374 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X315 VSS.t944 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 VSS.t943 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X316 VDPWR.t217 a_16027_11759# ringtest_0.x3.x2.GN2 VDPWR.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X317 VDPWR.t1119 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t25 VDPWR.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X318 VSS.t687 VDPWR.t1195 VSS.t686 VSS.t685 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X319 a_21395_6940# ringtest_0.x4.clknet_0_clk.t35 VSS.t664 VSS.t663 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X320 a_23949_6654# a_24045_6654# VDPWR.t54 VDPWR.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X321 VDPWR.t786 ringtest_0.x4.clknet_1_1__leaf_clk.t34 a_24361_5340# VDPWR.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X322 VDPWR.t193 a_23770_5308# ringtest_0.x4._18_ VDPWR.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X323 VSS.t976 a_22765_4478# ringtest_0.x4._14_ VSS.t975 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X324 VDPWR.t369 ringtest_0.ring_out.t10 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X325 VSS.t981 ringtest_0.x4._10_ a_22245_8054# VSS.t980 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X326 a_21675_10006# ringtest_0.x4.net2.t7 VSS.t921 VSS.t920 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X327 VSS.t147 a_22052_8875# a_21981_8976# VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X328 ringtest_0.x4.net9 a_25761_5058# VDPWR.t319 VDPWR.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X329 VDPWR.t675 VSS.t1157 VDPWR.t674 VDPWR.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X330 VSS.t758 a_19289_13081.t6 ringtest_0.drv_out.t7 VSS.t757 sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X331 VSS.t978 a_24968_5308# a_24926_5712# VSS.t977 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X332 VSS.t290 ui_in[1].t5 muxtest_0.x1.x1.nSEL1 VSS.t289 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X333 muxtest_0.x1.x3.GP1.t0 muxtest_0.x1.x3.GN1 VSS.t151 VSS.t150 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X334 a_16027_11759# a_16203_12091# a_16155_12151# VSS.t366 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X335 ringtest_0.x4.clknet_0_clk.t11 a_23879_6940# VSS.t634 VSS.t633 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X336 VDPWR.t48 ringtest_0.x4.net1 a_21049_8598# VDPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X337 VDPWR.t672 VSS.t1158 VDPWR.t671 VDPWR.t670 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X338 VSS.t690 VDPWR.t1196 VSS.t689 VSS.t688 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X339 VSS.t526 a_20318_32213# muxtest_0.x1.x3.GN4 VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X340 muxtest_0.x2.x1.nSEL0 ui_in[3].t3 VDPWR.t58 VDPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X341 a_16155_12151# ui_in[3].t4 VSS.t142 VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X342 a_26269_4612# ringtest_0.x4._15_ a_26173_4612# VSS.t574 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X343 VDPWR.t669 VSS.t1159 VDPWR.t668 VDPWR.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X344 VDPWR.t666 VSS.t1160 VDPWR.t665 VDPWR.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X345 VSS.t1037 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t8 VSS.t1036 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X346 a_25149_4220# ringtest_0.x4.net9 VDPWR.t298 VDPWR.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X347 a_22223_5712# a_21233_5340# a_22097_5334# VSS.t951 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X348 muxtest_0.x1.x3.GP4.t0 muxtest_0.x1.x3.GN4 VSS.t988 VSS.t987 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X349 VSS.t692 VDPWR.t1197 VSS.t691 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X350 VSS.t695 VDPWR.t1198 VSS.t694 VSS.t693 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X351 ringtest_0.x4.net5 a_22541_5058# VDPWR.t203 VDPWR.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X352 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR.t85 VDPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X353 VSS.t698 VDPWR.t1199 VSS.t697 VSS.t696 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X354 VSS.t287 ringtest_0.x4._11_.t9 ringtest_0.x4._01_ VSS.t286 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X355 a_22765_5308# ringtest_0.x4._16_.t3 a_23151_5334# VDPWR.t771 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X356 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP1.t4 muxtest_0.R7R8.t4 VDPWR.t1035 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X357 a_25977_4220# ringtest_0.x4._22_ VDPWR.t1052 VDPWR.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X358 a_25083_4790# ringtest_0.x4._07_ VDPWR.t1161 VDPWR.t1160 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 VSS.t701 VDPWR.t1200 VSS.t700 VSS.t699 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X360 VDPWR.t663 VSS.t1161 VDPWR.t662 VDPWR.t661 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X361 a_22983_5654# ringtest_0.x4._16_.t4 ringtest_0.x4._04_ VSS.t659 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X362 VSS.t704 VDPWR.t1201 VSS.t703 VSS.t702 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X363 VDPWR.t60 ui_in[3].t5 ringtest_0.x3.x1.nSEL0 VDPWR.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X364 a_23879_6940# ringtest_0.drv_out.t20 VDPWR.t1020 VDPWR.t1019 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X365 a_22164_4362# ringtest_0.x4._16_.t5 VSS.t1114 VSS.t1113 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X366 a_25168_5156# a_24729_4790# a_25083_4790# VSS.t316 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X367 VDPWR.t660 VSS.t1162 VDPWR.t659 VDPWR.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X368 VSS.t1019 a_22392_5990# a_22350_5878# VSS.t1018 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X369 VDPWR.t756 ringtest_0.x4._20_ a_23809_4790# VDPWR.t755 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X370 muxtest_0.x2.nselect2 VDPWR.t1202 VSS.t706 VSS.t705 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X371 a_21780_8964# a_21465_8830# VSS.t972 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X372 ringtest_0.x4._11_.t1 a_22245_8054# VSS.t567 VSS.t566 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X373 a_26895_3867# ringtest_0.x4.net9 VDPWR.t296 VDPWR.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X374 a_24715_5334# ringtest_0.x4._06_ VSS.t120 VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X375 VSS.t708 VDPWR.t1203 VSS.t707 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X376 VDPWR.t99 ringtest_0.x4._11_.t10 a_23899_5334# VDPWR.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X377 VDPWR.t1117 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t24 VDPWR.t1116 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X378 VDPWR.t332 a_25421_6641# ringtest_0.x4._05_ VDPWR.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X379 muxtest_0.x1.x3.GP3 muxtest_0.x1.x3.GN3 VSS.t837 VSS.t836 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X380 muxtest_0.x1.x4.A muxtest_0.x1.x5.GN ua[3].t3 VDPWR.t119 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X381 ua[2].t2 muxtest_0.x2.x2.GP1.t5 ua[3].t5 VDPWR.t315 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X382 ua[0].t0 muxtest_0.x2.x2.GN2 ua[2].t0 VSS.t354 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X383 a_25294_4790# a_24895_4790# a_25168_5156# VSS.t649 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X384 a_21863_4790# ringtest_0.x4._03_ VDPWR.t251 VDPWR.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X385 VDPWR.t657 VSS.t1163 VDPWR.t656 VDPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X386 VDPWR.t79 a_21007_3867# ringtest_0.x4.counter[0] VDPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X387 VSS.t711 VDPWR.t1204 VSS.t710 VSS.t709 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X388 a_21948_5156# a_21509_4790# a_21863_4790# VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X389 VSS.t714 VDPWR.t1205 VSS.t713 VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X390 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.ring_out.t11 VDPWR.t371 VDPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X391 VSS.t744 ringtest_0.x4.net11 a_27491_4566# VSS.t743 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X392 ringtest_0.x4.net11 a_27233_5058# VSS.t1112 VSS.t1111 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X393 ringtest_0.x4._21_ a_23809_4790# VDPWR.t33 VDPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X394 VSS.t349 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X395 VSS.t716 VDPWR.t1206 ringtest_0.x3.nselect2 VSS.t715 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X396 VDPWR.t919 ringtest_0.x4._01_ a_22399_8976# VDPWR.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X397 VDPWR.t417 a_23879_6940# ringtest_0.x4.clknet_0_clk.t27 VDPWR.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X398 a_25149_4220# ringtest_0.x4.net6.t6 a_25547_4612# VSS.t1000 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X399 ringtest_0.x4.net8 a_25393_5308# VSS.t603 VSS.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X400 VSS.t844 a_21425_9686# ringtest_0.x4._00_ VSS.t843 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X401 VSS.t589 a_25336_4902# a_25294_4790# VSS.t588 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X402 VDPWR.t415 a_23879_6940# ringtest_0.x4.clknet_0_clk.t26 VDPWR.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X403 ua[2].t8 muxtest_0.x2.x2.GP4.t4 muxtest_0.R7R8.t5 VDPWR.t762 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X404 a_22139_5878# ringtest_0.x4._04_ VSS.t955 VSS.t954 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X405 ringtest_0.x3.x2.GP2.t2 ringtest_0.x3.x2.GN2 VDPWR.t879 VDPWR.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X406 ringtest_0.x4.clknet_0_clk.t10 a_23879_6940# VSS.t632 VSS.t631 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X407 a_25977_4220# ringtest_0.x4.net10 a_26375_4612# VSS.t774 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X408 VSS.t719 VDPWR.t1207 VSS.t718 VSS.t717 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X409 VSS.t553 a_25421_6641# ringtest_0.x4._05_ VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X410 VDPWR.t969 ringtest_0.x4._24_ a_26749_6422# VDPWR.t968 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X411 VSS.t610 ringtest_0.x4.clknet_1_0__leaf_clk.t34 a_21785_5878# VSS.t609 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X412 VSS.t775 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 VDPWR.t820 a_19289_13081.t7 ringtest_0.drv_out.t17 VDPWR.t819 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X414 a_22021_4220# a_22164_4362# VDPWR.t266 VDPWR.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X415 VDPWR.t843 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR.t842 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X416 VSS.t781 VDPWR.t1208 VSS.t780 VSS.t779 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X417 VDPWR.t101 ringtest_0.x4._11_.t11 a_23809_4790# VDPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X418 ua[3].t11 muxtest_0.x2.x2.GN1 ua[2].t15 VSS.t1126 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X419 VDPWR.t655 VSS.t1164 VDPWR.t654 VDPWR.t653 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X420 a_19242_32347# ui_in[0].t4 VSS.t1059 VSS.t1058 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X421 muxtest_0.x1.x3.GP2.t1 muxtest_0.x1.x3.GN2 VSS.t346 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X422 ringtest_0.x4.clknet_1_0__leaf_clk.t7 a_21395_6940# VSS.t1035 VSS.t1034 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X423 VSS.t941 ringtest_0.x4._24_ a_26839_6788# VSS.t940 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X424 VDPWR.t391 ringtest_0.x4.clknet_1_0__leaf_clk.t35 a_21785_5878# VDPWR.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X425 VSS.t760 a_19289_13081.t8 ringtest_0.drv_out.t6 VSS.t759 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X426 VDPWR.t652 VSS.t1165 VDPWR.t651 VDPWR.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X427 ringtest_0.x4.net11 a_27233_5058# VDPWR.t1144 VDPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X428 muxtest_0.x2.x1.nSEL1 ui_in[4].t4 VDPWR.t115 VDPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X429 a_15575_12017# ringtest_0.x3.x1.nSEL0 a_15749_12123# VSS.t966 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X430 a_25083_4790# ringtest_0.x4._07_ VSS.t1120 VSS.t1119 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X431 VDPWR.t111 a_19666_31955# muxtest_0.x1.x3.GN3 VDPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X432 VSS.t939 ringtest_0.x4._14_ ringtest_0.x4._02_ VSS.t938 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 muxtest_0.R1R2.t2 ua[0].t4 VSS.t467 sky130_fd_pr__res_high_po_1p41 l=1.75
X434 VSS.t784 VDPWR.t1209 VSS.t783 VSS.t782 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X435 VSS.t630 a_23879_6940# ringtest_0.x4.clknet_0_clk.t9 VSS.t629 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X436 VSS.t670 ringtest_0.x4.clknet_1_1__leaf_clk.t35 a_24729_4790# VSS.t669 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X437 a_26808_5308# a_26640_5334# VSS.t756 VSS.t755 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X438 VDPWR.t1115 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t23 VDPWR.t1114 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X439 VDPWR.t649 VSS.t1166 VDPWR.t648 VDPWR.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X440 VDPWR.t647 VSS.t1167 VDPWR.t646 VDPWR.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X441 VSS.t787 VDPWR.t1210 VSS.t786 VSS.t785 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X442 VSS.t790 VDPWR.t1211 VSS.t789 VSS.t788 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X443 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP4.t4 muxtest_0.R4R5.t2 VDPWR.t956 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X444 VDPWR.t873 ringtest_0.x4.net4 a_21591_6128# VDPWR.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X445 a_21055_5334# ringtest_0.x4._13_ VDPWR.t877 VDPWR.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X446 VDPWR.t288 a_11845_23906# muxtest_0.x2.x2.GN1 VDPWR.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X447 VSS.t865 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X448 VDPWR.t645 VSS.t1168 VDPWR.t644 VDPWR.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X449 a_21395_6940# ringtest_0.x4.clknet_0_clk.t36 VSS.t666 VSS.t665 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X450 VDPWR.t800 ringtest_0.x4.net8 a_25149_4220# VDPWR.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X451 ringtest_0.drv_out.t16 a_19289_13081.t9 VDPWR.t822 VDPWR.t821 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X452 VDPWR.t889 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR.t888 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X453 VDPWR.t642 VSS.t1169 VDPWR.t641 VDPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X454 a_25168_5156# a_24895_4790# a_25083_4790# VDPWR.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X455 VDPWR.t787 ringtest_0.x4.clknet_1_1__leaf_clk.t36 a_26201_5340# VDPWR.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X456 VDPWR.t1028 ringtest_0.x4.net6.t7 a_22795_5334# VDPWR.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X457 a_25364_5878# ringtest_0.x4.clknet_0_clk.t37 VDPWR.t782 VDPWR.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X458 a_21863_4790# ringtest_0.x4._03_ VSS.t471 VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X459 ringtest_0.x3.nselect2 VDPWR.t1212 VSS.t792 VSS.t791 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X460 a_23949_6654# a_24045_6654# VSS.t138 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X461 a_23529_6422# a_23349_6422# VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X462 a_25055_3867# ringtest_0.x4.net7 VSS.t402 VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X463 a_26555_4790# ringtest_0.x4._09_ VDPWR.t264 VDPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X464 a_22795_5334# a_22765_5308# ringtest_0.x4._04_ VDPWR.t991 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X465 VDPWR.t982 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP4.t3 VDPWR.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X466 VSS.t795 VDPWR.t1213 VSS.t794 VSS.t793 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X467 VDPWR.t255 ringtest_0.drv_out.t21 a_23879_6940# VDPWR.t254 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X468 ringtest_0.x4._24_ a_26627_4246# VSS.t98 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X469 a_26640_5156# a_26201_4790# a_26555_4790# VSS.t318 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X470 a_21675_9686# ringtest_0.x4.net2.t8 VDPWR.t937 VDPWR.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X471 VDPWR.t27 a_22052_9116# a_21981_9142# VDPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X472 VDPWR.t899 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR.t898 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X473 VSS.t465 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X474 VDPWR.t639 VSS.t1170 VDPWR.t638 VDPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X475 a_27303_4246# ringtest_0.x4._23_ VDPWR.t389 VDPWR.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X476 a_21948_5156# a_21675_4790# a_21863_4790# VDPWR.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X477 a_13675_24012# ui_in[3].t6 VSS.t1005 VSS.t1004 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X478 VSS.t798 VDPWR.t1214 VSS.t797 VSS.t796 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X479 VSS.t801 VDPWR.t1215 VSS.t800 VSS.t799 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X480 VSS.t804 VDPWR.t1216 VSS.t803 VSS.t802 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X481 a_26766_4790# a_26367_4790# a_26640_5156# VSS.t323 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X482 VSS.t337 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X483 VDPWR.t636 VSS.t1171 VDPWR.t635 VDPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X484 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk.t37 VSS.t483 VSS.t482 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X485 VDPWR.t1097 ui_in[2].t2 muxtest_0.x1.x5.GN VDPWR.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X486 a_26721_4246# ringtest_0.x4._15_ VDPWR.t353 VDPWR.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X487 VSS.t125 a_22295_3867# ringtest_0.x4.counter[2] VSS.t124 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X488 VSS.t485 ringtest_0.x4.clknet_1_1__leaf_clk.t38 a_24361_5340# VSS.t484 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X489 VSS.t502 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X490 VSS.t1096 ringtest_0.x4._05_ a_24883_6800# VSS.t1095 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X491 VDPWR.t376 a_25336_4902# a_25263_5156# VDPWR.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X492 a_20318_32213# ui_in[0].t5 VDPWR.t1092 VDPWR.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X493 VSS.t1011 a_16579_11759# ringtest_0.x3.x2.GN3 VSS.t1010 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X494 ringtest_0.counter7.t2 ringtest_0.x3.x2.GN4 ua[1].t5 VSS.t382 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X495 VDPWR.t634 VSS.t1172 VDPWR.t633 VDPWR.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X496 a_23879_6940# ringtest_0.drv_out.t22 VDPWR.t257 VDPWR.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X497 a_26808_5308# a_26640_5334# VDPWR.t818 VDPWR.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X498 ringtest_0.x4.clknet_1_1__leaf_clk.t10 a_25364_5878# VSS.t1083 VSS.t1082 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X499 a_26095_6788# ringtest_0.x4.net7 a_26007_6788# VSS.t400 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X500 ringtest_0.x4._07_ a_24699_6200# VDPWR.t367 VDPWR.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14575 ps=1.335 w=1 l=0.15
X501 a_21840_5308# a_21672_5334# VSS.t496 VSS.t495 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X502 a_15749_12123# ringtest_0.x3.x1.nSEL1 VSS.t729 VSS.t728 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X503 VSS.t807 VDPWR.t1217 VSS.t806 VSS.t805 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X504 VSS.t573 ringtest_0.x4._15_ a_26201_6788# VSS.t572 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X505 VDPWR.t808 ringtest_0.x4.net11 a_27489_3702# VDPWR.t807 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X506 VSS.t370 a_26808_4902# a_26766_4790# VSS.t369 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X507 VDPWR.t632 VSS.t1173 VDPWR.t631 VDPWR.t630 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X508 a_25263_5156# a_24729_4790# a_25168_5156# VDPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X509 VSS.t353 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2.t0 VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X510 ua[2].t9 muxtest_0.x2.x2.GP4.t5 muxtest_0.R7R8.t6 VDPWR.t763 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X511 VSS.t628 a_23879_6940# ringtest_0.x4.clknet_0_clk.t8 VSS.t627 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X512 VSS.t809 VDPWR.t1218 VSS.t808 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X513 a_21375_3867# ringtest_0.x4.net3.t5 VSS.t647 VSS.t646 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X514 VDPWR.t292 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X515 VSS.t812 VDPWR.t1219 VSS.t811 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X516 ringtest_0.x4._15_ a_23381_4584# VDPWR.t847 VDPWR.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X517 VDPWR.t64 a_24135_3867# ringtest_0.x4.counter[4] VDPWR.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X518 VDPWR.t393 ringtest_0.x4.clknet_1_0__leaf_clk.t36 a_21233_5340# VDPWR.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X519 muxtest_0.x1.x1.nSEL1 ui_in[1].t6 VSS.t292 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X520 ringtest_0.ring_out.t3 ringtest_0.x3.x2.GN1 ua[1].t8 VSS.t527 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X521 ringtest_0.x4._10_ a_21785_8054# VDPWR.t95 VDPWR.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X522 ua[1].t3 ringtest_0.x3.x2.GP3 ringtest_0.counter3.t1 VDPWR.t50 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X523 a_22164_4362# ringtest_0.x4._16_.t6 VDPWR.t1147 VDPWR.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X524 a_23467_4584# ringtest_0.x4.net4 a_23381_4584# VSS.t854 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X525 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP2.t6 muxtest_0.R2R3.t1 VDPWR.t68 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X526 VSS.t668 ringtest_0.x4.clknet_0_clk.t38 a_21395_6940# VSS.t667 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X527 VDPWR.t629 VSS.t1174 VDPWR.t628 VDPWR.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X528 VSS.t175 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X529 a_24685_6788# a_24465_6800# VSS.t406 VSS.t405 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X530 VDPWR.t626 VSS.t1175 VDPWR.t625 VDPWR.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X531 VDPWR.t859 ui_in[6].t0 ringtest_0.ring_out.t7 VDPWR.t858 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X532 VSS.t814 VDPWR.t1220 VSS.t813 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X533 VSS.t817 VDPWR.t1221 VSS.t816 VSS.t815 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X534 VSS.t1033 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t6 VSS.t1032 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X535 VDPWR.t1050 ringtest_0.x4._22_ a_26721_4246# VDPWR.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X536 VSS.t645 ringtest_0.x4._20_ a_23963_4790# VSS.t644 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X537 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP1.t5 muxtest_0.R7R8.t3 VDPWR.t1036 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X538 a_22695_8304# ringtest_0.x4._12_ ringtest_0.x4._01_ VDPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X539 ringtest_0.x4._17_ a_25925_6788# VDPWR.t263 VDPWR.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X540 muxtest_0.x2.x2.GP4.t2 muxtest_0.x2.x2.GN4 VDPWR.t980 VDPWR.t979 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X541 ringtest_0.x4.clknet_0_clk.t7 a_23879_6940# VSS.t626 VSS.t625 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X542 a_26555_4790# ringtest_0.x4._09_ VSS.t481 VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X543 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VSS.t778 VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X544 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR.t897 VDPWR.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X545 ringtest_0.x4.clknet_1_1__leaf_clk.t22 a_25364_5878# VDPWR.t1113 VDPWR.t1112 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X546 VDPWR.t935 ringtest_0.x4.net2.t9 a_21785_8054# VDPWR.t934 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X547 a_27169_6641# ringtest_0.x4._25_ VDPWR.t901 VDPWR.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X548 a_24317_4942# ringtest_0.x4.net8 VDPWR.t798 VDPWR.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X549 ringtest_0.x4._16_.t0 a_23381_4818# VSS.t1094 VSS.t828 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X550 ringtest_0.drv_out.t15 a_19289_13081.t10 VDPWR.t824 VDPWR.t823 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X551 muxtest_0.R5R6.t4 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A VSS.t835 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X552 muxtest_0.R4R5.t0 muxtest_0.R3R4.t4 VSS.t371 sky130_fd_pr__res_high_po_1p41 l=1.75
X553 VSS.t1099 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 VSS.t1098 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X554 a_21845_8816# ringtest_0.x4.clknet_1_0__leaf_clk.t37 VSS.t761 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X555 a_27815_3867# ringtest_0.x4.net10 VSS.t773 VSS.t772 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X556 a_21561_9116# a_21845_9116# a_21780_9142# VSS.t308 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X557 a_21840_5308# a_21672_5334# VDPWR.t272 VDPWR.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X558 muxtest_0.x1.x5.GN ui_in[2].t3 VDPWR.t1099 VDPWR.t1098 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X559 VSS.t933 a_12297_23648# muxtest_0.x2.x2.GN2 VSS.t932 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X560 VDPWR.t988 ringtest_0.x3.x1.nSEL0 a_15575_12017# VDPWR.t987 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X561 ringtest_0.x4.clknet_1_0__leaf_clk.t5 a_21395_6940# VSS.t1031 VSS.t1030 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X562 VSS.t404 a_25149_4220# ringtest_0.x4._22_ VSS.t403 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X563 VDPWR.t211 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP4.t3 VDPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X564 VDPWR.t623 VSS.t1176 VDPWR.t622 VDPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X565 a_21561_8830# a_21845_8816# a_21780_8964# VSS.t308 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X566 VDPWR.t621 VSS.t1177 VDPWR.t620 VDPWR.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X567 VSS.t819 VDPWR.t1222 VSS.t818 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X568 VDPWR.t618 VSS.t1178 VDPWR.t617 VDPWR.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X569 VSS.t159 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X570 VSS.t508 a_18662_32213# muxtest_0.x1.x3.GN1 VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X571 VDPWR.t1165 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1.t3 VDPWR.t1164 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X572 VDPWR.t615 VSS.t1179 VDPWR.t614 VDPWR.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X573 VSS.t822 VDPWR.t1223 VSS.t821 VSS.t820 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X574 VDPWR.t31 a_13025_23980# a_12849_23648# VDPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X575 a_21507_9686# ringtest_0.x4.net1 a_21425_9686# VDPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X576 VDPWR.t612 VSS.t1180 VDPWR.t611 VDPWR.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X577 VSS.t825 VDPWR.t1224 VSS.t824 VSS.t823 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X578 a_24045_6654# a_24329_6640# a_24264_6788# VSS.t963 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X579 VSS.t937 ringtest_0.x4._14_ a_22390_4566# VSS.t936 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X580 a_25719_4790# a_24729_4790# a_25593_5156# VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X581 a_17405_12123# ui_in[3].t7 VSS.t1007 VSS.t1006 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X582 VDPWR.t609 VSS.t1181 VDPWR.t608 VDPWR.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X583 ringtest_0.counter3.t4 ringtest_0.x3.x2.GN3 ua[1].t15 VSS.t1097 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X584 a_27169_6641# ringtest_0.x4._25_ VSS.t878 VSS.t877 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X585 ringtest_0.drv_out.t5 a_19289_13081.t11 VSS.t561 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X586 ringtest_0.x3.x1.nSEL0 ui_in[3].t8 VDPWR.t1032 VDPWR.t1031 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X587 VSS.t827 VDPWR.t1225 VSS.t826 VSS.t815 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X588 VDPWR.t413 a_23879_6940# ringtest_0.x4.clknet_0_clk.t25 VDPWR.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X589 VSS.t235 VDPWR.t1226 VSS.t234 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X590 ringtest_0.x4._00_ ringtest_0.x4.net1 a_21675_10006# VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X591 VDPWR.t1149 ringtest_0.x4._16_.t7 a_24763_6143# VDPWR.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.129 ps=1.18 w=0.42 l=0.15
X592 VSS.t238 VDPWR.t1227 VSS.t237 VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X593 a_21803_8598# a_21465_8830# VDPWR.t997 VDPWR.t996 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X594 a_22457_5156# a_21675_4790# a_22373_5156# VDPWR.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X595 a_18836_32319# muxtest_0.x1.x1.nSEL1 VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X596 VSS.t241 VDPWR.t1228 VSS.t240 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X597 VDPWR.t607 VSS.t1182 VDPWR.t606 VDPWR.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X598 a_25364_5878# ringtest_0.x4.clknet_0_clk.t39 VDPWR.t774 VDPWR.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X599 VDPWR.t340 a_19289_13081.t12 ringtest_0.drv_out.t14 VDPWR.t339 sky130_fd_pr__pfet_01v8 ad=2.79 pd=18.62 as=1.485 ps=9.33 w=9 l=0.15
X600 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP3 muxtest_0.R5R6.t1 VDPWR.t122 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X601 muxtest_0.R4R5.t5 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A VSS.t986 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X602 ringtest_0.x4.net6.t0 a_22817_6146# VSS.t750 VSS.t749 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X603 a_24986_5878# ringtest_0.x4._22_ a_24763_6143# VSS.t1015 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.1092 ps=1.36 w=0.42 l=0.15
X604 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP4.t5 muxtest_0.R4R5.t1 VDPWR.t957 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X605 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk.t38 VDPWR.t826 VDPWR.t825 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X606 a_24287_6422# a_23949_6654# VDPWR.t380 VDPWR.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X607 VDPWR.t201 a_26808_4902# a_26735_5156# VDPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X608 a_26640_5334# a_26201_5340# a_26555_5334# VSS.t655 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X609 VSS.t864 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2.t1 VSS.t863 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X610 VDPWR.t259 ringtest_0.drv_out.t23 a_23879_6940# VDPWR.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X611 a_23837_5878# ringtest_0.x4._17_ VSS.t1108 VSS.t1107 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X612 ringtest_0.ring_out.t8 ui_in[6].t1 VDPWR.t861 VDPWR.t860 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X613 VDPWR.t137 a_21845_8816# a_21852_8720# VDPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X614 ringtest_0.x4.net4 a_22265_5308# VSS.t387 VSS.t386 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X615 VSS.t1009 ui_in[3].t9 a_13025_23980# VSS.t1008 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X616 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP4.t6 ua[0].t6 VDPWR.t958 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X617 VDPWR.t604 VSS.t1183 VDPWR.t603 VDPWR.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X618 VDPWR.t601 VSS.t1184 VDPWR.t600 VDPWR.t599 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X619 a_13501_23906# ui_in[3].t10 VDPWR.t1034 VDPWR.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X620 VSS.t244 VDPWR.t1229 VSS.t243 VSS.t242 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X621 a_26735_5156# a_26201_4790# a_26640_5156# VDPWR.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X622 VSS.t247 VDPWR.t1230 VSS.t246 VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X623 VDPWR.t598 VSS.t1185 VDPWR.t597 VDPWR.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X624 VSS.t377 a_17231_12017# ringtest_0.x3.x2.GN4 VSS.t376 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X625 ringtest_0.x4.clknet_0_clk.t6 a_23879_6940# VSS.t624 VSS.t623 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X626 VSS.t250 VDPWR.t1231 VSS.t249 VSS.t248 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X627 a_26766_5712# a_26367_5340# a_26640_5334# VSS.t974 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X628 VDPWR.t595 VSS.t1186 VDPWR.t594 VDPWR.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X629 a_21981_8976# a_21845_8816# a_21561_8830# VDPWR.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X630 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VSS.t500 VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X631 a_26007_6788# ringtest_0.x4.net6.t8 a_25925_6788# VSS.t1001 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X632 VDPWR.t593 VSS.t1187 VDPWR.t592 VDPWR.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X633 VDPWR.t363 ringtest_0.x4._21_ a_24070_5852# VDPWR.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.1176 ps=1.4 w=0.42 l=0.15
X634 VSS.t537 a_25761_5058# a_25719_4790# VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X635 VDPWR.t19 a_12473_23980# a_12297_23648# VDPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X636 a_15575_12017# ringtest_0.x3.x1.nSEL1 VDPWR.t793 VDPWR.t792 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X637 ringtest_0.x4.clknet_0_clk.t24 a_23879_6940# VDPWR.t411 VDPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X638 VSS.t253 VDPWR.t1232 VSS.t252 VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X639 a_24465_6800# a_24329_6640# a_24045_6654# VDPWR.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X640 VSS.t487 ringtest_0.x4.clknet_1_1__leaf_clk.t39 a_26201_5340# VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X641 VDPWR.t1111 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t21 VDPWR.t1110 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X642 VDPWR.t591 VSS.t1188 VDPWR.t590 VDPWR.t589 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X643 ringtest_0.x4._06_ a_24004_6128# VSS.t983 VSS.t982 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X644 VDPWR.t588 VSS.t1189 VDPWR.t587 VDPWR.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X645 ringtest_0.x4.net6.t1 a_22817_6146# VDPWR.t811 VDPWR.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X646 VSS.t834 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 VSS.t833 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X647 VSS.t255 VDPWR.t1233 VSS.t254 VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X648 ringtest_0.x4.clknet_1_0__leaf_clk.t4 a_21395_6940# VSS.t1029 VSS.t1028 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X649 ringtest_0.x4.clknet_1_1__leaf_clk.t9 a_25364_5878# VSS.t1081 VSS.t1080 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X650 muxtest_0.x2.x2.GP1.t2 muxtest_0.x2.x2.GN1 VDPWR.t1163 VDPWR.t1162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X651 VSS.t622 a_23879_6940# ringtest_0.x4.clknet_0_clk.t5 VSS.t621 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X652 VDPWR.t905 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR.t904 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X653 muxtest_0.R1R2.t5 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A VSS.t832 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X654 VSS.t258 VDPWR.t1234 VSS.t257 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X655 a_27065_5334# a_26201_5340# a_26808_5308# VDPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X656 VSS.t107 a_12849_23648# muxtest_0.x2.x2.GN3 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X657 VDPWR.t374 a_25977_4220# ringtest_0.x4._23_ VDPWR.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X658 VDPWR.t765 muxtest_0.x1.x1.nSEL0 a_18662_32213# VDPWR.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X659 a_23349_6422# ringtest_0.x4._17_ VSS.t1106 VSS.t1105 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X660 ringtest_0.x4.clknet_1_1__leaf_clk.t20 a_25364_5878# VDPWR.t1109 VDPWR.t1108 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X661 a_21675_4790# a_21509_4790# VDPWR.t335 VDPWR.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X662 a_21672_5334# a_21233_5340# a_21587_5334# VSS.t950 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X663 a_22765_4478# ringtest_0.x4.net4 a_22939_4584# VSS.t853 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X664 VSS.t296 ui_in[4].t5 a_12473_23980# VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X665 VSS.t1027 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t3 VSS.t1026 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X666 VDPWR.t585 VSS.t1190 VDPWR.t584 VDPWR.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X667 a_25441_4612# ringtest_0.x4.net8 a_25345_4612# VSS.t734 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X668 a_27149_5156# a_26367_4790# a_27065_5156# VDPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VSS.t336 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X670 VSS.t971 a_21465_8830# ringtest_0.x4.net3.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X671 muxtest_0.R2R3.t3 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A VSS.t344 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X672 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR.t887 VDPWR.t886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X673 a_22224_6244# a_21785_5878# a_22139_5878# VSS.t327 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X674 a_25055_3867# ringtest_0.x4.net7 VDPWR.t224 VDPWR.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X675 VSS.t601 a_25393_5308# a_25351_5712# VSS.t600 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X676 a_21798_5712# a_21399_5340# a_21672_5334# VSS.t516 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X677 muxtest_0.R7R8.t0 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A VSS.t149 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X678 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP2.t7 muxtest_0.R2R3.t0 VDPWR.t69 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X679 VDPWR.t582 VSS.t1191 VDPWR.t581 VDPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X680 VDPWR.t93 a_24763_6143# a_24699_6200# VDPWR.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.0672 ps=0.74 w=0.42 l=0.15
X681 VDPWR.t191 a_24536_6699# a_24465_6800# VDPWR.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X682 VDPWR.t830 a_27233_5308# a_27149_5334# VDPWR.t829 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X683 VSS.t261 VDPWR.t1235 VSS.t260 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X684 VSS.t343 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2.t0 VSS.t342 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X685 VDPWR.t342 a_19289_13081.t13 ringtest_0.drv_out.t13 VDPWR.t341 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X686 a_22350_5878# a_21951_5878# a_22224_6244# VSS.t739 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X687 VSS.t399 ringtest_0.x4.net7 a_23770_5308# VSS.t398 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X688 VSS.t763 ringtest_0.x4.clknet_1_0__leaf_clk.t39 a_21233_5340# VSS.t762 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X689 ringtest_0.x4.clknet_1_0__leaf_clk.t2 a_21395_6940# VSS.t1025 VSS.t1024 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X690 VDPWR.t117 ui_in[4].t6 muxtest_0.x2.x1.nSEL1 VDPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X691 a_19289_13081.t0 ringtest_0.ring_out.t12 VSS.t583 VSS.t582 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X692 VDPWR.t579 VSS.t1192 VDPWR.t578 VDPWR.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X693 VDPWR.t776 ringtest_0.x4.clknet_0_clk.t40 a_25364_5878# VDPWR.t775 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X694 ringtest_0.x4.counter[9] a_27489_3702# VSS.t285 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X695 ringtest_0.x4.clknet_1_1__leaf_clk.t8 a_25364_5878# VSS.t1079 VSS.t1078 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X696 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR.t311 VDPWR.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X697 a_17231_12017# ui_in[3].t11 VDPWR.t909 VDPWR.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X698 VDPWR.t576 VSS.t1193 VDPWR.t575 VDPWR.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X699 VSS.t263 VDPWR.t1236 VSS.t262 VSS.t205 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X700 VDPWR.t39 a_22295_3867# ringtest_0.x4.counter[2] VDPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X701 VDPWR.t573 VSS.t1194 VDPWR.t572 VDPWR.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X702 a_22765_5308# ringtest_0.x4.net6.t9 VSS.t1003 VSS.t1002 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X703 ua[3].t1 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A VSS.t298 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X704 VSS.t620 a_23879_6940# ringtest_0.x4.clknet_0_clk.t4 VSS.t619 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X705 ua[2].t7 muxtest_0.x2.x2.GP2.t4 ua[0].t3 VDPWR.t761 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X706 a_22097_5334# a_21233_5340# a_21840_5308# VDPWR.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X707 muxtest_0.R3R4.t8 muxtest_0.x2.x2.GN3 ua[2].t10 VSS.t942 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X708 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR.t903 VDPWR.t902 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X709 VSS.t266 VDPWR.t1237 VSS.t265 VSS.t264 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X710 VDPWR.t409 a_23879_6940# ringtest_0.x4.clknet_0_clk.t23 VDPWR.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X711 ringtest_0.x4._19_ a_23529_6422# VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X712 a_23381_4584# ringtest_0.x4.net4 VDPWR.t871 VDPWR.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X713 VSS.t652 a_25593_5156# a_25761_5058# VSS.t651 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X714 a_22139_5878# ringtest_0.x4._04_ VDPWR.t978 VDPWR.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X715 muxtest_0.x2.x1.nSEL0 ui_in[3].t12 VSS.t884 VSS.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X716 VSS.t269 VDPWR.t1238 VSS.t268 VSS.t267 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X717 a_21375_3867# ringtest_0.x4.net3.t6 VDPWR.t758 VDPWR.t757 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X718 a_24317_4942# ringtest_0.x4.net6.t10 VDPWR.t1030 VDPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X719 VDPWR.t197 a_16203_12091# a_16027_11759# VDPWR.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X720 VDPWR.t103 ringtest_0.x4._11_.t12 a_22695_8304# VDPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X721 ringtest_0.x4.clknet_1_0__leaf_clk.t26 a_21395_6940# VDPWR.t1076 VDPWR.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X722 VSS.t272 VDPWR.t1239 VSS.t271 VSS.t270 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X723 VSS.t524 a_26895_3867# ringtest_0.counter7.t4 VSS.t523 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X724 ua[1].t2 ringtest_0.x3.x2.GP3 ringtest_0.counter3.t0 VDPWR.t49 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X725 VSS.t275 VDPWR.t1240 VSS.t274 VSS.t273 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X726 VSS.t1023 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t1 VSS.t1022 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X727 ua[2].t4 muxtest_0.x2.x2.GP3 muxtest_0.R3R4.t2 VDPWR.t281 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X728 VDPWR.t570 VSS.t1195 VDPWR.t569 VDPWR.t568 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X729 VDPWR.t567 VSS.t1196 VDPWR.t566 VDPWR.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X730 VSS.t278 VDPWR.t1241 VSS.t277 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X731 a_26367_4790# a_26201_4790# VDPWR.t148 VDPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X732 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR.t247 VDPWR.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X733 a_24545_5878# ringtest_0.x4.net9 VSS.t520 VSS.t519 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X734 muxtest_0.R6R7.t2 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A VSS.t341 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X735 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP3 muxtest_0.R5R6.t0 VDPWR.t121 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X736 a_24968_5308# a_24800_5334# VSS.t310 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X737 VDPWR.t213 a_22265_5308# a_22181_5334# VDPWR.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X738 a_13501_23906# ui_in[4].t7 a_13675_24012# VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X739 VSS.t886 ui_in[3].t13 ringtest_0.x3.x1.nSEL0 VSS.t885 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X740 VDPWR.t378 a_23949_6654# ringtest_0.x4.net7 VDPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X741 VSS.t280 VDPWR.t1242 VSS.t279 VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X742 VDPWR.t564 VSS.t1197 VDPWR.t563 VDPWR.t562 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X743 VSS.t571 ringtest_0.x4._15_ a_23467_4818# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X744 VDPWR.t1074 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t25 VDPWR.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X745 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VSS.t157 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X746 VSS.t996 ui_in[4].t8 a_16203_12091# VSS.t995 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X747 VDPWR.t561 VSS.t1198 VDPWR.t560 VDPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X748 VSS.t283 VDPWR.t1243 VSS.t282 VSS.t281 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X749 VDPWR.t107 ui_in[1].t7 a_20318_32213# VDPWR.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X750 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP4.t7 ua[0].t5 VDPWR.t959 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X751 a_24004_6128# a_24070_5852# a_23837_5878# VSS.t533 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X752 VDPWR.t769 a_25593_5156# a_25761_5058# VDPWR.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X753 a_22373_5156# a_21675_4790# a_22116_4902# VSS.t559 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X754 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR.t280 VDPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X755 a_21465_9294# a_21561_9116# VSS.t882 VSS.t881 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X756 VDPWR.t1107 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t19 VDPWR.t1106 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X757 ua[3].t0 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A VSS.t298 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X758 a_23932_6128# ringtest_0.x4.net8 VDPWR.t796 VDPWR.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X759 a_23399_3867# ringtest_0.x4.net5 VSS.t300 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X760 a_27815_3867# ringtest_0.x4.net10 VDPWR.t836 VDPWR.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X761 ringtest_0.x4.clknet_1_1__leaf_clk.t7 a_25364_5878# VSS.t1077 VSS.t1076 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X762 VSS.t7 a_13501_23906# muxtest_0.x2.x2.GN4 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X763 VDPWR.t66 a_22052_8875# a_21981_8976# VDPWR.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X764 VDPWR.t558 VSS.t1199 VDPWR.t557 VDPWR.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X765 ringtest_0.x3.x2.GP4.t2 ringtest_0.x3.x2.GN4 VDPWR.t209 VDPWR.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X766 VDPWR.t913 ringtest_0.x4._11_.t13 a_26721_4246# VDPWR.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X767 a_23899_5654# ringtest_0.x4._15_ VSS.t570 VSS.t569 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X768 ringtest_0.x3.x2.GP2.t0 ringtest_0.x3.x2.GN2 VSS.t862 VSS.t861 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X769 VDPWR.t189 a_19114_31955# muxtest_0.x1.x3.GN2 VDPWR.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X770 VDPWR.t243 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.ring_out.t2 VDPWR.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X771 VDPWR.t1022 ui_in[4].t9 ringtest_0.x3.x1.nSEL1 VDPWR.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X772 VDPWR.t555 VSS.t1200 VDPWR.t554 VDPWR.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X773 a_24800_5334# a_24361_5340# a_24715_5334# VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X774 VSS.t409 VDPWR.t1244 VSS.t408 VSS.t407 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X775 VSS.t1021 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t0 VSS.t1020 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X776 a_23381_4818# ringtest_0.x4._11_.t14 VDPWR.t915 VDPWR.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X777 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR.t91 VDPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X778 a_21561_9116# a_21852_9416# a_21803_9508# VDPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X779 VSS.t777 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VSS.t497 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X780 VSS.t1075 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t6 VSS.t1074 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X781 a_24968_5308# a_24800_5334# VDPWR.t139 VDPWR.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X782 a_24926_5712# a_24527_5340# a_24800_5334# VSS.t754 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X783 VDPWR.t552 VSS.t1201 VDPWR.t551 VDPWR.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X784 VSS.t565 a_22245_8054# ringtest_0.x4._11_.t0 VSS.t564 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X785 a_21132_8918# ringtest_0.x4.net1 VSS.t131 VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X786 ringtest_0.x4._09_ a_27273_4220# VSS.t333 VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X787 a_24551_4790# ringtest_0.x4.net7 a_24479_4790# VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X788 VSS.t412 VDPWR.t1245 VSS.t411 VSS.t410 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X789 muxtest_0.x2.x1.nSEL1 ui_in[4].t10 VSS.t998 VSS.t997 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X790 ua[0].t7 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A VSS.t985 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X791 VDPWR.t961 a_16755_12091# a_16579_11759# VDPWR.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X792 a_27273_4220# ringtest_0.x4._23_ a_27659_4246# VDPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X793 VDPWR.t791 a_24317_4942# ringtest_0.x4._20_ VDPWR.t790 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X794 VSS.t767 a_27233_5308# a_27191_5712# VSS.t766 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X795 ua[2].t6 muxtest_0.x2.x2.GP2.t5 ua[0].t2 VDPWR.t760 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X796 VSS.t415 VDPWR.t1246 VSS.t414 VSS.t413 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X797 ringtest_0.x4.clknet_0_clk.t22 a_23879_6940# VDPWR.t407 VDPWR.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X798 a_22733_6244# a_21951_5878# a_22649_6244# VDPWR.t803 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X799 VDPWR.t549 VSS.t1202 VDPWR.t548 VDPWR.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X800 VDPWR.t547 VSS.t1203 VDPWR.t546 VDPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X801 a_27273_4220# ringtest_0.x4.net11 VSS.t742 VSS.t741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X802 VDPWR.t1140 a_25225_5334# a_25393_5308# VDPWR.t1139 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X803 a_25225_5334# a_24527_5340# a_24968_5308# VSS.t753 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X804 a_22111_10993# ui_in[5].t0 VDPWR.t1088 VDPWR.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X805 VDPWR.t1072 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t24 VDPWR.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X806 VDPWR.t544 VSS.t1204 VDPWR.t543 VDPWR.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X807 VDPWR.t45 ringtest_0.x4.net1 a_21785_8054# VDPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X808 a_27065_5156# a_26367_4790# a_26808_4902# VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X809 VSS.t868 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X810 a_17231_12017# ui_in[4].t11 a_17405_12123# VSS.t999 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X811 ringtest_0.x4._12_ ringtest_0.x4.net3.t7 a_21049_8598# VDPWR.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X812 a_25225_5334# a_24361_5340# a_24968_5308# VDPWR.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X813 VDPWR.t541 VSS.t1205 VDPWR.t540 VDPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X814 VDPWR.t538 VSS.t1206 VDPWR.t537 VDPWR.t536 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X815 VDPWR.t995 a_21465_8830# ringtest_0.x4.net3.t1 VDPWR.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X816 VSS.t418 VDPWR.t1247 VSS.t417 VSS.t416 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X817 muxtest_0.R5R6.t3 muxtest_0.R4R5.t3 VSS.t643 sky130_fd_pr__res_high_po_1p41 l=1.75
X818 ringtest_0.drv_out.t12 a_19289_13081.t14 VDPWR.t344 VDPWR.t343 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=2.79 ps=18.62 w=9 l=0.15
X819 VDPWR.t999 a_22765_4478# ringtest_0.x4._14_ VDPWR.t998 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X820 VSS.t389 a_16027_11759# ringtest_0.x3.x2.GN2 VSS.t388 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X821 VSS.t888 ui_in[3].t14 a_16755_12091# VSS.t887 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X822 VSS.t421 VDPWR.t1248 VSS.t420 VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X823 VSS.t960 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP4.t1 VSS.t959 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X824 VDPWR.t869 ringtest_0.x4.net4 a_22765_4478# VDPWR.t868 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X825 a_22074_4790# a_21675_4790# a_21948_5156# VSS.t558 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X826 a_21780_9142# a_21465_9294# VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X827 a_24763_6143# ringtest_0.x4._22_ VDPWR.t1048 VDPWR.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.20925 ps=1.345 w=0.42 l=0.15
X828 VSS.t424 VDPWR.t1249 VSS.t423 VSS.t422 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X829 ringtest_0.x4.clknet_1_0__leaf_clk.t23 a_21395_6940# VDPWR.t1070 VDPWR.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X830 ringtest_0.ring_out.t1 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR.t241 VDPWR.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X831 VSS.t876 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VSS.t873 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X832 a_23809_4790# ringtest_0.x4._15_ VDPWR.t351 VDPWR.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X833 VDPWR.t535 VSS.t1207 VDPWR.t534 VDPWR.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X834 VSS.t427 VDPWR.t1250 VSS.t426 VSS.t425 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X835 VSS.t458 muxtest_0.R7R8.t2 VSS.t457 sky130_fd_pr__res_high_po_1p41 l=1.75
X836 VSS.t429 VDPWR.t1251 VSS.t428 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X837 VDPWR.t533 VSS.t1208 VDPWR.t532 VDPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X838 a_22052_9116# a_21845_9116# a_22228_9508# VDPWR.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X839 a_22939_4584# ringtest_0.x4._11_.t15 VSS.t890 VSS.t889 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X840 VSS.t849 a_22116_4902# a_22074_4790# VSS.t848 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X841 ringtest_0.x4.clknet_1_1__leaf_clk.t18 a_25364_5878# VDPWR.t1105 VDPWR.t1104 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X842 VDPWR.t1024 ui_in[4].t12 a_13501_23906# VDPWR.t1023 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X843 a_22228_9508# a_21981_9142# VDPWR.t169 VDPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X844 VSS.t1061 ui_in[2].t4 muxtest_0.x1.x5.GN VSS.t1060 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X845 VDPWR.t382 a_25393_5308# a_25309_5334# VDPWR.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X846 a_24895_4790# a_24729_4790# VSS.t314 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X847 VSS.t385 a_22265_5308# a_22223_5712# VSS.t384 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X848 VSS.t1073 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t5 VSS.t1072 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X849 VSS.t432 VDPWR.t1252 VSS.t431 VSS.t430 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X850 VDPWR.t985 a_24329_6640# a_24336_6544# VDPWR.t984 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X851 VSS.t434 VDPWR.t1253 VSS.t433 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X852 muxtest_0.R7R8.t7 muxtest_0.x2.x2.GN4 ua[2].t12 VSS.t958 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X853 a_26555_5334# ringtest_0.x4._08_ VDPWR.t12 VDPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X854 a_19290_32287# ui_in[1].t8 VDPWR.t109 VDPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X855 muxtest_0.R6R7.t4 muxtest_0.R5R6.t2 VSS.t371 sky130_fd_pr__res_high_po_1p41 l=1.75
X856 VSS.t498 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VSS.t497 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X857 VDPWR.t530 VSS.t1209 VDPWR.t529 VDPWR.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X858 a_26627_4246# ringtest_0.x4.net10 VSS.t771 VSS.t770 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X859 VSS.t436 VDPWR.t1254 VSS.t435 VSS.t242 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X860 a_22775_5878# a_21785_5878# a_22649_6244# VSS.t326 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X861 VSS.t439 VDPWR.t1255 VSS.t438 VSS.t437 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X862 a_22795_5334# ringtest_0.x4._16_.t8 VDPWR.t1151 VDPWR.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X863 ringtest_0.x4._13_ ringtest_0.x4._11_.t16 VSS.t892 VSS.t891 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X864 VSS.t512 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X865 VSS.t591 a_23949_6654# ringtest_0.x4.net7 VSS.t590 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X866 VDPWR.t778 ringtest_0.x4.clknet_0_clk.t41 a_25364_5878# VDPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X867 a_26367_5340# a_26201_5340# VDPWR.t770 VDPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X868 VDPWR.t780 ringtest_0.x4.clknet_0_clk.t42 a_21395_6940# VDPWR.t779 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X869 ringtest_0.drv_out.t4 a_19289_13081.t15 VSS.t563 VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X870 ua[1].t12 ringtest_0.x3.x2.GP1.t4 ringtest_0.ring_out.t6 VDPWR.t1012 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X871 VSS.t365 ringtest_0.x4._18_ a_23619_6788# VSS.t364 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X872 VSS.t441 VDPWR.t1256 VSS.t440 VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X873 a_12849_23648# ui_in[4].t13 VDPWR.t925 VDPWR.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X874 ringtest_0.x4.clknet_1_1__leaf_clk.t4 a_25364_5878# VSS.t1071 VSS.t1070 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X875 VDPWR.t527 VSS.t1210 VDPWR.t526 VDPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X876 a_26640_5156# a_26367_4790# a_26555_4790# VDPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X877 muxtest_0.R3R4.t0 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A VSS.t148 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X878 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP1.t6 muxtest_0.R3R4.t6 VDPWR.t1037 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X879 VSS.t444 VDPWR.t1257 VSS.t443 VSS.t442 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X880 VSS.t447 VDPWR.t1258 VSS.t446 VSS.t445 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X881 VDPWR.t524 VSS.t1211 VDPWR.t523 VDPWR.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X882 a_22399_9142# a_21852_9416# a_22052_9116# VDPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X883 VDPWR.t43 ringtest_0.x4.net1 a_21675_9686# VDPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X884 ringtest_0.x4.counter[9] a_27489_3702# VDPWR.t97 VDPWR.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X885 VSS.t110 ringtest_0.x4.clknet_1_0__leaf_clk.t40 a_21509_4790# VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X886 a_22392_5990# a_22224_6244# VSS.t914 VSS.t913 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X887 muxtest_0.x1.x1.nSEL0 ui_in[0].t6 VDPWR.t234 VDPWR.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X888 a_17377_14114# ui_in[6].t2 ringtest_0.ring_out.t9 VSS.t845 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X889 ua[1].t13 ringtest_0.x3.x2.GP2.t4 ringtest_0.drv_out.t19 VDPWR.t1093 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X890 VDPWR.t806 ringtest_0.x4.net11 a_27303_4246# VDPWR.t805 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X891 muxtest_0.x2.x2.GP4.t0 muxtest_0.x2.x2.GN4 VSS.t957 VSS.t956 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X892 muxtest_0.R2R3.t4 muxtest_0.R1R2.t3 VSS.t551 sky130_fd_pr__res_high_po_1p41 l=1.75
X893 VSS.t173 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X894 ringtest_0.x4.clknet_1_0__leaf_clk.t22 a_21395_6940# VDPWR.t1068 VDPWR.t1067 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X895 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VSS.t875 VSS.t871 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X896 ringtest_0.x4.clknet_0_clk.t3 a_23879_6940# VSS.t618 VSS.t617 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X897 VDPWR.t222 ringtest_0.x4.net7 a_24317_4942# VDPWR.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X898 VSS.t748 a_22817_6146# a_22775_5878# VSS.t747 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X899 VSS.t450 VDPWR.t1259 VSS.t449 VSS.t448 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X900 VDPWR.t301 a_26895_3867# ringtest_0.counter7.t5 VDPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X901 VSS.t874 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VSS.t873 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X902 VDPWR.t521 VSS.t1212 VDPWR.t520 VDPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X903 VDPWR.t1005 ringtest_0.x4._10_ a_22245_8054# VDPWR.t1004 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X904 VSS.t1104 a_25225_5334# a_25393_5308# VSS.t1103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X905 a_21587_5334# ringtest_0.x4._02_ VDPWR.t10 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X906 muxtest_0.x1.x5.GN ui_in[2].t5 VSS.t661 VSS.t660 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X907 a_25336_4902# a_25168_5156# VSS.t506 VSS.t505 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X908 VSS.t1069 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t3 VSS.t1068 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X909 VSS.t381 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP4.t1 VSS.t380 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X910 VDPWR.t1103 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t17 VDPWR.t1102 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X911 VSS.t453 VDPWR.t1260 VSS.t452 VSS.t451 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X912 ringtest_0.x4.clknet_0_clk.t21 a_23879_6940# VDPWR.t405 VDPWR.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X913 VSS.t1125 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1.t1 VSS.t1124 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X914 ringtest_0.drv_out.t2 ringtest_0.x3.x2.GN2 ua[1].t11 VSS.t860 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X915 VSS.t129 ringtest_0.x4.net1 a_21939_8054# VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X916 a_21399_5340# a_21233_5340# VDPWR.t975 VDPWR.t974 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X917 muxtest_0.x1.x5.A ui_in[2].t6 ua[3].t6 VDPWR.t772 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X918 a_19289_13081.t1 ringtest_0.ring_out.t13 VDPWR.t373 VDPWR.t372 sky130_fd_pr__pfet_01v8 ad=2.61 pd=18.58 as=2.61 ps=18.58 w=9 l=0.15
X919 VDPWR.t518 VSS.t1213 VDPWR.t517 VDPWR.t516 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X920 a_12297_23648# ui_in[3].t15 VDPWR.t911 VDPWR.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X921 a_25345_4612# ringtest_0.x4.net9 VSS.t518 VSS.t517 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X922 VSS.t456 VDPWR.t1261 VSS.t455 VSS.t454 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X923 VSS.t183 VDPWR.t1262 VSS.t182 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X924 VDPWR.t1066 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t21 VDPWR.t1065 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X925 VSS.t186 VDPWR.t1263 VSS.t185 VSS.t184 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X926 ringtest_0.x3.x1.nSEL0 ui_in[3].t16 VSS.t840 VSS.t839 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X927 a_25547_4612# ringtest_0.x4.net7 a_25441_4612# VSS.t396 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X928 VDPWR.t865 a_22116_4902# a_22043_5156# VDPWR.t864 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X929 VDPWR.t927 ui_in[4].t14 a_17231_12017# VDPWR.t926 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X930 VDPWR.t386 ringtest_0.x4._23_ a_26569_6422# VDPWR.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X931 VDPWR.t321 a_27065_5334# a_27233_5308# VDPWR.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X932 a_27065_5334# a_26367_5340# a_26808_5308# VSS.t973 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X933 ringtest_0.x4._02_ ringtest_0.x4._14_ a_21055_5334# VDPWR.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X934 VDPWR.t515 VSS.t1214 VDPWR.t514 VDPWR.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X935 a_26173_4612# ringtest_0.x4._22_ VSS.t1014 VSS.t1013 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X936 VSS.t294 a_19666_31955# muxtest_0.x1.x3.GN3 VSS.t293 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X937 ringtest_0.x3.x1.nSEL1 ui_in[4].t15 VDPWR.t929 VDPWR.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X938 a_26375_4612# ringtest_0.x4._11_.t17 a_26269_4612# VSS.t893 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X939 VSS.t189 VDPWR.t1264 VSS.t188 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X940 VSS.t192 VDPWR.t1265 VSS.t191 VSS.t190 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X941 a_22043_5156# a_21509_4790# a_21948_5156# VDPWR.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X942 VSS.t534 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X943 a_26749_6422# a_26569_6422# VDPWR.t867 VDPWR.t866 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X944 a_23770_5308# ringtest_0.x4.net6.t11 a_23993_5654# VSS.t542 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X945 VSS.t103 a_22052_9116# a_21981_9142# VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X946 a_23399_3867# ringtest_0.x4.net5 VDPWR.t125 VDPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X947 VSS.t195 VDPWR.t1266 VSS.t194 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X948 ringtest_0.ring_out.t0 ui_in[6].t3 a_17377_14114# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X949 VDPWR.t261 a_15575_12017# ringtest_0.x3.x2.GN1 VDPWR.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X950 ringtest_0.x4._11_.t2 a_22245_8054# VDPWR.t347 VDPWR.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X951 ringtest_0.x4._02_ ringtest_0.x4._13_ VSS.t858 VSS.t857 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X952 ringtest_0.x4.clknet_1_0__leaf_clk.t20 a_21395_6940# VDPWR.t1064 VDPWR.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X953 muxtest_0.x1.x4.A muxtest_0.x1.x5.GN ua[3].t2 VDPWR.t119 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X954 VSS.t469 a_22021_4220# ringtest_0.x4._03_ VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X955 VSS.t489 ringtest_0.x4.clknet_1_1__leaf_clk.t40 a_26201_4790# VSS.t488 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X956 VDPWR.t512 VSS.t1215 VDPWR.t511 VDPWR.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X957 VDPWR.t509 VSS.t1216 VDPWR.t508 VDPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X958 VDPWR.t506 VSS.t1217 VDPWR.t505 VDPWR.t504 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X959 a_23879_6940# ringtest_0.drv_out.t24 VSS.t475 VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X960 ringtest_0.x4._24_ a_26627_4246# VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X961 a_25593_5156# a_24729_4790# a_25336_4902# VDPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X962 a_22111_10993# ui_in[5].t1 VSS.t1053 VSS.t1052 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X963 a_21395_6940# ringtest_0.x4.clknet_0_clk.t43 VDPWR.t1153 VDPWR.t1152 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X964 VDPWR.t245 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X965 ua[3].t10 muxtest_0.x2.x2.GN1 ua[2].t14 VSS.t1123 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X966 ringtest_0.drv_out.t1 ringtest_0.x3.x2.GN2 ua[1].t10 VSS.t859 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X967 VSS.t896 ringtest_0.x4._01_ a_22399_8976# VSS.t338 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X968 a_25336_4902# a_25168_5156# VDPWR.t284 VDPWR.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X969 VSS.t1067 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t2 VSS.t1066 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X970 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VSS.t872 VSS.t871 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X971 VSS.t198 VDPWR.t1267 VSS.t197 VSS.t196 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X972 VDPWR.t794 a_26808_5308# a_26735_5334# VDPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X973 ringtest_0.x4.clknet_0_clk.t20 a_23879_6940# VDPWR.t403 VDPWR.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X974 VDPWR.t278 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X975 VDPWR.t503 VSS.t1218 VDPWR.t502 VDPWR.t501 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X976 muxtest_0.x2.x2.GP1.t0 muxtest_0.x2.x2.GN1 VSS.t1122 VSS.t1121 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X977 a_21465_9294# a_21561_9116# VDPWR.t907 VDPWR.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X978 VDPWR.t500 VSS.t1219 VDPWR.t499 VDPWR.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X979 ringtest_0.x4._21_ a_23809_4790# VSS.t118 VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X980 VSS.t880 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VSS.t584 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X981 VSS.t201 VDPWR.t1268 VSS.t200 VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X982 VSS.t616 a_23879_6940# ringtest_0.x4.clknet_0_clk.t2 VSS.t615 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X983 muxtest_0.R3R4.t7 muxtest_0.R2R3.t5 VSS.t643 sky130_fd_pr__res_high_po_1p41 l=1.75
X984 VDPWR.t1062 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t19 VDPWR.t1061 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X985 a_23891_4790# ringtest_0.x4._11_.t18 a_23809_4790# VSS.t894 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X986 VDPWR.t497 VSS.t1220 VDPWR.t496 VDPWR.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X987 VDPWR.t37 a_22097_5334# a_22265_5308# VDPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X988 a_22097_5334# a_21399_5340# a_21840_5308# VSS.t515 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X989 ua[3].t7 ui_in[2].t7 muxtest_0.x1.x4.A VSS.t662 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X990 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR.t290 VDPWR.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X991 VSS.t916 a_25055_3867# ringtest_0.x4.counter[5] VSS.t915 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X992 VSS.t204 VDPWR.t1269 VSS.t203 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X993 VDPWR.t317 a_25761_5058# a_25677_5156# VDPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X994 a_26735_5334# a_26201_5340# a_26640_5334# VDPWR.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X995 ua[1].t4 ringtest_0.x3.x2.GP1.t5 ringtest_0.ring_out.t5 VDPWR.t118 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X996 VSS.t614 a_23879_6940# ringtest_0.x4.clknet_0_clk.t1 VSS.t613 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X997 ringtest_0.x4._25_ a_26749_6422# VSS.t492 VSS.t491 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X998 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk.t41 VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X999 VSS.t473 a_19289_13081.t16 ringtest_0.drv_out.t3 VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1000 VDPWR.t494 VSS.t1221 VDPWR.t493 VDPWR.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1001 a_22201_8964# a_21981_8976# VSS.t979 VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1002 VSS.t207 VDPWR.t1270 VSS.t206 VSS.t205 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1003 VSS.t210 VDPWR.t1271 VSS.t209 VSS.t208 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1004 VSS.t213 VDPWR.t1272 VSS.t212 VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1005 a_24135_3867# ringtest_0.x4.net6.t12 VSS.t544 VSS.t543 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1006 a_26808_4902# a_26640_5156# VSS.t368 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1007 a_22499_4790# a_21509_4790# a_22373_5156# VSS.t554 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1008 a_12849_23648# a_13025_23980# a_12977_24040# VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1009 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VSS.t867 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1010 VDPWR.t89 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1011 a_22765_4478# ringtest_0.x4._11_.t19 VDPWR.t917 VDPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1012 VDPWR.t491 VSS.t1222 VDPWR.t490 VDPWR.t489 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1013 a_19842_32287# ui_in[0].t7 VDPWR.t236 VDPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X1014 a_11845_23906# muxtest_0.x2.x1.nSEL0 a_12019_24012# VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1015 VDPWR.t488 VSS.t1223 VDPWR.t487 VDPWR.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1016 VDPWR.t485 VSS.t1224 VDPWR.t484 VDPWR.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1017 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR.t181 VDPWR.t180 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1018 VDPWR.t482 VSS.t1225 VDPWR.t481 VDPWR.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1019 VDPWR.t323 ringtest_0.x4.clknet_1_1__leaf_clk.t41 a_24729_4790# VDPWR.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1020 a_26367_5340# a_26201_5340# VSS.t654 VSS.t653 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1021 VDPWR.t479 VSS.t1226 VDPWR.t478 VDPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1022 a_24715_5334# ringtest_0.x4._06_ VDPWR.t35 VDPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1023 muxtest_0.R4R5.t4 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A VSS.t984 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X1024 a_23619_6788# a_23349_6422# a_23529_6422# VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1025 VSS.t1065 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t1 VSS.t1064 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1026 VSS.t918 ui_in[4].t16 muxtest_0.x2.x1.nSEL1 VSS.t917 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1027 a_21049_8598# ringtest_0.x4.net2.t10 VDPWR.t933 VDPWR.t932 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X1028 VSS.t216 VDPWR.t1273 VSS.t215 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1029 VSS.t931 a_21375_3867# ringtest_0.x4.counter[1] VSS.t930 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1030 VSS.t219 VDPWR.t1274 VSS.t218 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1031 VSS.t541 a_27065_5334# a_27233_5308# VSS.t540 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1032 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR.t839 VDPWR.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1033 VSS.t577 ringtest_0.x4._21_ a_24070_5852# VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1034 a_24527_5340# a_24361_5340# VDPWR.t82 VDPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1035 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP1.t7 muxtest_0.R3R4.t5 VDPWR.t345 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1036 VDPWR.t965 a_12297_23648# muxtest_0.x2.x2.GN2 VDPWR.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1037 a_27149_5334# a_26367_5340# a_27065_5334# VDPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1038 VDPWR.t230 a_25149_4220# ringtest_0.x4._22_ VDPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X1039 a_21767_5334# a_21233_5340# a_21672_5334# VDPWR.t973 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1040 VSS.t307 a_21845_8816# a_21852_8720# VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1041 VSS.t222 VDPWR.t1275 VSS.t221 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1042 ringtest_0.x4.clknet_0_clk.t19 a_23879_6940# VDPWR.t401 VDPWR.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1043 a_25364_5878# ringtest_0.x4.clknet_0_clk.t44 VSS.t1118 VSS.t1117 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1044 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VSS.t879 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1045 VDPWR.t325 ringtest_0.x4.net6.t13 a_25149_4220# VDPWR.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1046 VDPWR.t75 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1047 VSS.t225 VDPWR.t1276 VSS.t224 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1048 VSS.t373 a_22541_5058# a_22499_4790# VSS.t372 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1049 VDPWR.t476 VSS.t1227 VDPWR.t475 VDPWR.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1050 VSS.t595 ringtest_0.drv_out.t25 a_23879_6940# VSS.t594 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1051 a_22486_4246# ringtest_0.x4._14_ a_22021_4220# VDPWR.t966 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1052 VSS.t363 a_23770_5308# ringtest_0.x4._18_ VSS.t362 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1053 VDPWR.t834 ringtest_0.x4.net10 a_25977_4220# VDPWR.t833 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1054 a_12297_23648# a_12473_23980# a_12425_24040# VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1055 VSS.t585 ringtest_0.ring_out.t14 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VSS.t584 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1056 ua[1].t0 ringtest_0.x3.x2.GP4.t5 ringtest_0.counter7.t0 VDPWR.t1095 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1057 VDPWR.t307 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1.t3 VDPWR.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1058 ringtest_0.x4.clknet_1_0__leaf_clk.t18 a_21395_6940# VDPWR.t1060 VDPWR.t1059 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1059 a_24536_6699# a_24336_6544# a_24685_6788# VSS.t765 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1060 VDPWR.t473 VSS.t1228 VDPWR.t472 VDPWR.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1061 VSS.t227 VDPWR.t1277 VSS.t226 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1062 a_12425_24040# ui_in[3].t17 VSS.t842 VSS.t841 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X1063 VDPWR.t955 a_27169_6641# ringtest_0.x4._08_ VDPWR.t954 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1064 VDPWR.t303 a_20318_32213# muxtest_0.x1.x3.GN4 VDPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1065 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR.t883 VDPWR.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1066 VDPWR.t399 a_23879_6940# ringtest_0.x4.clknet_0_clk.t18 VDPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1067 a_24536_6699# a_24329_6640# a_24712_6422# VDPWR.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X1068 VSS.t312 a_27815_3867# ringtest_0.x4.counter[8] VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1069 muxtest_0.R1R2.t4 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A VSS.t831 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X1070 ua[1].t7 ringtest_0.x3.x2.GP2.t5 ringtest_0.drv_out.t0 VDPWR.t239 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1071 a_25421_6641# ringtest_0.x4._19_ VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1072 VDPWR.t470 VSS.t1229 VDPWR.t469 VDPWR.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1073 a_23879_6940# ringtest_0.drv_out.t26 VSS.t597 VSS.t596 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1074 a_21399_5340# a_21233_5340# VSS.t949 VSS.t948 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1075 VSS.t361 a_24536_6699# a_24465_6800# VSS.t360 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1076 a_24883_6800# a_24329_6640# a_24536_6699# VSS.t962 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1077 muxtest_0.x2.x2.GP3 muxtest_0.x2.x2.GN3 VDPWR.t972 VDPWR.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1078 a_21395_6940# ringtest_0.x4.clknet_0_clk.t45 VDPWR.t1155 VDPWR.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1079 a_26201_6788# ringtest_0.x4._11_.t20 a_26095_6788# VSS.t895 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1080 VSS.t329 a_22649_6244# a_22817_6146# VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1081 VSS.t229 VDPWR.t1278 VSS.t228 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1082 ringtest_0.x4._07_ a_24699_6200# VSS.t581 VSS.t580 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.098625 ps=0.98 w=0.65 l=0.15
X1083 VDPWR.t164 a_21845_9116# a_21852_9416# VDPWR.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1084 a_24712_6422# a_24465_6800# VDPWR.t232 VDPWR.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1085 VDPWR.t854 ui_in[3].t18 muxtest_0.x2.x1.nSEL0 VDPWR.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1086 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VSS.t171 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1087 VSS.t1116 ringtest_0.x4._16_.t9 a_22765_5308# VSS.t1115 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1088 VSS.t122 a_22097_5334# a_22265_5308# VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1089 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP3 muxtest_0.R1R2.t0 VDPWR.t120 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1090 a_16579_11759# ui_in[4].t17 VDPWR.t931 VDPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X1091 VDPWR.t467 VSS.t1230 VDPWR.t466 VDPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1092 VSS.t928 a_27169_6641# ringtest_0.x4._08_ VSS.t927 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1093 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR.t274 VDPWR.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1094 muxtest_0.R2R3.t2 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A VSS.t340 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X1095 a_25421_6641# ringtest_0.x4._19_ VSS.t95 VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1096 VDPWR.t41 a_22111_10993# ringtest_0.x4.net1 VDPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1097 ringtest_0.drv_out.t11 a_19289_13081.t17 VDPWR.t253 VDPWR.t252 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X1098 ringtest_0.x3.x2.GP4.t0 ringtest_0.x3.x2.GN4 VSS.t379 VSS.t378 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1099 a_21561_8830# a_21852_8720# a_21803_8598# VDPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1100 VDPWR.t464 VSS.t1231 VDPWR.t463 VDPWR.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1101 a_23993_5654# ringtest_0.x4._11_.t21 a_23899_5654# VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1102 VDPWR.t461 VSS.t1232 VDPWR.t460 VDPWR.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1103 VSS.t935 ui_in[1].t9 a_19290_32287# VSS.t934 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1104 a_17377_14114# ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VSS.t464 VSS.t463 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1105 VSS.t167 ui_in[4].t18 ringtest_0.x3.x1.nSEL1 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1106 a_24883_6800# a_24336_6544# a_24536_6699# VDPWR.t827 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X1107 VDPWR.t238 ui_in[0].t8 muxtest_0.x1.x1.nSEL0 VDPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1108 a_18662_32213# muxtest_0.x1.x1.nSEL1 VDPWR.t62 VDPWR.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1109 VDPWR.t458 VSS.t1233 VDPWR.t457 VDPWR.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1110 VDPWR.t455 VSS.t1234 VDPWR.t454 VDPWR.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1111 VDPWR.t158 a_22649_6244# a_22817_6146# VDPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1112 VDPWR.t452 VSS.t1235 VDPWR.t451 VDPWR.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1113 VSS.t1110 a_27233_5058# a_27191_4790# VSS.t1109 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1114 VDPWR.t29 a_12849_23648# muxtest_0.x2.x2.GN3 VDPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1115 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.ring_out.t15 VSS.t105 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1116 ringtest_0.x4.clknet_1_1__leaf_clk.t0 a_25364_5878# VSS.t1063 VSS.t1062 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1117 a_24699_6200# a_24763_6143# a_24545_5878# VSS.t178 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1118 muxtest_0.x2.x2.GP2.t2 muxtest_0.x2.x2.GN2 VDPWR.t185 VDPWR.t184 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1119 ringtest_0.x3.x2.GP1.t2 ringtest_0.x3.x2.GN1 VDPWR.t305 VDPWR.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1120 ringtest_0.x4.clknet_1_1__leaf_clk.t16 a_25364_5878# VDPWR.t1101 VDPWR.t1100 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1121 VDPWR.t146 muxtest_0.x2.x1.nSEL0 a_11845_23906# VDPWR.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1122 a_21951_5878# a_21785_5878# VSS.t325 VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1123 VSS.t494 a_22373_5156# a_22541_5058# VSS.t493 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1124 VDPWR.t449 VSS.t1236 VDPWR.t448 VDPWR.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1125 a_25975_3867# ringtest_0.x4.net8 VSS.t733 VSS.t732 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1126 a_21981_9142# a_21852_9416# a_21561_9116# VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1127 VSS.t232 VDPWR.t1279 VSS.t231 VSS.t230 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1128 VDPWR.t397 a_23879_6940# ringtest_0.x4.clknet_0_clk.t17 VDPWR.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1129 VSS.t18 VDPWR.t1280 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1130 a_21981_8976# a_21852_8720# a_21561_8830# VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1131 VDPWR.t446 VSS.t1237 VDPWR.t445 VDPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1132 a_22319_6244# a_21785_5878# a_22224_6244# VDPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1133 VDPWR.t71 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1.t2 VDPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1134 VSS.t21 VDPWR.t1281 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1135 VDPWR.t990 a_19290_32287# a_19114_31955# VDPWR.t989 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1136 VSS.t24 VDPWR.t1282 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1137 VDPWR.t443 VSS.t1238 VDPWR.t442 VDPWR.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1138 VSS.t27 VDPWR.t1283 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1139 a_21951_5878# a_21785_5878# VDPWR.t154 VDPWR.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1140 ringtest_0.x4._06_ a_24004_6128# VDPWR.t1007 VDPWR.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.18575 ps=1.415 w=1 l=0.15
X1141 VDPWR.t1001 a_24968_5308# a_24895_5334# VDPWR.t1000 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1142 a_24465_6800# a_24336_6544# a_24045_6654# VSS.t764 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1143 VDPWR.t440 VSS.t1239 VDPWR.t439 VDPWR.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1144 a_22390_4566# a_22164_4362# a_22021_4220# VSS.t490 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1145 VDPWR.t1157 ringtest_0.x4.clknet_0_clk.t46 a_21395_6940# VDPWR.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1146 VDPWR.t195 ringtest_0.x4._18_ a_23529_6422# VDPWR.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1147 VDPWR.t1009 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP4.t2 VDPWR.t1008 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1148 a_12977_24040# ui_in[4].t19 VSS.t169 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X1149 VDPWR.t437 VSS.t1240 VDPWR.t436 VDPWR.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1150 ringtest_0.x4._10_ a_21785_8054# VSS.t180 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1151 VSS.t612 a_23879_6940# ringtest_0.x4.clknet_0_clk.t0 VSS.t611 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1152 a_23963_4790# ringtest_0.x4._15_ a_23891_4790# VSS.t568 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1153 VDPWR.t1058 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t17 VDPWR.t1057 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1154 VSS.t30 VDPWR.t1284 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1155 a_24895_5334# a_24361_5340# a_24800_5334# VDPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1156 a_23770_5308# ringtest_0.x4.net7 a_23899_5334# VDPWR.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1157 a_22399_9142# a_21845_9116# a_22052_9116# VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1158 a_21867_8054# ringtest_0.x4.net2.t11 a_21785_8054# VSS.t919 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1159 VDPWR.t434 VSS.t1241 VDPWR.t433 VDPWR.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1160 ringtest_0.x4._04_ a_22765_5308# VSS.t969 VSS.t968 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1161 VSS.t33 VDPWR.t1285 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1162 ringtest_0.x4.clknet_0_clk.t16 a_23879_6940# VDPWR.t395 VDPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1163 a_25364_5878# ringtest_0.x4.clknet_0_clk.t47 VSS.t546 VSS.t545 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1164 a_22399_8976# a_21845_8816# a_22052_8875# VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1165 a_20492_32319# ui_in[0].t9 VSS.t460 VSS.t459 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1166 ringtest_0.x3.x2.GP3 ringtest_0.x3.x2.GN3 VDPWR.t1137 VDPWR.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1167 VDPWR.t270 a_22373_5156# a_22541_5058# VDPWR.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1168 VDPWR.t431 VSS.t1242 VDPWR.t430 VDPWR.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1169 a_22052_8875# a_21845_8816# a_22228_8598# VDPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X1170 a_22228_8598# a_21981_8976# VDPWR.t1003 VDPWR.t1002 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1171 ringtest_0.x4._01_ ringtest_0.x4._12_ VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1172 VSS.t599 ringtest_0.drv_out.t27 a_23879_6940# VSS.t598 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1173 ringtest_0.x4._16_.t1 a_23381_4818# VDPWR.t1133 VDPWR.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1174 a_23151_5334# ringtest_0.x4.net6.t14 VDPWR.t327 VDPWR.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1175 VDPWR.t944 VDPWR.t942 muxtest_0.x2.nselect2 VDPWR.t943 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1176 VSS.t510 a_11845_23906# muxtest_0.x2.x2.GN1 VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1177 a_22295_3867# ringtest_0.x4.net4 VSS.t852 VSS.t851 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1178 VDPWR.t428 VSS.t1243 VDPWR.t427 VDPWR.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1179 a_13025_23980# ui_in[3].t19 VDPWR.t856 VDPWR.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X1180 VSS.t462 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B a_17377_14114# VSS.t461 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1181 VSS.t36 VDPWR.t1286 VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1182 VDPWR.t923 a_25055_3867# ringtest_0.x4.counter[5] VDPWR.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1183 VSS.t953 ringtest_0.x4.net6.t15 a_22983_5654# VSS.t952 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1184 VDPWR.t970 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 VDPWR.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1185 ringtest_0.x4.clknet_1_0__leaf_clk.t16 a_21395_6940# VDPWR.t1056 VDPWR.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 ringtest_0.x4.net2.n14 ringtest_0.x4.net2.t1 315.034
R1 ringtest_0.x4.net2.t0 ringtest_0.x4.net2.n14 265.769
R2 ringtest_0.x4.net2 ringtest_0.x4.net2.t0 262.318
R3 ringtest_0.x4.net2.n4 ringtest_0.x4.net2.t5 260.322
R4 ringtest_0.x4.net2.n9 ringtest_0.x4.net2.t10 241.536
R5 ringtest_0.x4.net2.n0 ringtest_0.x4.net2.t8 212.081
R6 ringtest_0.x4.net2.n1 ringtest_0.x4.net2.t3 212.081
R7 ringtest_0.x4.net2.n6 ringtest_0.x4.net2.t9 183.505
R8 ringtest_0.x4.net2.n4 ringtest_0.x4.net2.t2 175.169
R9 ringtest_0.x4.net2.n9 ringtest_0.x4.net2.t6 169.237
R10 ringtest_0.x4.net2.n10 ringtest_0.x4.net2.n9 159.952
R11 ringtest_0.x4.net2.n7 ringtest_0.x4.net2.n6 153.863
R12 ringtest_0.x4.net2.n3 ringtest_0.x4.net2.n2 152.698
R13 ringtest_0.x4.net2.n5 ringtest_0.x4.net2.n4 152
R14 ringtest_0.x4.net2.n0 ringtest_0.x4.net2.t7 139.78
R15 ringtest_0.x4.net2.n1 ringtest_0.x4.net2.t4 139.78
R16 ringtest_0.x4.net2.n6 ringtest_0.x4.net2.t11 114.532
R17 ringtest_0.x4.net2.n2 ringtest_0.x4.net2.n0 37.246
R18 ringtest_0.x4.net2.n8 ringtest_0.x4.net2.n5 34.4715
R19 ringtest_0.x4.net2.n2 ringtest_0.x4.net2.n1 24.1005
R20 ringtest_0.x4.net2.n12 ringtest_0.x4.net2.n3 18.9449
R21 ringtest_0.x4.net2.n13 ringtest_0.x4.net2.n12 14.916
R22 ringtest_0.x4.net2.n11 ringtest_0.x4.net2.n10 13.8005
R23 ringtest_0.x4.net2 ringtest_0.x4.net2.n7 10.8927
R24 ringtest_0.x4.net2.n14 ringtest_0.x4.net2.n13 8.72777
R25 ringtest_0.x4.net2.n8 ringtest_0.x4.net2 6.07742
R26 ringtest_0.x4.net2.n10 ringtest_0.x4.net2 3.33963
R27 ringtest_0.x4.net2.n10 ringtest_0.x4.net2 3.29747
R28 ringtest_0.x4.net2 ringtest_0.x4.net2.n13 3.29747
R29 ringtest_0.x4.net2.n11 ringtest_0.x4.net2.n8 3.19006
R30 ringtest_0.x4.net2.n3 ringtest_0.x4.net2 1.97868
R31 ringtest_0.x4.net2.n7 ringtest_0.x4.net2 1.97868
R32 ringtest_0.x4.net2.n5 ringtest_0.x4.net2 1.55726
R33 ringtest_0.x4.net2.n12 ringtest_0.x4.net2.n11 1.38649
R34 VSS.n3406 VSS.n64 4.7454e+06
R35 VSS.n318 VSS.n65 4.7454e+06
R36 VSS.n3406 VSS.n65 3.52e+06
R37 VSS.n360 VSS.n64 3.52e+06
R38 VSS.n3212 VSS.n173 3.3176e+06
R39 VSS.n3281 VSS.n3280 3.3176e+06
R40 VSS.n378 VSS.n376 2.347e+06
R41 VSS.n376 VSS.n64 2.3386e+06
R42 VSS.n3191 VSS.n173 2.3386e+06
R43 VSS.n3281 VSS.n3250 2.3386e+06
R44 VSS.n321 VSS.n66 2.15447e+06
R45 VSS.n3250 VSS.n3249 2.1446e+06
R46 VSS.n3192 VSS.n3191 2.1446e+06
R47 VSS.n3283 VSS.n3234 1.86572e+06
R48 VSS.n303 VSS.n65 1.2338e+06
R49 VSS.n334 VSS.n65 1.18072e+06
R50 VSS.n310 VSS.n309 1.1798e+06
R51 VSS.n3284 VSS.n3232 1.1798e+06
R52 VSS.n3229 VSS.n176 1.1798e+06
R53 VSS.n311 VSS.n310 1.17976e+06
R54 VSS.n3284 VSS.n3233 1.17976e+06
R55 VSS.n3229 VSS.n3228 1.17976e+06
R56 VSS.n376 VSS.t152 1.17724e+06
R57 VSS.n3250 VSS.t378 1.17707e+06
R58 VSS.n3191 VSS.t956 1.17707e+06
R59 VSS.n3405 VSS.t845 1.0027e+06
R60 VSS.n3077 VSS.n224 573621
R61 VSS.n323 VSS.n318 396385
R62 VSS.n362 VSS.n360 396385
R63 VSS.n3214 VSS.n3212 396385
R64 VSS.n3280 VSS.n3279 396385
R65 VSS.n318 VSS.n317 391216
R66 VSS.n360 VSS.n359 391216
R67 VSS.n3280 VSS.n3251 391216
R68 VSS.n3212 VSS.n3211 391216
R69 VSS.n3283 VSS.n3282 293853
R70 VSS.n3405 VSS.n66 291597
R71 VSS.n3290 VSS.n3289 86912.4
R72 VSS.n3290 VSS.n66 81673.6
R73 VSS.n3235 VSS.n67 72143.6
R74 VSS.n310 VSS.n172 66245.4
R75 VSS.n3061 VSS.n224 61252.6
R76 VSS.n3081 VSS.n172 52488.3
R77 VSS.n3289 VSS.n3288 52128.6
R78 VSS.n3394 VSS.n3393 38301.6
R79 VSS VSS.n175 35992.3
R80 VSS.n3407 VSS.n63 35421.6
R81 VSS.n3395 VSS.n3394 29605.7
R82 VSS.n3288 VSS.n173 29419.1
R83 VSS.n3288 VSS.n172 29145.5
R84 VSS.n399 VSS 25742.3
R85 VSS.n2394 VSS 23608
R86 VSS.n3404 VSS.n67 18854
R87 VSS.n3288 VSS.n3287 17410.5
R88 VSS.n341 VSS.n222 16580.9
R89 VSS.n2394 VSS.t757 13977.5
R90 VSS VSS.n173 13964.9
R91 VSS.n3231 VSS.n174 13854.2
R92 VSS.n369 VSS.n341 13333.2
R93 VSS.n3289 VSS.n74 13232.9
R94 VSS.n379 VSS.n371 11744.7
R95 VSS.n383 VSS.n371 11744.7
R96 VSS.n379 VSS.n372 11744.7
R97 VSS.n383 VSS.n372 11744.7
R98 VSS.n358 VSS.n346 11744.7
R99 VSS.n354 VSS.n346 11744.7
R100 VSS.n358 VSS.n348 11744.7
R101 VSS.n354 VSS.n348 11744.7
R102 VSS.n396 VSS.n282 11744.7
R103 VSS.n396 VSS.n388 11744.7
R104 VSS.n388 VSS.n280 11744.7
R105 VSS.n282 VSS.n280 11744.7
R106 VSS.n335 VSS.n284 11744.7
R107 VSS.n339 VSS.n284 11744.7
R108 VSS.n335 VSS.n285 11744.7
R109 VSS.n339 VSS.n285 11744.7
R110 VSS.n316 VSS.n293 11744.7
R111 VSS.n312 VSS.n293 11744.7
R112 VSS.n316 VSS.n294 11744.7
R113 VSS.n312 VSS.n294 11744.7
R114 VSS.n304 VSS.n298 11744.7
R115 VSS.n308 VSS.n298 11744.7
R116 VSS.n304 VSS.n299 11744.7
R117 VSS.n308 VSS.n299 11744.7
R118 VSS.n320 VSS.n291 11744.7
R119 VSS.n320 VSS.n292 11744.7
R120 VSS.n324 VSS.n292 11744.7
R121 VSS.n324 VSS.n291 11744.7
R122 VSS.n363 VSS.n342 11744.7
R123 VSS.n367 VSS.n342 11744.7
R124 VSS.n363 VSS.n343 11744.7
R125 VSS.n367 VSS.n343 11744.7
R126 VSS.n3248 VSS.n3236 11744.7
R127 VSS.n3243 VSS.n3236 11744.7
R128 VSS.n3248 VSS.n3238 11744.7
R129 VSS.n3243 VSS.n3238 11744.7
R130 VSS.n3266 VSS.n3263 11744.7
R131 VSS.n3266 VSS.n3264 11744.7
R132 VSS.n3268 VSS.n3263 11744.7
R133 VSS.n3268 VSS.n3264 11744.7
R134 VSS.n206 VSS.n197 11744.7
R135 VSS.n206 VSS.n199 11744.7
R136 VSS.n199 VSS.n196 11744.7
R137 VSS.n197 VSS.n196 11744.7
R138 VSS.n3210 VSS.n177 11744.7
R139 VSS.n3227 VSS.n177 11744.7
R140 VSS.n3210 VSS.n178 11744.7
R141 VSS.n3227 VSS.n178 11744.7
R142 VSS.n3194 VSS.n185 11744.7
R143 VSS.n3194 VSS.n186 11744.7
R144 VSS.n3196 VSS.n185 11744.7
R145 VSS.n3196 VSS.n186 11744.7
R146 VSS.n3215 VSS.n3204 11744.7
R147 VSS.n3215 VSS.n3208 11744.7
R148 VSS.n3205 VSS.n3204 11744.7
R149 VSS.n3208 VSS.n3205 11744.7
R150 VSS.n3391 VSS.n75 11744.7
R151 VSS.n3391 VSS.n76 11744.7
R152 VSS.n75 VSS.n73 11744.7
R153 VSS.n76 VSS.n73 11744.7
R154 VSS.n3278 VSS.n3252 11744.7
R155 VSS.n3278 VSS.n3254 11744.7
R156 VSS.n3257 VSS.n3252 11744.7
R157 VSS.n3257 VSS.n3254 11744.7
R158 VSS.n3076 VSS.n225 11744.7
R159 VSS.n3072 VSS.n226 11744.7
R160 VSS.n3076 VSS.n226 11744.7
R161 VSS.n3059 VSS.n3057 11744.7
R162 VSS.n3063 VSS.n3057 11744.7
R163 VSS.n3060 VSS.n3059 11744.7
R164 VSS.n3063 VSS.n3060 11744.7
R165 VSS.n370 VSS.n369 9554.71
R166 VSS.n3396 VSS.n3395 9243.96
R167 VSS.n3082 VSS.n3081 8452.32
R168 VSS.n3078 VSS.n222 7337.33
R169 VSS.n323 VSS.t989 7088.89
R170 VSS.t985 VSS.n321 7088.89
R171 VSS.n362 VSS.t984 7088.89
R172 VSS.n368 VSS.t986 7088.89
R173 VSS.n3214 VSS.t958 7088.89
R174 VSS.t961 VSS.n174 7088.89
R175 VSS.n3279 VSS.t382 7088.89
R176 VSS.t383 VSS.n3234 7088.89
R177 VSS.n303 VSS.t340 6925.66
R178 VSS.n309 VSS.t344 6925.66
R179 VSS.n317 VSS.t831 6925.66
R180 VSS.n311 VSS.t832 6925.66
R181 VSS.n3249 VSS.t860 6925.66
R182 VSS.t859 VSS.n3232 6925.66
R183 VSS.t1097 VSS.n3251 6925.66
R184 VSS.t1100 VSS.n3233 6925.66
R185 VSS.t357 VSS.n3192 6925.66
R186 VSS.t354 VSS.n176 6925.66
R187 VSS.n3211 VSS.t942 6925.66
R188 VSS.n3228 VSS.t947 6925.66
R189 VSS.n359 VSS.t838 6925.66
R190 VSS.t835 VSS.n283 6925.66
R191 VSS.n378 VSS.t341 6925.66
R192 VSS.n384 VSS.t347 6925.66
R193 VSS.n3081 VSS.t959 6843.4
R194 VSS.t989 VSS.n322 6733.33
R195 VSS.n322 VSS.t985 6733.33
R196 VSS.t984 VSS.n361 6733.33
R197 VSS.n361 VSS.t986 6733.33
R198 VSS.t958 VSS.n3213 6733.33
R199 VSS.n3213 VSS.t961 6733.33
R200 VSS.n3253 VSS.t382 6733.33
R201 VSS.n3253 VSS.t383 6733.33
R202 VSS.t340 VSS.n302 6578.29
R203 VSS.n302 VSS.t344 6578.29
R204 VSS.n297 VSS.t831 6578.29
R205 VSS.t832 VSS.n297 6578.29
R206 VSS.n3237 VSS.t860 6578.29
R207 VSS.n3237 VSS.t859 6578.29
R208 VSS.n3267 VSS.t1097 6578.29
R209 VSS.n3267 VSS.t1100 6578.29
R210 VSS.n3195 VSS.t357 6578.29
R211 VSS.n3195 VSS.t354 6578.29
R212 VSS.t942 VSS.n3209 6578.29
R213 VSS.n3209 VSS.t947 6578.29
R214 VSS.n347 VSS.t838 6578.29
R215 VSS.n347 VSS.t835 6578.29
R216 VSS.t341 VSS.n377 6578.29
R217 VSS.n377 VSS.t347 6578.29
R218 VSS.n334 VSS.t155 6418.9
R219 VSS.n340 VSS.t148 6418.9
R220 VSS.t155 VSS.n333 6096.95
R221 VSS.n333 VSS.t148 6096.95
R222 VSS.n386 VSS.n385 5782.24
R223 VSS.n385 VSS.n370 5742.37
R224 VSS.n479 VSS.n423 5452.27
R225 VSS.n479 VSS.n470 5452.27
R226 VSS.n423 VSS.n421 5452.27
R227 VSS.n470 VSS.n421 5452.27
R228 VSS.n467 VSS.n428 5452.27
R229 VSS.n459 VSS.n428 5452.27
R230 VSS.n467 VSS.n429 5452.27
R231 VSS.n459 VSS.n429 5452.27
R232 VSS.n489 VSS.n402 5452.27
R233 VSS.n419 VSS.n402 5452.27
R234 VSS.n489 VSS.n403 5452.27
R235 VSS.n419 VSS.n403 5452.27
R236 VSS.n434 VSS.n425 5452.27
R237 VSS.n461 VSS.n434 5452.27
R238 VSS.n437 VSS.n425 5452.27
R239 VSS.n461 VSS.n437 5452.27
R240 VSS.n413 VSS.n400 5452.27
R241 VSS.n416 VSS.n413 5452.27
R242 VSS.n414 VSS.n400 5452.27
R243 VSS.n416 VSS.n414 5452.27
R244 VSS.n439 VSS.n427 5452.27
R245 VSS.n458 VSS.n439 5452.27
R246 VSS.n440 VSS.n427 5452.27
R247 VSS.n458 VSS.n440 5452.27
R248 VSS.n481 VSS.n410 5452.27
R249 VSS.n411 VSS.n410 5452.27
R250 VSS.n481 VSS.n480 5452.27
R251 VSS.n480 VSS.n411 5452.27
R252 VSS.n451 VSS.n449 5452.27
R253 VSS.n453 VSS.n449 5452.27
R254 VSS.n452 VSS.n451 5452.27
R255 VSS.n453 VSS.n452 5452.27
R256 VSS.n2392 VSS.n1001 5434.88
R257 VSS.n2392 VSS.n1003 5434.88
R258 VSS.n1003 VSS.n1000 5434.88
R259 VSS.n1001 VSS.n1000 5434.88
R260 VSS.n3230 VSS.n3229 5417.76
R261 VSS.n3082 VSS.n3080 5047.41
R262 VSS VSS.t810 4888.89
R263 VSS.n3080 VSS.n3079 4736.53
R264 VSS.t810 VSS 4408.43
R265 VSS.n385 VSS.n384 4081.58
R266 VSS.n370 VSS.n283 4038.16
R267 VSS.t46 VSS.t37 3877.39
R268 VSS.t820 VSS.t43 3877.39
R269 VSS.n310 VSS.n222 3666.67
R270 VSS.n1010 VSS.n1007 3464.88
R271 VSS.n1013 VSS.n1007 3464.88
R272 VSS.n1010 VSS.n1008 3464.88
R273 VSS.n1013 VSS.n1008 3464.88
R274 VSS.n3230 VSS.n175 3363.82
R275 VSS VSS.t696 3346.36
R276 VSS.t430 VSS 3346.36
R277 VSS.t902 VSS 3346.36
R278 VSS.t276 VSS 3346.36
R279 VSS VSS.t281 3346.36
R280 VSS VSS.t208 3346.36
R281 VSS VSS.t73 3346.36
R282 VSS.n3062 VSS.n3061 3340.87
R283 VSS.n3078 VSS.n3077 3323.88
R284 VSS.n198 VSS.n175 3119.26
R285 VSS.t845 VSS.n3404 3111.89
R286 VSS.t34 VSS.t793 3101.92
R287 VSS.t451 VSS.t779 3101.92
R288 VSS.t782 VSS.t823 3101.92
R289 VSS.n386 VSS.n224 2996.82
R290 VSS.n2031 VSS 2973.14
R291 VSS.n3284 VSS.n3283 2937.79
R292 VSS.n172 VSS.n66 2904
R293 VSS.n369 VSS.n368 2881.39
R294 VSS VSS.t259 2857.47
R295 VSS VSS.t52 2857.47
R296 VSS.t422 VSS 2857.47
R297 VSS.t25 VSS 2857.47
R298 VSS.t40 VSS 2857.47
R299 VSS VSS.t688 2857.47
R300 VSS.n3285 VSS.n3284 2647.82
R301 VSS.n341 VSS.n340 2595.64
R302 VSS.n399 VSS.n398 2555.51
R303 VSS.n1222 VSS 2552.48
R304 VSS.t1024 VSS.t28 2495.02
R305 VSS.n2037 VSS 2469.73
R306 VSS VSS.t58 2452.87
R307 VSS VSS.t217 2452.87
R308 VSS.t815 VSS.t236 2326.44
R309 VSS.t79 VSS.t193 2326.44
R310 VSS.t242 VSS.t85 2326.44
R311 VSS VSS.t248 2081.99
R312 VSS.t425 VSS 2081.99
R313 VSS.n3079 VSS.n223 2065.3
R314 VSS.n198 VSS.t1123 2053.05
R315 VSS.n3285 VSS.n3231 2012.27
R316 VSS.n207 VSS.t1123 1950.07
R317 VSS.n2036 VSS.t64 1938.7
R318 VSS.t1126 VSS.n207 1926.65
R319 VSS.n2035 VSS.n1222 1896.67
R320 VSS.n2035 VSS.n2034 1896.67
R321 VSS.n2034 VSS.n2033 1896.67
R322 VSS.n2033 VSS.n2032 1896.67
R323 VSS.n2032 VSS.n2031 1896.67
R324 VSS.t248 VSS 1812.26
R325 VSS VSS.t34 1795.4
R326 VSS.t779 VSS 1795.4
R327 VSS VSS.t782 1795.4
R328 VSS VSS.t410 1795.4
R329 VSS.n3406 VSS.n3405 1791.03
R330 VSS VSS.t897 1786.97
R331 VSS.t245 VSS 1786.97
R332 VSS VSS.t205 1786.97
R333 VSS VSS.t70 1702.68
R334 VSS VSS.n1368 1677.39
R335 VSS.t2 VSS.t881 1593.1
R336 VSS.t766 VSS.t540 1593.1
R337 VSS.t493 VSS.t372 1593.1
R338 VSS.t306 VSS.t338 1584.67
R339 VSS.t491 VSS.t927 1584.67
R340 VSS.t117 VSS.t187 1567.82
R341 VSS.t696 VSS.t211 1550.96
R342 VSS.t259 VSS.t430 1550.96
R343 VSS.t52 VSS.t902 1550.96
R344 VSS.t843 VSS.t132 1550.96
R345 VSS.t413 VSS.t276 1550.96
R346 VSS.t281 VSS.t785 1550.96
R347 VSS.t208 VSS.t25 1550.96
R348 VSS.t73 VSS.t40 1550.96
R349 VSS.t688 VSS.t245 1550.96
R350 VSS.n3084 VSS.t6 1550.96
R351 VSS.n3083 VSS.n3080 1530.43
R352 VSS VSS.t442 1502.01
R353 VSS.n491 VSS.n399 1445.53
R354 VSS.t332 VSS.t549 1416.09
R355 VSS VSS.t233 1407.66
R356 VSS.t256 VSS 1407.66
R357 VSS VSS.t671 1407.66
R358 VSS.t31 VSS 1407.66
R359 VSS.t828 VSS 1407.66
R360 VSS VSS.t419 1407.66
R361 VSS VSS.t251 1399.23
R362 VSS.t572 VSS.t478 1399.23
R363 VSS.t4 VSS 1390.8
R364 VSS.t211 VSS 1306.51
R365 VSS.t793 VSS 1306.51
R366 VSS VSS.t88 1306.51
R367 VSS.t897 VSS 1306.51
R368 VSS VSS.t413 1306.51
R369 VSS VSS.t451 1306.51
R370 VSS.t64 VSS 1306.51
R371 VSS.t264 VSS 1306.51
R372 VSS.t785 VSS 1306.51
R373 VSS.t823 VSS 1306.51
R374 VSS.t273 VSS 1306.51
R375 VSS VSS.t220 1306.51
R376 VSS.t28 VSS 1306.51
R377 VSS VSS.t49 1306.51
R378 VSS.t205 VSS 1306.51
R379 VSS.n2938 VSS.n522 1294.86
R380 VSS.t1054 VSS 1289.66
R381 VSS VSS.t887 1289.66
R382 VSS.t1008 VSS 1289.66
R383 VSS VSS.t1119 1272.8
R384 VSS.n3463 VSS.t525 1229.99
R385 VSS.n3421 VSS.n3408 1198.25
R386 VSS.n3462 VSS.n3461 1198.25
R387 VSS.n3368 VSS.n86 1198.25
R388 VSS.n113 VSS.n112 1198.25
R389 VSS.n71 VSS.n68 1198.25
R390 VSS.n3403 VSS.n3402 1198.25
R391 VSS.n1420 VSS.n1419 1198.25
R392 VSS.n1931 VSS.n1917 1198.25
R393 VSS.n2030 VSS.n2029 1198.25
R394 VSS.n2498 VSS.n2395 1198.25
R395 VSS.n2986 VSS.n2985 1198.25
R396 VSS.n2988 VSS.n2987 1198.25
R397 VSS.n2036 VSS.n581 1196.22
R398 VSS.n2038 VSS.n2037 1196.22
R399 VSS.n3464 VSS.n3463 1194.5
R400 VSS.n3190 VSS.n3189 1194.5
R401 VSS.n3094 VSS.n219 1194.5
R402 VSS.n3085 VSS.n3084 1194.5
R403 VSS.n3316 VSS.n72 1194.5
R404 VSS.n2236 VSS.n2225 1194.5
R405 VSS.n2224 VSS.n2223 1194.5
R406 VSS.n2725 VSS.n731 1194.5
R407 VSS.n2790 VSS.n693 1194.5
R408 VSS.n1500 VSS.n1368 1194.5
R409 VSS.n2594 VSS.n842 1194.5
R410 VSS.n1661 VSS.n1581 1194.5
R411 VSS.n1916 VSS.n1915 1194.5
R412 VSS.t576 VSS.t398 1188.51
R413 VSS.n3446 VSS.n38 1171.32
R414 VSS.n3175 VSS.n208 1171.32
R415 VSS.n95 VSS.n94 1171.32
R416 VSS.n1916 VSS.t651 1146.36
R417 VSS VSS.t843 1137.93
R418 VSS.n3393 VSS.n3392 1105.32
R419 VSS.t768 VSS 1104.21
R420 VSS.t948 VSS 1078.93
R421 VSS.t720 VSS.t735 1078.93
R422 VSS.t644 VSS.t117 1078.93
R423 VSS.t286 VSS 1070.5
R424 VSS.t179 VSS 1036.78
R425 VSS.t478 VSS 1036.78
R426 VSS.n491 VSS.n490 1032.02
R427 VSS VSS.t422 1019.92
R428 VSS VSS.t46 1019.92
R429 VSS VSS.t820 1019.92
R430 VSS.t220 VSS 1019.92
R431 VSS.t334 VSS.t102 1003.07
R432 VSS.t606 VSS 1003.07
R433 VSS.t846 VSS.t848 1003.07
R434 VSS.n2173 VSS.n2172 999.607
R435 VSS.n2142 VSS.n2141 999.607
R436 VSS.n2680 VSS.n2679 999.607
R437 VSS.t92 VSS.t617 960.92
R438 VSS.t747 VSS.t659 952.49
R439 VSS.t338 VSS.t305 944.062
R440 VSS.t480 VSS.t318 944.062
R441 VSS.t555 VSS.t470 944.062
R442 VSS VSS.n2224 927.203
R443 VSS.n731 VSS 927.203
R444 VSS.n3463 VSS 918.774
R445 VSS VSS.t507 918.774
R446 VSS VSS.n70 918.774
R447 VSS.t236 VSS 918.774
R448 VSS.n2225 VSS 918.774
R449 VSS.t233 VSS 918.774
R450 VSS VSS.t79 918.774
R451 VSS.t251 VSS 918.774
R452 VSS.t85 VSS 918.774
R453 VSS VSS.n693 918.774
R454 VSS VSS.t256 918.774
R455 VSS.t671 VSS 918.774
R456 VSS VSS.t31 918.774
R457 VSS.t190 VSS 918.774
R458 VSS.t419 VSS 918.774
R459 VSS VSS.n72 918.774
R460 VSS.t476 VSS 918.774
R461 VSS.n3084 VSS 918.774
R462 VSS.t509 VSS 918.774
R463 VSS.t303 VSS.t828 910.346
R464 VSS.t6 VSS.t1004 910.346
R465 VSS.n1419 VSS 901.917
R466 VSS.n1917 VSS 901.917
R467 VSS.t100 VSS.t308 893.487
R468 VSS.t740 VSS.t326 893.487
R469 VSS.n1432 VSS.n1431 870.4
R470 VSS.n1222 VSS 851.341
R471 VSS VSS.n2035 851.341
R472 VSS.t102 VSS.t100 851.341
R473 VSS.n2034 VSS 851.341
R474 VSS.n2033 VSS 851.341
R475 VSS.n2032 VSS 851.341
R476 VSS.t495 VSS.t515 851.341
R477 VSS.n2031 VSS 851.341
R478 VSS VSS.t854 851.341
R479 VSS VSS.n3082 851.341
R480 VSS.t578 VSS.t164 842.913
R481 VSS.n3080 VSS.n222 839.237
R482 VSS.t305 VSS.t101 834.484
R483 VSS.t101 VSS.t334 834.484
R484 VSS.t754 VSS.t162 834.484
R485 VSS.t569 VSS.t362 834.484
R486 VSS.t739 VSS.t1018 834.484
R487 VSS.t950 VSS.t516 834.484
R488 VSS.t316 VSS.t649 834.484
R489 VSS.t293 VSS.t751 826.054
R490 VSS.t358 VSS.t1058 826.054
R491 VSS.t940 VSS.t491 826.054
R492 VSS.t214 VSS.t99 826.054
R493 VSS.t490 VSS.t846 826.054
R494 VSS.t113 VSS.t1010 826.054
R495 VSS.t141 VSS.t388 826.054
R496 VSS.t168 VSS.t106 826.054
R497 VSS.t841 VSS.t932 826.054
R498 VSS.t895 VSS.t572 809.196
R499 VSS.t1119 VSS.t403 809.196
R500 VSS.n314 VSS.n313 807.013
R501 VSS.n307 VSS.n306 807.013
R502 VSS.n319 VSS.n290 807.013
R503 VSS.n338 VSS.n337 807.013
R504 VSS.n382 VSS.n381 807.013
R505 VSS.n356 VSS.n355 807.013
R506 VSS.n366 VSS.n365 807.013
R507 VSS.n204 VSS.n203 807.013
R508 VSS.t796 VSS 805.538
R509 VSS.t308 VSS.t2 800.766
R510 VSS.t980 VSS.t566 800.766
R511 VSS.t656 VSS.t766 800.766
R512 VSS.t319 VSS.t1109 800.766
R513 VSS.t289 VSS.t934 792.337
R514 VSS.t564 VSS.t802 792.337
R515 VSS.t400 VSS.t230 792.337
R516 VSS.t995 VSS.t166 792.337
R517 VSS.t295 VSS.t917 792.337
R518 VSS.n315 VSS.n314 785.722
R519 VSS.n306 VSS.n305 785.722
R520 VSS.n325 VSS.n290 785.722
R521 VSS.n337 VSS.n336 785.722
R522 VSS.n381 VSS.n380 785.722
R523 VSS.n357 VSS.n356 785.722
R524 VSS.n365 VSS.n364 785.722
R525 VSS.n203 VSS.n202 785.722
R526 VSS.t936 VSS.t559 783.909
R527 VSS.t410 VSS.t425 775.48
R528 VSS.n3074 VSS.n3073 767.294
R529 VSS.n3058 VSS.n3056 767.294
R530 VSS.n313 VSS.n296 763.106
R531 VSS.n307 VSS.n300 763.106
R532 VSS.n319 VSS.n289 763.106
R533 VSS.n338 VSS.n286 763.106
R534 VSS.n382 VSS.n373 763.106
R535 VSS.n355 VSS.n353 763.106
R536 VSS.n366 VSS.n344 763.106
R537 VSS.n205 VSS.n204 763.106
R538 VSS.n3073 VSS.n3070 763.106
R539 VSS.n3058 VSS.n3055 763.106
R540 VSS.n394 VSS.n393 763.09
R541 VSS.n3245 VSS.n3244 763.09
R542 VSS.n3269 VSS.n3262 763.09
R543 VSS.n3226 VSS.n3225 763.09
R544 VSS.n3207 VSS.n3206 763.09
R545 VSS.n3197 VSS.n184 763.09
R546 VSS.n3389 VSS.n3388 763.09
R547 VSS.n3259 VSS.n3258 763.09
R548 VSS.t1105 VSS.t214 758.621
R549 VSS.t1113 VSS.t558 758.621
R550 VSS.t922 VSS.t130 750.192
R551 VSS.n296 VSS.n295 748.977
R552 VSS.n301 VSS.n300 748.977
R553 VSS.n332 VSS.n286 748.977
R554 VSS.n345 VSS.n344 748.977
R555 VSS.n326 VSS.n289 748.977
R556 VSS.n375 VSS.n373 748.977
R557 VSS.n353 VSS.n352 748.977
R558 VSS.n205 VSS.n201 748.977
R559 VSS.t927 VSS.t877 741.763
R560 VSS.t1001 VSS.t400 741.763
R561 VSS.t1068 VSS.t973 741.763
R562 VSS.t893 VSS.t774 741.763
R563 VSS.n393 VSS.n392 732.236
R564 VSS.n3246 VSS.n3245 732.236
R565 VSS.n3270 VSS.n3269 732.236
R566 VSS.n3225 VSS.n3224 732.236
R567 VSS.n3207 VSS.n3202 732.236
R568 VSS.n3198 VSS.n3197 732.236
R569 VSS.n3388 VSS.n3387 732.236
R570 VSS.n3276 VSS.n3259 732.236
R571 VSS.t992 VSS.t922 724.904
R572 VSS.t474 VSS.t594 724.904
R573 VSS.t619 VSS.t641 724.904
R574 VSS.t625 VSS.t621 724.904
R575 VSS.t639 VSS.t637 724.904
R576 VSS.t635 VSS.t639 724.904
R577 VSS.t667 VSS.t663 724.904
R578 VSS.t663 VSS.t726 724.904
R579 VSS.t726 VSS.t665 724.904
R580 VSS.t665 VSS.t1036 724.904
R581 VSS.t1036 VSS.t1042 724.904
R582 VSS.t1046 VSS.t1050 724.904
R583 VSS.t1050 VSS.t1040 724.904
R584 VSS.t1040 VSS.t1044 724.904
R585 VSS.t1044 VSS.t1048 724.904
R586 VSS.t1048 VSS.t1038 724.904
R587 VSS.t1022 VSS.t1028 724.904
R588 VSS.t1028 VSS.t1032 724.904
R589 VSS.t1032 VSS.t1034 724.904
R590 VSS.t1034 VSS.t1026 724.904
R591 VSS.t1026 VSS.t1030 724.904
R592 VSS.t1030 VSS.t1020 724.904
R593 VSS.t1076 VSS.t1072 724.904
R594 VSS.t1070 VSS.t1066 724.904
R595 VSS.t1082 VSS.t1084 724.904
R596 VSS.t724 VSS.t1117 724.904
R597 VSS.t1117 VSS.t722 724.904
R598 VSS.t538 VSS.t1013 724.904
R599 VSS.t598 VSS.t552 716.476
R600 VSS.t1092 VSS.t196 716.476
R601 VSS.t398 VSS.t533 716.476
R602 VSS.t542 VSS.t1107 716.476
R603 VSS.n3392 VSS.n74 709.47
R604 VSS.t660 VSS.t1060 708.047
R605 VSS.t291 VSS.t289 708.047
R606 VSS.t0 VSS.t1056 708.047
R607 VSS.t143 VSS.t648 708.047
R608 VSS.n3395 VSS.n70 708.047
R609 VSS.t104 VSS.t584 708.047
R610 VSS.t156 VSS.t158 708.047
R611 VSS.t350 VSS.t348 708.047
R612 VSS.t170 VSS.t172 708.047
R613 VSS.t176 VSS.t174 708.047
R614 VSS.t513 VSS.t511 708.047
R615 VSS.t499 VSS.t497 708.047
R616 VSS.t503 VSS.t501 708.047
R617 VSS.t871 VSS.t873 708.047
R618 VSS.n3291 VSS.n3290 708.047
R619 VSS.t132 VSS.t920 708.047
R620 VSS.t920 VSS.t923 708.047
R621 VSS.t923 VSS.t133 708.047
R622 VSS.t111 VSS.t306 708.047
R623 VSS.t881 VSS.t4 708.047
R624 VSS.t8 VSS.t286 708.047
R625 VSS.t566 VSS.t564 708.047
R626 VSS.t519 VSS.t578 708.047
R627 VSS.t1002 VSS.t1115 708.047
R628 VSS.t954 VSS.t951 708.047
R629 VSS.t891 VSS.t855 708.047
R630 VSS.t762 VSS.t948 708.047
R631 VSS.t857 VSS.t938 708.047
R632 VSS.t743 VSS.t741 708.047
R633 VSS.t488 VSS.t320 708.047
R634 VSS.t669 VSS.t313 708.047
R635 VSS.t854 VSS.t303 708.047
R636 VSS.t556 VSS.t109 708.047
R637 VSS.n3394 VSS.n72 708.047
R638 VSS.t715 VSS.t791 708.047
R639 VSS.t166 VSS.t115 708.047
R640 VSS.t885 VSS.t839 708.047
R641 VSS.t966 VSS.t728 708.047
R642 VSS.t680 VSS.t705 708.047
R643 VSS.t917 VSS.t997 708.047
R644 VSS.t139 VSS.t883 708.047
R645 VSS.t317 VSS.t547 708.047
R646 VSS.t405 VSS.t631 699.617
R647 VSS.t617 VSS.t590 691.188
R648 VSS.t709 VSS.t768 691.188
R649 VSS.t600 VSS.t545 691.188
R650 VSS.t468 VSS 682.76
R651 VSS.n208 VSS.t717 681.482
R652 VSS.n94 VSS.t805 681.482
R653 VSS.t613 VSS.t137 674.331
R654 VSS.t1084 VSS 674.331
R655 VSS.t178 VSS.t119 674.331
R656 VSS.t586 VSS.t538 674.331
R657 VSS.t850 VSS.t940 657.471
R658 VSS.t99 VSS.t364 657.471
R659 VSS.t386 VSS.t740 657.471
R660 VSS.t1016 VSS.t322 657.471
R661 VSS VSS.t61 649.043
R662 VSS.t952 VSS.t749 640.614
R663 VSS.t659 VSS.t328 640.614
R664 VSS.n3291 VSS 632.184
R665 VSS VSS.t815 632.184
R666 VSS.n2224 VSS 632.184
R667 VSS.n2225 VSS 632.184
R668 VSS.t193 VSS 632.184
R669 VSS.n2037 VSS 632.184
R670 VSS VSS.n2036 632.184
R671 VSS VSS.t242 632.184
R672 VSS VSS.n731 632.184
R673 VSS VSS.n693 632.184
R674 VSS.t70 VSS 632.184
R675 VSS.n1368 VSS 632.184
R676 VSS.t592 VSS.t611 632.184
R677 VSS.n1419 VSS 632.184
R678 VSS.t58 VSS 632.184
R679 VSS.t1088 VSS.t602 632.184
R680 VSS VSS.n842 632.184
R681 VSS.t217 VSS 632.184
R682 VSS.n1917 VSS 632.184
R683 VSS.t1066 VSS.t14 623.755
R684 VSS.t1062 VSS.t755 615.327
R685 VSS.n1581 VSS.t1088 615.327
R686 VSS.t1090 VSS.t1103 615.327
R687 VSS.t91 VSS.t737 615.327
R688 VSS.t994 VSS.t128 606.898
R689 VSS.t919 VSS.t994 606.898
R690 VSS.t82 VSS.t1024 606.898
R691 VSS.t655 VSS.t1080 606.898
R692 VSS.t397 VSS.t330 606.898
R693 VSS.t735 VSS.t397 606.898
R694 VSS.t568 VSS.t644 606.898
R695 VSS.t894 VSS.t568 606.898
R696 VSS.t889 VSS.t374 606.898
R697 VSS.t239 VSS.n38 606.351
R698 VSS.n70 VSS.n69 599.125
R699 VSS.n3292 VSS.n3291 599.125
R700 VSS.t641 VSS.t964 598.467
R701 VSS.t968 VSS.t747 598.467
R702 VSS.t575 VSS.t367 598.467
R703 VSS.t734 VSS.t505 598.467
R704 VSS.t301 VSS.t554 598.467
R705 VSS.t765 VSS.t627 590.038
R706 VSS VSS.t850 581.61
R707 VSS.t615 VSS.t482 581.61
R708 VSS VSS.t857 581.61
R709 VSS.t608 VSS.t1111 573.181
R710 VSS.n3061 VSS.n175 570.136
R711 VSS VSS.t660 564.751
R712 VSS VSS.t0 564.751
R713 VSS.t648 VSS 564.751
R714 VSS.n398 VSS 564.751
R715 VSS VSS.t104 564.751
R716 VSS VSS.t156 564.751
R717 VSS VSS.t350 564.751
R718 VSS VSS.t170 564.751
R719 VSS VSS.t176 564.751
R720 VSS VSS.t513 564.751
R721 VSS VSS.t499 564.751
R722 VSS VSS.t503 564.751
R723 VSS VSS.t871 564.751
R724 VSS.n2394 VSS 564.751
R725 VSS.n2394 VSS 564.751
R726 VSS.t128 VSS 564.751
R727 VSS.n2394 VSS 564.751
R728 VSS.n2394 VSS 564.751
R729 VSS.t327 VSS.t384 564.751
R730 VSS.n2394 VSS 564.751
R731 VSS VSS.t853 564.751
R732 VSS.n2394 VSS 564.751
R733 VSS.t791 VSS 564.751
R734 VSS.t839 VSS 564.751
R735 VSS VSS.t966 564.751
R736 VSS.n3393 VSS 564.751
R737 VSS.t297 VSS 564.751
R738 VSS.t705 VSS 564.751
R739 VSS.t883 VSS 564.751
R740 VSS VSS.t317 564.751
R741 VSS.t459 VSS.t525 563.702
R742 VSS VSS.t980 556.322
R743 VSS.t963 VSS.t633 556.322
R744 VSS.t396 VSS.t650 556.322
R745 VSS VSS.t919 547.894
R746 VSS VSS.t606 547.894
R747 VSS VSS.t1001 547.894
R748 VSS VSS.t1105 547.894
R749 VSS.t309 VSS.t657 547.894
R750 VSS.t362 VSS 547.894
R751 VSS.t324 VSS.t495 547.894
R752 VSS VSS.t894 547.894
R753 VSS VSS.t8 539.465
R754 VSS VSS.t416 539.465
R755 VSS.t907 VSS 531.034
R756 VSS.t37 VSS 531.034
R757 VSS.t43 VSS 531.034
R758 VSS VSS.t223 531.034
R759 VSS.t685 VSS.t126 526.468
R760 VSS.t184 VSS.t143 522.606
R761 VSS VSS.t92 522.606
R762 VSS.t1086 VSS 522.606
R763 VSS.t728 VSS.t799 522.606
R764 VSS.n3083 VSS.t297 522.606
R765 VSS.t547 VSS.t712 522.606
R766 VSS VSS.t179 514.177
R767 VSS.t121 VSS.t913 514.177
R768 VSS VSS.t480 514.177
R769 VSS.t1015 VSS.t754 505.748
R770 VSS VSS.t12 505.748
R771 VSS.t55 VSS.t1046 497.318
R772 VSS.t974 VSS.t1064 497.318
R773 VSS VSS.t889 497.318
R774 VSS.t1018 VSS.t121 488.889
R775 VSS VSS.t967 480.461
R776 VSS.t962 VSS.t623 480.461
R777 VSS.t1074 VSS.t653 480.461
R778 VSS.t164 VSS 480.461
R779 VSS VSS.t536 480.461
R780 VSS.t366 VSS 480.461
R781 VSS.t96 VSS 480.461
R782 VSS VSS.t677 473.495
R783 VSS VSS.t19 473.495
R784 VSS VSS.t674 473.495
R785 VSS.n2395 VSS.t693 465.17
R786 VSS VSS.t598 463.603
R787 VSS.t623 VSS.t1095 463.603
R788 VSS.t629 VSS.t360 463.603
R789 VSS.t717 VSS 459.26
R790 VSS.t805 VSS 459.26
R791 VSS.t657 VSS.t977 455.173
R792 VSS.t869 VSS.t324 455.173
R793 VSS VSS.t319 455.173
R794 VSS.t318 VSS.t770 455.173
R795 VSS VSS.t656 446.743
R796 VSS.t973 VSS 446.743
R797 VSS VSS.t753 446.743
R798 VSS VSS.t604 446.743
R799 VSS.t536 VSS.n1916 446.743
R800 VSS VSS.t315 446.743
R801 VSS.t288 VSS.t459 438.435
R802 VSS VSS.t576 438.315
R803 VSS VSS.t1022 429.885
R804 VSS.t323 VSS.t1012 429.885
R805 VSS.t649 VSS.t517 429.885
R806 VSS.t677 VSS 426.228
R807 VSS.t19 VSS 426.228
R808 VSS.t674 VSS 426.228
R809 VSS VSS.t685 426.228
R810 VSS.n3231 VSS.n3230 406.803
R811 VSS VSS.t486 404.599
R812 VSS VSS.t609 404.599
R813 VSS VSS.t762 404.599
R814 VSS.t369 VSS.t575 404.599
R815 VSS.t1012 VSS.t369 404.599
R816 VSS.t588 VSS.t734 404.599
R817 VSS.t517 VSS.t588 404.599
R818 VSS VSS.t669 404.599
R819 VSS.t975 VSS.t493 404.599
R820 VSS.t109 VSS 404.599
R821 VSS.t530 VSS.n74 403.983
R822 VSS.t507 VSS.t184 387.74
R823 VSS.t764 VSS.t629 387.74
R824 VSS.t730 VSS.t1062 387.74
R825 VSS.t799 VSS.t476 387.74
R826 VSS.t712 VSS.t509 387.74
R827 VSS.n281 VSS 384.901
R828 VSS.t693 VSS 380.899
R829 VSS.t770 VSS.t323 379.31
R830 VSS.t1013 VSS 379.31
R831 VSS.t470 VSS.t190 370.882
R832 VSS VSS.t943 370.37
R833 VSS.t1124 VSS 370.37
R834 VSS VSS.t1098 370.37
R835 VSS.t531 VSS 370.37
R836 VSS.n2030 VSS.t437 361.798
R837 VSS.n415 VSS.n407 354.26
R838 VSS.n415 VSS.n406 354.26
R839 VSS.n418 VSS.n405 354.26
R840 VSS.n418 VSS.n417 354.26
R841 VSS.n478 VSS.n477 354.26
R842 VSS.n477 VSS.n476 354.26
R843 VSS.n445 VSS.n408 354.26
R844 VSS.n466 VSS.n430 354.26
R845 VSS.n466 VSS.n465 354.26
R846 VSS.n435 VSS.n432 354.26
R847 VSS.n436 VSS.n435 354.26
R848 VSS.n443 VSS.n442 354.26
R849 VSS.n444 VSS.n443 354.26
R850 VSS.n2391 VSS.n1004 353.13
R851 VSS.n2391 VSS.n2390 353.13
R852 VSS.n2539 VSS.n947 352
R853 VSS VSS.t288 349.704
R854 VSS VSS.t682 341.574
R855 VSS VSS.t67 341.574
R856 VSS VSS.t448 341.574
R857 VSS.t830 VSS.n3462 337.166
R858 VSS.t633 VSS.t764 337.166
R859 VSS.t1064 VSS.t730 337.166
R860 VSS.t753 VSS 337.166
R861 VSS.n112 VSS.t929 337.166
R862 VSS.t108 VSS.n219 337.166
R863 VSS.n3190 VSS.n187 334.815
R864 VSS.n93 VSS.n86 334.815
R865 VSS.n2390 VSS.n2389 330.486
R866 VSS.t977 VSS.t1015 328.736
R867 VSS.t1115 VSS 328.736
R868 VSS.t604 VSS 328.736
R869 VSS.n3075 VSS.n3074 325.502
R870 VSS.n3064 VSS.n3056 325.502
R871 VSS.t910 VSS 325.171
R872 VSS.n2388 VSS.n1004 324.425
R873 VSS VSS.t270 323.541
R874 VSS.n3462 VSS.t751 320.307
R875 VSS.t315 VSS 320.307
R876 VSS.n112 VSS.t113 320.307
R877 VSS.n219 VSS.t168 320.307
R878 VSS.t313 VSS 311.877
R879 VSS.n3075 VSS.n3069 308.137
R880 VSS.n3065 VSS.n3064 308.137
R881 VSS.n3206 VSS.n3203 304.553
R882 VSS.n3258 VSS.n3256 304.553
R883 VSS.n395 VSS.n394 304.553
R884 VSS.n3244 VSS.n3242 304.553
R885 VSS.n3265 VSS.n3262 304.553
R886 VSS.n3193 VSS.n184 304.553
R887 VSS.n3226 VSS.n179 304.553
R888 VSS.n3390 VSS.n3389 304.553
R889 VSS.t364 VSS 303.449
R890 VSS.t163 VSS 303.449
R891 VSS.t374 VSS.t975 303.449
R892 VSS.n3287 VSS.n3286 299.892
R893 VSS VSS.t830 295.019
R894 VSS.t505 VSS.t396 295.019
R895 VSS VSS.t556 295.019
R896 VSS.t929 VSS 295.019
R897 VSS VSS.t108 295.019
R898 VSS.n1008 VSS.n1005 292.5
R899 VSS.t582 VSS.n1008 292.5
R900 VSS.n1007 VSS.n1006 292.5
R901 VSS.t582 VSS.n1007 292.5
R902 VSS VSS.t992 286.591
R903 VSS.t1038 VSS 286.591
R904 VSS VSS.t574 286.591
R905 VSS.n637 VSS.t993 281.25
R906 VSS.t584 VSS 278.161
R907 VSS.t158 VSS 278.161
R908 VSS.t348 VSS 278.161
R909 VSS.t172 VSS 278.161
R910 VSS.t174 VSS 278.161
R911 VSS.t511 VSS 278.161
R912 VSS.t497 VSS 278.161
R913 VSS.t501 VSS 278.161
R914 VSS.t873 VSS 278.161
R915 VSS.n387 VSS.t154 277.575
R916 VSS.t682 VSS 277.529
R917 VSS.t437 VSS 277.529
R918 VSS.t67 VSS 277.529
R919 VSS.t448 VSS 277.529
R920 VSS.n1168 VSS.t1211 276.531
R921 VSS.n1204 VSS.t1191 276.531
R922 VSS.n747 VSS.t1192 276.531
R923 VSS.t270 VSS 276.274
R924 VSS VSS.t910 276.274
R925 VSS.n533 VSS.t134 275.293
R926 VSS.n2593 VSS.t1116 275.293
R927 VSS.n1845 VSS.t605 275.293
R928 VSS VSS.t667 269.733
R929 VSS.t162 VSS.t178 269.733
R930 VSS.t384 VSS.t739 269.733
R931 VSS.n2105 VSS.t1201 269.488
R932 VSS.n2889 VSS.t1162 269.445
R933 VSS.n395 VSS.n389 266.349
R934 VSS.n3242 VSS.n3239 266.349
R935 VSS.n3265 VSS.n3260 266.349
R936 VSS.n3193 VSS.n182 266.349
R937 VSS.n3222 VSS.n179 266.349
R938 VSS.n3217 VSS.n3203 266.349
R939 VSS.n3390 VSS.n77 266.349
R940 VSS.n3256 VSS.n3255 266.349
R941 VSS.n561 VSS.t1232 265.317
R942 VSS.n819 VSS.t1152 265.317
R943 VSS.n1152 VSS.t1157 265.298
R944 VSS.n732 VSS.t1203 265.298
R945 VSS.t149 VSS.n397 263.652
R946 VSS.n397 VSS.t154 263.652
R947 VSS.n1172 VSS.t1167 262.784
R948 VSS.n1173 VSS.t1151 262.784
R949 VSS.n1175 VSS.t1172 262.784
R950 VSS.n2171 VSS.t1212 262.784
R951 VSS.n548 VSS.t1166 262.784
R952 VSS.n549 VSS.t1131 262.784
R953 VSS.n1185 VSS.t1206 262.784
R954 VSS.n1187 VSS.t1238 262.784
R955 VSS.n1188 VSS.t1146 262.784
R956 VSS.n1197 VSS.t1178 262.784
R957 VSS.n612 VSS.t1183 262.784
R958 VSS.n613 VSS.t1214 262.784
R959 VSS.n2842 VSS.t1187 262.784
R960 VSS.n2844 VSS.t1190 262.784
R961 VSS.n751 VSS.t1207 262.784
R962 VSS.n752 VSS.t1210 262.784
R963 VSS.n754 VSS.t1149 262.784
R964 VSS.n2678 VSS.t1155 262.784
R965 VSS.n1320 VSS.t1171 262.784
R966 VSS.n1321 VSS.t1175 262.784
R967 VSS.n806 VSS.t1150 262.784
R968 VSS.n807 VSS.t1156 262.784
R969 VSS.n1538 VSS.t1138 262.784
R970 VSS.n1540 VSS.t1144 262.784
R971 VSS.n883 VSS.t1237 262.784
R972 VSS.n884 VSS.t1243 262.784
R973 VSS.n1292 VSS.t1222 262.784
R974 VSS.n1837 VSS.t1227 262.784
R975 VSS.n966 VSS.t1202 262.784
R976 VSS.n967 VSS.t1208 262.784
R977 VSS.n2207 VSS.t1229 262.719
R978 VSS.n2269 VSS.t1196 262.719
R979 VSS.n1132 VSS.t1180 262.719
R980 VSS.n1150 VSS.t1230 262.719
R981 VSS.n2241 VSS.t1193 262.719
R982 VSS.n2945 VSS.t1234 262.719
R983 VSS.n2945 VSS.t1164 262.719
R984 VSS.n1220 VSS.t1198 262.719
R985 VSS.n2075 VSS.t1127 262.719
R986 VSS.n2063 VSS.t1160 262.719
R987 VSS.n2898 VSS.t1165 262.719
R988 VSS.n2840 VSS.t1188 262.719
R989 VSS.n2817 VSS.t1173 262.719
R990 VSS.n2714 VSS.t1169 262.719
R991 VSS.n712 VSS.t1128 262.719
R992 VSS.n2754 VSS.t1241 262.719
R993 VSS.n696 VSS.t1168 262.719
R994 VSS.n2784 VSS.t1133 262.719
R995 VSS.n2635 VSS.t1141 262.719
R996 VSS.n1353 VSS.t1221 262.719
R997 VSS.n1502 VSS.t1145 262.719
R998 VSS.n1251 VSS.t1215 262.719
R999 VSS.n2349 VSS.t1181 262.719
R1000 VSS.n497 VSS.t1176 262.719
R1001 VSS.n1104 VSS.t1143 262.719
R1002 VSS.n275 VSS.t1177 262.719
R1003 VSS.t934 VSS 261.303
R1004 VSS VSS.t111 261.303
R1005 VSS.t94 VSS 261.303
R1006 VSS.t1095 VSS.t619 261.303
R1007 VSS.t49 VSS 261.303
R1008 VSS.t580 VSS.t309 261.303
R1009 VSS.t223 VSS 261.303
R1010 VSS.t741 VSS 261.303
R1011 VSS.t97 VSS 261.303
R1012 VSS.t774 VSS 261.303
R1013 VSS.t1000 VSS 261.303
R1014 VSS.t330 VSS 261.303
R1015 VSS VSS.t995 261.303
R1016 VSS VSS.t295 261.303
R1017 VSS.t160 VSS.t76 260.675
R1018 VSS.n1664 VSS.t1220 259.082
R1019 VSS.n1926 VSS.t1135 259.082
R1020 VSS.n2542 VSS.t1216 259.082
R1021 VSS.n1745 VSS.t1186 259.082
R1022 VSS.n2438 VSS.t1163 259.082
R1023 VSS.n2354 VSS.t1235 259.082
R1024 VSS.n1061 VSS.t1223 259.082
R1025 VSS.n3037 VSS.t1242 259.082
R1026 VSS.n245 VSS.t1233 259.082
R1027 VSS.n447 VSS.n446 255.839
R1028 VSS.n446 VSS.n445 253.365
R1029 VSS.t802 VSS 252.875
R1030 VSS.t360 VSS.t625 252.875
R1031 VSS VSS.t580 252.875
R1032 VSS.t609 VSS.t869 252.875
R1033 VSS.t938 VSS 252.875
R1034 VSS.n648 VSS.t3 251
R1035 VSS.n648 VSS.t972 251
R1036 VSS.n2587 VSS.t748 251
R1037 VSS.n916 VSS.t385 251
R1038 VSS.n1286 VSS.t1110 251
R1039 VSS.n2559 VSS.t373 251
R1040 VSS.t943 VSS.t945 248.889
R1041 VSS.t355 VSS.t352 248.889
R1042 VSS.t1121 VSS.t1124 248.889
R1043 VSS.t1098 VSS.t1101 248.889
R1044 VSS.t861 VSS.t863 248.889
R1045 VSS.t528 VSS.t531 248.889
R1046 VSS.n1460 VSS.t593 245.82
R1047 VSS.n1704 VSS.t767 245.82
R1048 VSS.n1599 VSS.t601 245.82
R1049 VSS.n1914 VSS.t537 245.82
R1050 VSS VSS.t702 244.445
R1051 VSS.t88 VSS 244.445
R1052 VSS VSS.t273 244.445
R1053 VSS.t267 VSS 244.445
R1054 VSS.t627 VSS.t962 244.445
R1055 VSS.t416 VSS 244.445
R1056 VSS.t22 VSS 244.445
R1057 VSS VSS.t454 244.445
R1058 VSS.n663 VSS.t339 243.028
R1059 VSS.n663 VSS.t896 243.028
R1060 VSS.n1631 VSS.t120 243.028
R1061 VSS.n911 VSS.t955 243.028
R1062 VSS.n1242 VSS.t1120 243.028
R1063 VSS.n1882 VSS.t481 243.028
R1064 VSS.n1447 VSS.t618 242.067
R1065 VSS.n1556 VSS.t1069 242.067
R1066 VSS VSS.t202 241.573
R1067 VSS.n1495 VSS.t595 240.948
R1068 VSS.n1642 VSS.t546 240.948
R1069 VSS.n16 VSS.t935 240.575
R1070 VSS.n110 VSS.t996 240.575
R1071 VSS.n1393 VSS.t1096 238.675
R1072 VSS.n1678 VSS.t15 238.675
R1073 VSS.n875 VSS.t13 238.675
R1074 VSS.n2543 VSS.t471 238.675
R1075 VSS.n803 VSS.t1025 238.44
R1076 VSS VSS.t16 238.202
R1077 VSS.n7 VSS.t1055 237.327
R1078 VSS.n3098 VSS.t296 237.327
R1079 VSS.n3088 VSS.t1009 237.327
R1080 VSS.n3320 VSS.t888 237.327
R1081 VSS.n1438 VSS.t1106 237.327
R1082 VSS.n1515 VSS.t607 237.327
R1083 VSS.t653 VSS.t1070 236.016
R1084 VSS.t982 VSS 236.016
R1085 VSS.t951 VSS.t327 236.016
R1086 VSS.n2816 VSS.t565 235.607
R1087 VSS.n1971 VSS.n1970 234.667
R1088 VSS.n1624 VSS.t399 230.977
R1089 VSS.n1866 VSS.t771 230.977
R1090 VSS.n621 VSS.t131 229.833
R1091 VSS.n1612 VSS.n1611 228.294
R1092 VSS.n943 VSS.n942 228.294
R1093 VSS.t788 VSS 228.09
R1094 VSS.t1042 VSS.t55 227.587
R1095 VSS.t1080 VSS.t974 227.587
R1096 VSS.t486 VSS.t1074 227.587
R1097 VSS VSS.t484 227.587
R1098 VSS.n2043 VSS.t47 227.256
R1099 VSS.n1431 VSS.t668 226.708
R1100 VSS.n3144 VSS.t797 225.427
R1101 VSS.n3169 VSS.t718 225.427
R1102 VSS.n3089 VSS.t455 225.427
R1103 VSS.n3108 VSS.t713 225.427
R1104 VSS.n1014 VSS.n1006 225.13
R1105 VSS.n1009 VSS.n1006 225.13
R1106 VSS.t445 VSS.t181 224.931
R1107 VSS.n1715 VSS.t1139 224.196
R1108 VSS.n1124 VSS.t1137 224.102
R1109 VSS.n717 VSS.t1197 224.102
R1110 VSS.n2791 VSS.t42 223.282
R1111 VSS.n1449 VSS.n1413 222.691
R1112 VSS VSS.n3190 222.222
R1113 VSS.n208 VSS 222.222
R1114 VSS VSS.n86 222.222
R1115 VSS.n94 VSS 222.222
R1116 VSS.n690 VSS.t1132 221.972
R1117 VSS.n845 VSS.n843 221.804
R1118 VSS.t152 VSS.t150 221.451
R1119 VSS.n839 VSS.t1218 220.952
R1120 VSS.n840 VSS.t1224 220.952
R1121 VSS.n692 VSS.t221 219.972
R1122 VSS.n628 VSS.n626 218.506
R1123 VSS.n628 VSS.n627 218.506
R1124 VSS.n1709 VSS.n1551 218.506
R1125 VSS.n1656 VSS.n1585 218.506
R1126 VSS.n918 VSS.n853 218.506
R1127 VSS.n1853 VSS.n1288 218.506
R1128 VSS.n1891 VSS.n1890 218.506
R1129 VSS.n934 VSS.n933 218.506
R1130 VSS.n57 VSS.t1184 218.308
R1131 VSS.n3436 VSS.t1205 218.308
R1132 VSS.n25 VSS.t1240 218.308
R1133 VSS.n9 VSS.t1185 218.308
R1134 VSS.n212 VSS.t1159 218.308
R1135 VSS.n3167 VSS.t1154 218.308
R1136 VSS.n221 VSS.t1147 218.308
R1137 VSS.n3107 VSS.t1213 218.308
R1138 VSS.n3302 VSS.t1209 218.308
R1139 VSS.n98 VSS.t1161 218.308
R1140 VSS.n3322 VSS.t1142 218.308
R1141 VSS.n3346 VSS.t1195 218.308
R1142 VSS.n555 VSS.t1129 218.308
R1143 VSS.n619 VSS.t1179 218.308
R1144 VSS.n2883 VSS.t1130 218.308
R1145 VSS.n813 VSS.t1148 218.308
R1146 VSS.n1440 VSS.t1136 218.308
R1147 VSS.n1844 VSS.t1219 218.308
R1148 VSS.n1811 VSS.t1239 218.308
R1149 VSS.n996 VSS.t1134 218.308
R1150 VSS.n1604 VSS.n1603 218.13
R1151 VSS.n1133 VSS.t903 217.977
R1152 VSS.n1123 VSS.t431 217.977
R1153 VSS.n2761 VSS.t74 217.977
R1154 VSS.n2740 VSS.t209 217.977
R1155 VSS.n2217 VSS.t795 217.953
R1156 VSS.n730 VSS.t825 217.953
R1157 VSS.n2261 VSS.t261 217.892
R1158 VSS.n2759 VSS.t27 217.892
R1159 VSS.n212 VSS.t798 217.78
R1160 VSS.n3167 VSS.t719 217.78
R1161 VSS.n221 VSS.t456 217.78
R1162 VSS.n3107 VSS.t714 217.78
R1163 VSS.n1340 VSS.t249 216.933
R1164 VSS.n1125 VSS.t89 216.589
R1165 VSS.n718 VSS.t274 216.589
R1166 VSS.n2802 VSS.t803 216.579
R1167 VSS.n1549 VSS.t710 215.992
R1168 VSS.n1124 VSS.t90 214.487
R1169 VSS.n717 VSS.t275 214.487
R1170 VSS.n8 VSS.t704 214.456
R1171 VSS.n3 VSS.t703 214.456
R1172 VSS.n58 VSS.t701 214.456
R1173 VSS.n42 VSS.t700 214.456
R1174 VSS.n3437 VSS.t241 214.456
R1175 VSS.n40 VSS.t240 214.456
R1176 VSS.n26 VSS.t186 214.456
R1177 VSS.n32 VSS.t185 214.456
R1178 VSS.n81 VSS.t201 214.456
R1179 VSS.n3305 VSS.t200 214.456
R1180 VSS.n99 VSS.t807 214.456
R1181 VSS.n97 VSS.t806 214.456
R1182 VSS.n3345 VSS.t801 214.456
R1183 VSS.n3341 VSS.t800 214.456
R1184 VSS.n3323 VSS.t24 214.456
R1185 VSS.n115 VSS.t23 214.456
R1186 VSS.n554 VSS.t909 214.456
R1187 VSS.n554 VSS.t899 214.456
R1188 VSS.n546 VSS.t898 214.456
R1189 VSS.n525 VSS.t908 214.456
R1190 VSS.n521 VSS.t819 214.456
R1191 VSS.n2227 VSS.t818 214.456
R1192 VSS.n521 VSS.t812 214.456
R1193 VSS.n2227 VSS.t811 214.456
R1194 VSS.n2226 VSS.t54 214.456
R1195 VSS.n1151 VSS.t904 214.456
R1196 VSS.n1140 VSS.t53 214.456
R1197 VSS.n2263 VSS.t432 214.456
R1198 VSS.n2277 VSS.t260 214.456
R1199 VSS.n1157 VSS.t794 214.456
R1200 VSS.n2214 VSS.t36 214.456
R1201 VSS.n1158 VSS.t213 214.456
R1202 VSS.n2185 VSS.t35 214.456
R1203 VSS.n2178 VSS.t698 214.456
R1204 VSS.n1171 VSS.t212 214.456
R1205 VSS.n1171 VSS.t697 214.456
R1206 VSS.n1172 VSS.t827 214.456
R1207 VSS.n1172 VSS.t826 214.456
R1208 VSS.n1173 VSS.t817 214.456
R1209 VSS.n1173 VSS.t816 214.456
R1210 VSS.n1175 VSS.t255 214.456
R1211 VSS.n1175 VSS.t254 214.456
R1212 VSS.n2171 VSS.t238 214.456
R1213 VSS.n2171 VSS.t237 214.456
R1214 VSS.n548 VSS.t235 214.456
R1215 VSS.n548 VSS.t234 214.456
R1216 VSS.n549 VSS.t814 214.456
R1217 VSS.n549 VSS.t813 214.456
R1218 VSS.n2892 VSS.t822 214.456
R1219 VSS.n577 VSS.t44 214.456
R1220 VSS.n2064 VSS.t821 214.456
R1221 VSS.n576 VSS.t39 214.456
R1222 VSS.n2069 VSS.t48 214.456
R1223 VSS.n2060 VSS.t38 214.456
R1224 VSS.n2082 VSS.t424 214.456
R1225 VSS.n2099 VSS.t453 214.456
R1226 VSS.n2039 VSS.t423 214.456
R1227 VSS.n2117 VSS.t452 214.456
R1228 VSS.n1221 VSS.t781 214.456
R1229 VSS.n1216 VSS.t415 214.456
R1230 VSS.n2131 VSS.t780 214.456
R1231 VSS.n1200 VSS.t278 214.456
R1232 VSS.n1198 VSS.t414 214.456
R1233 VSS.n1198 VSS.t277 214.456
R1234 VSS.n1185 VSS.t195 214.456
R1235 VSS.n1185 VSS.t194 214.456
R1236 VSS.n1187 VSS.t429 214.456
R1237 VSS.n1187 VSS.t428 214.456
R1238 VSS.n1188 VSS.t692 214.456
R1239 VSS.n1188 VSS.t691 214.456
R1240 VSS.n1197 VSS.t81 214.456
R1241 VSS.n1197 VSS.t80 214.456
R1242 VSS.n2882 VSS.t66 214.456
R1243 VSS.n582 VSS.t65 214.456
R1244 VSS.n2882 VSS.t45 214.456
R1245 VSS.n618 VSS.t266 214.456
R1246 VSS.n610 VSS.t265 214.456
R1247 VSS.n612 VSS.t280 214.456
R1248 VSS.n612 VSS.t279 214.456
R1249 VSS.n613 VSS.t253 214.456
R1250 VSS.n613 VSS.t252 214.456
R1251 VSS.n2785 VSS.t75 214.456
R1252 VSS.n2764 VSS.t41 214.456
R1253 VSS.n690 VSS.t222 214.456
R1254 VSS.n680 VSS.t804 214.456
R1255 VSS.n2829 VSS.t246 214.456
R1256 VSS.n2841 VSS.t690 214.456
R1257 VSS.n2836 VSS.t689 214.456
R1258 VSS.n2841 VSS.t247 214.456
R1259 VSS.n2842 VSS.t708 214.456
R1260 VSS.n2842 VSS.t707 214.456
R1261 VSS.n2844 VSS.t258 214.456
R1262 VSS.n2844 VSS.t257 214.456
R1263 VSS.n710 VSS.t210 214.456
R1264 VSS.n2742 VSS.t26 214.456
R1265 VSS.n736 VSS.t824 214.456
R1266 VSS.n2721 VSS.t784 214.456
R1267 VSS.n737 VSS.t787 214.456
R1268 VSS.n2692 VSS.t783 214.456
R1269 VSS.n2685 VSS.t283 214.456
R1270 VSS.n750 VSS.t786 214.456
R1271 VSS.n750 VSS.t282 214.456
R1272 VSS.n751 VSS.t244 214.456
R1273 VSS.n751 VSS.t243 214.456
R1274 VSS.n752 VSS.t436 214.456
R1275 VSS.n752 VSS.t435 214.456
R1276 VSS.n754 VSS.t906 214.456
R1277 VSS.n754 VSS.t905 214.456
R1278 VSS.n2678 VSS.t87 214.456
R1279 VSS.n2678 VSS.t86 214.456
R1280 VSS.n1320 VSS.t72 214.456
R1281 VSS.n1320 VSS.t71 214.456
R1282 VSS.n1321 VSS.t809 214.456
R1283 VSS.n1321 VSS.t808 214.456
R1284 VSS.n1439 VSS.t216 214.456
R1285 VSS.n1418 VSS.t215 214.456
R1286 VSS.n2628 VSS.t57 214.456
R1287 VSS.n1429 VSS.t56 214.456
R1288 VSS.n781 VSS.t83 214.456
R1289 VSS.n812 VSS.t30 214.456
R1290 VSS.n804 VSS.t29 214.456
R1291 VSS.n812 VSS.t84 214.456
R1292 VSS.n806 VSS.t901 214.456
R1293 VSS.n806 VSS.t900 214.456
R1294 VSS.n807 VSS.t673 214.456
R1295 VSS.n807 VSS.t672 214.456
R1296 VSS.n1370 VSS.t232 214.456
R1297 VSS.n1516 VSS.t231 214.456
R1298 VSS.n1361 VSS.t269 214.456
R1299 VSS.n1313 VSS.t268 214.456
R1300 VSS.n1346 VSS.t250 214.456
R1301 VSS.n879 VSS.t418 214.456
R1302 VSS.n877 VSS.t417 214.456
R1303 VSS.n1663 VSS.t198 214.456
R1304 VSS.n1578 VSS.t197 214.456
R1305 VSS.n1700 VSS.t711 214.456
R1306 VSS.n1715 VSS.t51 214.456
R1307 VSS.n1541 VSS.t50 214.456
R1308 VSS.n1538 VSS.t227 214.456
R1309 VSS.n1538 VSS.t226 214.456
R1310 VSS.n1540 VSS.t60 214.456
R1311 VSS.n1540 VSS.t59 214.456
R1312 VSS.n839 VSS.t263 214.456
R1313 VSS.n839 VSS.t262 214.456
R1314 VSS.n840 VSS.t207 214.456
R1315 VSS.n840 VSS.t206 214.456
R1316 VSS.n883 VSS.t434 214.456
R1317 VSS.n883 VSS.t433 214.456
R1318 VSS.n884 VSS.t33 214.456
R1319 VSS.n884 VSS.t32 214.456
R1320 VSS.n971 VSS.t427 214.456
R1321 VSS.n963 VSS.t426 214.456
R1322 VSS.n971 VSS.t412 214.456
R1323 VSS.n960 VSS.t411 214.456
R1324 VSS.n2541 VSS.t192 214.456
R1325 VSS.n944 VSS.t191 214.456
R1326 VSS.n1925 VSS.t63 214.456
R1327 VSS.n1918 VSS.t62 214.456
R1328 VSS.n1945 VSS.t189 214.456
R1329 VSS.n1968 VSS.t188 214.456
R1330 VSS.n1843 VSS.t225 214.456
R1331 VSS.n1290 VSS.t224 214.456
R1332 VSS.n1292 VSS.t229 214.456
R1333 VSS.n1292 VSS.t228 214.456
R1334 VSS.n1837 VSS.t219 214.456
R1335 VSS.n1837 VSS.t218 214.456
R1336 VSS.n966 VSS.t441 214.456
R1337 VSS.n966 VSS.t440 214.456
R1338 VSS.n967 VSS.t421 214.456
R1339 VSS.n967 VSS.t420 214.456
R1340 VSS.n2437 VSS.t78 214.456
R1341 VSS.n2435 VSS.t77 214.456
R1342 VSS.n2417 VSS.t450 214.456
R1343 VSS.n2416 VSS.t449 214.456
R1344 VSS.n2474 VSS.t695 214.456
R1345 VSS.n2397 VSS.t694 214.456
R1346 VSS.n997 VSS.t18 214.456
R1347 VSS.n2509 VSS.t17 214.456
R1348 VSS.n1996 VSS.t69 214.456
R1349 VSS.n1995 VSS.t68 214.456
R1350 VSS.n1227 VSS.t439 214.456
R1351 VSS.n1225 VSS.t438 214.456
R1352 VSS.n1781 VSS.t684 214.456
R1353 VSS.n1780 VSS.t683 214.456
R1354 VSS.n1810 VSS.t204 214.456
R1355 VSS.n1763 VSS.t203 214.456
R1356 VSS.n1741 VSS.t790 214.456
R1357 VSS.n1746 VSS.t789 214.456
R1358 VSS.n240 VSS.t447 214.456
R1359 VSS.n246 VSS.t446 214.456
R1360 VSS.n3036 VSS.t183 214.456
R1361 VSS.n3039 VSS.t182 214.456
R1362 VSS.n258 VSS.t271 214.456
R1363 VSS.n3021 VSS.t272 214.456
R1364 VSS.n277 VSS.t679 214.456
R1365 VSS.n271 VSS.t678 214.456
R1366 VSS.n1060 VSS.t409 214.456
R1367 VSS.n1059 VSS.t408 214.456
R1368 VSS.n1098 VSS.t21 214.456
R1369 VSS.n1075 VSS.t20 214.456
R1370 VSS.n495 VSS.t676 214.456
R1371 VSS.n1080 VSS.t675 214.456
R1372 VSS.n1039 VSS.t911 214.456
R1373 VSS.n1032 VSS.t912 214.456
R1374 VSS.n2350 VSS.t687 214.456
R1375 VSS.n2338 VSS.t686 214.456
R1376 VSS.n2353 VSS.t444 214.456
R1377 VSS.n2351 VSS.t443 214.456
R1378 VSS.n1009 VSS.n1005 214.409
R1379 VSS.n1015 VSS.n1014 213.911
R1380 VSS.n3401 VSS.n3400 212.78
R1381 VSS.n1631 VSS.n1608 212.317
R1382 VSS.t311 VSS.t284 211.237
R1383 VSS.t853 VSS 210.728
R1384 VSS.n3287 VSS.t530 209.996
R1385 VSS.n2601 VSS.n836 207.965
R1386 VSS.n937 VSS.n936 207.965
R1387 VSS.n1373 VSS.n1372 206.909
R1388 VSS.n3286 VSS.n3285 206.876
R1389 VSS.n1671 VSS.n1670 205.971
R1390 VSS.n1466 VSS.n1396 205.899
R1391 VSS.n1469 VSS.n1468 205.899
R1392 VSS.n1398 VSS.n1397 205.481
R1393 VSS.n1572 VSS.n1571 205.481
R1394 VSS.n2626 VSS.n2625 205.385
R1395 VSS.n1449 VSS.n1412 204.692
R1396 VSS.n1476 VSS.n1475 204.692
R1397 VSS.n48 VSS.n44 204.457
R1398 VSS.n3310 VSS.n3309 204.457
R1399 VSS.n1939 VSS.n1937 204.457
R1400 VSS.n1939 VSS.n1938 204.457
R1401 VSS.n1921 VSS.n1919 204.457
R1402 VSS.n2823 VSS.n2822 204.201
R1403 VSS.n1249 VSS.n1248 204.201
R1404 VSS.n1263 VSS.n1262 204.201
R1405 VSS.n1425 VSS.n1422 202.724
R1406 VSS.n772 VSS.n771 202.724
R1407 VSS.n1484 VSS.n1387 202.724
R1408 VSS.n1655 VSS.n1586 202.724
R1409 VSS.n1598 VSS.n1597 202.724
R1410 VSS VSS.t1092 202.299
R1411 VSS.t326 VSS.t968 202.299
R1412 VSS.t855 VSS.t950 202.299
R1413 VSS.t372 VSS.t301 202.299
R1414 VSS.n780 VSS.n779 201.458
R1415 VSS.n1575 VSS.n1574 201.458
R1416 VSS.n1459 VSS.n1400 201.129
R1417 VSS.n2618 VSS.n784 201.129
R1418 VSS.n2620 VSS.n783 201.129
R1419 VSS.n1680 VSS.n1573 201.129
R1420 VSS.n2084 VSS.n2083 200.692
R1421 VSS.n1702 VSS.n1701 200.692
R1422 VSS.n2479 VSS.n2478 200.692
R1423 VSS.n3023 VSS.n3022 200.692
R1424 VSS.n2327 VSS.n2326 200.692
R1425 VSS.n2599 VSS.n838 200.516
R1426 VSS.n1285 VSS.n1284 200.516
R1427 VSS.n793 VSS.n792 200.508
R1428 VSS.n774 VSS.n773 200.508
R1429 VSS.n2634 VSS.n776 200.508
R1430 VSS.n1392 VSS.n1391 200.508
R1431 VSS.n1560 VSS.n1559 200.508
R1432 VSS.n1665 VSS.n1580 200.508
R1433 VSS.n1583 VSS.n1582 200.508
R1434 VSS.n3460 VSS.n15 200.231
R1435 VSS.n3452 VSS.n21 200.231
R1436 VSS.n3329 VSS.n3328 200.231
R1437 VSS.n108 VSS.n107 200.231
R1438 VSS.n1446 VSS.n1416 200.231
R1439 VSS.n845 VSS.n844 200.127
R1440 VSS.n1851 VSS.n1850 200.127
R1441 VSS.n30 VSS.n24 200.105
R1442 VSS.n3109 VSS.n3106 200.105
R1443 VSS.n3138 VSS.n214 200.105
R1444 VSS.n3348 VSS.n3343 200.105
R1445 VSS.n599 VSS.n597 199.739
R1446 VSS.n599 VSS.n598 199.739
R1447 VSS.n1494 VSS.n1374 199.739
R1448 VSS.n1629 VSS.n1610 199.739
R1449 VSS.n1272 VSS.n1271 199.739
R1450 VSS.n1823 VSS.n1758 199.739
R1451 VSS.n1818 VSS.n1762 199.739
R1452 VSS.n1805 VSS.n1767 199.739
R1453 VSS.n1784 VSS.n1783 199.739
R1454 VSS.n1992 VSS.n1991 199.739
R1455 VSS.n2519 VSS.n990 199.739
R1456 VSS.n999 VSS.n998 199.739
R1457 VSS.n2413 VSS.n2412 199.739
R1458 VSS.n2421 VSS.n2420 199.739
R1459 VSS.n2444 VSS.n2434 199.739
R1460 VSS.n1031 VSS.n1030 199.739
R1461 VSS.n682 VSS.n681 199.662
R1462 VSS.n657 VSS.n655 199.53
R1463 VSS.n657 VSS.n656 199.53
R1464 VSS.n1470 VSS.n1467 199.53
R1465 VSS.n1637 VSS.n1605 199.53
R1466 VSS.n917 VSS.n854 199.53
R1467 VSS.n1241 VSS.n1240 199.53
R1468 VSS.n1865 VSS.n1864 199.53
R1469 VSS.n940 VSS.n939 199.53
R1470 VSS.t956 VSS 198.519
R1471 VSS.t945 VSS 198.519
R1472 VSS VSS.t355 198.519
R1473 VSS VSS.t1121 198.519
R1474 VSS.t378 VSS 198.519
R1475 VSS.t1101 VSS 198.519
R1476 VSS VSS.t861 198.519
R1477 VSS VSS.t528 198.519
R1478 VSS VSS.n38 197.724
R1479 VSS.n3101 VSS.n3100 197.476
R1480 VSS.n3095 VSS.n218 197.476
R1481 VSS.n1359 VSS.n1307 197.476
R1482 VSS.n536 VSS.n535 196.831
R1483 VSS.n1694 VSS.n1558 196.589
R1484 VSS.n909 VSS.n859 196.589
R1485 VSS.n1352 VSS.n1310 196.442
R1486 VSS.n1483 VSS.n1388 196.442
R1487 VSS.n1673 VSS.n1577 196.442
R1488 VSS.n861 VSS.n860 196.442
R1489 VSS.n890 VSS.n878 196.442
R1490 VSS.n308 VSS.n307 195
R1491 VSS.n309 VSS.n308 195
R1492 VSS.n305 VSS.n304 195
R1493 VSS.n304 VSS.n303 195
R1494 VSS.n313 VSS.n312 195
R1495 VSS.n312 VSS.n311 195
R1496 VSS.n316 VSS.n315 195
R1497 VSS.n317 VSS.n316 195
R1498 VSS.n320 VSS.n319 195
R1499 VSS.n321 VSS.n320 195
R1500 VSS.n325 VSS.n324 195
R1501 VSS.n324 VSS.n323 195
R1502 VSS.n367 VSS.n366 195
R1503 VSS.n368 VSS.n367 195
R1504 VSS.n364 VSS.n363 195
R1505 VSS.n363 VSS.n362 195
R1506 VSS.n339 VSS.n338 195
R1507 VSS.n340 VSS.n339 195
R1508 VSS.n336 VSS.n335 195
R1509 VSS.n335 VSS.n334 195
R1510 VSS.n391 VSS.n282 195
R1511 VSS.n282 VSS.n281 195
R1512 VSS.n3244 VSS.n3243 195
R1513 VSS.n3243 VSS.n3232 195
R1514 VSS.n3248 VSS.n3247 195
R1515 VSS.n3249 VSS.n3248 195
R1516 VSS.n3264 VSS.n3262 195
R1517 VSS.n3264 VSS.n3233 195
R1518 VSS.n3263 VSS.n3261 195
R1519 VSS.n3263 VSS.n3251 195
R1520 VSS.n3206 VSS.n3205 195
R1521 VSS.n3205 VSS.n174 195
R1522 VSS.n3216 VSS.n3215 195
R1523 VSS.n3215 VSS.n3214 195
R1524 VSS.n186 VSS.n184 195
R1525 VSS.n186 VSS.n176 195
R1526 VSS.n185 VSS.n183 195
R1527 VSS.n3192 VSS.n185 195
R1528 VSS.n3227 VSS.n3226 195
R1529 VSS.n3228 VSS.n3227 195
R1530 VSS.n3210 VSS.n180 195
R1531 VSS.n3211 VSS.n3210 195
R1532 VSS.n3389 VSS.n76 195
R1533 VSS.n3286 VSS.n76 195
R1534 VSS.n202 VSS.n197 195
R1535 VSS.n197 VSS.n187 195
R1536 VSS.n204 VSS.n199 195
R1537 VSS.n199 VSS.n198 195
R1538 VSS.n3258 VSS.n3257 195
R1539 VSS.n3257 VSS.n3234 195
R1540 VSS.n3278 VSS.n3277 195
R1541 VSS.n3279 VSS.n3278 195
R1542 VSS.n3386 VSS.n75 195
R1543 VSS.n93 VSS.n75 195
R1544 VSS.n355 VSS.n354 195
R1545 VSS.n354 VSS.n283 195
R1546 VSS.n358 VSS.n357 195
R1547 VSS.n359 VSS.n358 195
R1548 VSS.n383 VSS.n382 195
R1549 VSS.n384 VSS.n383 195
R1550 VSS.n380 VSS.n379 195
R1551 VSS.n379 VSS.n378 195
R1552 VSS.n394 VSS.n388 195
R1553 VSS.n388 VSS.n387 195
R1554 VSS.n3074 VSS.n226 195
R1555 VSS.n226 VSS.t298 195
R1556 VSS.n3070 VSS.n225 195
R1557 VSS.n3060 VSS.n3056 195
R1558 VSS.t662 VSS.n3060 195
R1559 VSS.n3057 VSS.n3055 195
R1560 VSS.t662 VSS.n3057 195
R1561 VSS.n398 VSS.t149 194.406
R1562 VSS.t913 VSS.t386 193.87
R1563 VSS.t367 VSS.t1016 193.87
R1564 VSS.n2057 VSS.n2055 190.399
R1565 VSS.n1555 VSS.n1552 190.399
R1566 VSS.n2477 VSS.n2476 190.399
R1567 VSS.n263 VSS.n261 190.399
R1568 VSS.n2325 VSS.n2324 190.399
R1569 VSS.n1970 VSS.n1244 189.268
R1570 VSS.n947 VSS.n946 189.201
R1571 VSS.n3071 VSS.n225 188.968
R1572 VSS.t515 VSS.t954 185.441
R1573 VSS.t650 VSS.t1000 185.441
R1574 VSS.t1004 VSS.n3083 185.441
R1575 VSS.n438 VSS.t699 179.556
R1576 VSS.t523 VSS 177.529
R1577 VSS.t915 VSS 177.529
R1578 VSS.t145 VSS 177.529
R1579 VSS.t124 VSS 177.529
R1580 VSS.t930 VSS 177.529
R1581 VSS.t1058 VSS 177.012
R1582 VSS.t737 VSS.t569 177.012
R1583 VSS.t1109 VSS.t332 177.012
R1584 VSS.t322 VSS.t97 177.012
R1585 VSS VSS.t141 177.012
R1586 VSS VSS.t841 177.012
R1587 VSS.t150 VSS 176.633
R1588 VSS.n398 VSS 176.633
R1589 VSS.n3072 VSS.n3071 174.41
R1590 VSS.t202 VSS 174.157
R1591 VSS.t16 VSS 174.157
R1592 VSS.t611 VSS.t963 168.583
R1593 VSS.t484 VSS.t982 168.583
R1594 VSS.n387 VSS.n386 163.297
R1595 VSS.n3429 VSS.t991 162.471
R1596 VSS.n3424 VSS.t834 162.471
R1597 VSS.n3420 VSS.t343 162.471
R1598 VSS.n3415 VSS.t153 162.471
R1599 VSS.n3455 VSS.t290 162.471
R1600 VSS.n3376 VSS.t381 162.471
R1601 VSS.n3371 VSS.t1099 162.471
R1602 VSS.n3367 VSS.t864 162.471
R1603 VSS.n3362 VSS.t532 162.471
R1604 VSS.n3334 VSS.t167 162.471
R1605 VSS.n2986 VSS 162.179
R1606 VSS.n127 VSS.t880 162.022
R1607 VSS.n132 VSS.t337 162.022
R1608 VSS.n137 VSS.t349 162.022
R1609 VSS.n142 VSS.t868 162.022
R1610 VSS.n147 VSS.t865 162.022
R1611 VSS.n152 VSS.t512 162.022
R1612 VSS.n157 VSS.t777 162.022
R1613 VSS.n162 VSS.t775 162.022
R1614 VSS.n167 VSS.t876 162.022
R1615 VSS.n131 VSS.t105 162.022
R1616 VSS.n136 VSS.t157 162.022
R1617 VSS.n141 VSS.t466 162.022
R1618 VSS.n146 VSS.t171 162.022
R1619 VSS.n151 VSS.t177 162.022
R1620 VSS.n156 VSS.t535 162.022
R1621 VSS.n161 VSS.t500 162.022
R1622 VSS.n166 VSS.t504 162.022
R1623 VSS.n171 VSS.t872 162.022
R1624 VSS.n3460 VSS.t1061 160.046
R1625 VSS.n3452 VSS.t1057 160.046
R1626 VSS.n3329 VSS.t716 160.046
R1627 VSS.n108 VSS.t886 160.046
R1628 VSS.n127 VSS.t585 160.017
R1629 VSS.n132 VSS.t159 160.017
R1630 VSS.n137 VSS.t465 160.017
R1631 VSS.n142 VSS.t173 160.017
R1632 VSS.n147 VSS.t175 160.017
R1633 VSS.n152 VSS.t534 160.017
R1634 VSS.n157 VSS.t498 160.017
R1635 VSS.n162 VSS.t502 160.017
R1636 VSS.n167 VSS.t874 160.017
R1637 VSS.n60 VSS.t988 160.017
R1638 VSS.n3422 VSS.t837 160.017
R1639 VSS.n3411 VSS.t346 160.017
R1640 VSS.n39 VSS.t151 160.017
R1641 VSS.n3453 VSS.t292 160.017
R1642 VSS.n22 VSS.t1 160.017
R1643 VSS.n83 VSS.t379 160.017
R1644 VSS.n3369 VSS.t1102 160.017
R1645 VSS.n89 VSS.t862 160.017
R1646 VSS.n3360 VSS.t529 160.017
R1647 VSS.n3336 VSS.t116 160.017
R1648 VSS.n3353 VSS.t840 160.017
R1649 VSS.n131 VSS.t879 160.017
R1650 VSS.n136 VSS.t336 160.017
R1651 VSS.n141 VSS.t351 160.017
R1652 VSS.n146 VSS.t867 160.017
R1653 VSS.n151 VSS.t866 160.017
R1654 VSS.n156 VSS.t514 160.017
R1655 VSS.n161 VSS.t778 160.017
R1656 VSS.n166 VSS.t776 160.017
R1657 VSS.n171 VSS.t875 160.017
R1658 VSS.n16 VSS.t661 158.534
R1659 VSS.n110 VSS.t792 158.534
R1660 VSS.t10 VSS.n2030 157.304
R1661 VSS.n2395 VSS.t135 157.304
R1662 VSS.n3146 VSS.t960 157.291
R1663 VSS.n3148 VSS.t944 157.291
R1664 VSS.n191 VSS.t353 157.291
R1665 VSS.n192 VSS.t1125 157.291
R1666 VSS.n3097 VSS.t681 157.291
R1667 VSS.n3124 VSS.t918 157.291
R1668 VSS.n3117 VSS.t140 157.291
R1669 VSS.n3156 VSS.t957 155.286
R1670 VSS.n3150 VSS.t946 155.286
R1671 VSS.n3184 VSS.t356 155.286
R1672 VSS.n3178 VSS.t1122 155.286
R1673 VSS.n3129 VSS.t706 155.286
R1674 VSS.n3122 VSS.t998 155.286
R1675 VSS.n3115 VSS.t884 155.286
R1676 VSS.n904 VSS.t856 154.131
R1677 VSS.n2814 VSS.t9 152.381
R1678 VSS.n874 VSS.t892 152.381
R1679 VSS.n882 VSS.t939 152.381
R1680 VSS.n2085 VSS.n2084 152
R1681 VSS.n1703 VSS.n1702 152
R1682 VSS.n2478 VSS.n2411 152
R1683 VSS.n2326 VSS.n1034 152
R1684 VSS.n3024 VSS.n3023 152
R1685 VSS.n2803 VSS.t287 150.101
R1686 VSS.n882 VSS.t858 150.101
R1687 VSS.n2987 VSS.t407 149.954
R1688 VSS VSS.n3403 144.951
R1689 VSS.n848 VSS.t969 144.886
R1690 VSS.n1858 VSS.t333 144.886
R1691 VSS.t482 VSS.t596 143.296
R1692 VSS VSS.n842 143.296
R1693 VSS.t61 VSS 143.296
R1694 VSS.n474 VSS.n473 139.727
R1695 VSS.t662 VSS.n223 137.912
R1696 VSS.n3062 VSS.t662 137.912
R1697 VSS.t123 VSS 135.415
R1698 VSS.t631 VSS.t765 134.867
R1699 VSS.t1111 VSS.t743 134.867
R1700 VSS.t549 VSS.t608 134.867
R1701 VSS.t403 VSS.t316 134.867
R1702 VSS.n71 VSS.t376 133.507
R1703 VSS.t964 VSS.t615 126.438
R1704 VSS.n522 VSS.t844 124.688
R1705 VSS.n431 VSS.n430 123.882
R1706 VSS.t76 VSS 122.472
R1707 VSS.n879 VSS.t1231 121.927
R1708 VSS.n2417 VSS.t1228 121.927
R1709 VSS.n1996 VSS.t1158 121.927
R1710 VSS.n1227 VSS.t1225 121.927
R1711 VSS.n1781 VSS.t1170 121.927
R1712 VSS VSS.t1126 121.481
R1713 VSS VSS.t527 121.481
R1714 VSS.n3079 VSS.n3078 120.984
R1715 VSS.n3077 VSS.n3076 118.285
R1716 VSS.t596 VSS 118.008
R1717 VSS.t1020 VSS.t82 118.008
R1718 VSS.t1072 VSS.t655 118.008
R1719 VSS.t574 VSS.t488 118.008
R1720 VSS.n452 VSS.n448 117.001
R1721 VSS.n452 VSS.t467 117.001
R1722 VSS.n449 VSS.n447 117.001
R1723 VSS.n449 VSS.t467 117.001
R1724 VSS.n480 VSS.n412 117.001
R1725 VSS.n480 VSS.t551 117.001
R1726 VSS.n410 VSS.n408 117.001
R1727 VSS.t551 VSS.n410 117.001
R1728 VSS.n444 VSS.n440 117.001
R1729 VSS.n440 VSS.t643 117.001
R1730 VSS.n442 VSS.n439 117.001
R1731 VSS.t643 VSS.n439 117.001
R1732 VSS.n414 VSS.n407 117.001
R1733 VSS.n414 VSS.t371 117.001
R1734 VSS.n413 VSS.n406 117.001
R1735 VSS.n413 VSS.t371 117.001
R1736 VSS.n437 VSS.n436 117.001
R1737 VSS.t643 VSS.n437 117.001
R1738 VSS.n434 VSS.n432 117.001
R1739 VSS.t643 VSS.n434 117.001
R1740 VSS.n405 VSS.n403 117.001
R1741 VSS.t371 VSS.n403 117.001
R1742 VSS.n417 VSS.n402 117.001
R1743 VSS.t371 VSS.n402 117.001
R1744 VSS.n465 VSS.n429 117.001
R1745 VSS.t643 VSS.n429 117.001
R1746 VSS.n430 VSS.n428 117.001
R1747 VSS.t643 VSS.n428 117.001
R1748 VSS.n476 VSS.n421 117.001
R1749 VSS.t457 VSS.n421 117.001
R1750 VSS.n479 VSS.n478 117.001
R1751 VSS.t457 VSS.n479 117.001
R1752 VSS.n972 VSS.t1200 116.734
R1753 VSS.n1347 VSS.t1189 116.734
R1754 VSS.n1978 VSS.n1977 114.377
R1755 VSS.n1509 VSS.n1365 110.349
R1756 VSS.n1889 VSS.n1270 110.349
R1757 VSS.t755 VSS.t1068 109.579
R1758 VSS.n1581 VSS.t1086 109.579
R1759 VSS.t1103 VSS.t724 109.579
R1760 VSS.t545 VSS.t163 109.579
R1761 VSS.t554 VSS.t936 109.579
R1762 VSS.n1365 VSS.t573 108.505
R1763 VSS.n1977 VSS.t518 108.505
R1764 VSS.n1270 VSS.t1014 108.505
R1765 VSS VSS.t380 106.942
R1766 VSS.t463 VSS.t999 102.992
R1767 VSS.t461 VSS.t1006 102.992
R1768 VSS.n2178 VSS.t1140 102.353
R1769 VSS.n1200 VSS.t1226 102.353
R1770 VSS.n2685 VSS.t1199 102.353
R1771 VSS.n2822 VSS.t129 101.43
R1772 VSS.n1248 VSS.t736 101.43
R1773 VSS.n1262 VSS.t645 101.43
R1774 VSS.t230 VSS.t895 101.15
R1775 VSS.t14 VSS.t1076 101.15
R1776 VSS.n2850 VSS.t1182 99.7825
R1777 VSS.n964 VSS.t1204 99.7825
R1778 VSS.t772 VSS.t311 98.8769
R1779 VSS.t284 VSS.t745 98.8769
R1780 VSS.t521 VSS.t523 98.8769
R1781 VSS.t732 VSS.t10 98.8769
R1782 VSS.t401 VSS.t915 98.8769
R1783 VSS.t543 VSS.t145 98.8769
R1784 VSS.t299 VSS.t135 98.8769
R1785 VSS.t851 VSS.t124 98.8769
R1786 VSS.t646 VSS.t930 98.8769
R1787 VSS.t925 VSS.t160 98.8769
R1788 VSS.t637 VSS.t592 92.7208
R1789 VSS.t1078 VSS 92.7208
R1790 VSS.t602 VSS.t1090 92.7208
R1791 VSS.t533 VSS.t542 92.7208
R1792 VSS.t1107 VSS.t91 92.7208
R1793 VSS VSS.t555 92.7208
R1794 VSS.n476 VSS.n475 89.224
R1795 VSS.n465 VSS.n464 89.224
R1796 VSS.n463 VSS.n432 89.224
R1797 VSS.n436 VSS.n433 89.224
R1798 VSS.n442 VSS.n441 89.224
R1799 VSS.n456 VSS.n444 89.224
R1800 VSS.t181 VSS 88.8318
R1801 VSS.t407 VSS 88.8318
R1802 VSS.n455 VSS.n447 88.4711
R1803 VSS.t352 VSS.n187 85.9264
R1804 VSS.t863 VSS.n93 85.9264
R1805 VSS.n483 VSS.n408 84.7064
R1806 VSS.t967 VSS.t291 84.2917
R1807 VSS.t133 VSS.t907 84.2917
R1808 VSS.t115 VSS.t366 84.2917
R1809 VSS.t997 VSS.t96 84.2917
R1810 VSS VSS.t788 84.2702
R1811 VSS.n3282 VSS 83.8426
R1812 VSS.n484 VSS.n407 80.1887
R1813 VSS.n486 VSS.n406 80.1887
R1814 VSS.n487 VSS.n405 80.1887
R1815 VSS.n417 VSS.n404 80.1887
R1816 VSS.n2394 VSS 76.6073
R1817 VSS.t848 VSS.t1113 75.8626
R1818 VSS VSS.n2394 75.2814
R1819 VSS.n655 VSS.t103 74.8666
R1820 VSS.n656 VSS.t147 74.8666
R1821 VSS.n1467 VSS.t361 74.8666
R1822 VSS.n1558 VSS.t756 74.8666
R1823 VSS.n1605 VSS.t310 74.8666
R1824 VSS.n854 VSS.t914 74.8666
R1825 VSS.n859 VSS.t496 74.8666
R1826 VSS.n1240 VSS.t506 74.8666
R1827 VSS.n1864 VSS.t368 74.8666
R1828 VSS.n939 VSS.t847 74.8666
R1829 VSS.n24 VSS.t144 72.8576
R1830 VSS.n44 VSS.t460 72.8576
R1831 VSS.n3106 VSS.t548 72.8576
R1832 VSS.n214 VSS.t1005 72.8576
R1833 VSS.n3309 VSS.t1007 72.8576
R1834 VSS.n3343 VSS.t729 72.8576
R1835 VSS.n1937 VSS.t571 72.8576
R1836 VSS.n1938 VSS.t304 72.8576
R1837 VSS.n1919 VSS.t890 72.8576
R1838 VSS.t643 VSS.n426 72.7469
R1839 VSS.n460 VSS.t467 72.7469
R1840 VSS.t126 VSS.t1052 71.7175
R1841 VSS.t745 VSS 70.787
R1842 VSS.t959 VSS.t796 67.6928
R1843 VSS.t749 VSS.t1002 67.4335
R1844 VSS.t328 VSS.t952 67.4335
R1845 VSS.t320 VSS.t893 67.4335
R1846 VSS.n422 VSS.t371 66.396
R1847 VSS.t457 VSS.n420 66.396
R1848 VSS.n482 VSS.n409 64.8307
R1849 VSS.n3077 VSS.t298 61.6916
R1850 VSS VSS.t445 61.1229
R1851 VSS VSS.n2986 61.1229
R1852 VSS.n1002 VSS.n63 59.6152
R1853 VSS.n1011 VSS.n63 59.6152
R1854 VSS.t558 VSS.t468 59.0043
R1855 VSS.n451 VSS.n450 58.7133
R1856 VSS.n15 VSS.t752 58.5719
R1857 VSS.n21 VSS.t1059 58.5719
R1858 VSS.n3100 VSS.t842 58.5719
R1859 VSS.n218 VSS.t169 58.5719
R1860 VSS.n3328 VSS.t114 58.5719
R1861 VSS.n107 VSS.t142 58.5719
R1862 VSS.n1416 VSS.t365 58.5719
R1863 VSS.n1307 VSS.t941 58.5719
R1864 VSS.n3404 VSS.t123 57.2177
R1865 VSS.t999 VSS.t461 57.2177
R1866 VSS.n3394 VSS.n71 57.2177
R1867 VSS VSS.n492 56.2331
R1868 VSS.n391 VSS.n389 54.2123
R1869 VSS.n3247 VSS.n3239 54.2123
R1870 VSS.n3261 VSS.n3260 54.2123
R1871 VSS.n3222 VSS.n180 54.2123
R1872 VSS.n3217 VSS.n3216 54.2123
R1873 VSS.n183 VSS.n182 54.2123
R1874 VSS.n3386 VSS.n77 54.2123
R1875 VSS.n3277 VSS.n3255 54.2123
R1876 VSS.n1004 VSS.n1001 53.1823
R1877 VSS.n1001 VSS.t757 53.1823
R1878 VSS.n2390 VSS.n1003 53.1823
R1879 VSS.n1003 VSS.n1002 53.1823
R1880 VSS.n1014 VSS.n1013 53.1823
R1881 VSS.n1013 VSS.n1012 53.1823
R1882 VSS.n1010 VSS.n1009 53.1823
R1883 VSS.n1011 VSS.n1010 53.1823
R1884 VSS.n681 VSS.t567 52.8576
R1885 VSS.n454 VSS.n448 51.7522
R1886 VSS.t1060 VSS.t293 50.5752
R1887 VSS.t1056 VSS.t358 50.5752
R1888 VSS.t137 VSS.t635 50.5752
R1889 VSS VSS.t1078 50.5752
R1890 VSS.t1010 VSS.t715 50.5752
R1891 VSS.t388 VSS.t885 50.5752
R1892 VSS.t106 VSS.t680 50.5752
R1893 VSS.t932 VSS.t139 50.5752
R1894 VSS.n1002 VSS.t560 50.3004
R1895 VSS.t582 VSS.n1011 49.0584
R1896 VSS.n1012 VSS.t582 49.0584
R1897 VSS.n2389 VSS.n1000 48.7505
R1898 VSS.n2393 VSS.n1000 48.7505
R1899 VSS.n2392 VSS.n2391 48.7505
R1900 VSS.n2393 VSS.n2392 48.7505
R1901 VSS.n1603 VSS.t658 48.5719
R1902 VSS.t380 VSS.n3281 47.9103
R1903 VSS.n1611 VSS.t577 47.1434
R1904 VSS.n942 VSS.t1114 47.1434
R1905 VSS.t699 VSS 44.7453
R1906 VSS.n50 VSS 43.9579
R1907 VSS.n3140 VSS 43.9579
R1908 VSS.n3308 VSS 43.9579
R1909 VSS.n475 VSS.n474 42.1089
R1910 VSS.n488 VSS.n404 42.1089
R1911 VSS.n488 VSS.n487 42.1089
R1912 VSS.n486 VSS.n485 42.1089
R1913 VSS.n485 VSS.n484 42.1089
R1914 VSS.n483 VSS.n482 42.1089
R1915 VSS.n3403 VSS.t376 41.9598
R1916 VSS.n655 VSS.t335 40.0005
R1917 VSS.n656 VSS.t979 40.0005
R1918 VSS.n681 VSS.t981 40.0005
R1919 VSS.n1400 VSS.t638 40.0005
R1920 VSS.n1400 VSS.t640 40.0005
R1921 VSS.n784 VSS.t1035 40.0005
R1922 VSS.n784 VSS.t1027 40.0005
R1923 VSS.n783 VSS.t1029 40.0005
R1924 VSS.n783 VSS.t1033 40.0005
R1925 VSS.n792 VSS.t1031 40.0005
R1926 VSS.n792 VSS.t1021 40.0005
R1927 VSS.n1422 VSS.t664 40.0005
R1928 VSS.n1422 VSS.t727 40.0005
R1929 VSS.n771 VSS.t666 40.0005
R1930 VSS.n771 VSS.t1037 40.0005
R1931 VSS.n773 VSS.t1043 40.0005
R1932 VSS.n773 VSS.t1047 40.0005
R1933 VSS.n776 VSS.t1051 40.0005
R1934 VSS.n776 VSS.t1041 40.0005
R1935 VSS.n779 VSS.t1045 40.0005
R1936 VSS.n779 VSS.t1049 40.0005
R1937 VSS.n2625 VSS.t1039 40.0005
R1938 VSS.n1396 VSS.t626 40.0005
R1939 VSS.n1397 VSS.t634 40.0005
R1940 VSS.n1397 VSS.t612 40.0005
R1941 VSS.n1412 VSS.t636 40.0005
R1942 VSS.n1412 VSS.t614 40.0005
R1943 VSS.n1467 VSS.t406 40.0005
R1944 VSS.n1468 VSS.t632 40.0005
R1945 VSS.n1468 VSS.t622 40.0005
R1946 VSS.n1475 VSS.t624 40.0005
R1947 VSS.n1475 VSS.t628 40.0005
R1948 VSS.n1391 VSS.t642 40.0005
R1949 VSS.n1391 VSS.t620 40.0005
R1950 VSS.n1387 VSS.t597 40.0005
R1951 VSS.n1387 VSS.t616 40.0005
R1952 VSS.n1372 VSS.t475 40.0005
R1953 VSS.n1372 VSS.t599 40.0005
R1954 VSS.n1559 VSS.t1063 40.0005
R1955 VSS.n1559 VSS.t1065 40.0005
R1956 VSS.n1558 VSS.t731 40.0005
R1957 VSS.n1571 VSS.t1081 40.0005
R1958 VSS.n1571 VSS.t1073 40.0005
R1959 VSS.n1573 VSS.t1077 40.0005
R1960 VSS.n1573 VSS.t1067 40.0005
R1961 VSS.n1574 VSS.t1075 40.0005
R1962 VSS.n1670 VSS.t1079 40.0005
R1963 VSS.n1670 VSS.t1085 40.0005
R1964 VSS.n1580 VSS.t1083 40.0005
R1965 VSS.n1580 VSS.t1093 40.0005
R1966 VSS.n1582 VSS.t1087 40.0005
R1967 VSS.n1582 VSS.t1089 40.0005
R1968 VSS.n1586 VSS.t1091 40.0005
R1969 VSS.n1586 VSS.t725 40.0005
R1970 VSS.n1597 VSS.t1118 40.0005
R1971 VSS.n1597 VSS.t723 40.0005
R1972 VSS.n1605 VSS.t978 40.0005
R1973 VSS.n854 VSS.t1019 40.0005
R1974 VSS.n859 VSS.t870 40.0005
R1975 VSS.n1240 VSS.t589 40.0005
R1976 VSS.n1864 VSS.t370 40.0005
R1977 VSS.n939 VSS.t849 40.0005
R1978 VSS.n484 VSS.n483 39.4771
R1979 VSS.n1365 VSS.t479 38.7697
R1980 VSS.n838 VSS.t363 38.7697
R1981 VSS.n1977 VSS.t404 38.7697
R1982 VSS.n1284 VSS.t98 38.7697
R1983 VSS.n1270 VSS.t587 38.7697
R1984 VSS.n597 VSS.t112 38.5719
R1985 VSS.n597 VSS.t331 38.5719
R1986 VSS.n598 VSS.t761 38.5719
R1987 VSS.n598 VSS.t307 38.5719
R1988 VSS.n2625 VSS.t1023 38.5719
R1989 VSS.n1396 VSS.t630 38.5719
R1990 VSS.n1388 VSS.t483 38.5719
R1991 VSS.n1388 VSS.t965 38.5719
R1992 VSS.n1574 VSS.t1071 38.5719
R1993 VSS.n1577 VSS.t654 38.5719
R1994 VSS.n1577 VSS.t487 38.5719
R1995 VSS.n1608 VSS.t520 38.5719
R1996 VSS.n1608 VSS.t579 38.5719
R1997 VSS.n1610 VSS.t165 38.5719
R1998 VSS.n1610 VSS.t485 38.5719
R1999 VSS.n860 VSS.t325 38.5719
R2000 VSS.n860 VSS.t610 38.5719
R2001 VSS.n878 VSS.t949 38.5719
R2002 VSS.n878 VSS.t763 38.5719
R2003 VSS.n1244 VSS.t314 38.5719
R2004 VSS.n1244 VSS.t670 38.5719
R2005 VSS.n1271 VSS.t321 38.5719
R2006 VSS.n1271 VSS.t489 38.5719
R2007 VSS.n946 VSS.t557 38.5719
R2008 VSS.n946 VSS.t110 38.5719
R2009 VSS.n3407 VSS.t342 38.3944
R2010 VSS VSS.t990 36.085
R2011 VSS VSS.t833 36.085
R2012 VSS.n1611 VSS.t983 35.4291
R2013 VSS.n942 VSS.t469 35.4291
R2014 VSS.n487 VSS.n486 35.2902
R2015 VSS.n464 VSS.n431 34.659
R2016 VSS.n463 VSS.n462 34.659
R2017 VSS.n462 VSS.n433 34.659
R2018 VSS.n457 VSS.n441 34.659
R2019 VSS.n457 VSS.n456 34.659
R2020 VSS.n455 VSS.n454 34.659
R2021 VSS.n1478 VSS.n1477 34.6358
R2022 VSS.n50 VSS.n49 34.6358
R2023 VSS.n47 VSS.n2 34.6358
R2024 VSS.n3161 VSS.n3145 34.6358
R2025 VSS.n3161 VSS.n3160 34.6358
R2026 VSS.n3155 VSS.n3154 34.6358
R2027 VSS.n3189 VSS.n188 34.6358
R2028 VSS.n3189 VSS.n189 34.6358
R2029 VSS.n3183 VSS.n3182 34.6358
R2030 VSS.n3177 VSS.n3176 34.6358
R2031 VSS.n3176 VSS.n195 34.6358
R2032 VSS.n3170 VSS.n195 34.6358
R2033 VSS.n3140 VSS.n3139 34.6358
R2034 VSS.n3137 VSS.n215 34.6358
R2035 VSS.n3085 VSS.n215 34.6358
R2036 VSS.n3087 VSS.n3085 34.6358
R2037 VSS.n3090 VSS.n220 34.6358
R2038 VSS.n3094 VSS.n220 34.6358
R2039 VSS.n3114 VSS.n3103 34.6358
R2040 VSS.n3110 VSS.n3103 34.6358
R2041 VSS.n3311 VSS.n3308 34.6358
R2042 VSS.n3315 VSS.n3299 34.6358
R2043 VSS.n636 VSS.n629 34.6358
R2044 VSS.n654 VSS.n602 34.6358
R2045 VSS.n650 VSS.n602 34.6358
R2046 VSS.n650 VSS.n649 34.6358
R2047 VSS.n662 VSS.n600 34.6358
R2048 VSS.n658 VSS.n600 34.6358
R2049 VSS.n1459 VSS.n1401 34.6358
R2050 VSS.n1474 VSS.n1394 34.6358
R2051 VSS.n1482 VSS.n1389 34.6358
R2052 VSS.n1658 VSS.n1657 34.6358
R2053 VSS.n1654 VSS.n1587 34.6358
R2054 VSS.n1641 VSS.n1601 34.6358
R2055 VSS.n1636 VSS.n1635 34.6358
R2056 VSS.n1635 VSS.n1606 34.6358
R2057 VSS.n2602 VSS.n835 34.6358
R2058 VSS.n920 VSS.n919 34.6358
R2059 VSS.n915 VSS.n857 34.6358
R2060 VSS.n903 VSS.n863 34.6358
R2061 VSS.n1936 VSS.n1935 34.6358
R2062 VSS.n1935 VSS.n1267 34.6358
R2063 VSS.n1940 VSS.n1265 34.6358
R2064 VSS.n1913 VSS.n1896 34.6358
R2065 VSS.n1904 VSS.n1896 34.6358
R2066 VSS.n1905 VSS.n1904 34.6358
R2067 VSS.n1888 VSS.n1887 34.6358
R2068 VSS.n1915 VSS.n1268 34.6358
R2069 VSS.n2555 VSS.n2554 34.6358
R2070 VSS.n2554 VSS.n2553 34.6358
R2071 VSS.n2549 VSS.n2548 34.6358
R2072 VSS.n1822 VSS.n1760 34.6358
R2073 VSS.n1804 VSS.n1768 34.6358
R2074 VSS.n2007 VSS.n2006 34.6358
R2075 VSS.n2518 VSS.n991 34.6358
R2076 VSS.n2468 VSS.n2467 34.6358
R2077 VSS.n2449 VSS.n2448 34.6358
R2078 VSS.n2448 VSS.n2432 34.6358
R2079 VSS.n1042 VSS.n493 34.6358
R2080 VSS.n2057 VSS.t1236 34.2973
R2081 VSS.n1555 VSS.t1194 34.2973
R2082 VSS.n2477 VSS.t1174 34.2973
R2083 VSS.n263 VSS.t1217 34.2973
R2084 VSS.n2325 VSS.t1153 34.2973
R2085 VSS.n3157 VSS.n3156 33.8829
R2086 VSS.n3151 VSS.n3150 33.8829
R2087 VSS.n3185 VSS.n3184 33.8829
R2088 VSS.n3179 VSS.n3178 33.8829
R2089 VSS.n3130 VSS.n3129 33.8829
R2090 VSS.n3123 VSS.n3122 33.8829
R2091 VSS.n3116 VSS.n3115 33.8829
R2092 VSS.n1673 VSS.n1672 33.8829
R2093 VSS.n905 VSS.n861 33.8829
R2094 VSS.t590 VSS.t613 33.717
R2095 VSS.t722 VSS.t600 33.717
R2096 VSS.t119 VSS.t519 33.717
R2097 VSS.t516 VSS 33.717
R2098 VSS.t12 VSS.t891 33.717
R2099 VSS.t651 VSS.t586 33.717
R2100 VSS.n1310 VSS.t878 33.462
R2101 VSS.n1310 VSS.t928 33.462
R2102 VSS.n1374 VSS.t95 33.462
R2103 VSS.n1374 VSS.t553 33.462
R2104 VSS.n1758 VSS.t773 33.462
R2105 VSS.n1758 VSS.t312 33.462
R2106 VSS.n1762 VSS.t285 33.462
R2107 VSS.n1762 VSS.t746 33.462
R2108 VSS.n1767 VSS.t522 33.462
R2109 VSS.n1767 VSS.t524 33.462
R2110 VSS.n1783 VSS.t733 33.462
R2111 VSS.n1783 VSS.t11 33.462
R2112 VSS.n1991 VSS.t402 33.462
R2113 VSS.n1991 VSS.t916 33.462
R2114 VSS.n990 VSS.t544 33.462
R2115 VSS.n990 VSS.t146 33.462
R2116 VSS.n998 VSS.t300 33.462
R2117 VSS.n998 VSS.t136 33.462
R2118 VSS.n2412 VSS.t852 33.462
R2119 VSS.n2412 VSS.t125 33.462
R2120 VSS.n2420 VSS.t647 33.462
R2121 VSS.n2420 VSS.t931 33.462
R2122 VSS.n2434 VSS.t926 33.462
R2123 VSS.n2434 VSS.t161 33.462
R2124 VSS.n1030 VSS.t1053 33.462
R2125 VSS.n1030 VSS.t127 33.462
R2126 VSS.n3157 VSS.n3146 33.1299
R2127 VSS.n3151 VSS.n3148 33.1299
R2128 VSS.n3185 VSS.n191 33.1299
R2129 VSS.n3179 VSS.n192 33.1299
R2130 VSS.n3095 VSS.n3094 33.1299
R2131 VSS.n3130 VSS.n3097 33.1299
R2132 VSS.n3124 VSS.n3123 33.1299
R2133 VSS.n3121 VSS.n3101 33.1299
R2134 VSS.n3117 VSS.n3116 33.1299
R2135 VSS.n492 VSS.n491 32.9096
R2136 VSS.n2383 VSS.t561 32.8043
R2137 VSS.n1018 VSS.t758 32.8043
R2138 VSS VSS.t772 32.5848
R2139 VSS VSS.t521 32.5848
R2140 VSS VSS.t732 32.5848
R2141 VSS VSS.t401 32.5848
R2142 VSS VSS.t543 32.5848
R2143 VSS VSS.t299 32.5848
R2144 VSS VSS.t851 32.5848
R2145 VSS VSS.t646 32.5848
R2146 VSS VSS.t925 32.5848
R2147 VSS.n1603 VSS.t581 32.5719
R2148 VSS.n454 VSS.n453 32.5005
R2149 VSS.n453 VSS.n438 32.5005
R2150 VSS.n451 VSS.n426 32.5005
R2151 VSS.n445 VSS.n411 32.5005
R2152 VSS.n424 VSS.n411 32.5005
R2153 VSS.n482 VSS.n481 32.5005
R2154 VSS.n481 VSS.n401 32.5005
R2155 VSS.n458 VSS.n457 32.5005
R2156 VSS.n460 VSS.n458 32.5005
R2157 VSS.n443 VSS.n427 32.5005
R2158 VSS.n468 VSS.n427 32.5005
R2159 VSS.n416 VSS.n415 32.5005
R2160 VSS.n420 VSS.n416 32.5005
R2161 VSS.n485 VSS.n400 32.5005
R2162 VSS.n490 VSS.n400 32.5005
R2163 VSS.n462 VSS.n461 32.5005
R2164 VSS.n461 VSS.n460 32.5005
R2165 VSS.n435 VSS.n425 32.5005
R2166 VSS.n468 VSS.n425 32.5005
R2167 VSS.n419 VSS.n418 32.5005
R2168 VSS.n420 VSS.n419 32.5005
R2169 VSS.n489 VSS.n488 32.5005
R2170 VSS.n490 VSS.n489 32.5005
R2171 VSS.n459 VSS.n431 32.5005
R2172 VSS.n460 VSS.n459 32.5005
R2173 VSS.n467 VSS.n466 32.5005
R2174 VSS.n468 VSS.n467 32.5005
R2175 VSS.n477 VSS.n470 32.5005
R2176 VSS.n470 VSS.n469 32.5005
R2177 VSS.n474 VSS.n423 32.5005
R2178 VSS.n423 VSS.n422 32.5005
R2179 VSS.n441 VSS.n433 32.4928
R2180 VSS.n3125 VSS.n3098 32.377
R2181 VSS.n628 VSS.n604 32.377
R2182 VSS.n1854 VSS.n1853 32.377
R2183 VSS.n1891 VSS.n1268 32.377
R2184 VSS.n2560 VSS.n934 32.377
R2185 VSS.n1678 VSS.n1677 32.377
R2186 VSS.n1889 VSS.n1888 31.624
R2187 VSS.n648 VSS.n604 31.2476
R2188 VSS.n2588 VSS.n2587 31.2476
R2189 VSS.n1854 VSS.n1286 31.2476
R2190 VSS.n2560 VSS.n2559 31.2476
R2191 VSS.n456 VSS.n455 30.9174
R2192 VSS.n478 VSS.n473 30.8711
R2193 VSS.n392 VSS.n391 30.8711
R2194 VSS.n3247 VSS.n3246 30.8711
R2195 VSS.n3270 VSS.n3261 30.8711
R2196 VSS.n3224 VSS.n180 30.8711
R2197 VSS.n3216 VSS.n3202 30.8711
R2198 VSS.n3198 VSS.n183 30.8711
R2199 VSS.n3387 VSS.n3386 30.8711
R2200 VSS.n3277 VSS.n3276 30.8711
R2201 VSS.n658 VSS.n657 30.8711
R2202 VSS.n1637 VSS.n1636 30.8711
R2203 VSS.n1979 VSS.n1241 30.8711
R2204 VSS.n1867 VSS.n1865 30.8711
R2205 VSS.n475 VSS.n404 30.7444
R2206 VSS.n1570 VSS.n1560 30.4946
R2207 VSS.n1624 VSS.n835 30.4946
R2208 VSS.n1867 VSS.n1866 30.4946
R2209 VSS.n2377 VSS.t583 30.3424
R2210 VSS.n1461 VSS.n1460 30.1181
R2211 VSS.n1681 VSS.n1680 30.1181
R2212 VSS.n1600 VSS.n1599 30.1181
R2213 VSS.n1914 VSS.n1913 30.1181
R2214 VSS.n3402 VSS.n3401 29.8168
R2215 VSS.t392 VSS.t472 29.8079
R2216 VSS.t472 VSS.t562 29.8079
R2217 VSS.t394 VSS.t759 29.8079
R2218 VSS.t390 VSS.t394 29.8079
R2219 VSS.t560 VSS.t390 29.8079
R2220 VSS.n1465 VSS.n1398 29.7417
R2221 VSS.n2593 VSS.n2592 29.3652
R2222 VSS.n1449 VSS.n1448 28.9887
R2223 VSS.n464 VSS.n463 28.259
R2224 VSS.n1485 VSS.n1484 27.8593
R2225 VSS.n1655 VSS.n1654 27.8593
R2226 VSS.n663 VSS.n662 27.4829
R2227 VSS.n1631 VSS.n1606 27.4829
R2228 VSS.n2599 VSS.n2598 27.4829
R2229 VSS.n917 VSS.n916 27.4829
R2230 VSS.n911 VSS.n857 27.4829
R2231 VSS.n1978 VSS.n1976 27.4829
R2232 VSS.n1976 VSS.n1242 27.4829
R2233 VSS.n1859 VSS.n1285 27.4829
R2234 VSS.n1882 VSS.n1273 27.4829
R2235 VSS.n1485 VSS.n1373 27.1064
R2236 VSS.n3446 VSS.n3445 26.9246
R2237 VSS.n3359 VSS.n95 26.9246
R2238 VSS.n1625 VSS.n1612 26.7299
R2239 VSS.n2337 VSS.n2336 26.6009
R2240 VSS.n1944 VSS.n1265 26.314
R2241 VSS.n2383 VSS.n2382 26.1653
R2242 VSS.n2385 VSS.n2384 26.1653
R2243 VSS.n1018 VSS.n1017 26.1653
R2244 VSS.n469 VSS.n468 25.9813
R2245 VSS.n2822 VSS.t180 25.9346
R2246 VSS.n1248 VSS.t721 25.9346
R2247 VSS.n1262 VSS.t118 25.9346
R2248 VSS.n3235 VSS.t199 25.8199
R2249 VSS.n1662 VSS.n1661 25.7355
R2250 VSS.n1924 VSS.n1922 25.7355
R2251 VSS.n2548 VSS.n2547 25.7355
R2252 VSS.n1824 VSS.n1757 25.7355
R2253 VSS.n2443 VSS.n2442 25.7355
R2254 VSS.n3464 VSS.n2 25.6926
R2255 VSS.n3316 VSS.n3315 25.6926
R2256 VSS.n1817 VSS.n1816 25.6926
R2257 VSS.n1809 VSS.n1765 25.6926
R2258 VSS.n1779 VSS.n1768 25.6926
R2259 VSS.n2006 VSS.n1993 25.6926
R2260 VSS.n2510 VSS.n991 25.6926
R2261 VSS.n2504 VSS.n2503 25.6926
R2262 VSS.n2467 VSS.n2414 25.6926
R2263 VSS.n1043 VSS.n1042 25.6926
R2264 VSS.n637 VSS.n636 25.6005
R2265 VSS.n1677 VSS.n1575 25.6005
R2266 VSS.n15 VSS.t294 25.4291
R2267 VSS.n21 VSS.t359 25.4291
R2268 VSS.n3100 VSS.t933 25.4291
R2269 VSS.n218 VSS.t107 25.4291
R2270 VSS.n3328 VSS.t1011 25.4291
R2271 VSS.n107 VSS.t389 25.4291
R2272 VSS.n1416 VSS.t93 25.4291
R2273 VSS.n1307 VSS.t492 25.4291
R2274 VSS.t130 VSS.t264 25.2879
R2275 VSS.t621 VSS.t405 25.2879
R2276 VSS.t559 VSS.t490 25.2879
R2277 VSS.n3429 VSS.n3428 25.224
R2278 VSS.n3428 VSS.n60 25.224
R2279 VSS.n3424 VSS.n3423 25.224
R2280 VSS.n3423 VSS.n3422 25.224
R2281 VSS.n3420 VSS.n3419 25.224
R2282 VSS.n3419 VSS.n3411 25.224
R2283 VSS.n3415 VSS.n3414 25.224
R2284 VSS.n3414 VSS.n39 25.224
R2285 VSS.n3455 VSS.n3454 25.224
R2286 VSS.n3454 VSS.n3453 25.224
R2287 VSS.n3451 VSS.n22 25.224
R2288 VSS.n3376 VSS.n3375 25.224
R2289 VSS.n3375 VSS.n83 25.224
R2290 VSS.n3371 VSS.n3370 25.224
R2291 VSS.n3370 VSS.n3369 25.224
R2292 VSS.n3367 VSS.n3366 25.224
R2293 VSS.n3366 VSS.n89 25.224
R2294 VSS.n3362 VSS.n3361 25.224
R2295 VSS.n3361 VSS.n3360 25.224
R2296 VSS.n3335 VSS.n3334 25.224
R2297 VSS.n3336 VSS.n3335 25.224
R2298 VSS.n3353 VSS.n3340 25.224
R2299 VSS.n127 VSS.n125 25.224
R2300 VSS.n131 VSS.n125 25.224
R2301 VSS.n132 VSS.n124 25.224
R2302 VSS.n136 VSS.n124 25.224
R2303 VSS.n137 VSS.n123 25.224
R2304 VSS.n141 VSS.n123 25.224
R2305 VSS.n142 VSS.n122 25.224
R2306 VSS.n146 VSS.n122 25.224
R2307 VSS.n147 VSS.n121 25.224
R2308 VSS.n151 VSS.n121 25.224
R2309 VSS.n152 VSS.n120 25.224
R2310 VSS.n156 VSS.n120 25.224
R2311 VSS.n157 VSS.n119 25.224
R2312 VSS.n161 VSS.n119 25.224
R2313 VSS.n162 VSS.n118 25.224
R2314 VSS.n166 VSS.n118 25.224
R2315 VSS.n167 VSS.n117 25.224
R2316 VSS.n171 VSS.n117 25.224
R2317 VSS.n1572 VSS.n1570 25.224
R2318 VSS.n1681 VSS.n1572 25.224
R2319 VSS.n2473 VSS.n2472 24.9894
R2320 VSS.n2332 VSS.n2331 24.9894
R2321 VSS.n3144 VSS.n3143 24.9767
R2322 VSS.n3169 VSS.n3168 24.9767
R2323 VSS.n3108 VSS.n3105 24.9767
R2324 VSS.n2881 VSS.n585 24.968
R2325 VSS.n3400 VSS.t464 24.9236
R2326 VSS.n3400 VSS.t462 24.9236
R2327 VSS.n535 VSS.t921 24.9236
R2328 VSS.n535 VSS.t924 24.9236
R2329 VSS.n627 VSS.t970 24.9236
R2330 VSS.n627 VSS.t971 24.9236
R2331 VSS.n626 VSS.t882 24.9236
R2332 VSS.n626 VSS.t5 24.9236
R2333 VSS.n1413 VSS.t138 24.9236
R2334 VSS.n1413 VSS.t591 24.9236
R2335 VSS.n1551 VSS.t769 24.9236
R2336 VSS.n1551 VSS.t541 24.9236
R2337 VSS.n1585 VSS.t603 24.9236
R2338 VSS.n1585 VSS.t1104 24.9236
R2339 VSS.n836 VSS.t1108 24.9236
R2340 VSS.n836 VSS.t738 24.9236
R2341 VSS.n838 VSS.t570 24.9236
R2342 VSS.n844 VSS.t1003 24.9236
R2343 VSS.n844 VSS.t953 24.9236
R2344 VSS.n843 VSS.t750 24.9236
R2345 VSS.n843 VSS.t329 24.9236
R2346 VSS.n853 VSS.t387 24.9236
R2347 VSS.n853 VSS.t122 24.9236
R2348 VSS.n1850 VSS.t742 24.9236
R2349 VSS.n1850 VSS.t744 24.9236
R2350 VSS.n1288 VSS.t1112 24.9236
R2351 VSS.n1288 VSS.t550 24.9236
R2352 VSS.n1284 VSS.t1017 24.9236
R2353 VSS.n1890 VSS.t539 24.9236
R2354 VSS.n1890 VSS.t652 24.9236
R2355 VSS.n933 VSS.t375 24.9236
R2356 VSS.n933 VSS.t494 24.9236
R2357 VSS.n936 VSS.t302 24.9236
R2358 VSS.n936 VSS.t937 24.9236
R2359 VSS VSS.t463 24.7946
R2360 VSS.n1695 VSS.n1694 24.4711
R2361 VSS.n910 VSS.n909 24.4711
R2362 VSS.n2602 VSS.n2601 24.4711
R2363 VSS.n905 VSS.n904 24.4711
R2364 VSS.n904 VSS.n903 24.4711
R2365 VSS.n2555 VSS.n937 24.4711
R2366 VSS.t990 VSS.t987 24.2493
R2367 VSS.t833 VSS.t836 24.2493
R2368 VSS.t342 VSS.t345 24.2493
R2369 VSS.n3459 VSS.n16 24.0946
R2370 VSS.n3330 VSS.n110 24.0946
R2371 VSS.n281 VSS.t239 23.7273
R2372 VSS.n2594 VSS.n841 23.7181
R2373 VSS.n1328 VSS.n1314 23.7181
R2374 VSS.n1339 VSS.n1314 23.7181
R2375 VSS.n1433 VSS.n1420 23.7181
R2376 VSS.n1433 VSS.n1432 23.7181
R2377 VSS.n1642 VSS.n1641 23.7181
R2378 VSS.n2598 VSS.n841 23.7181
R2379 VSS.n2586 VSS.n848 23.7181
R2380 VSS.n920 VSS.n848 23.7181
R2381 VSS.n1931 VSS.n1267 23.7181
R2382 VSS.n1859 VSS.n1858 23.7181
R2383 VSS.n1789 VSS.n1788 23.7181
R2384 VSS.n2029 VSS.n1223 23.7181
R2385 VSS.n2012 VSS.n2011 23.7181
R2386 VSS.n1999 VSS.n989 23.7181
R2387 VSS.n2499 VSS.n2498 23.7181
R2388 VSS.n2460 VSS.n2459 23.7181
R2389 VSS.n2985 VSS.n493 23.7181
R2390 VSS.t1052 VSS 23.6345
R2391 VSS.n876 VSS.n875 23.4338
R2392 VSS.n1392 VSS.n1389 23.3417
R2393 VSS.n1658 VSS.n1583 23.3417
R2394 VSS.n450 VSS.n448 23.2076
R2395 VSS.n3176 VSS.n3175 23.1729
R2396 VSS.n664 VSS.n599 22.9652
R2397 VSS.n664 VSS.n663 22.9652
R2398 VSS.n1631 VSS.n1630 22.9652
R2399 VSS.n1630 VSS.n1629 22.9652
R2400 VSS.n2588 VSS.n845 22.9652
R2401 VSS.n911 VSS.n910 22.9652
R2402 VSS.n1972 VSS.n1242 22.9652
R2403 VSS.n1972 VSS.n1971 22.9652
R2404 VSS.n1852 VSS.n1851 22.9652
R2405 VSS.n1883 VSS.n1882 22.9652
R2406 VSS.n1883 VSS.n1272 22.9652
R2407 VSS.n943 VSS.n940 22.9652
R2408 VSS.n3282 VSS.n3235 22.9387
R2409 VSS.n3393 VSS.t527 22.8805
R2410 VSS.n1642 VSS.n1600 22.5887
R2411 VSS.n24 VSS.t508 22.3257
R2412 VSS.n44 VSS.t526 22.3257
R2413 VSS.n3106 VSS.t510 22.3257
R2414 VSS.n214 VSS.t7 22.3257
R2415 VSS.n3309 VSS.t377 22.3257
R2416 VSS.n3343 VSS.t477 22.3257
R2417 VSS.n1937 VSS.t1094 22.3257
R2418 VSS.n1938 VSS.t829 22.3257
R2419 VSS.n1919 VSS.t976 22.3257
R2420 VSS.n649 VSS.n648 22.2123
R2421 VSS.n2587 VSS.n2586 22.2123
R2422 VSS.n916 VSS.n915 22.2123
R2423 VSS.n2559 VSS.n2558 22.2123
R2424 VSS.n1824 VSS.n1823 22.2123
R2425 VSS.n1823 VSS.n1822 22.2123
R2426 VSS.n1818 VSS.n1760 22.2123
R2427 VSS.n1818 VSS.n1817 22.2123
R2428 VSS.n1805 VSS.n1765 22.2123
R2429 VSS.n1805 VSS.n1804 22.2123
R2430 VSS.n1788 VSS.n1784 22.2123
R2431 VSS.n1784 VSS.n1223 22.2123
R2432 VSS.n2011 VSS.n1992 22.2123
R2433 VSS.n2007 VSS.n1992 22.2123
R2434 VSS.n2519 VSS.n989 22.2123
R2435 VSS.n2519 VSS.n2518 22.2123
R2436 VSS.n2503 VSS.n999 22.2123
R2437 VSS.n2499 VSS.n999 22.2123
R2438 VSS.n2472 VSS.n2413 22.2123
R2439 VSS.n2468 VSS.n2413 22.2123
R2440 VSS.n2459 VSS.n2421 22.2123
R2441 VSS.n2449 VSS.n2421 22.2123
R2442 VSS.n2444 VSS.n2432 22.2123
R2443 VSS.n2444 VSS.n2443 22.2123
R2444 VSS.n2336 VSS.n1031 22.2123
R2445 VSS.n2332 VSS.n1031 22.2123
R2446 VSS.n446 VSS.n412 21.6752
R2447 VSS.n3408 VSS 21.6512
R2448 VSS.n3460 VSS.n3459 21.4593
R2449 VSS.n3452 VSS.n3451 21.4593
R2450 VSS.n3330 VSS.n3329 21.4593
R2451 VSS.n3340 VSS.n108 21.4593
R2452 VSS.n599 VSS.n585 21.4593
R2453 VSS.n1629 VSS.n1628 21.4593
R2454 VSS.n2592 VSS.n845 21.4593
R2455 VSS.n1979 VSS.n1978 21.4593
R2456 VSS.n1887 VSS.n1272 21.4593
R2457 VSS.n1699 VSS.n1556 20.8482
R2458 VSS.n1461 VSS.n1398 20.7064
R2459 VSS.n1449 VSS.n1401 20.7064
R2460 VSS.n3424 VSS.n60 20.3299
R2461 VSS.n3415 VSS.n3411 20.3299
R2462 VSS.n3371 VSS.n83 20.3299
R2463 VSS.n3362 VSS.n89 20.3299
R2464 VSS.t987 VSS 19.3418
R2465 VSS.t836 VSS 19.3418
R2466 VSS.t345 VSS 19.3418
R2467 VSS.n3430 VSS.n3429 19.2926
R2468 VSS.n3377 VSS.n3376 19.2926
R2469 VSS.n2394 VSS.t392 19.2511
R2470 VSS.t1006 VSS 19.0729
R2471 VSS.n3138 VSS.n3137 18.824
R2472 VSS.n132 VSS.n131 18.824
R2473 VSS.n137 VSS.n136 18.824
R2474 VSS.n142 VSS.n141 18.824
R2475 VSS.n147 VSS.n146 18.824
R2476 VSS.n152 VSS.n151 18.824
R2477 VSS.n157 VSS.n156 18.824
R2478 VSS.n162 VSS.n161 18.824
R2479 VSS.n167 VSS.n166 18.824
R2480 VSS.n2828 VSS.n2827 18.2791
R2481 VSS.n1517 VSS.n1362 18.2791
R2482 VSS.n1097 VSS.n1096 18.2791
R2483 VSS.n33 VSS.n22 17.7867
R2484 VSS.n3353 VSS.n3352 17.7867
R2485 VSS.n1074 VSS.n1055 17.7007
R2486 VSS.n2359 VSS.n2358 17.4137
R2487 VSS.n3421 VSS.n3420 17.3181
R2488 VSS.n3145 VSS.n3144 17.3181
R2489 VSS.n3170 VSS.n3169 17.3181
R2490 VSS.n3090 VSS.n3089 17.3181
R2491 VSS.n3368 VSS.n3367 17.3181
R2492 VSS.n1447 VSS.n1446 17.3181
R2493 VSS.n2233 VSS.n2232 17.195
R2494 VSS.n2792 VSS.n692 16.9936
R2495 VSS.n3020 VSS.n264 16.9545
R2496 VSS.n2600 VSS.n2599 16.9417
R2497 VSS.n1863 VSS.n1285 16.9417
R2498 VSS.t702 VSS.t1054 16.8587
R2499 VSS.t877 VSS.t267 16.8587
R2500 VSS.t540 VSS.t709 16.8587
R2501 VSS.t187 VSS.t720 16.8587
R2502 VSS.t887 VSS.t22 16.8587
R2503 VSS.t454 VSS.t1008 16.8587
R2504 VSS.n3040 VSS.n255 16.8353
R2505 VSS.n3035 VSS.n256 16.7924
R2506 VSS.n523 VSS.n522 16.763
R2507 VSS.n1012 VSS.n67 16.4566
R2508 VSS.n1466 VSS.n1465 16.1887
R2509 VSS.n1448 VSS.n1447 16.1887
R2510 VSS.n1695 VSS.n1556 16.1887
R2511 VSS.n3422 VSS.n3421 15.8123
R2512 VSS.n3445 VSS.n39 15.8123
R2513 VSS.n3139 VSS.n3138 15.8123
R2514 VSS.n3110 VSS.n3109 15.8123
R2515 VSS.n3369 VSS.n3368 15.8123
R2516 VSS.n3360 VSS.n3359 15.8123
R2517 VSS.n127 VSS.n69 15.8123
R2518 VSS.n3292 VSS.n171 15.8123
R2519 VSS.n1496 VSS.n1495 15.3963
R2520 VSS.n2985 VSS.n2984 15.3963
R2521 VSS.n2989 VSS.n2988 15.3963
R2522 VSS.n3089 VSS.n3088 15.0593
R2523 VSS.t562 VSS.n2393 14.9042
R2524 VSS.n2393 VSS.t759 14.9042
R2525 VSS.n1931 VSS.n1930 14.8179
R2526 VSS.n2988 VSS.n278 14.8179
R2527 VSS.n3445 VSS.n3444 14.775
R2528 VSS.n3461 VSS.n4 14.775
R2529 VSS.n3359 VSS.n92 14.775
R2530 VSS.n3324 VSS.n113 14.775
R2531 VSS.n617 VSS.n614 14.775
R2532 VSS.n1437 VSS.n1420 14.775
R2533 VSS.n1721 VSS.n1720 14.775
R2534 VSS.n1839 VSS.n1838 14.775
R2535 VSS.n2029 VSS.n2028 14.775
R2536 VSS.n2498 VSS.n2497 14.775
R2537 VSS.n2939 VSS.n2938 14.2735
R2538 VSS.n2540 VSS.n2539 14.065
R2539 VSS.n553 VSS.n550 14.0503
R2540 VSS.n2846 VSS.n2845 14.0503
R2541 VSS.n811 VSS.n808 14.0503
R2542 VSS.n1625 VSS.n1624 13.9299
R2543 VSS.n1866 VSS.n1273 13.9299
R2544 VSS.n970 VSS.n969 13.8859
R2545 VSS.n3455 VSS.n16 13.5534
R2546 VSS.n3334 VSS.n110 13.5534
R2547 VSS.n3396 VSS.n69 12.8005
R2548 VSS.n3396 VSS.n68 12.8005
R2549 VSS.n3402 VSS.n68 12.8005
R2550 VSS.n2172 VSS.n1174 12.8005
R2551 VSS.n2143 VSS.n2142 12.8005
R2552 VSS.n2679 VSS.n753 12.8005
R2553 VSS.n887 VSS.n886 12.8005
R2554 VSS.n1851 VSS.n1289 12.5161
R2555 VSS.n3070 VSS.n3069 12.424
R2556 VSS.n3065 VSS.n3055 12.424
R2557 VSS.n2792 VSS.n2791 12.1384
R2558 VSS.n1672 VSS.n1671 11.9309
R2559 VSS.n3143 VSS.n3142 11.3835
R2560 VSS.n1661 VSS.n1583 11.2946
R2561 VSS.n1858 VSS.n1286 11.2946
R2562 VSS.n53 VSS.n52 11.2844
R2563 VSS.n3307 VSS.n3306 11.2844
R2564 VSS.n306 VSS.n299 11.0382
R2565 VSS.n302 VSS.n299 11.0382
R2566 VSS.n300 VSS.n298 11.0382
R2567 VSS.n302 VSS.n298 11.0382
R2568 VSS.n314 VSS.n294 11.0382
R2569 VSS.n297 VSS.n294 11.0382
R2570 VSS.n296 VSS.n293 11.0382
R2571 VSS.n297 VSS.n293 11.0382
R2572 VSS.n291 VSS.n289 11.0382
R2573 VSS.n322 VSS.n291 11.0382
R2574 VSS.n292 VSS.n290 11.0382
R2575 VSS.n322 VSS.n292 11.0382
R2576 VSS.n365 VSS.n343 11.0382
R2577 VSS.n361 VSS.n343 11.0382
R2578 VSS.n344 VSS.n342 11.0382
R2579 VSS.n361 VSS.n342 11.0382
R2580 VSS.n337 VSS.n285 11.0382
R2581 VSS.n333 VSS.n285 11.0382
R2582 VSS.n286 VSS.n284 11.0382
R2583 VSS.n333 VSS.n284 11.0382
R2584 VSS.n3245 VSS.n3238 11.0382
R2585 VSS.n3238 VSS.n3237 11.0382
R2586 VSS.n3242 VSS.n3236 11.0382
R2587 VSS.n3237 VSS.n3236 11.0382
R2588 VSS.n3269 VSS.n3268 11.0382
R2589 VSS.n3268 VSS.n3267 11.0382
R2590 VSS.n3266 VSS.n3265 11.0382
R2591 VSS.n3267 VSS.n3266 11.0382
R2592 VSS.n3208 VSS.n3207 11.0382
R2593 VSS.n3213 VSS.n3208 11.0382
R2594 VSS.n3204 VSS.n3203 11.0382
R2595 VSS.n3213 VSS.n3204 11.0382
R2596 VSS.n3197 VSS.n3196 11.0382
R2597 VSS.n3196 VSS.n3195 11.0382
R2598 VSS.n3194 VSS.n3193 11.0382
R2599 VSS.n3195 VSS.n3194 11.0382
R2600 VSS.n3225 VSS.n178 11.0382
R2601 VSS.n3209 VSS.n178 11.0382
R2602 VSS.n179 VSS.n177 11.0382
R2603 VSS.n3209 VSS.n177 11.0382
R2604 VSS.n203 VSS.n196 11.0382
R2605 VSS.n207 VSS.n196 11.0382
R2606 VSS.n206 VSS.n205 11.0382
R2607 VSS.n207 VSS.n206 11.0382
R2608 VSS.n3259 VSS.n3254 11.0382
R2609 VSS.n3254 VSS.n3253 11.0382
R2610 VSS.n3256 VSS.n3252 11.0382
R2611 VSS.n3253 VSS.n3252 11.0382
R2612 VSS.n3388 VSS.n73 11.0382
R2613 VSS.n3392 VSS.n73 11.0382
R2614 VSS.n3391 VSS.n3390 11.0382
R2615 VSS.n3392 VSS.n3391 11.0382
R2616 VSS.n356 VSS.n348 11.0382
R2617 VSS.n348 VSS.n347 11.0382
R2618 VSS.n353 VSS.n346 11.0382
R2619 VSS.n347 VSS.n346 11.0382
R2620 VSS.n381 VSS.n372 11.0382
R2621 VSS.n377 VSS.n372 11.0382
R2622 VSS.n373 VSS.n371 11.0382
R2623 VSS.n377 VSS.n371 11.0382
R2624 VSS.n393 VSS.n280 11.0382
R2625 VSS.n397 VSS.n280 11.0382
R2626 VSS.n396 VSS.n395 11.0382
R2627 VSS.n397 VSS.n396 11.0382
R2628 VSS.n3076 VSS.n3075 11.0382
R2629 VSS.n3073 VSS.n3072 11.0382
R2630 VSS.n3064 VSS.n3063 11.0382
R2631 VSS.n3063 VSS.n3062 11.0382
R2632 VSS.n3059 VSS.n3058 11.0382
R2633 VSS.n3059 VSS.n223 11.0382
R2634 VSS.n2098 VSS.n2042 10.9091
R2635 VSS.n1431 VSS.n1430 10.8805
R2636 VSS.n471 VSS.t458 10.6509
R2637 VSS.n3066 VSS.n3065 10.6195
R2638 VSS.n3069 VSS.n3068 10.6189
R2639 VSS.n1340 VSS.n1339 10.5983
R2640 VSS.n657 VSS.n654 10.5417
R2641 VSS.n1470 VSS.n1466 10.5417
R2642 VSS.n1905 VSS.n1241 10.5417
R2643 VSS.n1865 VSS.n1863 10.5417
R2644 VSS.n2553 VSS.n940 10.5417
R2645 VSS.n392 VSS.n390 10.4476
R2646 VSS.n3246 VSS.n3241 10.4476
R2647 VSS.n3271 VSS.n3270 10.4476
R2648 VSS.n3224 VSS.n3223 10.4476
R2649 VSS.n3218 VSS.n3202 10.4476
R2650 VSS.n3199 VSS.n3198 10.4476
R2651 VSS.n3387 VSS.n3385 10.4476
R2652 VSS.n3276 VSS.n3275 10.4476
R2653 VSS.n3453 VSS.n3452 10.1652
R2654 VSS.n3336 VSS.n108 10.1652
R2655 VSS.n1495 VSS.n1494 10.1652
R2656 VSS.n1494 VSS.n1373 10.1652
R2657 VSS.n1694 VSS.n1693 10.1652
R2658 VSS.n2601 VSS.n2600 10.1652
R2659 VSS.n909 VSS.n908 10.1652
R2660 VSS.n2558 VSS.n937 10.1652
R2661 VSS.n637 VSS.n625 9.88085
R2662 VSS.n1747 VSS.n1746 9.7205
R2663 VSS.n247 VSS.n246 9.7205
R2664 VSS.n2437 VSS.n2436 9.71789
R2665 VSS.n2353 VSS.n2352 9.71789
R2666 VSS.n53 VSS.n42 9.70901
R2667 VSS.n3438 VSS.n3437 9.70901
R2668 VSS.n27 VSS.n26 9.70901
R2669 VSS.n3306 VSS.n3305 9.70901
R2670 VSS.n100 VSS.n99 9.70901
R2671 VSS.n3345 VSS.n3344 9.70901
R2672 VSS.n48 VSS.n47 9.41227
R2673 VSS.n3310 VSS.n3299 9.41227
R2674 VSS.n1637 VSS.n1604 9.41227
R2675 VSS.n1940 VSS.n1939 9.41227
R2676 VSS.n1921 VSS.n1920 9.41227
R2677 VSS.n2153 VSS.n1174 9.3031
R2678 VSS.n2143 VSS.n1182 9.3031
R2679 VSS.n2661 VSS.n753 9.3031
R2680 VSS.n1328 VSS.n1327 9.3031
R2681 VSS.n1721 VSS.n1535 9.3031
R2682 VSS.n1838 VSS.n1836 9.3031
R2683 VSS.n3447 VSS.n3446 9.3005
R2684 VSS.n3440 VSS.n3439 9.3005
R2685 VSS.n3442 VSS.n3441 9.3005
R2686 VSS.n3444 VSS.n3443 9.3005
R2687 VSS.n3445 VSS.n36 9.3005
R2688 VSS.n55 VSS.n54 9.3005
R2689 VSS.n56 VSS.n41 9.3005
R2690 VSS.n3431 VSS.n3430 9.3005
R2691 VSS.n3429 VSS.n59 9.3005
R2692 VSS.n3428 VSS.n3427 9.3005
R2693 VSS.n3426 VSS.n60 9.3005
R2694 VSS.n3425 VSS.n3424 9.3005
R2695 VSS.n3423 VSS.n61 9.3005
R2696 VSS.n3422 VSS.n62 9.3005
R2697 VSS.n3421 VSS.n3409 9.3005
R2698 VSS.n3420 VSS.n3410 9.3005
R2699 VSS.n3419 VSS.n3418 9.3005
R2700 VSS.n3417 VSS.n3411 9.3005
R2701 VSS.n3416 VSS.n3415 9.3005
R2702 VSS.n3414 VSS.n3413 9.3005
R2703 VSS.n3412 VSS.n39 9.3005
R2704 VSS.n29 VSS.n28 9.3005
R2705 VSS.n31 VSS.n23 9.3005
R2706 VSS.n34 VSS.n33 9.3005
R2707 VSS.n3461 VSS.n13 9.3005
R2708 VSS.n3460 VSS.n14 9.3005
R2709 VSS.n3459 VSS.n3458 9.3005
R2710 VSS.n3457 VSS.n16 9.3005
R2711 VSS.n3456 VSS.n3455 9.3005
R2712 VSS.n3454 VSS.n18 9.3005
R2713 VSS.n3453 VSS.n19 9.3005
R2714 VSS.n3452 VSS.n20 9.3005
R2715 VSS.n3451 VSS.n3450 9.3005
R2716 VSS.n35 VSS.n22 9.3005
R2717 VSS.n51 VSS.n50 9.3005
R2718 VSS.n49 VSS.n43 9.3005
R2719 VSS.n47 VSS.n46 9.3005
R2720 VSS.n45 VSS.n2 9.3005
R2721 VSS.n3465 VSS.n3464 9.3005
R2722 VSS.n6 VSS.n5 9.3005
R2723 VSS.n11 VSS.n10 9.3005
R2724 VSS.n12 VSS.n4 9.3005
R2725 VSS.n3111 VSS.n3110 9.3005
R2726 VSS.n3112 VSS.n3103 9.3005
R2727 VSS.n3141 VSS.n3140 9.3005
R2728 VSS.n3139 VSS.n213 9.3005
R2729 VSS.n3137 VSS.n3136 9.3005
R2730 VSS.n3135 VSS.n215 9.3005
R2731 VSS.n3085 VSS.n216 9.3005
R2732 VSS.n3087 VSS.n3086 9.3005
R2733 VSS.n3091 VSS.n3090 9.3005
R2734 VSS.n3092 VSS.n220 9.3005
R2735 VSS.n3094 VSS.n3093 9.3005
R2736 VSS.n3096 VSS.n217 9.3005
R2737 VSS.n3131 VSS.n3130 9.3005
R2738 VSS.n3128 VSS.n3127 9.3005
R2739 VSS.n3126 VSS.n3125 9.3005
R2740 VSS.n3123 VSS.n3099 9.3005
R2741 VSS.n3121 VSS.n3120 9.3005
R2742 VSS.n3119 VSS.n3118 9.3005
R2743 VSS.n3116 VSS.n3102 9.3005
R2744 VSS.n3114 VSS.n3113 9.3005
R2745 VSS.n3175 VSS.n3174 9.3005
R2746 VSS.n3171 VSS.n3170 9.3005
R2747 VSS.n3172 VSS.n195 9.3005
R2748 VSS.n3176 VSS.n194 9.3005
R2749 VSS.n3145 VSS.n211 9.3005
R2750 VSS.n3162 VSS.n3161 9.3005
R2751 VSS.n3160 VSS.n3159 9.3005
R2752 VSS.n3158 VSS.n3157 9.3005
R2753 VSS.n3155 VSS.n3147 9.3005
R2754 VSS.n3154 VSS.n3153 9.3005
R2755 VSS.n3152 VSS.n3151 9.3005
R2756 VSS.n3149 VSS.n188 9.3005
R2757 VSS.n3189 VSS.n3188 9.3005
R2758 VSS.n3187 VSS.n189 9.3005
R2759 VSS.n3186 VSS.n3185 9.3005
R2760 VSS.n3183 VSS.n190 9.3005
R2761 VSS.n3182 VSS.n3181 9.3005
R2762 VSS.n3180 VSS.n3179 9.3005
R2763 VSS.n3177 VSS.n193 9.3005
R2764 VSS.n3356 VSS.n95 9.3005
R2765 VSS.n102 VSS.n101 9.3005
R2766 VSS.n104 VSS.n103 9.3005
R2767 VSS.n105 VSS.n92 9.3005
R2768 VSS.n3359 VSS.n3358 9.3005
R2769 VSS.n3304 VSS.n3301 9.3005
R2770 VSS.n3303 VSS.n80 9.3005
R2771 VSS.n3378 VSS.n3377 9.3005
R2772 VSS.n3376 VSS.n82 9.3005
R2773 VSS.n3375 VSS.n3374 9.3005
R2774 VSS.n3373 VSS.n83 9.3005
R2775 VSS.n3372 VSS.n3371 9.3005
R2776 VSS.n3370 VSS.n84 9.3005
R2777 VSS.n3369 VSS.n85 9.3005
R2778 VSS.n3368 VSS.n87 9.3005
R2779 VSS.n3367 VSS.n88 9.3005
R2780 VSS.n3366 VSS.n3365 9.3005
R2781 VSS.n3364 VSS.n89 9.3005
R2782 VSS.n3363 VSS.n3362 9.3005
R2783 VSS.n3361 VSS.n90 9.3005
R2784 VSS.n3360 VSS.n91 9.3005
R2785 VSS.n3347 VSS.n3342 9.3005
R2786 VSS.n3350 VSS.n3349 9.3005
R2787 VSS.n3352 VSS.n3351 9.3005
R2788 VSS.n3308 VSS.n3300 9.3005
R2789 VSS.n3312 VSS.n3311 9.3005
R2790 VSS.n3313 VSS.n3299 9.3005
R2791 VSS.n3315 VSS.n3314 9.3005
R2792 VSS.n3317 VSS.n3316 9.3005
R2793 VSS.n3319 VSS.n3318 9.3005
R2794 VSS.n3321 VSS.n114 9.3005
R2795 VSS.n3325 VSS.n3324 9.3005
R2796 VSS.n3326 VSS.n113 9.3005
R2797 VSS.n3329 VSS.n3327 9.3005
R2798 VSS.n3331 VSS.n3330 9.3005
R2799 VSS.n3332 VSS.n110 9.3005
R2800 VSS.n3334 VSS.n3333 9.3005
R2801 VSS.n3335 VSS.n109 9.3005
R2802 VSS.n3337 VSS.n3336 9.3005
R2803 VSS.n3338 VSS.n108 9.3005
R2804 VSS.n3340 VSS.n3339 9.3005
R2805 VSS.n3354 VSS.n3353 9.3005
R2806 VSS.n3293 VSS.n3292 9.3005
R2807 VSS.n171 VSS.n170 9.3005
R2808 VSS.n3402 VSS.n3399 9.3005
R2809 VSS.n3398 VSS.n68 9.3005
R2810 VSS.n3397 VSS.n3396 9.3005
R2811 VSS.n126 VSS.n69 9.3005
R2812 VSS.n128 VSS.n127 9.3005
R2813 VSS.n129 VSS.n125 9.3005
R2814 VSS.n131 VSS.n130 9.3005
R2815 VSS.n133 VSS.n132 9.3005
R2816 VSS.n134 VSS.n124 9.3005
R2817 VSS.n136 VSS.n135 9.3005
R2818 VSS.n138 VSS.n137 9.3005
R2819 VSS.n139 VSS.n123 9.3005
R2820 VSS.n141 VSS.n140 9.3005
R2821 VSS.n143 VSS.n142 9.3005
R2822 VSS.n144 VSS.n122 9.3005
R2823 VSS.n146 VSS.n145 9.3005
R2824 VSS.n148 VSS.n147 9.3005
R2825 VSS.n149 VSS.n121 9.3005
R2826 VSS.n151 VSS.n150 9.3005
R2827 VSS.n153 VSS.n152 9.3005
R2828 VSS.n154 VSS.n120 9.3005
R2829 VSS.n156 VSS.n155 9.3005
R2830 VSS.n158 VSS.n157 9.3005
R2831 VSS.n159 VSS.n119 9.3005
R2832 VSS.n161 VSS.n160 9.3005
R2833 VSS.n163 VSS.n162 9.3005
R2834 VSS.n164 VSS.n118 9.3005
R2835 VSS.n166 VSS.n165 9.3005
R2836 VSS.n168 VSS.n167 9.3005
R2837 VSS.n169 VSS.n117 9.3005
R2838 VSS.n553 VSS.n552 9.3005
R2839 VSS.n556 VSS.n547 9.3005
R2840 VSS.n558 VSS.n557 9.3005
R2841 VSS.n560 VSS.n559 9.3005
R2842 VSS.n563 VSS.n562 9.3005
R2843 VSS.n545 VSS.n544 9.3005
R2844 VSS.n538 VSS.n537 9.3005
R2845 VSS.n527 VSS.n526 9.3005
R2846 VSS.n2932 VSS.n2931 9.3005
R2847 VSS.n2933 VSS.n524 9.3005
R2848 VSS.n2935 VSS.n2934 9.3005
R2849 VSS.n2937 VSS.n2936 9.3005
R2850 VSS.n2160 VSS.n1174 9.3005
R2851 VSS.n2156 VSS.n1174 9.3005
R2852 VSS.n2174 VSS.n2173 9.3005
R2853 VSS.n2176 VSS.n2175 9.3005
R2854 VSS.n2177 VSS.n1170 9.3005
R2855 VSS.n2181 VSS.n2180 9.3005
R2856 VSS.n2184 VSS.n2183 9.3005
R2857 VSS.n2186 VSS.n1167 9.3005
R2858 VSS.n2188 VSS.n2187 9.3005
R2859 VSS.n2201 VSS.n2200 9.3005
R2860 VSS.n2203 VSS.n2202 9.3005
R2861 VSS.n2205 VSS.n2204 9.3005
R2862 VSS.n2206 VSS.n1156 9.3005
R2863 VSS.n2209 VSS.n2208 9.3005
R2864 VSS.n2210 VSS.n1155 9.3005
R2865 VSS.n2212 VSS.n2211 9.3005
R2866 VSS.n2213 VSS.n1154 9.3005
R2867 VSS.n2216 VSS.n2215 9.3005
R2868 VSS.n2223 VSS.n2222 9.3005
R2869 VSS.n2221 VSS.n1153 9.3005
R2870 VSS.n2220 VSS.n2219 9.3005
R2871 VSS.n2219 VSS.n2218 9.3005
R2872 VSS.n2287 VSS.n2286 9.3005
R2873 VSS.n2286 VSS.n2285 9.3005
R2874 VSS.n2279 VSS.n2278 9.3005
R2875 VSS.n2276 VSS.n1127 9.3005
R2876 VSS.n2275 VSS.n2274 9.3005
R2877 VSS.n2273 VSS.n1128 9.3005
R2878 VSS.n2272 VSS.n2271 9.3005
R2879 VSS.n2270 VSS.n1129 9.3005
R2880 VSS.n2268 VSS.n2267 9.3005
R2881 VSS.n2266 VSS.n1130 9.3005
R2882 VSS.n2265 VSS.n2264 9.3005
R2883 VSS.n2262 VSS.n1131 9.3005
R2884 VSS.n1143 VSS.n1142 9.3005
R2885 VSS.n1147 VSS.n1146 9.3005
R2886 VSS.n2250 VSS.n2249 9.3005
R2887 VSS.n2248 VSS.n1139 9.3005
R2888 VSS.n2247 VSS.n2246 9.3005
R2889 VSS.n2245 VSS.n1148 9.3005
R2890 VSS.n2244 VSS.n2243 9.3005
R2891 VSS.n2242 VSS.n1149 9.3005
R2892 VSS.n2240 VSS.n2239 9.3005
R2893 VSS.n2238 VSS.n2237 9.3005
R2894 VSS.n2236 VSS.n2235 9.3005
R2895 VSS.n2234 VSS.n2233 9.3005
R2896 VSS.n2232 VSS.n2231 9.3005
R2897 VSS.n2230 VSS.n2229 9.3005
R2898 VSS.n2228 VSS.n513 9.3005
R2899 VSS.n517 VSS.n514 9.3005
R2900 VSS.n2952 VSS.n2951 9.3005
R2901 VSS.n2950 VSS.n2949 9.3005
R2902 VSS.n2948 VSS.n518 9.3005
R2903 VSS.n2947 VSS.n2946 9.3005
R2904 VSS.n2944 VSS.n519 9.3005
R2905 VSS.n2943 VSS.n2942 9.3005
R2906 VSS.n2941 VSS.n520 9.3005
R2907 VSS.n2940 VSS.n2939 9.3005
R2908 VSS.n2891 VSS.n580 9.3005
R2909 VSS.n2894 VSS.n2893 9.3005
R2910 VSS.n2895 VSS.n579 9.3005
R2911 VSS.n2897 VSS.n2896 9.3005
R2912 VSS.n2899 VSS.n578 9.3005
R2913 VSS.n2901 VSS.n2900 9.3005
R2914 VSS.n2903 VSS.n2902 9.3005
R2915 VSS.n583 VSS.n581 9.3005
R2916 VSS.n2888 VSS.n2887 9.3005
R2917 VSS.n2886 VSS.n2885 9.3005
R2918 VSS.n2884 VSS.n584 9.3005
R2919 VSS.n2881 VSS.n2880 9.3005
R2920 VSS.n599 VSS.n595 9.3005
R2921 VSS.n663 VSS.n596 9.3005
R2922 VSS.n638 VSS.n637 9.3005
R2923 VSS.n620 VSS.n611 9.3005
R2924 VSS.n617 VSS.n616 9.3005
R2925 VSS.n623 VSS.n622 9.3005
R2926 VSS.n625 VSS.n624 9.3005
R2927 VSS.n636 VSS.n635 9.3005
R2928 VSS.n631 VSS.n629 9.3005
R2929 VSS.n605 VSS.n604 9.3005
R2930 VSS.n648 VSS.n647 9.3005
R2931 VSS.n649 VSS.n603 9.3005
R2932 VSS.n651 VSS.n650 9.3005
R2933 VSS.n652 VSS.n602 9.3005
R2934 VSS.n654 VSS.n653 9.3005
R2935 VSS.n657 VSS.n601 9.3005
R2936 VSS.n659 VSS.n658 9.3005
R2937 VSS.n660 VSS.n600 9.3005
R2938 VSS.n662 VSS.n661 9.3005
R2939 VSS.n665 VSS.n664 9.3005
R2940 VSS.n593 VSS.n585 9.3005
R2941 VSS.n2905 VSS.n2904 9.3005
R2942 VSS.n2914 VSS.n2913 9.3005
R2943 VSS.n2916 VSS.n2915 9.3005
R2944 VSS.n2065 VSS.n575 9.3005
R2945 VSS.n2067 VSS.n2066 9.3005
R2946 VSS.n2144 VSS.n2143 9.3005
R2947 VSS.n2143 VSS.n1186 9.3005
R2948 VSS.n2141 VSS.n2140 9.3005
R2949 VSS.n2139 VSS.n2138 9.3005
R2950 VSS.n2137 VSS.n1199 9.3005
R2951 VSS.n2136 VSS.n2135 9.3005
R2952 VSS.n2133 VSS.n2132 9.3005
R2953 VSS.n2130 VSS.n2129 9.3005
R2954 VSS.n1212 VSS.n1205 9.3005
R2955 VSS.n1217 VSS.n1214 9.3005
R2956 VSS.n2119 VSS.n2118 9.3005
R2957 VSS.n2116 VSS.n1215 9.3005
R2958 VSS.n2115 VSS.n2114 9.3005
R2959 VSS.n2113 VSS.n1218 9.3005
R2960 VSS.n2112 VSS.n2111 9.3005
R2961 VSS.n2110 VSS.n1219 9.3005
R2962 VSS.n2109 VSS.n2108 9.3005
R2963 VSS.n2107 VSS.n2106 9.3005
R2964 VSS.n2040 VSS.n2038 9.3005
R2965 VSS.n2103 VSS.n2102 9.3005
R2966 VSS.n2101 VSS.n2100 9.3005
R2967 VSS.n2098 VSS.n2097 9.3005
R2968 VSS.n2044 VSS.n2043 9.3005
R2969 VSS.n2054 VSS.n2052 9.3005
R2970 VSS.n2087 VSS.n2086 9.3005
R2971 VSS.n2056 VSS.n2053 9.3005
R2972 VSS.n2081 VSS.n2080 9.3005
R2973 VSS.n2079 VSS.n2058 9.3005
R2974 VSS.n2078 VSS.n2077 9.3005
R2975 VSS.n2076 VSS.n2059 9.3005
R2976 VSS.n2074 VSS.n2073 9.3005
R2977 VSS.n2072 VSS.n2061 9.3005
R2978 VSS.n2071 VSS.n2070 9.3005
R2979 VSS.n2068 VSS.n2062 9.3005
R2980 VSS.n2788 VSS.n694 9.3005
R2981 VSS.n2787 VSS.n2786 9.3005
R2982 VSS.n2783 VSS.n695 9.3005
R2983 VSS.n2782 VSS.n2781 9.3005
R2984 VSS.n2780 VSS.n2779 9.3005
R2985 VSS.n2778 VSS.n697 9.3005
R2986 VSS.n2777 VSS.n2776 9.3005
R2987 VSS.n2775 VSS.n698 9.3005
R2988 VSS.n2763 VSS.n2762 9.3005
R2989 VSS.n2766 VSS.n2765 9.3005
R2990 VSS.n2790 VSS.n2789 9.3005
R2991 VSS.n2793 VSS.n2792 9.3005
R2992 VSS.n2801 VSS.n2800 9.3005
R2993 VSS.n2804 VSS.n2803 9.3005
R2994 VSS.n685 VSS.n684 9.3005
R2995 VSS.n2813 VSS.n2812 9.3005
R2996 VSS.n2815 VSS.n683 9.3005
R2997 VSS.n2819 VSS.n2818 9.3005
R2998 VSS.n2820 VSS.n682 9.3005
R2999 VSS.n2821 VSS 9.3005
R3000 VSS.n2825 VSS.n2824 9.3005
R3001 VSS.n2827 VSS.n2826 9.3005
R3002 VSS.n2828 VSS.n679 9.3005
R3003 VSS.n2831 VSS.n2830 9.3005
R3004 VSS.n2832 VSS.n678 9.3005
R3005 VSS.n2834 VSS.n2833 9.3005
R3006 VSS.n2835 VSS.n676 9.3005
R3007 VSS.n2864 VSS.n2863 9.3005
R3008 VSS.n2862 VSS.n2861 9.3005
R3009 VSS.n2854 VSS.n2837 9.3005
R3010 VSS.n2853 VSS.n2852 9.3005
R3011 VSS.n2851 VSS.n2839 9.3005
R3012 VSS.n2849 VSS.n2848 9.3005
R3013 VSS.n2847 VSS.n2846 9.3005
R3014 VSS.n2668 VSS.n753 9.3005
R3015 VSS.n2664 VSS.n753 9.3005
R3016 VSS.n2681 VSS.n2680 9.3005
R3017 VSS.n2683 VSS.n2682 9.3005
R3018 VSS.n2684 VSS.n749 9.3005
R3019 VSS.n2688 VSS.n2687 9.3005
R3020 VSS.n2691 VSS.n2690 9.3005
R3021 VSS.n2693 VSS.n746 9.3005
R3022 VSS.n2695 VSS.n2694 9.3005
R3023 VSS.n2708 VSS.n2707 9.3005
R3024 VSS.n2710 VSS.n2709 9.3005
R3025 VSS.n2712 VSS.n2711 9.3005
R3026 VSS.n2713 VSS.n735 9.3005
R3027 VSS.n2716 VSS.n2715 9.3005
R3028 VSS.n2717 VSS.n734 9.3005
R3029 VSS.n2719 VSS.n2718 9.3005
R3030 VSS.n2720 VSS.n733 9.3005
R3031 VSS.n2723 VSS.n2722 9.3005
R3032 VSS.n2725 VSS.n2724 9.3005
R3033 VSS.n2727 VSS.n2726 9.3005
R3034 VSS.n2729 VSS.n2728 9.3005
R3035 VSS.n2730 VSS.n2729 9.3005
R3036 VSS.n2739 VSS.n716 9.3005
R3037 VSS.n2739 VSS.n2738 9.3005
R3038 VSS.n2741 VSS.n715 9.3005
R3039 VSS.n2744 VSS.n2743 9.3005
R3040 VSS.n2745 VSS.n714 9.3005
R3041 VSS.n2747 VSS.n2746 9.3005
R3042 VSS.n2748 VSS.n713 9.3005
R3043 VSS.n2750 VSS.n2749 9.3005
R3044 VSS.n2752 VSS.n2751 9.3005
R3045 VSS.n2753 VSS.n711 9.3005
R3046 VSS.n2756 VSS.n2755 9.3005
R3047 VSS.n2758 VSS.n2757 9.3005
R3048 VSS.n1494 VSS.n1493 9.3005
R3049 VSS.n1482 VSS.n1481 9.3005
R3050 VSS.n1479 VSS.n1478 9.3005
R3051 VSS.n1446 VSS.n1445 9.3005
R3052 VSS.n1437 VSS.n1436 9.3005
R3053 VSS.n1426 VSS.n1421 9.3005
R3054 VSS.n1428 VSS.n1427 9.3005
R3055 VSS.n1424 VSS.n767 9.3005
R3056 VSS.n1423 VSS.n768 9.3005
R3057 VSS.n2642 VSS.n2641 9.3005
R3058 VSS.n2640 VSS.n2639 9.3005
R3059 VSS.n2638 VSS.n2637 9.3005
R3060 VSS.n2636 VSS.n775 9.3005
R3061 VSS.n2633 VSS.n2632 9.3005
R3062 VSS.n2631 VSS.n777 9.3005
R3063 VSS.n2630 VSS.n2629 9.3005
R3064 VSS.n2627 VSS.n778 9.3005
R3065 VSS.n2624 VSS.n2623 9.3005
R3066 VSS.n2622 VSS.n2621 9.3005
R3067 VSS.n2619 VSS.n782 9.3005
R3068 VSS.n2618 VSS.n2617 9.3005
R3069 VSS.n786 VSS.n785 9.3005
R3070 VSS.n801 VSS.n800 9.3005
R3071 VSS.n802 VSS.n791 9.3005
R3072 VSS.n821 VSS.n820 9.3005
R3073 VSS.n818 VSS.n817 9.3005
R3074 VSS.n816 VSS.n815 9.3005
R3075 VSS.n814 VSS.n805 9.3005
R3076 VSS.n811 VSS.n810 9.3005
R3077 VSS.n1434 VSS.n1433 9.3005
R3078 VSS.n1435 VSS.n1420 9.3005
R3079 VSS.n1441 VSS.n1417 9.3005
R3080 VSS.n1443 VSS.n1442 9.3005
R3081 VSS.n1444 VSS.n1415 9.3005
R3082 VSS.n1447 VSS.n1414 9.3005
R3083 VSS.n1448 VSS.n1411 9.3005
R3084 VSS.n1450 VSS.n1449 9.3005
R3085 VSS.n1403 VSS.n1401 9.3005
R3086 VSS.n1459 VSS.n1458 9.3005
R3087 VSS.n1462 VSS.n1461 9.3005
R3088 VSS.n1463 VSS.n1398 9.3005
R3089 VSS.n1465 VSS.n1464 9.3005
R3090 VSS.n1466 VSS.n1395 9.3005
R3091 VSS.n1471 VSS.n1470 9.3005
R3092 VSS.n1472 VSS.n1394 9.3005
R3093 VSS.n1474 VSS.n1473 9.3005
R3094 VSS.n1477 VSS.n1390 9.3005
R3095 VSS.n1480 VSS.n1389 9.3005
R3096 VSS.n1486 VSS.n1485 9.3005
R3097 VSS.n1386 VSS.n1373 9.3005
R3098 VSS.n1495 VSS.n1371 9.3005
R3099 VSS.n1497 VSS.n1496 9.3005
R3100 VSS.n1498 VSS.n1369 9.3005
R3101 VSS.n1500 VSS.n1499 9.3005
R3102 VSS.n1501 VSS.n1367 9.3005
R3103 VSS.n1504 VSS.n1503 9.3005
R3104 VSS.n1505 VSS.n1366 9.3005
R3105 VSS.n1507 VSS.n1506 9.3005
R3106 VSS.n1508 VSS.n1364 9.3005
R3107 VSS.n1511 VSS.n1510 9.3005
R3108 VSS.n1512 VSS.n1363 9.3005
R3109 VSS.n1514 VSS.n1513 9.3005
R3110 VSS.n1518 VSS.n1517 9.3005
R3111 VSS.n1328 VSS.n1318 9.3005
R3112 VSS.n1329 VSS.n1328 9.3005
R3113 VSS.n1337 VSS.n1314 9.3005
R3114 VSS.n1339 VSS.n1338 9.3005
R3115 VSS.n1342 VSS.n1341 9.3005
R3116 VSS.n1344 VSS.n1343 9.3005
R3117 VSS.n1345 VSS.n1312 9.3005
R3118 VSS.n1348 VSS.n1347 9.3005
R3119 VSS.n1349 VSS.n1311 9.3005
R3120 VSS.n1351 VSS.n1350 9.3005
R3121 VSS.n1352 VSS.n1309 9.3005
R3122 VSS.n1355 VSS.n1354 9.3005
R3123 VSS.n1356 VSS.n1308 9.3005
R3124 VSS.n1358 VSS.n1357 9.3005
R3125 VSS.n1360 VSS.n1303 9.3005
R3126 VSS.n1362 VSS.n1304 9.3005
R3127 VSS.n1722 VSS.n1721 9.3005
R3128 VSS.n1721 VSS.n1539 9.3005
R3129 VSS.n1720 VSS.n1719 9.3005
R3130 VSS.n1718 VSS.n1717 9.3005
R3131 VSS.n1712 VSS.n1711 9.3005
R3132 VSS.n1710 VSS.n1550 9.3005
R3133 VSS.n1708 VSS.n1707 9.3005
R3134 VSS.n1706 VSS.n1705 9.3005
R3135 VSS.n1554 VSS.n1553 9.3005
R3136 VSS.n1699 VSS.n1698 9.3005
R3137 VSS.n1697 VSS.n1556 9.3005
R3138 VSS.n1696 VSS.n1695 9.3005
R3139 VSS.n1693 VSS.n1692 9.3005
R3140 VSS.n1570 VSS.n1569 9.3005
R3141 VSS.n1572 VSS.n1566 9.3005
R3142 VSS.n1682 VSS.n1681 9.3005
R3143 VSS.n1679 VSS.n1567 9.3005
R3144 VSS.n1677 VSS.n1676 9.3005
R3145 VSS.n1675 VSS.n1674 9.3005
R3146 VSS.n1672 VSS.n1576 9.3005
R3147 VSS.n1669 VSS.n1668 9.3005
R3148 VSS.n1667 VSS.n1666 9.3005
R3149 VSS.n1662 VSS.n1579 9.3005
R3150 VSS.n1661 VSS.n1660 9.3005
R3151 VSS.n1659 VSS.n1658 9.3005
R3152 VSS.n1657 VSS.n1584 9.3005
R3153 VSS.n1654 VSS.n1653 9.3005
R3154 VSS.n1589 VSS.n1587 9.3005
R3155 VSS.n1600 VSS.n1596 9.3005
R3156 VSS.n1643 VSS.n1642 9.3005
R3157 VSS.n1641 VSS.n1640 9.3005
R3158 VSS.n1639 VSS.n1601 9.3005
R3159 VSS.n1638 VSS.n1637 9.3005
R3160 VSS.n1636 VSS.n1602 9.3005
R3161 VSS.n1635 VSS.n1634 9.3005
R3162 VSS.n1633 VSS.n1606 9.3005
R3163 VSS.n1632 VSS.n1631 9.3005
R3164 VSS.n1630 VSS.n1607 9.3005
R3165 VSS.n1629 VSS.n1609 9.3005
R3166 VSS.n1628 VSS.n1627 9.3005
R3167 VSS.n1626 VSS.n1625 9.3005
R3168 VSS.n1624 VSS.n1623 9.3005
R3169 VSS.n1615 VSS.n835 9.3005
R3170 VSS.n2603 VSS.n2602 9.3005
R3171 VSS.n2600 VSS.n834 9.3005
R3172 VSS.n2599 VSS.n837 9.3005
R3173 VSS.n2598 VSS.n2597 9.3005
R3174 VSS.n2595 VSS.n2594 9.3005
R3175 VSS.n2592 VSS.n2591 9.3005
R3176 VSS.n2590 VSS.n845 9.3005
R3177 VSS.n2589 VSS.n2588 9.3005
R3178 VSS.n2587 VSS.n847 9.3005
R3179 VSS.n2586 VSS.n2585 9.3005
R3180 VSS.n850 VSS.n848 9.3005
R3181 VSS.n921 VSS.n920 9.3005
R3182 VSS.n919 VSS.n852 9.3005
R3183 VSS.n917 VSS.n855 9.3005
R3184 VSS.n916 VSS.n856 9.3005
R3185 VSS.n915 VSS.n914 9.3005
R3186 VSS.n913 VSS.n857 9.3005
R3187 VSS.n912 VSS.n911 9.3005
R3188 VSS.n910 VSS.n858 9.3005
R3189 VSS.n908 VSS.n907 9.3005
R3190 VSS.n906 VSS.n905 9.3005
R3191 VSS.n904 VSS.n862 9.3005
R3192 VSS.n903 VSS.n902 9.3005
R3193 VSS.n865 VSS.n863 9.3005
R3194 VSS.n876 VSS.n872 9.3005
R3195 VSS.n892 VSS.n891 9.3005
R3196 VSS.n889 VSS.n873 9.3005
R3197 VSS.n887 VSS.n881 9.3005
R3198 VSS.n1838 VSS.n1294 9.3005
R3199 VSS.n1838 VSS.n1293 9.3005
R3200 VSS.n1840 VSS.n1839 9.3005
R3201 VSS.n1842 VSS.n1841 9.3005
R3202 VSS.n1847 VSS.n1846 9.3005
R3203 VSS.n1848 VSS.n1289 9.3005
R3204 VSS.n1851 VSS.n1849 9.3005
R3205 VSS.n1852 VSS.n1287 9.3005
R3206 VSS.n1855 VSS.n1854 9.3005
R3207 VSS.n1856 VSS.n1286 9.3005
R3208 VSS.n1858 VSS.n1857 9.3005
R3209 VSS.n1860 VSS.n1859 9.3005
R3210 VSS.n1861 VSS.n1285 9.3005
R3211 VSS.n1863 VSS.n1862 9.3005
R3212 VSS.n1865 VSS.n1282 9.3005
R3213 VSS.n1868 VSS.n1867 9.3005
R3214 VSS.n1866 VSS.n1274 9.3005
R3215 VSS.n1880 VSS.n1273 9.3005
R3216 VSS.n1882 VSS.n1881 9.3005
R3217 VSS.n1884 VSS.n1883 9.3005
R3218 VSS.n1885 VSS.n1272 9.3005
R3219 VSS.n1887 VSS.n1886 9.3005
R3220 VSS.n1888 VSS.n1269 9.3005
R3221 VSS.n1893 VSS.n1892 9.3005
R3222 VSS.n1894 VSS.n1268 9.3005
R3223 VSS.n1915 VSS.n1895 9.3005
R3224 VSS.n1913 VSS.n1912 9.3005
R3225 VSS.n1911 VSS.n1896 9.3005
R3226 VSS.n1904 VSS.n1897 9.3005
R3227 VSS.n1906 VSS.n1905 9.3005
R3228 VSS.n1241 VSS.n1238 9.3005
R3229 VSS.n1980 VSS.n1979 9.3005
R3230 VSS.n1978 VSS.n1239 9.3005
R3231 VSS.n1976 VSS.n1975 9.3005
R3232 VSS.n1974 VSS.n1242 9.3005
R3233 VSS.n1973 VSS.n1972 9.3005
R3234 VSS.n1246 VSS.n1243 9.3005
R3235 VSS.n1967 VSS.n1966 9.3005
R3236 VSS.n1965 VSS.n1245 9.3005
R3237 VSS.n1964 VSS.n1963 9.3005
R3238 VSS.n1962 VSS.n1247 9.3005
R3239 VSS.n1961 VSS.n1960 9.3005
R3240 VSS.n1959 VSS.n1958 9.3005
R3241 VSS.n1957 VSS.n1956 9.3005
R3242 VSS.n1264 VSS.n1253 9.3005
R3243 VSS.n1948 VSS.n1947 9.3005
R3244 VSS.n1946 VSS.n1261 9.3005
R3245 VSS.n1944 VSS.n1943 9.3005
R3246 VSS.n1942 VSS.n1265 9.3005
R3247 VSS.n1941 VSS.n1940 9.3005
R3248 VSS.n1936 VSS.n1266 9.3005
R3249 VSS.n1935 VSS.n1934 9.3005
R3250 VSS.n1933 VSS.n1267 9.3005
R3251 VSS.n1932 VSS.n1931 9.3005
R3252 VSS.n1930 VSS.n1929 9.3005
R3253 VSS.n1928 VSS.n1927 9.3005
R3254 VSS.n1924 VSS.n1923 9.3005
R3255 VSS.n1922 VSS.n929 9.3005
R3256 VSS.n1920 VSS.n930 9.3005
R3257 VSS.n2561 VSS.n2560 9.3005
R3258 VSS.n2559 VSS.n935 9.3005
R3259 VSS.n2558 VSS.n2557 9.3005
R3260 VSS.n2556 VSS.n2555 9.3005
R3261 VSS.n2554 VSS.n938 9.3005
R3262 VSS.n2553 VSS.n2552 9.3005
R3263 VSS.n2551 VSS.n940 9.3005
R3264 VSS.n2550 VSS.n2549 9.3005
R3265 VSS.n2548 VSS.n941 9.3005
R3266 VSS.n2547 VSS.n2546 9.3005
R3267 VSS.n2545 VSS.n2544 9.3005
R3268 VSS.n2540 VSS.n945 9.3005
R3269 VSS.n2538 VSS.n2537 9.3005
R3270 VSS.n961 VSS.n950 9.3005
R3271 VSS.n962 VSS.n958 9.3005
R3272 VSS.n978 VSS.n977 9.3005
R3273 VSS.n976 VSS.n959 9.3005
R3274 VSS.n975 VSS.n974 9.3005
R3275 VSS.n973 VSS.n972 9.3005
R3276 VSS.n970 VSS.n965 9.3005
R3277 VSS.n2440 VSS.n2439 9.3005
R3278 VSS.n2442 VSS.n2441 9.3005
R3279 VSS.n1744 VSS.n1742 9.3005
R3280 VSS.n1757 VSS.n1756 9.3005
R3281 VSS.n1825 VSS.n1824 9.3005
R3282 VSS.n1823 VSS.n1759 9.3005
R3283 VSS.n1822 VSS.n1821 9.3005
R3284 VSS.n1820 VSS.n1760 9.3005
R3285 VSS.n1819 VSS.n1818 9.3005
R3286 VSS.n1817 VSS.n1761 9.3005
R3287 VSS.n1816 VSS.n1815 9.3005
R3288 VSS.n1814 VSS.n1813 9.3005
R3289 VSS.n1812 VSS.n1764 9.3005
R3290 VSS.n1809 VSS.n1808 9.3005
R3291 VSS.n1807 VSS.n1765 9.3005
R3292 VSS.n1806 VSS.n1805 9.3005
R3293 VSS.n1804 VSS.n1803 9.3005
R3294 VSS.n1775 VSS.n1768 9.3005
R3295 VSS.n1779 VSS.n1777 9.3005
R3296 VSS.n1793 VSS.n1792 9.3005
R3297 VSS.n1791 VSS.n1778 9.3005
R3298 VSS.n1788 VSS.n1787 9.3005
R3299 VSS.n1786 VSS.n1784 9.3005
R3300 VSS.n1785 VSS.n1223 9.3005
R3301 VSS.n2029 VSS.n1224 9.3005
R3302 VSS.n2028 VSS.n2027 9.3005
R3303 VSS.n2026 VSS.n2025 9.3005
R3304 VSS.n2024 VSS.n2023 9.3005
R3305 VSS.n2012 VSS.n1229 9.3005
R3306 VSS.n2012 VSS.n1990 9.3005
R3307 VSS.n2013 VSS.n2012 9.3005
R3308 VSS.n2011 VSS.n2010 9.3005
R3309 VSS.n2009 VSS.n1992 9.3005
R3310 VSS.n2008 VSS.n2007 9.3005
R3311 VSS.n2006 VSS.n2005 9.3005
R3312 VSS.n2004 VSS.n1993 9.3005
R3313 VSS.n2003 VSS.n2002 9.3005
R3314 VSS.n2001 VSS.n1994 9.3005
R3315 VSS.n1997 VSS.n989 9.3005
R3316 VSS.n2520 VSS.n2519 9.3005
R3317 VSS.n2518 VSS.n2517 9.3005
R3318 VSS.n2512 VSS.n991 9.3005
R3319 VSS.n2511 VSS.n2510 9.3005
R3320 VSS.n2508 VSS.n995 9.3005
R3321 VSS.n2507 VSS.n2506 9.3005
R3322 VSS.n2505 VSS.n2504 9.3005
R3323 VSS.n2503 VSS.n2502 9.3005
R3324 VSS.n2501 VSS.n999 9.3005
R3325 VSS.n2500 VSS.n2499 9.3005
R3326 VSS.n2498 VSS.n2396 9.3005
R3327 VSS.n2497 VSS.n2496 9.3005
R3328 VSS.n2495 VSS.n2494 9.3005
R3329 VSS.n2493 VSS.n2398 9.3005
R3330 VSS.n2492 VSS.n2491 9.3005
R3331 VSS.n2407 VSS.n2399 9.3005
R3332 VSS.n2475 VSS.n2409 9.3005
R3333 VSS.n2481 VSS.n2480 9.3005
R3334 VSS.n2473 VSS.n2410 9.3005
R3335 VSS.n2472 VSS.n2471 9.3005
R3336 VSS.n2470 VSS.n2413 9.3005
R3337 VSS.n2469 VSS.n2468 9.3005
R3338 VSS.n2467 VSS.n2466 9.3005
R3339 VSS.n2465 VSS.n2414 9.3005
R3340 VSS.n2464 VSS.n2463 9.3005
R3341 VSS.n2462 VSS.n2415 9.3005
R3342 VSS.n2460 VSS.n2418 9.3005
R3343 VSS.n2459 VSS.n2458 9.3005
R3344 VSS.n2431 VSS.n2421 9.3005
R3345 VSS.n2450 VSS.n2449 9.3005
R3346 VSS.n2448 VSS.n2447 9.3005
R3347 VSS.n2446 VSS.n2432 9.3005
R3348 VSS.n2445 VSS.n2444 9.3005
R3349 VSS.n2443 VSS.n2433 9.3005
R3350 VSS.n244 VSS.n241 9.3005
R3351 VSS.n255 VSS.n254 9.3005
R3352 VSS.n3041 VSS.n3040 9.3005
R3353 VSS.n3038 VSS.n239 9.3005
R3354 VSS.n3035 VSS.n3034 9.3005
R3355 VSS.n3033 VSS.n256 9.3005
R3356 VSS.n3032 VSS.n3031 9.3005
R3357 VSS.n3030 VSS.n257 9.3005
R3358 VSS.n3029 VSS.n3028 9.3005
R3359 VSS.n3027 VSS.n259 9.3005
R3360 VSS.n3026 VSS.n3025 9.3005
R3361 VSS.n262 VSS.n260 9.3005
R3362 VSS.n3020 VSS.n3019 9.3005
R3363 VSS.n3018 VSS.n264 9.3005
R3364 VSS.n272 VSS.n265 9.3005
R3365 VSS.n3010 VSS.n3009 9.3005
R3366 VSS.n3008 VSS.n3007 9.3005
R3367 VSS.n3001 VSS.n273 9.3005
R3368 VSS.n3000 VSS.n2999 9.3005
R3369 VSS.n2998 VSS.n274 9.3005
R3370 VSS.n2997 VSS.n2996 9.3005
R3371 VSS.n2995 VSS.n2994 9.3005
R3372 VSS.n2993 VSS.n276 9.3005
R3373 VSS.n2992 VSS.n2991 9.3005
R3374 VSS.n2990 VSS.n2989 9.3005
R3375 VSS.n2988 VSS.n279 9.3005
R3376 VSS.n1058 VSS.n278 9.3005
R3377 VSS.n1063 VSS.n1062 9.3005
R3378 VSS.n1065 VSS.n1055 9.3005
R3379 VSS.n1074 VSS.n1073 9.3005
R3380 VSS.n1076 VSS.n1053 9.3005
R3381 VSS.n1113 VSS.n1112 9.3005
R3382 VSS.n1111 VSS.n1054 9.3005
R3383 VSS.n1110 VSS.n1109 9.3005
R3384 VSS.n1108 VSS.n1077 9.3005
R3385 VSS.n1107 VSS.n1106 9.3005
R3386 VSS.n1105 VSS.n1078 9.3005
R3387 VSS.n1103 VSS.n1102 9.3005
R3388 VSS.n1101 VSS.n1079 9.3005
R3389 VSS.n1100 VSS.n1099 9.3005
R3390 VSS.n1097 VSS 9.3005
R3391 VSS.n1096 VSS.n1095 9.3005
R3392 VSS.n1094 VSS.n1093 9.3005
R3393 VSS.n1092 VSS.n1091 9.3005
R3394 VSS.n1084 VSS.n1082 9.3005
R3395 VSS.n2972 VSS.n499 9.3005
R3396 VSS.n2974 VSS.n2973 9.3005
R3397 VSS.n2975 VSS.n498 9.3005
R3398 VSS.n2977 VSS.n2976 9.3005
R3399 VSS.n2979 VSS.n2978 9.3005
R3400 VSS.n2980 VSS.n496 9.3005
R3401 VSS.n2982 VSS.n2981 9.3005
R3402 VSS.n2984 VSS.n2983 9.3005
R3403 VSS.n2985 VSS.n494 9.3005
R3404 VSS.n1040 VSS.n493 9.3005
R3405 VSS.n1042 VSS.n1041 9.3005
R3406 VSS.n1044 VSS.n1043 9.3005
R3407 VSS.n2314 VSS.n2313 9.3005
R3408 VSS.n2316 VSS.n2315 9.3005
R3409 VSS.n1036 VSS.n1035 9.3005
R3410 VSS.n2322 VSS.n2321 9.3005
R3411 VSS.n2323 VSS.n1033 9.3005
R3412 VSS.n2329 VSS.n2328 9.3005
R3413 VSS.n2331 VSS.n2330 9.3005
R3414 VSS.n2333 VSS.n2332 9.3005
R3415 VSS.n2334 VSS.n1031 9.3005
R3416 VSS.n2336 VSS.n2335 9.3005
R3417 VSS.n2337 VSS.n1029 9.3005
R3418 VSS.n2340 VSS.n2339 9.3005
R3419 VSS.n2341 VSS.n1028 9.3005
R3420 VSS.n2343 VSS.n2342 9.3005
R3421 VSS.n2344 VSS.n1025 9.3005
R3422 VSS.n2371 VSS.n2370 9.3005
R3423 VSS.n2369 VSS.n2368 9.3005
R3424 VSS.n2366 VSS.n2345 9.3005
R3425 VSS.n2365 VSS.n2364 9.3005
R3426 VSS.n2363 VSS.n2348 9.3005
R3427 VSS.n2362 VSS.n2361 9.3005
R3428 VSS.n2360 VSS.n2359 9.3005
R3429 VSS.n2358 VSS.n2357 9.3005
R3430 VSS.n2356 VSS.n2355 9.3005
R3431 VSS.n1446 VSS.n1415 9.12791
R3432 VSS.n1477 VSS.n1476 9.03579
R3433 VSS.n1393 VSS.n1392 9.03579
R3434 VSS.n1674 VSS.n1575 9.03579
R3435 VSS.n2626 VSS.n2624 8.9684
R3436 VSS.n328 VSS.n327 8.44328
R3437 VSS.n350 VSS.n349 8.44328
R3438 VSS.n3220 VSS.n3219 8.44328
R3439 VSS.n3274 VSS.n3273 8.44328
R3440 VSS.t594 VSS.t94 8.42962
R3441 VSS.t552 VSS.t474 8.42962
R3442 VSS.t196 VSS.t1082 8.42962
R3443 VSS VSS.n3406 8.3721
R3444 VSS.n331 VSS.n330 8.33966
R3445 VSS.n3384 VSS.n3383 8.33966
R3446 VSS.n200 VSS.n181 8.31061
R3447 VSS.n3054 VSS.n227 8.30267
R3448 VSS.n918 VSS.n917 8.28285
R3449 VSS.n2223 VSS.n1153 8.23546
R3450 VSS.n2934 VSS.n2933 8.23546
R3451 VSS.n2933 VSS.n2932 8.23546
R3452 VSS.n2932 VSS.n526 8.23546
R3453 VSS.n562 VSS.n545 8.23546
R3454 VSS.n2830 VSS.n678 8.23546
R3455 VSS.n2834 VSS.n678 8.23546
R3456 VSS.n2803 VSS.n684 8.23546
R3457 VSS.n2813 VSS.n684 8.23546
R3458 VSS.n2821 VSS.n682 8.23546
R3459 VSS.n2824 VSS.n2821 8.23546
R3460 VSS.n2726 VSS.n2725 8.23546
R3461 VSS.n2619 VSS.n2618 8.23546
R3462 VSS.n2618 VSS.n785 8.23546
R3463 VSS.n802 VSS.n801 8.23546
R3464 VSS.n1424 VSS.n1423 8.23546
R3465 VSS.n2641 VSS.n2640 8.23546
R3466 VSS.n2637 VSS.n2636 8.23546
R3467 VSS.n2633 VSS.n777 8.23546
R3468 VSS.n1352 VSS.n1351 8.23546
R3469 VSS.n1354 VSS.n1352 8.23546
R3470 VSS.n1358 VSS.n1308 8.23546
R3471 VSS.n1514 VSS.n1363 8.23546
R3472 VSS.n1510 VSS.n1363 8.23546
R3473 VSS.n1508 VSS.n1507 8.23546
R3474 VSS.n1507 VSS.n1366 8.23546
R3475 VSS.n1503 VSS.n1366 8.23546
R3476 VSS.n1501 VSS.n1500 8.23546
R3477 VSS.n1500 VSS.n1369 8.23546
R3478 VSS.n1967 VSS.n1245 8.23546
R3479 VSS.n1963 VSS.n1245 8.23546
R3480 VSS.n1963 VSS.n1962 8.23546
R3481 VSS.n1962 VSS.n1961 8.23546
R3482 VSS.n1958 VSS.n1957 8.23546
R3483 VSS.n1947 VSS.n1264 8.23546
R3484 VSS.n1947 VSS.n1946 8.23546
R3485 VSS.n2339 VSS.n1028 8.23546
R3486 VSS.n2343 VSS.n1028 8.23546
R3487 VSS.n2344 VSS.n2343 8.23546
R3488 VSS.n2370 VSS.n2344 8.23546
R3489 VSS.n2370 VSS.n2369 8.23546
R3490 VSS.n2369 VSS.n2345 8.23546
R3491 VSS.n2364 VSS.n2363 8.23546
R3492 VSS.n2363 VSS.n2362 8.23546
R3493 VSS.n1093 VSS.n1092 8.23546
R3494 VSS.n1092 VSS.n1082 8.23546
R3495 VSS.n1082 VSS.n499 8.23546
R3496 VSS.n2974 VSS.n499 8.23546
R3497 VSS.n2975 VSS.n2974 8.23546
R3498 VSS.n2976 VSS.n2975 8.23546
R3499 VSS.n2980 VSS.n2979 8.23546
R3500 VSS.n2981 VSS.n2980 8.23546
R3501 VSS.n1112 VSS.n1076 8.23546
R3502 VSS.n1112 VSS.n1111 8.23546
R3503 VSS.n1111 VSS.n1110 8.23546
R3504 VSS.n1110 VSS.n1077 8.23546
R3505 VSS.n1106 VSS.n1077 8.23546
R3506 VSS.n1106 VSS.n1105 8.23546
R3507 VSS.n1103 VSS.n1079 8.23546
R3508 VSS.n1099 VSS.n1079 8.23546
R3509 VSS.n3009 VSS.n272 8.23546
R3510 VSS.n3009 VSS.n3008 8.23546
R3511 VSS.n3008 VSS.n273 8.23546
R3512 VSS.n2999 VSS.n273 8.23546
R3513 VSS.n2999 VSS.n2998 8.23546
R3514 VSS.n2998 VSS.n2997 8.23546
R3515 VSS.n2994 VSS.n2993 8.23546
R3516 VSS.n2993 VSS.n2992 8.23546
R3517 VSS.n2815 VSS.n2814 8.14595
R3518 VSS.n537 VSS.n536 8.05644
R3519 VSS.n329 VSS.n287 7.97888
R3520 VSS.n374 VSS.n228 7.97888
R3521 VSS.n3240 VSS.n78 7.97888
R3522 VSS.n3201 VSS.n3200 7.97888
R3523 VSS.n328 VSS.n288 7.97601
R3524 VSS.n351 VSS.n350 7.97601
R3525 VSS.n3273 VSS.n3272 7.97601
R3526 VSS.n3221 VSS.n3220 7.97601
R3527 VSS.n1470 VSS.n1469 7.90638
R3528 VSS.n1628 VSS.n1612 7.90638
R3529 VSS.n2549 VSS.n943 7.90638
R3530 VSS.n1360 VSS.n1359 7.78791
R3531 VSS.n1970 VSS.n1969 7.72113
R3532 VSS.n2236 VSS.n2226 7.6984
R3533 VSS.n2934 VSS.n525 7.6984
R3534 VSS.n2830 VSS.n2829 7.6984
R3535 VSS.n2818 VSS.n2816 7.6984
R3536 VSS.n2621 VSS.n781 7.6984
R3537 VSS.n1429 VSS.n1428 7.6984
R3538 VSS.n1428 VSS.n1425 7.6984
R3539 VSS.n2629 VSS.n2628 7.6984
R3540 VSS.n1361 VSS.n1360 7.6984
R3541 VSS.n1370 VSS.n1369 7.6984
R3542 VSS.n1968 VSS.n1967 7.6984
R3543 VSS.n1946 VSS.n1945 7.6984
R3544 VSS.n2339 VSS.n2338 7.6984
R3545 VSS.n2362 VSS.n2350 7.6984
R3546 VSS.n1093 VSS.n1080 7.6984
R3547 VSS.n2981 VSS.n495 7.6984
R3548 VSS.n1076 VSS.n1075 7.6984
R3549 VSS.n1099 VSS.n1098 7.6984
R3550 VSS.n272 VSS.n271 7.6984
R3551 VSS.n2992 VSS.n277 7.6984
R3552 VSS.n3144 VSS.n212 7.64725
R3553 VSS.n3169 VSS.n3167 7.64725
R3554 VSS.n3089 VSS.n221 7.64725
R3555 VSS.n3108 VSS.n3107 7.64725
R3556 VSS.n948 VSS.n947 7.6005
R3557 VSS.n1509 VSS.n1508 7.51938
R3558 VSS.n2824 VSS.n2823 7.34036
R3559 VSS.n1958 VSS.n1249 7.34036
R3560 VSS.n793 VSS.n785 7.25085
R3561 VSS.n1516 VSS.n1515 7.25085
R3562 VSS.n390 VSS.n227 7.16724
R3563 VSS.n3241 VSS.n3240 7.16724
R3564 VSS.n3272 VSS.n3271 7.16724
R3565 VSS.n3223 VSS.n3221 7.16724
R3566 VSS.n3219 VSS.n3218 7.16724
R3567 VSS.n3200 VSS.n3199 7.16724
R3568 VSS.n3385 VSS.n3384 7.16724
R3569 VSS.n3275 VSS.n3274 7.16724
R3570 VSS.n2620 VSS.n2619 7.16134
R3571 VSS.n3461 VSS.n3460 7.15344
R3572 VSS.n3329 VSS.n113 7.15344
R3573 VSS.n2237 VSS.n2236 7.11268
R3574 VSS.n2790 VSS.n694 7.11268
R3575 VSS.n537 VSS.n533 6.98232
R3576 VSS.n2835 VSS.n2834 6.88949
R3577 VSS.n1351 VSS.n1311 6.88949
R3578 VSS.n1423 VSS.n772 6.62428
R3579 VSS.n2286 VSS.n1125 6.61527
R3580 VSS.n2739 VSS.n718 6.61527
R3581 VSS.n2382 VSS.t395 6.6005
R3582 VSS.n2382 VSS.t391 6.6005
R3583 VSS.n2384 VSS.t563 6.6005
R3584 VSS.n2384 VSS.t760 6.6005
R3585 VSS.n1017 VSS.t393 6.6005
R3586 VSS.n1017 VSS.t473 6.6005
R3587 VSS.n2219 VSS.n1125 6.57117
R3588 VSS.n2729 VSS.n718 6.57117
R3589 VSS.n1714 VSS.n1549 6.57117
R3590 VSS.n1716 VSS.n1714 6.57117
R3591 VSS.n803 VSS.n802 6.53477
R3592 VSS.n3449 VSS.n3448 6.50373
R3593 VSS.n3104 VSS.n209 6.50373
R3594 VSS.n3357 VSS.n3355 6.50373
R3595 VSS.n49 VSS.n48 6.4005
R3596 VSS.n3311 VSS.n3310 6.4005
R3597 VSS.n1939 VSS.n1936 6.4005
R3598 VSS.n1922 VSS.n1921 6.4005
R3599 VSS.n56 VSS.n55 6.26433
R3600 VSS.n3441 VSS.n3440 6.26433
R3601 VSS.n3304 VSS.n3303 6.26433
R3602 VSS.n103 VSS.n102 6.26433
R3603 VSS.n1442 VSS.n1441 6.26433
R3604 VSS.n1711 VSS.n1710 6.26433
R3605 VSS.n1846 VSS.n1842 6.26433
R3606 VSS.n1813 VSS.n1812 6.26433
R3607 VSS.n1792 VSS.n1791 6.26433
R3608 VSS.n2025 VSS.n2024 6.26433
R3609 VSS.n2002 VSS.n2001 6.26433
R3610 VSS.n2508 VSS.n2507 6.26433
R3611 VSS.n2494 VSS.n2493 6.26433
R3612 VSS.n2493 VSS.n2492 6.26433
R3613 VSS.n2463 VSS.n2462 6.26433
R3614 VSS.n2315 VSS.n2314 6.26433
R3615 VSS.n2315 VSS.n1035 6.26433
R3616 VSS.n3031 VSS.n3030 6.26433
R3617 VSS.n3030 VSS.n3029 6.26433
R3618 VSS.n890 VSS.n889 6.12816
R3619 VSS.n622 VSS.n621 6.06007
R3620 VSS.n315 VSS.n295 6.05269
R3621 VSS.n305 VSS.n301 6.05269
R3622 VSS.n326 VSS.n325 6.05269
R3623 VSS.n336 VSS.n332 6.05269
R3624 VSS.n380 VSS.n375 6.05269
R3625 VSS.n357 VSS.n352 6.05269
R3626 VSS.n364 VSS.n345 6.05269
R3627 VSS.n202 VSS.n201 6.05269
R3628 VSS.n2202 VSS.n2201 6.02861
R3629 VSS.n2118 VSS.n1217 6.02861
R3630 VSS.n2068 VSS.n2067 6.02861
R3631 VSS.n2904 VSS.n2903 6.02861
R3632 VSS.n2709 VSS.n2708 6.02861
R3633 VSS.n1476 VSS.n1474 6.02403
R3634 VSS.n1484 VSS.n1483 6.02403
R3635 VSS.n1666 VSS.n1578 5.98311
R3636 VSS.n1927 VSS.n1918 5.98311
R3637 VSS.n2544 VSS.n944 5.98311
R3638 VSS.n1744 VSS.n1741 5.98311
R3639 VSS.n2439 VSS.n2435 5.98311
R3640 VSS.n2355 VSS.n2351 5.98311
R3641 VSS.n1062 VSS.n1059 5.98311
R3642 VSS.n3039 VSS.n3038 5.98311
R3643 VSS.n244 VSS.n240 5.98311
R3644 VSS.n55 VSS.n42 5.85582
R3645 VSS.n3441 VSS.n40 5.85582
R3646 VSS.n32 VSS.n31 5.85582
R3647 VSS.n6 VSS.n3 5.85582
R3648 VSS.n10 VSS.n7 5.85582
R3649 VSS.n3305 VSS.n3304 5.85582
R3650 VSS.n103 VSS.n97 5.85582
R3651 VSS.n3319 VSS.n115 5.85582
R3652 VSS.n3321 VSS.n3320 5.85582
R3653 VSS.n3349 VSS.n3341 5.85582
R3654 VSS.n622 VSS.n610 5.85582
R3655 VSS.n1442 VSS.n1418 5.85582
R3656 VSS.n1717 VSS.n1541 5.85582
R3657 VSS.n891 VSS.n877 5.85582
R3658 VSS.n1842 VSS.n1290 5.85582
R3659 VSS.n961 VSS.n960 5.85582
R3660 VSS.n1813 VSS.n1763 5.85582
R3661 VSS.n1792 VSS.n1780 5.85582
R3662 VSS.n2025 VSS.n1225 5.85582
R3663 VSS.n2002 VSS.n1995 5.85582
R3664 VSS.n2509 VSS.n2508 5.85582
R3665 VSS.n2494 VSS.n2397 5.85582
R3666 VSS.n2463 VSS.n2416 5.85582
R3667 VSS.n2314 VSS.n1039 5.85582
R3668 VSS.n3031 VSS.n258 5.85582
R3669 VSS.n2492 VSS.n2399 5.65809
R3670 VSS.n2322 VSS.n1035 5.65809
R3671 VSS.n3029 VSS.n259 5.65809
R3672 VSS.n2217 VSS.n1153 5.63966
R3673 VSS.n2803 VSS.n2802 5.63966
R3674 VSS.n2791 VSS.n2790 5.63966
R3675 VSS.n2726 VSS.n730 5.63966
R3676 VSS.n2890 VSS.n581 5.5878
R3677 VSS.n2640 VSS.n774 5.55015
R3678 VSS.n2104 VSS.n2038 5.48621
R3679 VSS.n2081 VSS.n2058 5.48128
R3680 VSS.n962 VSS.n961 5.37524
R3681 VSS.n2594 VSS.n2593 5.27109
R3682 VSS.n1709 VSS.n1708 5.24958
R3683 VSS.n1174 VSS.n1172 5.13108
R3684 VSS.n1174 VSS.n1173 5.13108
R3685 VSS.n2172 VSS.n1175 5.13108
R3686 VSS.n2172 VSS.n2171 5.13108
R3687 VSS.n550 VSS.n548 5.13108
R3688 VSS.n550 VSS.n549 5.13108
R3689 VSS.n2143 VSS.n1185 5.13108
R3690 VSS.n2143 VSS.n1187 5.13108
R3691 VSS.n2142 VSS.n1188 5.13108
R3692 VSS.n2142 VSS.n1197 5.13108
R3693 VSS.n614 VSS.n612 5.13108
R3694 VSS.n614 VSS.n613 5.13108
R3695 VSS.n2845 VSS.n2842 5.13108
R3696 VSS.n2845 VSS.n2844 5.13108
R3697 VSS.n753 VSS.n751 5.13108
R3698 VSS.n753 VSS.n752 5.13108
R3699 VSS.n2679 VSS.n754 5.13108
R3700 VSS.n2679 VSS.n2678 5.13108
R3701 VSS.n1328 VSS.n1320 5.13108
R3702 VSS.n1328 VSS.n1321 5.13108
R3703 VSS.n808 VSS.n806 5.13108
R3704 VSS.n808 VSS.n807 5.13108
R3705 VSS.n1721 VSS.n1538 5.13108
R3706 VSS.n1721 VSS.n1540 5.13108
R3707 VSS.n886 VSS.n883 5.13108
R3708 VSS.n886 VSS.n884 5.13108
R3709 VSS.n1838 VSS.n1292 5.13108
R3710 VSS.n1838 VSS.n1837 5.13108
R3711 VSS.n969 VSS.n966 5.13108
R3712 VSS.n969 VSS.n967 5.13108
R3713 VSS.n2629 VSS.n780 4.92358
R3714 VSS.n2987 VSS.n492 4.89029
R3715 VSS.n2084 VSS.n2057 4.85762
R3716 VSS.n1702 VSS.n1555 4.85762
R3717 VSS.n2478 VSS.n2477 4.85762
R3718 VSS.n3023 VSS.n263 4.85762
R3719 VSS.n2326 VSS.n2325 4.85762
R3720 VSS.n1927 VSS.n1926 4.8005
R3721 VSS.n1745 VSS.n1744 4.8005
R3722 VSS.n2439 VSS.n2438 4.8005
R3723 VSS.n2355 VSS.n2354 4.8005
R3724 VSS.n1062 VSS.n1061 4.8005
R3725 VSS.n3038 VSS.n3037 4.8005
R3726 VSS.n245 VSS.n244 4.8005
R3727 VSS.n3448 VSS.n36 4.788
R3728 VSS.n209 VSS.n194 4.788
R3729 VSS.n3358 VSS.n3357 4.788
R3730 VSS.n2261 VSS.n2260 4.72533
R3731 VSS.n2760 VSS.n2759 4.72533
R3732 VSS.n2187 VSS.n2186 4.67352
R3733 VSS.n2206 VSS.n2205 4.67352
R3734 VSS.n2208 VSS.n2206 4.67352
R3735 VSS.n2212 VSS.n1155 4.67352
R3736 VSS.n2213 VSS.n2212 4.67352
R3737 VSS.n2276 VSS.n2275 4.67352
R3738 VSS.n2275 VSS.n1128 4.67352
R3739 VSS.n2271 VSS.n1128 4.67352
R3740 VSS.n2271 VSS.n2270 4.67352
R3741 VSS.n2268 VSS.n1130 4.67352
R3742 VSS.n2249 VSS.n1147 4.67352
R3743 VSS.n2249 VSS.n2248 4.67352
R3744 VSS.n2248 VSS.n2247 4.67352
R3745 VSS.n2247 VSS.n1148 4.67352
R3746 VSS.n2243 VSS.n2242 4.67352
R3747 VSS.n2229 VSS.n2228 4.67352
R3748 VSS.n2228 VSS.n517 4.67352
R3749 VSS.n2951 VSS.n517 4.67352
R3750 VSS.n2951 VSS.n2950 4.67352
R3751 VSS.n2950 VSS.n518 4.67352
R3752 VSS.n2946 VSS.n518 4.67352
R3753 VSS.n2944 VSS.n2943 4.67352
R3754 VSS.n2943 VSS.n520 4.67352
R3755 VSS.n2130 VSS.n1205 4.67352
R3756 VSS.n2116 VSS.n2115 4.67352
R3757 VSS.n2115 VSS.n1218 4.67352
R3758 VSS.n2111 VSS.n2110 4.67352
R3759 VSS.n2110 VSS.n2109 4.67352
R3760 VSS.n2077 VSS.n2076 4.67352
R3761 VSS.n2074 VSS.n2061 4.67352
R3762 VSS.n2070 VSS.n2061 4.67352
R3763 VSS.n2915 VSS.n575 4.67352
R3764 VSS.n2915 VSS.n2914 4.67352
R3765 VSS.n2900 VSS.n2899 4.67352
R3766 VSS.n2897 VSS.n579 4.67352
R3767 VSS.n2893 VSS.n579 4.67352
R3768 VSS.n2694 VSS.n2693 4.67352
R3769 VSS.n2713 VSS.n2712 4.67352
R3770 VSS.n2715 VSS.n2713 4.67352
R3771 VSS.n2719 VSS.n734 4.67352
R3772 VSS.n2720 VSS.n2719 4.67352
R3773 VSS.n2743 VSS.n714 4.67352
R3774 VSS.n2747 VSS.n714 4.67352
R3775 VSS.n2748 VSS.n2747 4.67352
R3776 VSS.n2749 VSS.n2748 4.67352
R3777 VSS.n2753 VSS.n2752 4.67352
R3778 VSS.n2763 VSS.n698 4.67352
R3779 VSS.n2777 VSS.n698 4.67352
R3780 VSS.n2778 VSS.n2777 4.67352
R3781 VSS.n2779 VSS.n2778 4.67352
R3782 VSS.n2783 VSS.n2782 4.67352
R3783 VSS.n2286 VSS.n1123 4.63943
R3784 VSS.n2260 VSS.n1133 4.63943
R3785 VSS.n2740 VSS.n2739 4.63943
R3786 VSS.n2761 VSS.n2760 4.63943
R3787 VSS.n887 VSS.n880 4.62124
R3788 VSS.n2460 VSS.n2419 4.62124
R3789 VSS.n2260 VSS.n2259 4.62124
R3790 VSS.n2801 VSS.n2794 4.62124
R3791 VSS.n2760 VSS.n709 4.62124
R3792 VSS.n1714 VSS.n1713 4.62124
R3793 VSS.n2219 VSS.n2217 4.6085
R3794 VSS.n2729 VSS.n730 4.6085
R3795 VSS.n2262 VSS.n2261 4.60638
R3796 VSS.n2759 VSS.n2758 4.60638
R3797 VSS.n473 VSS.n472 4.5578
R3798 VSS.n2278 VSS.n1123 4.55559
R3799 VSS.n1142 VSS.n1133 4.55559
R3800 VSS.n2741 VSS.n2740 4.55559
R3801 VSS.n2765 VSS.n2761 4.55559
R3802 VSS.n1460 VSS.n1459 4.51815
R3803 VSS.n1469 VSS.n1394 4.51815
R3804 VSS.n1680 VSS.n1679 4.51815
R3805 VSS.n1656 VSS.n1655 4.51815
R3806 VSS.n1915 VSS.n1914 4.51815
R3807 VSS.n1046 VSS.n1045 4.51401
R3808 VSS.n2320 VSS.n2319 4.51401
R3809 VSS.n247 VSS.n243 4.51401
R3810 VSS.n3043 VSS.n3042 4.51401
R3811 VSS.n2570 VSS.n927 4.51401
R3812 VSS.n932 VSS.n931 4.51401
R3813 VSS.n1064 VSS.n1057 4.51401
R3814 VSS.n1115 VSS.n1114 4.51401
R3815 VSS.n2578 VSS.n846 4.51401
R3816 VSS.n2582 VSS.n922 4.51401
R3817 VSS.n1085 VSS.n1081 4.51401
R3818 VSS.n2971 VSS.n2970 4.51401
R3819 VSS.n2961 VSS.n511 4.51401
R3820 VSS.n516 VSS.n515 4.51401
R3821 VSS.n2290 VSS.n1120 4.51401
R3822 VSS VSS.n2284 4.51401
R3823 VSS.n2194 VSS.n1165 4.51401
R3824 VSS.n2199 VSS.n2198 4.51401
R3825 VSS.n2163 VSS.n2153 4.51401
R3826 VSS.n2169 VSS.n2168 4.51401
R3827 VSS.n2930 VSS.n2929 4.51401
R3828 VSS.n565 VSS.n564 4.51401
R3829 VSS.n2258 VSS.n2257 4.51401
R3830 VSS.n2252 VSS.n2251 4.51401
R3831 VSS.n1207 VSS.n1203 4.51401
R3832 VSS.n2121 VSS.n2120 4.51401
R3833 VSS.n2147 VSS.n1182 4.51401
R3834 VSS.n1195 VSS.n1194 4.51401
R3835 VSS.n646 VSS.n645 4.51401
R3836 VSS.n640 VSS.n639 4.51401
R3837 VSS.n587 VSS.n586 4.51401
R3838 VSS.n667 VSS.n666 4.51401
R3839 VSS.n2045 VSS.n2041 4.51401
R3840 VSS.n2089 VSS.n2088 4.51401
R3841 VSS.n2919 VSS.n572 4.51401
R3842 VSS.n2910 VSS.n2906 4.51401
R3843 VSS.n2701 VSS.n744 4.51401
R3844 VSS.n2706 VSS.n2705 4.51401
R3845 VSS.n2671 VSS.n2661 4.51401
R3846 VSS.n2676 VSS.n2675 4.51401
R3847 VSS.n2867 VSS.n674 4.51401
R3848 VSS.n2860 VSS.n2859 4.51401
R3849 VSS.n2797 VSS.n2795 4.51401
R3850 VSS.n2811 VSS.n2810 4.51401
R3851 VSS.n2733 VSS.n725 4.51401
R3852 VSS VSS.n2737 4.51401
R3853 VSS.n2769 VSS.n704 4.51401
R3854 VSS.n2774 VSS.n2773 4.51401
R3855 VSS.n1327 VSS.n1326 4.51401
R3856 VSS.n1336 VSS.n1335 4.51401
R3857 VSS.n2616 VSS.n2615 4.51401
R3858 VSS.n823 VSS.n822 4.51401
R3859 VSS.n2651 VSS.n765 4.51401
R3860 VSS.n770 VSS.n769 4.51401
R3861 VSS.n1383 VSS.n1381 4.51401
R3862 VSS.n1487 VSS 4.51401
R3863 VSS.n1527 VSS.n1301 4.51401
R3864 VSS.n1306 VSS.n1305 4.51401
R3865 VSS.n1407 VSS.n1399 4.51401
R3866 VSS.n1452 VSS.n1451 4.51401
R3867 VSS.n1257 VSS.n1250 4.51401
R3868 VSS.n1950 VSS.n1949 4.51401
R3869 VSS.n2523 VSS.n986 4.51401
R3870 VSS.n2514 VSS.n2513 4.51401
R3871 VSS.n1616 VSS.n1613 4.51401
R3872 VSS.n2605 VSS.n2604 4.51401
R3873 VSS.n1562 VSS.n1557 4.51401
R3874 VSS.n1684 VSS.n1683 4.51401
R3875 VSS.n1725 VSS.n1535 4.51401
R3876 VSS.n1548 VSS.n1547 4.51401
R3877 VSS.n866 VSS.n864 4.51401
R3878 VSS.n894 VSS.n893 4.51401
R3879 VSS.n1590 VSS.n1588 4.51401
R3880 VSS.n1645 VSS.n1644 4.51401
R3881 VSS.n1230 VSS.n1226 4.51401
R3882 VSS.n2015 VSS.n2014 4.51401
R3883 VSS.n1910 VSS.n1909 4.51401
R3884 VSS.n1982 VSS.n1981 4.51401
R3885 VSS.n1836 VSS.n1835 4.51401
R3886 VSS.n1735 VSS.n1291 4.51401
R3887 VSS.n951 VSS.n949 4.51401
R3888 VSS.n980 VSS.n979 4.51401
R3889 VSS.n1874 VSS.n1280 4.51401
R3890 VSS.n1879 VSS.n1878 4.51401
R3891 VSS.n1769 VSS.n1766 4.51401
R3892 VSS.n1795 VSS.n1794 4.51401
R3893 VSS.n1747 VSS.n1743 4.51401
R3894 VSS.n1827 VSS.n1826 4.51401
R3895 VSS.n2427 VSS.n2424 4.51401
R3896 VSS.n2452 VSS.n2451 4.51401
R3897 VSS.n2402 VSS.n2400 4.51401
R3898 VSS.n2483 VSS.n2482 4.51401
R3899 VSS.n2374 VSS.n1024 4.51401
R3900 VSS.n2367 VSS.n1022 4.51401
R3901 VSS.n3017 VSS.n3016 4.51401
R3902 VSS.n3006 VSS.n3005 4.51401
R3903 VSS.n3448 VSS.n3447 4.50726
R3904 VSS.n3174 VSS.n209 4.50726
R3905 VSS.n3357 VSS.n3356 4.50726
R3906 VSS.n534 VSS.n528 4.5005
R3907 VSS.n542 VSS.n541 4.5005
R3908 VSS.n543 VSS.n532 4.5005
R3909 VSS.n2162 VSS.n2161 4.5005
R3910 VSS.n2159 VSS.n2158 4.5005
R3911 VSS.n2155 VSS.n1176 4.5005
R3912 VSS.n2193 VSS.n2192 4.5005
R3913 VSS.n2191 VSS.n2190 4.5005
R3914 VSS.n1160 VSS.n1159 4.5005
R3915 VSS.n2289 VSS.n2288 4.5005
R3916 VSS.n2280 VSS.n1122 4.5005
R3917 VSS.n2283 VSS.n1126 4.5005
R3918 VSS.n2960 VSS.n2959 4.5005
R3919 VSS.n2958 VSS.n2957 4.5005
R3920 VSS.n2954 VSS.n2953 4.5005
R3921 VSS.n1141 VSS.n1134 4.5005
R3922 VSS.n1145 VSS.n1144 4.5005
R3923 VSS.n1138 VSS.n1137 4.5005
R3924 VSS.n2051 VSS.n2049 4.5005
R3925 VSS.n2879 VSS.n2878 4.5005
R3926 VSS.n592 VSS.n588 4.5005
R3927 VSS.n594 VSS.n591 4.5005
R3928 VSS.n630 VSS.n606 4.5005
R3929 VSS.n633 VSS.n632 4.5005
R3930 VSS.n634 VSS.n609 4.5005
R3931 VSS.n2146 VSS.n2145 4.5005
R3932 VSS.n1189 VSS.n1184 4.5005
R3933 VSS.n1193 VSS.n1192 4.5005
R3934 VSS.n2128 VSS.n2127 4.5005
R3935 VSS.n1208 VSS.n1206 4.5005
R3936 VSS.n1213 VSS.n1211 4.5005
R3937 VSS.n2096 VSS.n2095 4.5005
R3938 VSS.n2050 VSS.n2046 4.5005
R3939 VSS.n2918 VSS.n2917 4.5005
R3940 VSS.n2907 VSS.n574 4.5005
R3941 VSS.n2912 VSS.n2911 4.5005
R3942 VSS.n720 VSS.n719 4.5005
R3943 VSS.n2799 VSS.n2798 4.5005
R3944 VSS.n2806 VSS.n2805 4.5005
R3945 VSS.n689 VSS.n686 4.5005
R3946 VSS.n2866 VSS.n2865 4.5005
R3947 VSS.n2855 VSS.n677 4.5005
R3948 VSS.n2858 VSS.n2838 4.5005
R3949 VSS.n2670 VSS.n2669 4.5005
R3950 VSS.n2667 VSS.n2666 4.5005
R3951 VSS.n2663 VSS.n755 4.5005
R3952 VSS.n2700 VSS.n2699 4.5005
R3953 VSS.n2698 VSS.n2697 4.5005
R3954 VSS.n739 VSS.n738 4.5005
R3955 VSS.n2732 VSS.n2731 4.5005
R3956 VSS.n728 VSS.n727 4.5005
R3957 VSS.n2768 VSS.n2767 4.5005
R3958 VSS.n708 VSS.n707 4.5005
R3959 VSS.n700 VSS.n699 4.5005
R3960 VSS.n1382 VSS.n1375 4.5005
R3961 VSS.n1492 VSS.n1491 4.5005
R3962 VSS.n1378 VSS.n1376 4.5005
R3963 VSS.n2650 VSS.n2649 4.5005
R3964 VSS.n2648 VSS.n2647 4.5005
R3965 VSS.n2644 VSS.n2643 4.5005
R3966 VSS.n794 VSS.n787 4.5005
R3967 VSS.n799 VSS.n798 4.5005
R3968 VSS.n795 VSS.n790 4.5005
R3969 VSS.n1323 VSS.n1322 4.5005
R3970 VSS.n1331 VSS.n1330 4.5005
R3971 VSS.n1319 VSS.n1315 4.5005
R3972 VSS.n1526 VSS.n1525 4.5005
R3973 VSS.n1524 VSS.n1523 4.5005
R3974 VSS.n1520 VSS.n1519 4.5005
R3975 VSS.n1406 VSS.n1402 4.5005
R3976 VSS.n1457 VSS.n1456 4.5005
R3977 VSS.n1410 VSS.n1405 4.5005
R3978 VSS.n871 VSS.n869 4.5005
R3979 VSS.n1724 VSS.n1723 4.5005
R3980 VSS.n1542 VSS.n1537 4.5005
R3981 VSS.n1546 VSS.n1545 4.5005
R3982 VSS.n1691 VSS.n1690 4.5005
R3983 VSS.n1563 VSS.n1561 4.5005
R3984 VSS.n1568 VSS.n1565 4.5005
R3985 VSS.n1617 VSS.n1614 4.5005
R3986 VSS.n1622 VSS.n1621 4.5005
R3987 VSS.n833 VSS.n832 4.5005
R3988 VSS.n2577 VSS.n2576 4.5005
R3989 VSS.n2574 VSS.n849 4.5005
R3990 VSS.n2584 VSS.n2583 4.5005
R3991 VSS.n901 VSS.n900 4.5005
R3992 VSS.n870 VSS.n867 4.5005
R3993 VSS.n1652 VSS.n1651 4.5005
R3994 VSS.n1594 VSS.n1591 4.5005
R3995 VSS.n1595 VSS.n1593 4.5005
R3996 VSS.n957 VSS.n955 4.5005
R3997 VSS.n1296 VSS.n1295 4.5005
R3998 VSS.n1731 VSS.n1730 4.5005
R3999 VSS.n1734 VSS.n1733 4.5005
R4000 VSS.n1908 VSS.n1907 4.5005
R4001 VSS.n1903 VSS.n1902 4.5005
R4002 VSS.n1900 VSS.n1237 4.5005
R4003 VSS.n1256 VSS.n1252 4.5005
R4004 VSS.n1955 VSS.n1954 4.5005
R4005 VSS.n1260 VSS.n1255 4.5005
R4006 VSS.n2569 VSS.n2568 4.5005
R4007 VSS.n2567 VSS.n2566 4.5005
R4008 VSS.n2563 VSS.n2562 4.5005
R4009 VSS.n2536 VSS.n2535 4.5005
R4010 VSS.n956 VSS.n952 4.5005
R4011 VSS.n1873 VSS.n1872 4.5005
R4012 VSS.n1871 VSS.n1870 4.5005
R4013 VSS.n1283 VSS.n1275 4.5005
R4014 VSS.n2430 VSS.n2423 4.5005
R4015 VSS.n1749 VSS.n1748 4.5005
R4016 VSS.n1754 VSS.n1753 4.5005
R4017 VSS.n1755 VSS.n1740 4.5005
R4018 VSS.n1802 VSS.n1801 4.5005
R4019 VSS.n1774 VSS.n1770 4.5005
R4020 VSS.n1776 VSS.n1773 4.5005
R4021 VSS.n2022 VSS.n2021 4.5005
R4022 VSS.n1988 VSS.n1231 4.5005
R4023 VSS.n1989 VSS.n1987 4.5005
R4024 VSS.n2522 VSS.n2521 4.5005
R4025 VSS.n992 VSS.n988 4.5005
R4026 VSS.n2516 VSS.n2515 4.5005
R4027 VSS.n2426 VSS.n2425 4.5005
R4028 VSS.n2457 VSS.n2456 4.5005
R4029 VSS.n2490 VSS.n2489 4.5005
R4030 VSS.n2403 VSS.n2401 4.5005
R4031 VSS.n2408 VSS.n2406 4.5005
R4032 VSS.n2347 VSS.n2346 4.5005
R4033 VSS.n249 VSS.n248 4.5005
R4034 VSS.n252 VSS.n251 4.5005
R4035 VSS.n253 VSS.n238 4.5005
R4036 VSS.n1067 VSS.n1066 4.5005
R4037 VSS.n1072 VSS.n1071 4.5005
R4038 VSS.n1056 VSS.n1052 4.5005
R4039 VSS.n1086 VSS.n1083 4.5005
R4040 VSS.n1090 VSS.n1089 4.5005
R4041 VSS.n501 VSS.n500 4.5005
R4042 VSS.n2312 VSS.n2311 4.5005
R4043 VSS.n1047 VSS.n1038 4.5005
R4044 VSS.n2318 VSS.n2317 4.5005
R4045 VSS.n2373 VSS.n2372 4.5005
R4046 VSS.n1027 VSS.n1026 4.5005
R4047 VSS.n269 VSS.n266 4.5005
R4048 VSS.n3012 VSS.n3011 4.5005
R4049 VSS.n3002 VSS.n270 4.5005
R4050 VSS.n2389 VSS.n2388 4.4805
R4051 VSS.n2543 VSS.n2542 4.38311
R4052 VSS.n2186 VSS.n2185 4.36875
R4053 VSS.n2187 VSS.n1158 4.36875
R4054 VSS.n2205 VSS.n1157 4.36875
R4055 VSS.n2214 VSS.n2213 4.36875
R4056 VSS.n2277 VSS.n2276 4.36875
R4057 VSS.n2264 VSS.n2263 4.36875
R4058 VSS.n1147 VSS.n1140 4.36875
R4059 VSS.n2240 VSS.n1151 4.36875
R4060 VSS.n2229 VSS.n2227 4.36875
R4061 VSS.n521 VSS.n520 4.36875
R4062 VSS.n2131 VSS.n2130 4.36875
R4063 VSS.n1216 VSS.n1205 4.36875
R4064 VSS.n2117 VSS.n2116 4.36875
R4065 VSS.n2109 VSS.n1221 4.36875
R4066 VSS.n2077 VSS.n2060 4.36875
R4067 VSS.n2070 VSS.n2069 4.36875
R4068 VSS.n2914 VSS.n576 4.36875
R4069 VSS.n2900 VSS.n577 4.36875
R4070 VSS.n2893 VSS.n2892 4.36875
R4071 VSS.n2693 VSS.n2692 4.36875
R4072 VSS.n2694 VSS.n737 4.36875
R4073 VSS.n2712 VSS.n736 4.36875
R4074 VSS.n2721 VSS.n2720 4.36875
R4075 VSS.n2743 VSS.n2742 4.36875
R4076 VSS.n2755 VSS.n710 4.36875
R4077 VSS.n2764 VSS.n2763 4.36875
R4078 VSS.n2786 VSS.n2785 4.36875
R4079 VSS.n1717 VSS.n1716 4.28986
R4080 VSS.n1711 VSS.n1549 4.28986
R4081 VSS.n889 VSS.n888 4.28986
R4082 VSS.n1791 VSS.n1790 4.28986
R4083 VSS.n2024 VSS.n1228 4.28986
R4084 VSS.n2001 VSS.n2000 4.28986
R4085 VSS.n2462 VSS.n2461 4.28986
R4086 VSS.n1693 VSS.n1560 4.14168
R4087 VSS.n2818 VSS.n2817 4.11798
R4088 VSS.n2817 VSS.n682 4.11798
R4089 VSS.n2636 VSS.n2635 4.11798
R4090 VSS.n1354 VSS.n1353 4.11798
R4091 VSS.n1353 VSS.n1308 4.11798
R4092 VSS.n1503 VSS.n1502 4.11798
R4093 VSS.n1502 VSS.n1501 4.11798
R4094 VSS.n1957 VSS.n1251 4.11798
R4095 VSS.n2349 VSS.n2345 4.11798
R4096 VSS.n2364 VSS.n2349 4.11798
R4097 VSS.n2976 VSS.n497 4.11798
R4098 VSS.n2979 VSS.n497 4.11798
R4099 VSS.n1105 VSS.n1104 4.11798
R4100 VSS.n1104 VSS.n1103 4.11798
R4101 VSS.n2997 VSS.n275 4.11798
R4102 VSS.n2994 VSS.n275 4.11798
R4103 VSS.n2801 VSS.n691 4.09013
R4104 VSS.n888 VSS.n887 4.07323
R4105 VSS.n1790 VSS.n1789 4.07323
R4106 VSS.n2012 VSS.n1228 4.07323
R4107 VSS.n2000 VSS.n1999 4.07323
R4108 VSS.n2461 VSS.n2460 4.07323
R4109 VSS.n562 VSS.n561 4.03876
R4110 VSS.n820 VSS.n819 4.03876
R4111 VSS.n3053 VSS 4.02175
R4112 VSS.n230 VSS 4.02175
R4113 VSS.n3382 VSS 4.02175
R4114 VSS.n231 VSS 4.02175
R4115 VSS.n2223 VSS.n1152 3.97459
R4116 VSS.n2725 VSS.n732 3.97459
R4117 VSS.n2177 VSS.n2176 3.96548
R4118 VSS.n2180 VSS.n2177 3.96548
R4119 VSS.n557 VSS.n556 3.96548
R4120 VSS.n2138 VSS.n2137 3.96548
R4121 VSS.n2137 VSS.n2136 3.96548
R4122 VSS.n2885 VSS.n2884 3.96548
R4123 VSS.n2863 VSS.n2862 3.96548
R4124 VSS.n2862 VSS.n2837 3.96548
R4125 VSS.n2852 VSS.n2851 3.96548
R4126 VSS.n2684 VSS.n2683 3.96548
R4127 VSS.n2687 VSS.n2684 3.96548
R4128 VSS.n815 VSS.n814 3.96548
R4129 VSS.n1345 VSS.n1344 3.96548
R4130 VSS.n1347 VSS.n1345 3.96548
R4131 VSS.n841 VSS.n839 3.90948
R4132 VSS.n841 VSS.n840 3.90948
R4133 VSS.n390 VSS.n389 3.78485
R4134 VSS.n3241 VSS.n3239 3.78485
R4135 VSS.n3271 VSS.n3260 3.78485
R4136 VSS.n3223 VSS.n3222 3.78485
R4137 VSS.n3218 VSS.n3217 3.78485
R4138 VSS.n3199 VSS.n182 3.78485
R4139 VSS.n3385 VSS.n77 3.78485
R4140 VSS.n3275 VSS.n3255 3.78485
R4141 VSS.n2634 VSS.n2633 3.75994
R4142 VSS.n412 VSS.n409 3.75517
R4143 VSS.n2176 VSS.n1171 3.7069
R4144 VSS.n557 VSS.n546 3.7069
R4145 VSS.n2138 VSS.n1198 3.7069
R4146 VSS.n2885 VSS.n582 3.7069
R4147 VSS.n2100 VSS.n2039 3.7069
R4148 VSS.n2100 VSS.n2099 3.7069
R4149 VSS.n2863 VSS.n2836 3.7069
R4150 VSS.n2849 VSS.n2841 3.7069
R4151 VSS.n2683 VSS.n750 3.7069
R4152 VSS.n815 VSS.n804 3.7069
R4153 VSS.n1344 VSS.n1313 3.7069
R4154 VSS.n1347 VSS.n1346 3.7069
R4155 VSS.n1705 VSS.n1552 3.50735
R4156 VSS.n2476 VSS.n2475 3.50735
R4157 VSS.n2324 VSS.n2323 3.50735
R4158 VSS.n3025 VSS.n261 3.50735
R4159 VSS.n490 VSS.n401 3.46461
R4160 VSS.n422 VSS.n401 3.46461
R4161 VSS.t551 VSS.t371 3.46461
R4162 VSS.t551 VSS.t457 3.46461
R4163 VSS.n424 VSS.n420 3.46461
R4164 VSS.n469 VSS.n424 3.46461
R4165 VSS.n977 VSS.n976 3.44377
R4166 VSS.n976 VSS.n975 3.44377
R4167 VSS.n931 VSS.n924 3.43925
R4168 VSS.n2571 VSS.n2570 3.43925
R4169 VSS.n2582 VSS.n2581 3.43925
R4170 VSS.n2579 VSS.n2578 3.43925
R4171 VSS.n515 VSS.n508 3.43925
R4172 VSS.n2962 VSS.n2961 3.43925
R4173 VSS.n2284 VSS.n1117 3.43925
R4174 VSS.n2291 VSS.n2290 3.43925
R4175 VSS.n2198 VSS.n2197 3.43925
R4176 VSS.n2195 VSS.n2194 3.43925
R4177 VSS.n566 VSS.n565 3.43925
R4178 VSS.n2929 VSS.n2928 3.43925
R4179 VSS.n2253 VSS.n2252 3.43925
R4180 VSS.n2257 VSS.n2256 3.43925
R4181 VSS.n2122 VSS.n2121 3.43925
R4182 VSS.n2124 VSS.n1207 3.43925
R4183 VSS.n1194 VSS.n1180 3.43925
R4184 VSS.n2148 VSS.n2147 3.43925
R4185 VSS.n641 VSS.n640 3.43925
R4186 VSS.n645 VSS.n644 3.43925
R4187 VSS.n668 VSS.n667 3.43925
R4188 VSS.n2875 VSS.n587 3.43925
R4189 VSS.n2090 VSS.n2089 3.43925
R4190 VSS.n2092 VSS.n2045 3.43925
R4191 VSS.n2910 VSS.n569 3.43925
R4192 VSS.n2920 VSS.n2919 3.43925
R4193 VSS.n2705 VSS.n2704 3.43925
R4194 VSS.n2702 VSS.n2701 3.43925
R4195 VSS.n2675 VSS.n2674 3.43925
R4196 VSS.n2672 VSS.n2671 3.43925
R4197 VSS.n2859 VSS.n671 3.43925
R4198 VSS.n2868 VSS.n2867 3.43925
R4199 VSS.n2810 VSS.n2809 3.43925
R4200 VSS.n2797 VSS.n2796 3.43925
R4201 VSS.n2737 VSS.n2736 3.43925
R4202 VSS.n2734 VSS.n2733 3.43925
R4203 VSS.n2773 VSS.n2772 3.43925
R4204 VSS.n2770 VSS.n2769 3.43925
R4205 VSS.n824 VSS.n823 3.43925
R4206 VSS.n2615 VSS.n2614 3.43925
R4207 VSS.n769 VSS.n762 3.43925
R4208 VSS.n2652 VSS.n2651 3.43925
R4209 VSS.n1488 VSS.n1487 3.43925
R4210 VSS.n1384 VSS.n1383 3.43925
R4211 VSS.n1305 VSS.n1299 3.43925
R4212 VSS.n1528 VSS.n1527 3.43925
R4213 VSS.n1453 VSS.n1452 3.43925
R4214 VSS.n1408 VSS.n1407 3.43925
R4215 VSS.n1951 VSS.n1950 3.43925
R4216 VSS.n1258 VSS.n1257 3.43925
R4217 VSS.n2514 VSS.n984 3.43925
R4218 VSS.n2524 VSS.n2523 3.43925
R4219 VSS.n1685 VSS.n1684 3.43925
R4220 VSS.n1687 VSS.n1562 3.43925
R4221 VSS.n1547 VSS.n1533 3.43925
R4222 VSS.n1726 VSS.n1725 3.43925
R4223 VSS.n895 VSS.n894 3.43925
R4224 VSS.n897 VSS.n866 3.43925
R4225 VSS.n1646 VSS.n1645 3.43925
R4226 VSS.n1648 VSS.n1590 3.43925
R4227 VSS.n2016 VSS.n2015 3.43925
R4228 VSS.n2018 VSS.n1230 3.43925
R4229 VSS.n981 VSS.n980 3.43925
R4230 VSS.n2532 VSS.n951 3.43925
R4231 VSS.n1878 VSS.n1877 3.43925
R4232 VSS.n1875 VSS.n1874 3.43925
R4233 VSS.n1796 VSS.n1795 3.43925
R4234 VSS.n1798 VSS.n1769 3.43925
R4235 VSS.n2453 VSS.n2452 3.43925
R4236 VSS.n2428 VSS.n2427 3.43925
R4237 VSS.n2484 VSS.n2483 3.43925
R4238 VSS.n2486 VSS.n2402 3.43925
R4239 VSS.n3044 VSS.n3043 3.41839
R4240 VSS.n243 VSS.n242 3.41839
R4241 VSS.n3005 VSS.n3004 3.41636
R4242 VSS.n3016 VSS.n3015 3.41636
R4243 VSS.n1116 VSS.n1115 3.41624
R4244 VSS.n1057 VSS.n1050 3.41624
R4245 VSS.n2970 VSS.n2969 3.41605
R4246 VSS.n1085 VSS.n503 3.41605
R4247 VSS.n2168 VSS.n2167 3.41514
R4248 VSS.n1335 VSS.n1334 3.41514
R4249 VSS.n1736 VSS.n1735 3.41514
R4250 VSS.n250 VSS.n235 3.4105
R4251 VSS.n3045 VSS.n236 3.4105
R4252 VSS.n928 VSS.n926 3.4105
R4253 VSS.n2565 VSS.n2564 3.4105
R4254 VSS.n1069 VSS.n1068 3.4105
R4255 VSS.n1070 VSS.n1051 3.4105
R4256 VSS.n2575 VSS.n2573 3.4105
R4257 VSS.n923 VSS.n851 3.4105
R4258 VSS.n1087 VSS.n1048 3.4105
R4259 VSS.n1088 VSS.n502 3.4105
R4260 VSS.n512 VSS.n510 3.4105
R4261 VSS.n2956 VSS.n2955 3.4105
R4262 VSS.n1121 VSS.n1119 3.4105
R4263 VSS.n2282 VSS.n2281 3.4105
R4264 VSS.n1166 VSS.n1164 3.4105
R4265 VSS.n2189 VSS.n1161 3.4105
R4266 VSS.n2164 VSS.n2163 3.4105
R4267 VSS.n2154 VSS.n2152 3.4105
R4268 VSS.n2157 VSS.n1177 3.4105
R4269 VSS.n539 VSS.n529 3.4105
R4270 VSS.n540 VSS.n531 3.4105
R4271 VSS.n2255 VSS.n1135 3.4105
R4272 VSS.n2254 VSS.n1136 3.4105
R4273 VSS.n2126 VSS.n2125 3.4105
R4274 VSS.n1210 VSS.n1209 3.4105
R4275 VSS.n1183 VSS.n1181 3.4105
R4276 VSS.n1191 VSS.n1190 3.4105
R4277 VSS.n643 VSS.n607 3.4105
R4278 VSS.n642 VSS.n608 3.4105
R4279 VSS.n2877 VSS.n2876 3.4105
R4280 VSS.n590 VSS.n589 3.4105
R4281 VSS.n2094 VSS.n2093 3.4105
R4282 VSS.n2048 VSS.n2047 3.4105
R4283 VSS.n573 VSS.n571 3.4105
R4284 VSS.n2909 VSS.n2908 3.4105
R4285 VSS.n745 VSS.n743 3.4105
R4286 VSS.n2696 VSS.n740 3.4105
R4287 VSS.n2662 VSS.n2660 3.4105
R4288 VSS.n2665 VSS.n756 3.4105
R4289 VSS.n675 VSS.n673 3.4105
R4290 VSS.n2857 VSS.n2856 3.4105
R4291 VSS.n688 VSS.n687 3.4105
R4292 VSS.n2808 VSS.n2807 3.4105
R4293 VSS.n729 VSS.n724 3.4105
R4294 VSS.n726 VSS.n721 3.4105
R4295 VSS.n705 VSS.n703 3.4105
R4296 VSS.n706 VSS.n701 3.4105
R4297 VSS.n1326 VSS.n1325 3.4105
R4298 VSS.n1317 VSS.n1316 3.4105
R4299 VSS.n1333 VSS.n1332 3.4105
R4300 VSS.n796 VSS.n788 3.4105
R4301 VSS.n797 VSS.n789 3.4105
R4302 VSS.n766 VSS.n764 3.4105
R4303 VSS.n2646 VSS.n2645 3.4105
R4304 VSS.n1379 VSS.n1377 3.4105
R4305 VSS.n1490 VSS.n1489 3.4105
R4306 VSS.n1302 VSS.n1300 3.4105
R4307 VSS.n1522 VSS.n1521 3.4105
R4308 VSS.n1409 VSS.n1404 3.4105
R4309 VSS.n1455 VSS.n1454 3.4105
R4310 VSS.n1259 VSS.n1254 3.4105
R4311 VSS.n1953 VSS.n1952 3.4105
R4312 VSS.n987 VSS.n985 3.4105
R4313 VSS.n994 VSS.n993 3.4105
R4314 VSS.n2607 VSS.n2606 3.4105
R4315 VSS.n2607 VSS.n829 3.4105
R4316 VSS.n2606 VSS.n2605 3.4105
R4317 VSS.n1616 VSS.n829 3.4105
R4318 VSS.n1619 VSS.n1618 3.4105
R4319 VSS.n1620 VSS.n831 3.4105
R4320 VSS.n1689 VSS.n1688 3.4105
R4321 VSS.n1686 VSS.n1564 3.4105
R4322 VSS.n1536 VSS.n1534 3.4105
R4323 VSS.n1544 VSS.n1543 3.4105
R4324 VSS.n899 VSS.n898 3.4105
R4325 VSS.n896 VSS.n868 3.4105
R4326 VSS.n1650 VSS.n1649 3.4105
R4327 VSS.n1647 VSS.n1592 3.4105
R4328 VSS.n2020 VSS.n2019 3.4105
R4329 VSS.n1986 VSS.n1232 3.4105
R4330 VSS.n1984 VSS.n1983 3.4105
R4331 VSS.n1984 VSS.n1235 3.4105
R4332 VSS.n1983 VSS.n1982 3.4105
R4333 VSS.n1909 VSS.n1235 3.4105
R4334 VSS.n1899 VSS.n1898 3.4105
R4335 VSS.n1901 VSS.n1236 3.4105
R4336 VSS.n1835 VSS.n1834 3.4105
R4337 VSS.n1729 VSS.n1298 3.4105
R4338 VSS.n1732 VSS.n1728 3.4105
R4339 VSS.n2534 VSS.n2533 3.4105
R4340 VSS.n954 VSS.n953 3.4105
R4341 VSS.n1281 VSS.n1279 3.4105
R4342 VSS.n1869 VSS.n1276 3.4105
R4343 VSS.n1800 VSS.n1799 3.4105
R4344 VSS.n1772 VSS.n1771 3.4105
R4345 VSS.n1829 VSS.n1828 3.4105
R4346 VSS.n1829 VSS.n1738 3.4105
R4347 VSS.n1828 VSS.n1827 3.4105
R4348 VSS.n1743 VSS.n1738 3.4105
R4349 VSS.n1751 VSS.n1750 3.4105
R4350 VSS.n1752 VSS.n1739 3.4105
R4351 VSS.n2429 VSS.n2422 3.4105
R4352 VSS.n2455 VSS.n2454 3.4105
R4353 VSS.n2488 VSS.n2487 3.4105
R4354 VSS.n2405 VSS.n2404 3.4105
R4355 VSS.n2375 VSS.n2374 3.4105
R4356 VSS.n3014 VSS.n3013 3.4105
R4357 VSS.n3003 VSS.n268 3.4105
R4358 VSS.n2319 VSS.n1019 3.4105
R4359 VSS.n2305 VSS.n1046 3.4105
R4360 VSS.n2310 VSS.n2309 3.4105
R4361 VSS.n2308 VSS.n1037 3.4105
R4362 VSS.n2375 VSS.n1022 3.4105
R4363 VSS.n2375 VSS.n1021 3.4105
R4364 VSS.n2375 VSS.n1020 3.4105
R4365 VSS.n30 VSS.n29 3.40476
R4366 VSS.n3348 VSS.n3347 3.40476
R4367 VSS.n780 VSS.n777 3.31239
R4368 VSS.n1263 VSS.n1251 3.22288
R4369 VSS.n977 VSS.n963 3.21921
R4370 VSS.n972 VSS.n971 3.21921
R4371 VSS.n1703 VSS.n1554 3.2005
R4372 VSS.n2480 VSS.n2411 3.2005
R4373 VSS.n2328 VSS.n1034 3.2005
R4374 VSS.n3024 VSS.n262 3.2005
R4375 VSS.n57 VSS.n56 3.13241
R4376 VSS.n3440 VSS.n3436 3.13241
R4377 VSS.n29 VSS.n25 3.13241
R4378 VSS.n10 VSS.n9 3.13241
R4379 VSS.n3303 VSS.n3302 3.13241
R4380 VSS.n102 VSS.n98 3.13241
R4381 VSS.n3322 VSS.n3321 3.13241
R4382 VSS.n3347 VSS.n3346 3.13241
R4383 VSS.n620 VSS.n619 3.13241
R4384 VSS.n1441 VSS.n1440 3.13241
R4385 VSS.n1812 VSS.n1811 3.13241
R4386 VSS.n2507 VSS.n996 3.13241
R4387 VSS.n1016 VSS.n1015 3.1005
R4388 VSS.n2043 VSS.n2042 3.09945
R4389 VSS.n2215 VSS.n1152 3.05276
R4390 VSS.n2722 VSS.n732 3.05276
R4391 VSS.n551 VSS.n550 3.04861
R4392 VSS.n2172 VSS.n2170 3.04861
R4393 VSS.n615 VSS.n614 3.04861
R4394 VSS.n2142 VSS.n1196 3.04861
R4395 VSS.n2845 VSS.n2843 3.04861
R4396 VSS.n2679 VSS.n2677 3.04861
R4397 VSS.n809 VSS.n808 3.04861
R4398 VSS.n886 VSS.n885 3.04861
R4399 VSS.n969 VSS.n968 3.04861
R4400 VSS.n1789 VSS.n1782 3.04861
R4401 VSS.n1999 VSS.n1998 3.04861
R4402 VSS.n1892 VSS.n1889 3.01226
R4403 VSS.n1666 VSS.n1665 2.92224
R4404 VSS.n2802 VSS.n2801 2.92166
R4405 VSS.n3468 VSS.n3467 2.90519
R4406 VSS.n3071 VSS.t298 2.89674
R4407 VSS.n2180 VSS.n2179 2.88804
R4408 VSS.n2136 VSS.n1201 2.88804
R4409 VSS.n2687 VSS.n2686 2.88804
R4410 VSS.n3134 VSS.n3133 2.88636
R4411 VSS.n31 VSS.n30 2.86007
R4412 VSS.n3349 VSS.n3348 2.86007
R4413 VSS.n2179 VSS.n2178 2.79323
R4414 VSS.n1201 VSS.n1200 2.79323
R4415 VSS.n2686 VSS.n2685 2.79323
R4416 VSS.n561 VSS.n560 2.77203
R4417 VSS.n819 VSS.n818 2.77203
R4418 VSS.n58 VSS.n57 2.7239
R4419 VSS.n3437 VSS.n3436 2.7239
R4420 VSS.n26 VSS.n25 2.7239
R4421 VSS.n9 VSS.n8 2.7239
R4422 VSS.n3302 VSS.n81 2.7239
R4423 VSS.n99 VSS.n98 2.7239
R4424 VSS.n3323 VSS.n3322 2.7239
R4425 VSS.n3346 VSS.n3345 2.7239
R4426 VSS.n619 VSS.n618 2.7239
R4427 VSS.n1440 VSS.n1439 2.7239
R4428 VSS.n1844 VSS.n1843 2.7239
R4429 VSS.n1811 VSS.n1810 2.7239
R4430 VSS.n997 VSS.n996 2.7239
R4431 VSS.n2637 VSS.n774 2.68581
R4432 VSS.n3467 VSS.n3466 2.63717
R4433 VSS.n3298 VSS.n3297 2.63717
R4434 VSS.n1701 VSS.n1700 2.63064
R4435 VSS.n2479 VSS.n2474 2.63064
R4436 VSS.n2327 VSS.n1032 2.63064
R4437 VSS.n3022 VSS.n3021 2.63064
R4438 VSS.n3408 VSS.n3407 2.59858
R4439 VSS VSS.n229 2.56738
R4440 VSS.n2086 VSS.n2055 2.55412
R4441 VSS.n2938 VSS.n2937 2.50679
R4442 VSS.n1432 VSS.n1421 2.50679
R4443 VSS.n1971 VSS.n1243 2.50679
R4444 VSS.n692 VSS.n691 2.38348
R4445 VSS.n2208 VSS.n2207 2.33701
R4446 VSS.n2207 VSS.n1155 2.33701
R4447 VSS.n2270 VSS.n2269 2.33701
R4448 VSS.n2269 VSS.n2268 2.33701
R4449 VSS.n1132 VSS.n1130 2.33701
R4450 VSS.n2264 VSS.n1132 2.33701
R4451 VSS.n1150 VSS.n1148 2.33701
R4452 VSS.n2243 VSS.n1150 2.33701
R4453 VSS.n2242 VSS.n2241 2.33701
R4454 VSS.n2241 VSS.n2240 2.33701
R4455 VSS.n2946 VSS.n2945 2.33701
R4456 VSS.n2945 VSS.n2944 2.33701
R4457 VSS.n1220 VSS.n1218 2.33701
R4458 VSS.n2111 VSS.n1220 2.33701
R4459 VSS.n2076 VSS.n2075 2.33701
R4460 VSS.n2075 VSS.n2074 2.33701
R4461 VSS.n2063 VSS.n575 2.33701
R4462 VSS.n2899 VSS.n2898 2.33701
R4463 VSS.n2898 VSS.n2897 2.33701
R4464 VSS.n2715 VSS.n2714 2.33701
R4465 VSS.n2714 VSS.n734 2.33701
R4466 VSS.n2749 VSS.n712 2.33701
R4467 VSS.n2752 VSS.n712 2.33701
R4468 VSS.n2754 VSS.n2753 2.33701
R4469 VSS.n2755 VSS.n2754 2.33701
R4470 VSS.n2779 VSS.n696 2.33701
R4471 VSS.n2782 VSS.n696 2.33701
R4472 VSS.n2784 VSS.n2783 2.33701
R4473 VSS.n2786 VSS.n2784 2.33701
R4474 VSS.n2085 VSS.n2056 2.33067
R4475 VSS.n295 VSS.n288 2.3255
R4476 VSS.n301 VSS.n287 2.3255
R4477 VSS.n327 VSS.n326 2.3255
R4478 VSS.n332 VSS.n331 2.3255
R4479 VSS.n375 VSS.n374 2.3255
R4480 VSS.n352 VSS.n351 2.3255
R4481 VSS.n349 VSS.n345 2.3255
R4482 VSS.n201 VSS.n200 2.3255
R4483 VSS.n3088 VSS.n3087 2.25932
R4484 VSS.n3128 VSS.n3098 2.25932
R4485 VSS.n629 VSS.n628 2.25932
R4486 VSS.n1478 VSS.n1393 2.25932
R4487 VSS.n1679 VSS.n1678 2.25932
R4488 VSS.n1657 VSS.n1656 2.25932
R4489 VSS.n1598 VSS.n1587 2.25932
R4490 VSS.n1599 VSS.n1598 2.25932
R4491 VSS.n919 VSS.n918 2.25932
R4492 VSS.n1853 VSS.n1852 2.25932
R4493 VSS.n1892 VSS.n1891 2.25932
R4494 VSS.n1920 VSS.n934 2.25932
R4495 VSS.n2182 VSS.n1169 2.25312
R4496 VSS.n2134 VSS.n1202 2.25312
R4497 VSS.n2689 VSS.n748 2.25312
R4498 VSS.n2596 VSS.n841 2.25293
R4499 VSS.n3050 VSS.n3049 2.23999
R4500 VSS.n1169 VSS.n1168 2.2228
R4501 VSS.n1204 VSS.n1202 2.2228
R4502 VSS.n748 VSS.n747 2.2228
R4503 VSS.n1845 VSS.n1844 2.17922
R4504 VSS.n3295 VSS.n3294 2.14347
R4505 VSS.n1716 VSS.n1715 2.13383
R4506 VSS.n1125 VSS.n1124 2.11085
R4507 VSS.n718 VSS.n717 2.11085
R4508 VSS.n2851 VSS.n2850 2.06919
R4509 VSS.n3067 VSS.n3066 2.03479
R4510 VSS.n2064 VSS.n2063 2.03225
R4511 VSS.n556 VSS.n555 1.98299
R4512 VSS.n2884 VSS.n2883 1.98299
R4513 VSS.n2840 VSS.n2837 1.98299
R4514 VSS.n2852 VSS.n2840 1.98299
R4515 VSS.n814 VSS.n813 1.98299
R4516 VSS.n2539 VSS.n2538 1.97497
R4517 VSS.n2083 VSS.n2082 1.91571
R4518 VSS.n2850 VSS.n2849 1.8968
R4519 VSS.n875 VSS.n874 1.88285
R4520 VSS.n1665 VSS.n1664 1.87876
R4521 VSS.n975 VSS.n964 1.79699
R4522 VSS.n3068 VSS.n3067 1.77326
R4523 VSS.n2627 VSS.n2626 1.75824
R4524 VSS.n3435 VSS.n3434 1.753
R4525 VSS.n3433 VSS.n3432 1.753
R4526 VSS.n3166 VSS.n3165 1.753
R4527 VSS.n3164 VSS.n3163 1.753
R4528 VSS.n96 VSS.n79 1.753
R4529 VSS.n3380 VSS.n3379 1.753
R4530 VSS.n1671 VSS.n1669 1.7528
R4531 VSS.n555 VSS.n554 1.72441
R4532 VSS.n2883 VSS.n2882 1.72441
R4533 VSS.n813 VSS.n812 1.72441
R4534 VSS.n2307 VSS.n507 1.70468
R4535 VSS.n2306 VSS.n507 1.70468
R4536 VSS.n1832 VSS.n1736 1.70393
R4537 VSS.n1833 VSS.n1832 1.70393
R4538 VSS.n1334 VSS.n760 1.70393
R4539 VSS.n1324 VSS.n760 1.70393
R4540 VSS.n2167 VSS.n2166 1.70393
R4541 VSS.n2166 VSS.n2165 1.70393
R4542 VSS.n2969 VSS.n2968 1.70348
R4543 VSS.n2968 VSS.n503 1.70348
R4544 VSS.n2294 VSS.n1116 1.70338
R4545 VSS.n2294 VSS.n1050 1.70338
R4546 VSS.n3004 VSS.n267 1.70332
R4547 VSS.n3015 VSS.n267 1.70332
R4548 VSS.n3044 VSS.n237 1.70231
R4549 VSS.n242 VSS.n237 1.70231
R4550 VSS.n820 VSS.n803 1.7012
R4551 VSS.n2525 VSS.n984 1.69188
R4552 VSS.n2525 VSS.n2524 1.69188
R4553 VSS.n1951 VSS.n830 1.69188
R4554 VSS.n1258 VSS.n830 1.69188
R4555 VSS.n1453 VSS.n827 1.69188
R4556 VSS.n1408 VSS.n827 1.69188
R4557 VSS.n2772 VSS.n2771 1.69188
R4558 VSS.n2771 VSS.n2770 1.69188
R4559 VSS.n2921 VSS.n569 1.69188
R4560 VSS.n2921 VSS.n2920 1.69188
R4561 VSS.n2253 VSS.n504 1.69188
R4562 VSS.n2256 VSS.n504 1.69188
R4563 VSS.n2607 VSS.n828 1.69188
R4564 VSS.n2017 VSS.n2016 1.69188
R4565 VSS.n2018 VSS.n2017 1.69188
R4566 VSS.n1646 VSS.n1233 1.69188
R4567 VSS.n1648 VSS.n1233 1.69188
R4568 VSS.n1488 VSS.n1385 1.69188
R4569 VSS.n1385 VSS.n1384 1.69188
R4570 VSS.n2736 VSS.n2735 1.69188
R4571 VSS.n2735 VSS.n2734 1.69188
R4572 VSS.n2091 VSS.n2090 1.69188
R4573 VSS.n2092 VSS.n2091 1.69188
R4574 VSS.n2292 VSS.n1117 1.69188
R4575 VSS.n2292 VSS.n2291 1.69188
R4576 VSS.n1984 VSS.n1234 1.69188
R4577 VSS.n1797 VSS.n1796 1.69188
R4578 VSS.n1798 VSS.n1797 1.69188
R4579 VSS.n1877 VSS.n1876 1.69188
R4580 VSS.n1876 VSS.n1875 1.69188
R4581 VSS.n1685 VSS.n1277 1.69188
R4582 VSS.n1687 VSS.n1277 1.69188
R4583 VSS.n1529 VSS.n1299 1.69188
R4584 VSS.n1529 VSS.n1528 1.69188
R4585 VSS.n2704 VSS.n2703 1.69188
R4586 VSS.n2703 VSS.n2702 1.69188
R4587 VSS.n2123 VSS.n2122 1.69188
R4588 VSS.n2124 VSS.n2123 1.69188
R4589 VSS.n2197 VSS.n2196 1.69188
R4590 VSS.n2196 VSS.n2195 1.69188
R4591 VSS.n1727 VSS.n1533 1.69188
R4592 VSS.n1727 VSS.n1726 1.69188
R4593 VSS.n2674 VSS.n2673 1.69188
R4594 VSS.n2673 VSS.n2672 1.69188
R4595 VSS.n2149 VSS.n1180 1.69188
R4596 VSS.n2149 VSS.n2148 1.69188
R4597 VSS.n1829 VSS.n1737 1.69188
R4598 VSS.n2485 VSS.n2484 1.69188
R4599 VSS.n2486 VSS.n2485 1.69188
R4600 VSS.n2572 VSS.n924 1.69188
R4601 VSS.n2572 VSS.n2571 1.69188
R4602 VSS.n2581 VSS.n2580 1.69188
R4603 VSS.n2580 VSS.n2579 1.69188
R4604 VSS.n2653 VSS.n762 1.69188
R4605 VSS.n2653 VSS.n2652 1.69188
R4606 VSS.n2809 VSS.n669 1.69188
R4607 VSS.n2796 VSS.n669 1.69188
R4608 VSS.n2874 VSS.n668 1.69188
R4609 VSS.n2875 VSS.n2874 1.69188
R4610 VSS.n2963 VSS.n508 1.69188
R4611 VSS.n2963 VSS.n2962 1.69188
R4612 VSS.n2453 VSS.n982 1.69188
R4613 VSS.n2428 VSS.n982 1.69188
R4614 VSS.n2531 VSS.n981 1.69188
R4615 VSS.n2532 VSS.n2531 1.69188
R4616 VSS.n895 VSS.n825 1.69188
R4617 VSS.n897 VSS.n825 1.69188
R4618 VSS.n2613 VSS.n824 1.69188
R4619 VSS.n2614 VSS.n2613 1.69188
R4620 VSS.n2869 VSS.n671 1.69188
R4621 VSS.n2869 VSS.n2868 1.69188
R4622 VSS.n641 VSS.n567 1.69188
R4623 VSS.n644 VSS.n567 1.69188
R4624 VSS.n2927 VSS.n566 1.69188
R4625 VSS.n2928 VSS.n2927 1.69188
R4626 VSS.n972 VSS.n964 1.64728
R4627 VSS.n2641 VSS.n772 1.61169
R4628 VSS.n3401 VSS 1.54822
R4629 VSS.n3160 VSS.n3146 1.50638
R4630 VSS.n3154 VSS.n3148 1.50638
R4631 VSS.n191 VSS.n189 1.50638
R4632 VSS.n3182 VSS.n192 1.50638
R4633 VSS.n3096 VSS.n3095 1.50638
R4634 VSS.n3097 VSS.n3096 1.50638
R4635 VSS.n3125 VSS.n3124 1.50638
R4636 VSS.n3118 VSS.n3101 1.50638
R4637 VSS.n3118 VSS.n3117 1.50638
R4638 VSS.n3109 VSS.n3108 1.50638
R4639 VSS.n2891 VSS.n2890 1.47352
R4640 VSS.n3067 VSS.n3054 1.44312
R4641 VSS.n2106 VSS.n2105 1.34658
R4642 VSS.n3052 VSS.n229 1.3415
R4643 VSS.n691 VSS.n690 1.3283
R4644 VSS.n3051 VSS.n3050 1.31337
R4645 VSS.n2184 VSS.n1168 1.29527
R4646 VSS.n2132 VSS.n1204 1.29527
R4647 VSS.n2691 VSS.n747 1.29527
R4648 VSS.n545 VSS.n533 1.25365
R4649 VSS.n2104 VSS.n2103 1.25033
R4650 VSS.n17 VSS.n1 1.21169
R4651 VSS.n3133 VSS.n3132 1.21169
R4652 VSS.n3296 VSS.n111 1.21169
R4653 VSS.n1341 VSS.n1340 1.20723
R4654 VSS.n1664 VSS.n1663 1.18311
R4655 VSS.n1926 VSS.n1925 1.18311
R4656 VSS.n2542 VSS.n2541 1.18311
R4657 VSS.n1746 VSS.n1745 1.18311
R4658 VSS.n2438 VSS.n2437 1.18311
R4659 VSS.n2354 VSS.n2353 1.18311
R4660 VSS.n1061 VSS.n1060 1.18311
R4661 VSS.n3037 VSS.n3036 1.18311
R4662 VSS.n246 VSS.n245 1.18311
R4663 VSS.n450 VSS.n409 1.15795
R4664 VSS.n1701 VSS.n1554 1.14023
R4665 VSS.n2480 VSS.n2479 1.14023
R4666 VSS.n2328 VSS.n2327 1.14023
R4667 VSS.n3022 VSS.n262 1.14023
R4668 VSS.n1604 VSS.n1601 1.12991
R4669 VSS.n2889 VSS.n2888 1.12954
R4670 VSS.n2296 VSS 1.12383
R4671 VSS.n2295 VSS 1.11689
R4672 VSS.n2300 VSS 1.11689
R4673 VSS.n3050 VSS.n232 1.11056
R4674 VSS.n2299 VSS 1.07702
R4675 VSS.n2621 VSS.n2620 1.07463
R4676 VSS.n3469 VSS 1.06996
R4677 VSS.n3052 VSS.n3051 1.05425
R4678 VSS.n3433 VSS 1.00137
R4679 VSS.n2381 VSS.n2380 0.993972
R4680 VSS.n801 VSS.n793 0.985115
R4681 VSS.n1846 VSS.n1845 0.953691
R4682 VSS.n888 VSS.n879 0.952566
R4683 VSS.n1790 VSS.n1781 0.952566
R4684 VSS.n1228 VSS.n1227 0.952566
R4685 VSS.n2000 VSS.n1996 0.952566
R4686 VSS.n2461 VSS.n2417 0.952566
R4687 VSS.n472 VSS.n0 0.927421
R4688 VSS.n887 VSS.n882 0.899674
R4689 VSS.n1961 VSS.n1249 0.895605
R4690 VSS.n1264 VSS.n1263 0.895605
R4691 VSS.n2179 VSS.n1169 0.892621
R4692 VSS.n1202 VSS.n1201 0.892621
R4693 VSS.n2686 VSS.n748 0.892621
R4694 VSS.n2375 VSS.n1023 0.853
R4695 VSS.n2379 VSS.n2378 0.842928
R4696 VSS.n2475 VSS.n2411 0.833377
R4697 VSS.n2323 VSS.n1034 0.833377
R4698 VSS.n3025 VSS.n3024 0.833377
R4699 VSS.n2083 VSS.n2056 0.830425
R4700 VSS.n2054 VSS.n2042 0.798505
R4701 VSS.n2388 VSS.n2387 0.777453
R4702 VSS.n3434 VSS.n3433 0.761313
R4703 VSS.n3165 VSS.n3164 0.761313
R4704 VSS.n3380 VSS.n79 0.761313
R4705 VSS.n3156 VSS.n3155 0.753441
R4706 VSS.n3150 VSS.n188 0.753441
R4707 VSS.n3184 VSS.n3183 0.753441
R4708 VSS.n3178 VSS.n3177 0.753441
R4709 VSS.n3129 VSS.n3128 0.753441
R4710 VSS.n3122 VSS.n3121 0.753441
R4711 VSS.n3115 VSS.n3114 0.753441
R4712 VSS.n1483 VSS.n1482 0.753441
R4713 VSS.n1674 VSS.n1673 0.753441
R4714 VSS.n908 VSS.n861 0.753441
R4715 VSS.n1510 VSS.n1509 0.716584
R4716 VSS.n2086 VSS.n2085 0.606984
R4717 VSS.n468 VSS.n426 0.577852
R4718 VSS.t643 VSS.t467 0.577852
R4719 VSS.n460 VSS.n438 0.577852
R4720 VSS.n2233 VSS.n2226 0.537563
R4721 VSS.n2829 VSS.n2828 0.537563
R4722 VSS.n2816 VSS.n2815 0.537563
R4723 VSS.n2827 VSS.n680 0.537563
R4724 VSS.n2624 VSS.n781 0.537563
R4725 VSS.n1425 VSS.n1424 0.537563
R4726 VSS.n2628 VSS.n2627 0.537563
R4727 VSS.n1362 VSS.n1361 0.537563
R4728 VSS.n1517 VSS.n1516 0.537563
R4729 VSS.n1496 VSS.n1370 0.537563
R4730 VSS.n1945 VSS.n1944 0.537563
R4731 VSS.n2338 VSS.n2337 0.537563
R4732 VSS.n2359 VSS.n2350 0.537563
R4733 VSS.n1096 VSS.n1080 0.537563
R4734 VSS.n2984 VSS.n495 0.537563
R4735 VSS.n1075 VSS.n1074 0.537563
R4736 VSS.n1098 VSS.n1097 0.537563
R4737 VSS.n271 VSS.n264 0.537563
R4738 VSS.n2989 VSS.n277 0.537563
R4739 VSS.n1 VSS 0.531208
R4740 VSS.n3133 VSS 0.531208
R4741 VSS.n1708 VSS.n1552 0.526527
R4742 VSS.n1705 VSS.n1704 0.526527
R4743 VSS.n2476 VSS.n2399 0.526527
R4744 VSS.n2324 VSS.n2322 0.526527
R4745 VSS.n261 VSS.n259 0.526527
R4746 VSS.n1532 VSS.n1531 0.500125
R4747 VSS.n1831 VSS.n1830 0.500125
R4748 VSS.n1179 VSS.n1178 0.500125
R4749 VSS.n2151 VSS.n2150 0.500125
R4750 VSS.n759 VSS.n758 0.500125
R4751 VSS.n2659 VSS.n2658 0.500125
R4752 VSS.n3382 VSS.n3381 0.482665
R4753 VSS.n3049 VSS.n0 0.473674
R4754 VSS.n329 VSS.n328 0.467019
R4755 VSS.n350 VSS.n228 0.467019
R4756 VSS.n3220 VSS.n3201 0.467019
R4757 VSS.n3273 VSS.n78 0.467019
R4758 VSS.n3294 VSS 0.448179
R4759 VSS.n525 VSS.n523 0.448052
R4760 VSS.n1359 VSS.n1358 0.448052
R4761 VSS.n1515 VSS.n1514 0.448052
R4762 VSS.n232 VSS.n210 0.426643
R4763 VSS.n1669 VSS.n1578 0.417891
R4764 VSS.n1663 VSS.n1662 0.417891
R4765 VSS.n1930 VSS.n1918 0.417891
R4766 VSS.n1925 VSS.n1924 0.417891
R4767 VSS.n2547 VSS.n944 0.417891
R4768 VSS.n2544 VSS.n2543 0.417891
R4769 VSS.n2541 VSS.n2540 0.417891
R4770 VSS.n1757 VSS.n1741 0.417891
R4771 VSS.n2442 VSS.n2435 0.417891
R4772 VSS.n2358 VSS.n2351 0.417891
R4773 VSS.n1059 VSS.n278 0.417891
R4774 VSS.n1060 VSS.n1055 0.417891
R4775 VSS.n3040 VSS.n3039 0.417891
R4776 VSS.n3036 VSS.n3035 0.417891
R4777 VSS.n255 VSS.n240 0.417891
R4778 VSS.n2387 VSS.n1016 0.410656
R4779 VSS.n3430 VSS.n58 0.409011
R4780 VSS.n3444 VSS.n40 0.409011
R4781 VSS.n33 VSS.n32 0.409011
R4782 VSS.n3464 VSS.n3 0.409011
R4783 VSS.n7 VSS.n6 0.409011
R4784 VSS.n8 VSS.n4 0.409011
R4785 VSS.n3377 VSS.n81 0.409011
R4786 VSS.n97 VSS.n92 0.409011
R4787 VSS.n3316 VSS.n115 0.409011
R4788 VSS.n3320 VSS.n3319 0.409011
R4789 VSS.n3324 VSS.n3323 0.409011
R4790 VSS.n3352 VSS.n3341 0.409011
R4791 VSS.n625 VSS.n610 0.409011
R4792 VSS.n618 VSS.n617 0.409011
R4793 VSS.n1418 VSS.n1415 0.409011
R4794 VSS.n1720 VSS.n1541 0.409011
R4795 VSS.n1710 VSS.n1709 0.409011
R4796 VSS.n877 VSS.n876 0.409011
R4797 VSS.n1839 VSS.n1290 0.409011
R4798 VSS.n1843 VSS.n1289 0.409011
R4799 VSS.n1816 VSS.n1763 0.409011
R4800 VSS.n1810 VSS.n1809 0.409011
R4801 VSS.n1780 VSS.n1779 0.409011
R4802 VSS.n2028 VSS.n1225 0.409011
R4803 VSS.n1995 VSS.n1993 0.409011
R4804 VSS.n2510 VSS.n2509 0.409011
R4805 VSS.n2504 VSS.n997 0.409011
R4806 VSS.n2497 VSS.n2397 0.409011
R4807 VSS.n2416 VSS.n2414 0.409011
R4808 VSS.n1043 VSS.n1039 0.409011
R4809 VSS.n258 VSS.n256 0.409011
R4810 VSS.n2055 VSS.n2054 0.383542
R4811 VSS.n1834 VSS.n1297 0.381255
R4812 VSS.n2656 VSS.n702 0.3805
R4813 VSS.n670 VSS.n570 0.3805
R4814 VSS.n2923 VSS.n2922 0.3805
R4815 VSS.n2967 VSS.n2966 0.3805
R4816 VSS.n2527 VSS.n2526 0.3805
R4817 VSS.n2609 VSS.n2608 0.3805
R4818 VSS.n2293 VSS.n505 0.3805
R4819 VSS.n1118 VSS.n568 0.3805
R4820 VSS.n757 VSS.n722 0.3805
R4821 VSS.n2657 VSS.n723 0.3805
R4822 VSS.n1380 VSS.n826 0.3805
R4823 VSS.n1985 VSS.n983 0.3805
R4824 VSS.n1178 VSS.n1162 0.3805
R4825 VSS.n2150 VSS.n1163 0.3805
R4826 VSS.n758 VSS.n741 0.3805
R4827 VSS.n2658 VSS.n742 0.3805
R4828 VSS.n1531 VSS.n1530 0.3805
R4829 VSS.n1830 VSS.n1278 0.3805
R4830 VSS.n2965 VSS.n2964 0.3805
R4831 VSS.n2924 VSS.n509 0.3805
R4832 VSS.n2873 VSS.n2872 0.3805
R4833 VSS.n2655 VSS.n2654 0.3805
R4834 VSS.n2610 VSS.n763 0.3805
R4835 VSS.n2528 VSS.n925 0.3805
R4836 VSS.n761 VSS.n672 0.3805
R4837 VSS.n2871 VSS.n2870 0.3805
R4838 VSS.n2926 VSS.n2925 0.3805
R4839 VSS.n530 VSS.n506 0.3805
R4840 VSS.n2530 VSS.n2529 0.3805
R4841 VSS.n2612 VSS.n2611 0.3805
R4842 VSS.n874 VSS.n863 0.376971
R4843 uio_oe[7] VSS.n3491 0.371345
R4844 VSS VSS.n3295 0.366908
R4845 VSS.n3049 VSS.n3048 0.364419
R4846 VSS.n3297 VSS.n116 0.358995
R4847 VSS.n2823 VSS.n680 0.358542
R4848 VSS.n1430 VSS.n1429 0.358542
R4849 VSS.n2635 VSS.n2634 0.358542
R4850 VSS.n1969 VSS.n1243 0.358542
R4851 VSS.n1438 VSS.n1437 0.340926
R4852 VSS.n3048 VSS.n3047 0.335802
R4853 VSS.n3469 uo_out[0] 0.3295
R4854 VSS.n3470 uo_out[1] 0.3295
R4855 VSS.n3471 uo_out[2] 0.3295
R4856 VSS.n3472 uo_out[3] 0.3295
R4857 VSS.n3473 uo_out[4] 0.3295
R4858 VSS.n3474 uo_out[5] 0.3295
R4859 VSS.n3475 uo_out[6] 0.3295
R4860 VSS.n3476 uo_out[7] 0.3295
R4861 VSS.n3477 uio_out[0] 0.3295
R4862 VSS.n3478 uio_out[1] 0.3295
R4863 VSS.n3479 uio_out[2] 0.3295
R4864 VSS.n3480 uio_out[3] 0.3295
R4865 VSS.n3481 uio_out[4] 0.3295
R4866 VSS.n3482 uio_out[5] 0.3295
R4867 VSS.n3483 uio_out[6] 0.3295
R4868 VSS.n3484 uio_out[7] 0.3295
R4869 VSS.n3485 uio_oe[0] 0.3295
R4870 VSS.n3486 uio_oe[1] 0.3295
R4871 VSS.n3487 uio_oe[2] 0.3295
R4872 VSS.n3488 uio_oe[3] 0.3295
R4873 VSS.n3489 uio_oe[4] 0.3295
R4874 VSS.n3490 uio_oe[5] 0.3295
R4875 VSS.n3491 uio_oe[6] 0.3295
R4876 VSS.n1704 VSS.n1703 0.307349
R4877 VSS.n2185 VSS.n2184 0.305262
R4878 VSS.n2201 VSS.n1158 0.305262
R4879 VSS.n2202 VSS.n1157 0.305262
R4880 VSS.n2215 VSS.n2214 0.305262
R4881 VSS.n2278 VSS.n2277 0.305262
R4882 VSS.n2263 VSS.n2262 0.305262
R4883 VSS.n1142 VSS.n1140 0.305262
R4884 VSS.n2237 VSS.n1151 0.305262
R4885 VSS.n2232 VSS.n2227 0.305262
R4886 VSS.n2939 VSS.n521 0.305262
R4887 VSS.n2132 VSS.n2131 0.305262
R4888 VSS.n1217 VSS.n1216 0.305262
R4889 VSS.n2118 VSS.n2117 0.305262
R4890 VSS.n2106 VSS.n1221 0.305262
R4891 VSS.n2060 VSS.n2058 0.305262
R4892 VSS.n2069 VSS.n2068 0.305262
R4893 VSS.n2067 VSS.n2064 0.305262
R4894 VSS.n2904 VSS.n576 0.305262
R4895 VSS.n2903 VSS.n577 0.305262
R4896 VSS.n2892 VSS.n2891 0.305262
R4897 VSS.n2692 VSS.n2691 0.305262
R4898 VSS.n2708 VSS.n737 0.305262
R4899 VSS.n2709 VSS.n736 0.305262
R4900 VSS.n2722 VSS.n2721 0.305262
R4901 VSS.n2742 VSS.n2741 0.305262
R4902 VSS.n2758 VSS.n710 0.305262
R4903 VSS.n2765 VSS.n2764 0.305262
R4904 VSS.n2785 VSS.n694 0.305262
R4905 VSS.n2380 VSS.n2379 0.298799
R4906 VSS.n2182 VSS.n2181 0.298074
R4907 VSS.n2135 VSS.n2134 0.298074
R4908 VSS.n2689 VSS.n2688 0.298074
R4909 VSS.n471 VSS 0.286698
R4910 VSS.n1325 VSS.n1297 0.281546
R4911 VSS.n2164 VSS.n233 0.281132
R4912 VSS.n2302 VSS.n2301 0.278782
R4913 VSS VSS.n3468 0.268171
R4914 VSS.n1700 VSS.n1699 0.263514
R4915 VSS.n2474 VSS.n2473 0.263514
R4916 VSS.n2331 VSS.n1032 0.263514
R4917 VSS.n3021 VSS.n3020 0.263514
R4918 VSS.n3296 VSS 0.260439
R4919 VSS.n2173 VSS.n1171 0.259086
R4920 VSS.n560 VSS.n546 0.259086
R4921 VSS.n554 VSS.n553 0.259086
R4922 VSS.n2141 VSS.n1198 0.259086
R4923 VSS.n2888 VSS.n582 0.259086
R4924 VSS.n2882 VSS.n2881 0.259086
R4925 VSS.n2103 VSS.n2039 0.259086
R4926 VSS.n2099 VSS.n2098 0.259086
R4927 VSS.n2836 VSS.n2835 0.259086
R4928 VSS.n2846 VSS.n2841 0.259086
R4929 VSS.n2680 VSS.n750 0.259086
R4930 VSS.n818 VSS.n804 0.259086
R4931 VSS.n812 VSS.n811 0.259086
R4932 VSS.n1341 VSS.n1313 0.259086
R4933 VSS.n1346 VSS.n1311 0.259086
R4934 VSS.n1015 VSS.n1005 0.2565
R4935 VSS.n3467 VSS.n1 0.249698
R4936 VSS.n1782 VSS.n1778 0.239381
R4937 VSS.n1998 VSS.n1994 0.239381
R4938 VSS VSS.n2596 0.237784
R4939 VSS.n2379 VSS.n116 0.23574
R4940 VSS.n963 VSS.n962 0.225061
R4941 VSS.n971 VSS.n970 0.225061
R4942 VSS.n2380 VSS.n2376 0.224703
R4943 VSS.n2297 VSS.n237 0.218753
R4944 VSS.n621 VSS.n620 0.204755
R4945 VSS.n2538 VSS.n948 0.204755
R4946 VSS.n960 VSS.n948 0.204755
R4947 VSS.n2596 VSS 0.200023
R4948 VSS VSS.n2182 0.199635
R4949 VSS.n2134 VSS 0.199635
R4950 VSS VSS.n2689 0.199635
R4951 VSS.n231 VSS.n181 0.198729
R4952 VSS.n2298 VSS.n2297 0.196532
R4953 VSS.n1049 VSS.n234 0.196532
R4954 VSS.n2301 VSS.n2300 0.195539
R4955 VSS.n3054 VSS.n3053 0.194976
R4956 VSS.n2082 VSS.n2081 0.192021
R4957 VSS.n3047 VSS.n234 0.18942
R4958 VSS.n2376 VSS.n1019 0.184476
R4959 VSS.n330 VSS.n230 0.1838
R4960 VSS.n3383 VSS.n3382 0.1838
R4961 VSS.n2419 VSS.n2415 0.180304
R4962 VSS.n885 VSS 0.17983
R4963 VSS.n968 VSS 0.17983
R4964 VSS.n536 VSS.n526 0.179521
R4965 VSS.n1430 VSS.n1421 0.179521
R4966 VSS.n1969 VSS.n1968 0.179521
R4967 VSS VSS.n551 0.179485
R4968 VSS VSS.n615 0.179485
R4969 VSS.n2843 VSS 0.179485
R4970 VSS VSS.n809 0.179485
R4971 VSS.n2305 VSS.n2304 0.175416
R4972 VSS.n2387 VSS.n2386 0.173577
R4973 VSS.n2607 VSS.n830 0.1603
R4974 VSS.n1984 VSS.n1233 0.1603
R4975 VSS.n1876 VSS.n1277 0.1603
R4976 VSS.n1832 VSS.n1727 0.1603
R4977 VSS.n2580 VSS.n2572 0.1603
R4978 VSS.n2531 VSS.n825 0.1603
R4979 VSS.n2608 VSS.n827 0.159712
R4980 VSS.n1385 VSS.n1380 0.159712
R4981 VSS.n1530 VSS.n1529 0.159712
R4982 VSS.n1532 VSS.n760 0.159712
R4983 VSS.n2653 VSS.n763 0.159712
R4984 VSS.n2613 VSS.n2612 0.159712
R4985 VSS.n2259 VSS 0.158169
R4986 VSS VSS.n709 0.158169
R4987 VSS.n2794 VSS 0.158169
R4988 VSS VSS.n880 0.156867
R4989 VSS.n2424 VSS.n2419 0.151658
R4990 VSS.n2170 VSS.n2169 0.143027
R4991 VSS.n1196 VSS.n1195 0.143027
R4992 VSS.n2677 VSS.n2676 0.143027
R4993 VSS.n2170 VSS 0.14207
R4994 VSS.n551 VSS 0.14207
R4995 VSS VSS.n1196 0.14207
R4996 VSS.n615 VSS 0.14207
R4997 VSS.n2677 VSS 0.14207
R4998 VSS.n2843 VSS 0.14207
R4999 VSS.n809 VSS 0.14207
R5000 VSS VSS.n1782 0.14207
R5001 VSS.n1998 VSS 0.14207
R5002 VSS.n885 VSS 0.141725
R5003 VSS.n968 VSS 0.141725
R5004 VSS.n1297 VSS.n233 0.141676
R5005 VSS.n3111 VSS.n3105 0.141672
R5006 VSS.n3143 VSS.n211 0.141672
R5007 VSS.n2967 VSS.n504 0.137387
R5008 VSS.n2293 VSS.n2292 0.137387
R5009 VSS.n2196 VSS.n1162 0.137387
R5010 VSS.n2166 VSS.n1179 0.137387
R5011 VSS.n2964 VSS.n2963 0.137387
R5012 VSS.n2927 VSS.n530 0.137387
R5013 VSS.n891 VSS.n890 0.13667
R5014 VSS.n2526 VSS.n2525 0.126812
R5015 VSS.n2017 VSS.n1985 0.126812
R5016 VSS.n1797 VSS.n1278 0.126812
R5017 VSS.n1831 VSS.n1829 0.126812
R5018 VSS.n2485 VSS.n925 0.126812
R5019 VSS.n2530 VSS.n982 0.126812
R5020 VSS.n2105 VSS.n2104 0.126617
R5021 VSS.n2771 VSS.n702 0.125637
R5022 VSS.n2735 VSS.n723 0.125637
R5023 VSS.n2703 VSS.n742 0.125637
R5024 VSS.n2673 VSS.n2659 0.125637
R5025 VSS.n2654 VSS.n669 0.125637
R5026 VSS.n2869 VSS.n672 0.125637
R5027 VSS.n3447 VSS.n37 0.1255
R5028 VSS.n3174 VSS.n3173 0.1255
R5029 VSS.n3356 VSS.n106 0.1255
R5030 VSS.n3297 VSS.n3296 0.122556
R5031 VSS.n3105 VSS 0.121778
R5032 VSS.n3168 VSS 0.121778
R5033 VSS.n2890 VSS.n2889 0.120632
R5034 VSS.n1713 VSS 0.120408
R5035 VSS.n54 VSS.n53 0.120292
R5036 VSS.n54 VSS.n41 0.120292
R5037 VSS.n3427 VSS.n59 0.120292
R5038 VSS.n3427 VSS.n3426 0.120292
R5039 VSS.n3425 VSS.n61 0.120292
R5040 VSS.n62 VSS.n61 0.120292
R5041 VSS.n3418 VSS.n3410 0.120292
R5042 VSS.n3418 VSS.n3417 0.120292
R5043 VSS.n3416 VSS.n3413 0.120292
R5044 VSS.n3413 VSS.n3412 0.120292
R5045 VSS.n3443 VSS.n3442 0.120292
R5046 VSS.n3439 VSS.n3438 0.120292
R5047 VSS.n51 VSS.n43 0.120292
R5048 VSS.n46 VSS.n43 0.120292
R5049 VSS.n46 VSS.n45 0.120292
R5050 VSS.n12 VSS.n11 0.120292
R5051 VSS.n3456 VSS.n18 0.120292
R5052 VSS.n19 VSS.n18 0.120292
R5053 VSS.n3450 VSS.n20 0.120292
R5054 VSS.n34 VSS.n23 0.120292
R5055 VSS.n28 VSS.n23 0.120292
R5056 VSS.n28 VSS.n27 0.120292
R5057 VSS.n3141 VSS.n213 0.120292
R5058 VSS.n3136 VSS.n213 0.120292
R5059 VSS.n3136 VSS.n3135 0.120292
R5060 VSS.n3092 VSS.n3091 0.120292
R5061 VSS.n3126 VSS.n3099 0.120292
R5062 VSS.n3120 VSS.n3099 0.120292
R5063 VSS.n3119 VSS.n3102 0.120292
R5064 VSS.n3112 VSS.n3111 0.120292
R5065 VSS.n3159 VSS.n3158 0.120292
R5066 VSS.n3158 VSS.n3147 0.120292
R5067 VSS.n3153 VSS.n3152 0.120292
R5068 VSS.n3152 VSS.n3149 0.120292
R5069 VSS.n3187 VSS.n3186 0.120292
R5070 VSS.n3186 VSS.n190 0.120292
R5071 VSS.n3181 VSS.n3180 0.120292
R5072 VSS.n3180 VSS.n193 0.120292
R5073 VSS.n3172 VSS.n3171 0.120292
R5074 VSS.n3306 VSS.n3301 0.120292
R5075 VSS.n3301 VSS.n80 0.120292
R5076 VSS.n3374 VSS.n82 0.120292
R5077 VSS.n3374 VSS.n3373 0.120292
R5078 VSS.n3372 VSS.n84 0.120292
R5079 VSS.n85 VSS.n84 0.120292
R5080 VSS.n3365 VSS.n88 0.120292
R5081 VSS.n3365 VSS.n3364 0.120292
R5082 VSS.n3363 VSS.n90 0.120292
R5083 VSS.n91 VSS.n90 0.120292
R5084 VSS.n105 VSS.n104 0.120292
R5085 VSS.n101 VSS.n100 0.120292
R5086 VSS.n3312 VSS.n3300 0.120292
R5087 VSS.n3313 VSS.n3312 0.120292
R5088 VSS.n3314 VSS.n3313 0.120292
R5089 VSS.n3325 VSS.n114 0.120292
R5090 VSS.n3333 VSS.n109 0.120292
R5091 VSS.n3337 VSS.n109 0.120292
R5092 VSS.n3339 VSS.n3338 0.120292
R5093 VSS.n3351 VSS.n3350 0.120292
R5094 VSS.n3350 VSS.n3342 0.120292
R5095 VSS.n3344 VSS.n3342 0.120292
R5096 VSS.n2175 VSS.n2174 0.120292
R5097 VSS.n2175 VSS.n1170 0.120292
R5098 VSS.n2181 VSS.n1170 0.120292
R5099 VSS.n2204 VSS.n2203 0.120292
R5100 VSS.n2204 VSS.n1156 0.120292
R5101 VSS.n2209 VSS.n1156 0.120292
R5102 VSS.n2210 VSS.n2209 0.120292
R5103 VSS.n2211 VSS.n2210 0.120292
R5104 VSS.n2211 VSS.n1154 0.120292
R5105 VSS.n2216 VSS.n1154 0.120292
R5106 VSS.n2279 VSS.n1127 0.120292
R5107 VSS.n2274 VSS.n1127 0.120292
R5108 VSS.n2274 VSS.n2273 0.120292
R5109 VSS.n2273 VSS.n2272 0.120292
R5110 VSS.n2272 VSS.n1129 0.120292
R5111 VSS.n2267 VSS.n1129 0.120292
R5112 VSS.n2267 VSS.n2266 0.120292
R5113 VSS.n2266 VSS.n2265 0.120292
R5114 VSS.n2265 VSS.n1131 0.120292
R5115 VSS.n2250 VSS.n1139 0.120292
R5116 VSS.n2246 VSS.n1139 0.120292
R5117 VSS.n2246 VSS.n2245 0.120292
R5118 VSS.n2245 VSS.n2244 0.120292
R5119 VSS.n2244 VSS.n1149 0.120292
R5120 VSS.n2239 VSS.n1149 0.120292
R5121 VSS.n2239 VSS.n2238 0.120292
R5122 VSS.n2231 VSS.n2230 0.120292
R5123 VSS.n2949 VSS.n2948 0.120292
R5124 VSS.n2948 VSS.n2947 0.120292
R5125 VSS.n2947 VSS.n519 0.120292
R5126 VSS.n2942 VSS.n519 0.120292
R5127 VSS.n2942 VSS.n2941 0.120292
R5128 VSS.n2941 VSS.n2940 0.120292
R5129 VSS.n2936 VSS.n2935 0.120292
R5130 VSS.n2935 VSS.n524 0.120292
R5131 VSS.n2931 VSS.n524 0.120292
R5132 VSS.n559 VSS.n558 0.120292
R5133 VSS.n558 VSS.n547 0.120292
R5134 VSS.n552 VSS.n547 0.120292
R5135 VSS.n2140 VSS.n2139 0.120292
R5136 VSS.n2139 VSS.n1199 0.120292
R5137 VSS.n2135 VSS.n1199 0.120292
R5138 VSS.n2119 VSS.n1215 0.120292
R5139 VSS.n2114 VSS.n1215 0.120292
R5140 VSS.n2114 VSS.n2113 0.120292
R5141 VSS.n2113 VSS.n2112 0.120292
R5142 VSS.n2112 VSS.n1219 0.120292
R5143 VSS.n2108 VSS.n1219 0.120292
R5144 VSS.n2108 VSS.n2107 0.120292
R5145 VSS.n2102 VSS.n2101 0.120292
R5146 VSS.n2087 VSS.n2053 0.120292
R5147 VSS.n2080 VSS.n2053 0.120292
R5148 VSS.n2079 VSS.n2078 0.120292
R5149 VSS.n2078 VSS.n2059 0.120292
R5150 VSS.n2073 VSS.n2059 0.120292
R5151 VSS.n2073 VSS.n2072 0.120292
R5152 VSS.n2072 VSS.n2071 0.120292
R5153 VSS.n2071 VSS.n2062 0.120292
R5154 VSS.n2066 VSS.n2065 0.120292
R5155 VSS.n2902 VSS.n2901 0.120292
R5156 VSS.n2901 VSS.n578 0.120292
R5157 VSS.n2896 VSS.n578 0.120292
R5158 VSS.n2896 VSS.n2895 0.120292
R5159 VSS.n2895 VSS.n2894 0.120292
R5160 VSS.n2894 VSS.n580 0.120292
R5161 VSS.n2887 VSS.n2886 0.120292
R5162 VSS.n2886 VSS.n584 0.120292
R5163 VSS.n665 VSS.n596 0.120292
R5164 VSS.n661 VSS.n596 0.120292
R5165 VSS.n661 VSS.n660 0.120292
R5166 VSS.n660 VSS.n659 0.120292
R5167 VSS.n659 VSS.n601 0.120292
R5168 VSS.n653 VSS.n601 0.120292
R5169 VSS.n653 VSS.n652 0.120292
R5170 VSS.n652 VSS.n651 0.120292
R5171 VSS.n651 VSS.n603 0.120292
R5172 VSS.n647 VSS.n603 0.120292
R5173 VSS.n624 VSS.n623 0.120292
R5174 VSS.n623 VSS.n611 0.120292
R5175 VSS.n2682 VSS.n2681 0.120292
R5176 VSS.n2682 VSS.n749 0.120292
R5177 VSS.n2688 VSS.n749 0.120292
R5178 VSS.n2711 VSS.n2710 0.120292
R5179 VSS.n2711 VSS.n735 0.120292
R5180 VSS.n2716 VSS.n735 0.120292
R5181 VSS.n2717 VSS.n2716 0.120292
R5182 VSS.n2718 VSS.n2717 0.120292
R5183 VSS.n2718 VSS.n733 0.120292
R5184 VSS.n2723 VSS.n733 0.120292
R5185 VSS.n2744 VSS.n715 0.120292
R5186 VSS.n2745 VSS.n2744 0.120292
R5187 VSS.n2746 VSS.n2745 0.120292
R5188 VSS.n2746 VSS.n713 0.120292
R5189 VSS.n2750 VSS.n713 0.120292
R5190 VSS.n2751 VSS.n2750 0.120292
R5191 VSS.n2751 VSS.n711 0.120292
R5192 VSS.n2756 VSS.n711 0.120292
R5193 VSS.n2757 VSS.n2756 0.120292
R5194 VSS.n2776 VSS.n2775 0.120292
R5195 VSS.n2776 VSS.n697 0.120292
R5196 VSS.n2780 VSS.n697 0.120292
R5197 VSS.n2781 VSS.n2780 0.120292
R5198 VSS.n2781 VSS.n695 0.120292
R5199 VSS.n2787 VSS.n695 0.120292
R5200 VSS.n2788 VSS.n2787 0.120292
R5201 VSS.n2819 VSS.n683 0.120292
R5202 VSS.n2820 VSS.n2819 0.120292
R5203 VSS VSS.n2820 0.120292
R5204 VSS.n2826 VSS.n2825 0.120292
R5205 VSS.n2831 VSS.n679 0.120292
R5206 VSS.n2832 VSS.n2831 0.120292
R5207 VSS.n2854 VSS.n2853 0.120292
R5208 VSS.n2853 VSS.n2839 0.120292
R5209 VSS.n2848 VSS.n2839 0.120292
R5210 VSS.n2848 VSS.n2847 0.120292
R5211 VSS.n1343 VSS.n1342 0.120292
R5212 VSS.n1343 VSS.n1312 0.120292
R5213 VSS.n1348 VSS.n1312 0.120292
R5214 VSS.n1349 VSS.n1348 0.120292
R5215 VSS.n1355 VSS.n1309 0.120292
R5216 VSS.n1357 VSS.n1356 0.120292
R5217 VSS.n1512 VSS.n1511 0.120292
R5218 VSS.n1511 VSS.n1364 0.120292
R5219 VSS.n1506 VSS.n1364 0.120292
R5220 VSS.n1506 VSS.n1505 0.120292
R5221 VSS.n1505 VSS.n1504 0.120292
R5222 VSS.n1504 VSS.n1367 0.120292
R5223 VSS.n1498 VSS.n1497 0.120292
R5224 VSS.n1481 VSS.n1480 0.120292
R5225 VSS.n1480 VSS.n1479 0.120292
R5226 VSS.n1479 VSS.n1390 0.120292
R5227 VSS.n1473 VSS.n1390 0.120292
R5228 VSS.n1473 VSS.n1472 0.120292
R5229 VSS.n1472 VSS.n1471 0.120292
R5230 VSS.n1471 VSS.n1395 0.120292
R5231 VSS.n1464 VSS.n1395 0.120292
R5232 VSS.n1464 VSS.n1463 0.120292
R5233 VSS.n1463 VSS.n1462 0.120292
R5234 VSS.n1450 VSS.n1411 0.120292
R5235 VSS.n1444 VSS.n1443 0.120292
R5236 VSS.n1443 VSS.n1417 0.120292
R5237 VSS.n1436 VSS.n1417 0.120292
R5238 VSS.n2639 VSS.n2638 0.120292
R5239 VSS.n2638 VSS.n775 0.120292
R5240 VSS.n2632 VSS.n775 0.120292
R5241 VSS.n2632 VSS.n2631 0.120292
R5242 VSS.n2631 VSS.n2630 0.120292
R5243 VSS.n2630 VSS.n778 0.120292
R5244 VSS.n2623 VSS.n2622 0.120292
R5245 VSS.n2622 VSS.n782 0.120292
R5246 VSS.n2617 VSS.n782 0.120292
R5247 VSS.n817 VSS.n816 0.120292
R5248 VSS.n816 VSS.n805 0.120292
R5249 VSS.n810 VSS.n805 0.120292
R5250 VSS.n1719 VSS.n1718 0.120292
R5251 VSS.n1712 VSS.n1550 0.120292
R5252 VSS.n1707 VSS.n1550 0.120292
R5253 VSS.n1707 VSS.n1706 0.120292
R5254 VSS.n1706 VSS.n1553 0.120292
R5255 VSS.n1698 VSS.n1553 0.120292
R5256 VSS.n1697 VSS.n1696 0.120292
R5257 VSS.n1682 VSS.n1567 0.120292
R5258 VSS.n1676 VSS.n1567 0.120292
R5259 VSS.n1676 VSS.n1675 0.120292
R5260 VSS.n1675 VSS.n1576 0.120292
R5261 VSS.n1668 VSS.n1667 0.120292
R5262 VSS.n1667 VSS.n1579 0.120292
R5263 VSS.n1659 VSS.n1584 0.120292
R5264 VSS.n1639 VSS.n1638 0.120292
R5265 VSS.n1638 VSS.n1602 0.120292
R5266 VSS.n1634 VSS.n1602 0.120292
R5267 VSS.n1634 VSS.n1633 0.120292
R5268 VSS.n1633 VSS.n1632 0.120292
R5269 VSS.n1632 VSS.n1607 0.120292
R5270 VSS.n2603 VSS.n834 0.120292
R5271 VSS.n837 VSS.n834 0.120292
R5272 VSS.n2591 VSS.n2590 0.120292
R5273 VSS.n2590 VSS.n2589 0.120292
R5274 VSS.n921 VSS.n852 0.120292
R5275 VSS.n855 VSS.n852 0.120292
R5276 VSS.n856 VSS.n855 0.120292
R5277 VSS.n914 VSS.n856 0.120292
R5278 VSS.n914 VSS.n913 0.120292
R5279 VSS.n913 VSS.n912 0.120292
R5280 VSS.n912 VSS.n858 0.120292
R5281 VSS.n907 VSS.n858 0.120292
R5282 VSS.n907 VSS.n906 0.120292
R5283 VSS.n892 VSS.n873 0.120292
R5284 VSS.n1841 VSS.n1840 0.120292
R5285 VSS.n1849 VSS.n1287 0.120292
R5286 VSS.n1855 VSS.n1287 0.120292
R5287 VSS.n1856 VSS.n1855 0.120292
R5288 VSS.n1857 VSS.n1856 0.120292
R5289 VSS.n1862 VSS.n1861 0.120292
R5290 VSS.n1885 VSS.n1884 0.120292
R5291 VSS.n1886 VSS.n1885 0.120292
R5292 VSS.n1893 VSS.n1269 0.120292
R5293 VSS.n1894 VSS.n1893 0.120292
R5294 VSS.n1980 VSS.n1239 0.120292
R5295 VSS.n1975 VSS.n1239 0.120292
R5296 VSS.n1974 VSS.n1973 0.120292
R5297 VSS.n1966 VSS.n1246 0.120292
R5298 VSS.n1964 VSS.n1247 0.120292
R5299 VSS.n1960 VSS.n1247 0.120292
R5300 VSS.n1960 VSS.n1959 0.120292
R5301 VSS.n1948 VSS.n1261 0.120292
R5302 VSS.n1943 VSS.n1261 0.120292
R5303 VSS.n1942 VSS.n1941 0.120292
R5304 VSS.n1941 VSS.n1266 0.120292
R5305 VSS.n1934 VSS.n1266 0.120292
R5306 VSS.n1934 VSS.n1933 0.120292
R5307 VSS.n2557 VSS.n935 0.120292
R5308 VSS.n2557 VSS.n2556 0.120292
R5309 VSS.n2556 VSS.n938 0.120292
R5310 VSS.n2552 VSS.n938 0.120292
R5311 VSS.n2552 VSS.n2551 0.120292
R5312 VSS.n2551 VSS.n2550 0.120292
R5313 VSS.n2550 VSS.n941 0.120292
R5314 VSS.n2546 VSS.n2545 0.120292
R5315 VSS.n2545 VSS.n945 0.120292
R5316 VSS.n978 VSS.n959 0.120292
R5317 VSS.n974 VSS.n959 0.120292
R5318 VSS.n974 VSS.n973 0.120292
R5319 VSS.n973 VSS.n965 0.120292
R5320 VSS.n1821 VSS.n1759 0.120292
R5321 VSS.n1820 VSS.n1819 0.120292
R5322 VSS.n1819 VSS.n1761 0.120292
R5323 VSS.n1815 VSS.n1814 0.120292
R5324 VSS.n1814 VSS.n1764 0.120292
R5325 VSS.n1808 VSS.n1764 0.120292
R5326 VSS.n1793 VSS.n1778 0.120292
R5327 VSS.n1786 VSS.n1785 0.120292
R5328 VSS.n2027 VSS.n2026 0.120292
R5329 VSS.n2009 VSS.n2008 0.120292
R5330 VSS.n2004 VSS.n2003 0.120292
R5331 VSS.n2003 VSS.n1994 0.120292
R5332 VSS.n2511 VSS.n995 0.120292
R5333 VSS.n2506 VSS.n995 0.120292
R5334 VSS.n2506 VSS.n2505 0.120292
R5335 VSS.n2501 VSS.n2500 0.120292
R5336 VSS.n2496 VSS.n2495 0.120292
R5337 VSS.n2495 VSS.n2398 0.120292
R5338 VSS.n2481 VSS.n2410 0.120292
R5339 VSS.n2470 VSS.n2469 0.120292
R5340 VSS.n2465 VSS.n2464 0.120292
R5341 VSS.n2464 VSS.n2415 0.120292
R5342 VSS.n2445 VSS.n2433 0.120292
R5343 VSS.n2441 VSS.n2440 0.120292
R5344 VSS.n2440 VSS.n2436 0.120292
R5345 VSS.n3041 VSS.n239 0.120292
R5346 VSS.n3034 VSS.n239 0.120292
R5347 VSS.n3033 VSS.n3032 0.120292
R5348 VSS.n3032 VSS.n257 0.120292
R5349 VSS.n3028 VSS.n257 0.120292
R5350 VSS.n3028 VSS.n3027 0.120292
R5351 VSS.n3027 VSS.n3026 0.120292
R5352 VSS.n3026 VSS.n260 0.120292
R5353 VSS.n3019 VSS.n260 0.120292
R5354 VSS.n3001 VSS.n3000 0.120292
R5355 VSS.n3000 VSS.n274 0.120292
R5356 VSS.n2996 VSS.n274 0.120292
R5357 VSS.n2996 VSS.n2995 0.120292
R5358 VSS.n2995 VSS.n276 0.120292
R5359 VSS.n2991 VSS.n276 0.120292
R5360 VSS.n2991 VSS.n2990 0.120292
R5361 VSS.n1063 VSS.n1058 0.120292
R5362 VSS.n1113 VSS.n1054 0.120292
R5363 VSS.n1109 VSS.n1054 0.120292
R5364 VSS.n1109 VSS.n1108 0.120292
R5365 VSS.n1108 VSS.n1107 0.120292
R5366 VSS.n1107 VSS.n1078 0.120292
R5367 VSS.n1102 VSS.n1078 0.120292
R5368 VSS.n1102 VSS.n1101 0.120292
R5369 VSS.n1101 VSS.n1100 0.120292
R5370 VSS.n1100 VSS 0.120292
R5371 VSS.n1095 VSS.n1094 0.120292
R5372 VSS.n2973 VSS.n2972 0.120292
R5373 VSS.n2973 VSS.n498 0.120292
R5374 VSS.n2977 VSS.n498 0.120292
R5375 VSS.n2978 VSS.n2977 0.120292
R5376 VSS.n2978 VSS.n496 0.120292
R5377 VSS.n2982 VSS.n496 0.120292
R5378 VSS.n2983 VSS.n2982 0.120292
R5379 VSS.n1041 VSS.n1040 0.120292
R5380 VSS.n2321 VSS.n1033 0.120292
R5381 VSS.n2329 VSS.n1033 0.120292
R5382 VSS.n2330 VSS.n2329 0.120292
R5383 VSS.n2335 VSS.n2334 0.120292
R5384 VSS.n2340 VSS.n1029 0.120292
R5385 VSS.n2341 VSS.n2340 0.120292
R5386 VSS.n2342 VSS.n2341 0.120292
R5387 VSS.n2366 VSS.n2365 0.120292
R5388 VSS.n2365 VSS.n2348 0.120292
R5389 VSS.n2361 VSS.n2348 0.120292
R5390 VSS.n2361 VSS.n2360 0.120292
R5391 VSS.n2357 VSS.n2356 0.120292
R5392 VSS.n2356 VSS.n2352 0.120292
R5393 VSS.n1531 VSS.n826 0.120125
R5394 VSS.n2609 VSS.n826 0.120125
R5395 VSS.n2610 VSS.n2609 0.120125
R5396 VSS.n2611 VSS.n2610 0.120125
R5397 VSS.n1830 VSS.n983 0.120125
R5398 VSS.n2527 VSS.n983 0.120125
R5399 VSS.n2528 VSS.n2527 0.120125
R5400 VSS.n2529 VSS.n2528 0.120125
R5401 VSS.n1178 VSS.n505 0.120125
R5402 VSS.n2966 VSS.n505 0.120125
R5403 VSS.n2966 VSS.n2965 0.120125
R5404 VSS.n2965 VSS.n506 0.120125
R5405 VSS.n2150 VSS.n568 0.120125
R5406 VSS.n2923 VSS.n568 0.120125
R5407 VSS.n2924 VSS.n2923 0.120125
R5408 VSS.n2925 VSS.n2924 0.120125
R5409 VSS.n758 VSS.n757 0.120125
R5410 VSS.n757 VSS.n670 0.120125
R5411 VSS.n2872 VSS.n670 0.120125
R5412 VSS.n2872 VSS.n2871 0.120125
R5413 VSS.n2658 VSS.n2657 0.120125
R5414 VSS.n2657 VSS.n2656 0.120125
R5415 VSS.n2656 VSS.n2655 0.120125
R5416 VSS.n2655 VSS.n761 0.120125
R5417 VSS.n116 VSS 0.114397
R5418 VSS.n330 VSS.n329 0.113648
R5419 VSS.n3383 VSS.n78 0.113648
R5420 VSS.n229 VSS 0.11275
R5421 VSS.n130 VSS.n129 0.111077
R5422 VSS.n135 VSS.n134 0.111077
R5423 VSS.n140 VSS.n139 0.111077
R5424 VSS.n145 VSS.n144 0.111077
R5425 VSS.n150 VSS.n149 0.111077
R5426 VSS.n155 VSS.n154 0.111077
R5427 VSS.n160 VSS.n159 0.111077
R5428 VSS.n165 VSS.n164 0.111077
R5429 VSS.n170 VSS.n169 0.111077
R5430 VSS.n2795 VSS.n2794 0.109992
R5431 VSS.n2304 VSS.n2303 0.10744
R5432 VSS.n2922 VSS.n2921 0.103312
R5433 VSS.n2091 VSS.n1118 0.103312
R5434 VSS.n2123 VSS.n1163 0.103312
R5435 VSS.n2151 VSS.n2149 0.103312
R5436 VSS.n2874 VSS.n509 0.103312
R5437 VSS.n2926 VSS.n567 0.103312
R5438 VSS.n1513 VSS.n1306 0.102062
R5439 VSS.n1683 VSS.n1682 0.102062
R5440 VSS.n1880 VSS.n1879 0.102062
R5441 VSS.n1794 VSS.n1793 0.102062
R5442 VSS.n3006 VSS.n3001 0.102062
R5443 VSS.n11 VSS 0.0981562
R5444 VSS.n3091 VSS 0.0981562
R5445 VSS VSS.n114 0.0981562
R5446 VSS.n2203 VSS 0.0981562
R5447 VSS.n2222 VSS 0.0981562
R5448 VSS.n2235 VSS 0.0981562
R5449 VSS.n2936 VSS 0.0981562
R5450 VSS VSS.n2119 0.0981562
R5451 VSS.n2040 VSS 0.0981562
R5452 VSS.n2066 VSS 0.0981562
R5453 VSS.n2902 VSS 0.0981562
R5454 VSS.n583 VSS 0.0981562
R5455 VSS.n2710 VSS 0.0981562
R5456 VSS.n2724 VSS 0.0981562
R5457 VSS.n2789 VSS 0.0981562
R5458 VSS VSS.n679 0.0981562
R5459 VSS VSS.n1309 0.0981562
R5460 VSS.n1481 VSS 0.0981562
R5461 VSS.n1427 VSS 0.0981562
R5462 VSS.n2623 VSS 0.0981562
R5463 VSS.n1627 VSS 0.0981562
R5464 VSS.n1848 VSS 0.0981562
R5465 VSS.n1884 VSS 0.0981562
R5466 VSS VSS.n1964 0.0981562
R5467 VSS.n1923 VSS 0.0981562
R5468 VSS.n279 VSS 0.0981562
R5469 VSS.n1095 VSS 0.0981562
R5470 VSS VSS.n494 0.0981562
R5471 VSS.n2357 VSS 0.0981562
R5472 VSS.n2949 VSS.n516 0.0968542
R5473 VSS.n666 VSS.n665 0.0968542
R5474 VSS.n2812 VSS.n2811 0.0968542
R5475 VSS.n2639 VSS.n770 0.0968542
R5476 VSS VSS.n1639 0.0968542
R5477 VSS.n1861 VSS 0.0968542
R5478 VSS.n2482 VSS.n2481 0.0968542
R5479 VSS.n2321 VSS.n2320 0.0968542
R5480 VSS.n1759 VSS 0.0955521
R5481 VSS VSS.n1806 0.0955521
R5482 VSS VSS.n1786 0.0955521
R5483 VSS VSS.n2009 0.0955521
R5484 VSS VSS.n2501 0.0955521
R5485 VSS VSS.n2470 0.0955521
R5486 VSS VSS.n2445 0.0955521
R5487 VSS.n2334 VSS 0.0955521
R5488 VSS.n2311 VSS.n1046 0.0950946
R5489 VSS.n2319 VSS.n2318 0.0950946
R5490 VSS.n249 VSS.n243 0.0950946
R5491 VSS.n3043 VSS.n238 0.0950946
R5492 VSS.n2570 VSS.n2569 0.0950946
R5493 VSS.n2563 VSS.n931 0.0950946
R5494 VSS.n1067 VSS.n1057 0.0950946
R5495 VSS.n1115 VSS.n1052 0.0950946
R5496 VSS.n2578 VSS.n2577 0.0950946
R5497 VSS.n2583 VSS.n2582 0.0950946
R5498 VSS.n1086 VSS.n1085 0.0950946
R5499 VSS.n2970 VSS.n501 0.0950946
R5500 VSS.n2961 VSS.n2960 0.0950946
R5501 VSS.n2954 VSS.n515 0.0950946
R5502 VSS.n2290 VSS.n2289 0.0950946
R5503 VSS.n2284 VSS.n2283 0.0950946
R5504 VSS.n2194 VSS.n2193 0.0950946
R5505 VSS.n2198 VSS.n1160 0.0950946
R5506 VSS.n2163 VSS.n2162 0.0950946
R5507 VSS.n2168 VSS.n1176 0.0950946
R5508 VSS.n2929 VSS.n528 0.0950946
R5509 VSS.n565 VSS.n532 0.0950946
R5510 VSS.n2257 VSS.n1134 0.0950946
R5511 VSS.n2252 VSS.n1137 0.0950946
R5512 VSS.n2127 VSS.n1207 0.0950946
R5513 VSS.n2121 VSS.n1211 0.0950946
R5514 VSS.n2147 VSS.n2146 0.0950946
R5515 VSS.n1194 VSS.n1193 0.0950946
R5516 VSS.n645 VSS.n606 0.0950946
R5517 VSS.n640 VSS.n609 0.0950946
R5518 VSS.n2878 VSS.n587 0.0950946
R5519 VSS.n667 VSS.n591 0.0950946
R5520 VSS.n2095 VSS.n2045 0.0950946
R5521 VSS.n2089 VSS.n2049 0.0950946
R5522 VSS.n2919 VSS.n2918 0.0950946
R5523 VSS.n2911 VSS.n2910 0.0950946
R5524 VSS.n2701 VSS.n2700 0.0950946
R5525 VSS.n2705 VSS.n739 0.0950946
R5526 VSS.n2671 VSS.n2670 0.0950946
R5527 VSS.n2675 VSS.n755 0.0950946
R5528 VSS.n2867 VSS.n2866 0.0950946
R5529 VSS.n2859 VSS.n2858 0.0950946
R5530 VSS.n2798 VSS.n2797 0.0950946
R5531 VSS.n2810 VSS.n686 0.0950946
R5532 VSS.n2733 VSS.n2732 0.0950946
R5533 VSS.n2737 VSS.n720 0.0950946
R5534 VSS.n2769 VSS.n2768 0.0950946
R5535 VSS.n2773 VSS.n700 0.0950946
R5536 VSS.n1326 VSS.n1323 0.0950946
R5537 VSS.n1335 VSS.n1315 0.0950946
R5538 VSS.n2615 VSS.n787 0.0950946
R5539 VSS.n823 VSS.n790 0.0950946
R5540 VSS.n2651 VSS.n2650 0.0950946
R5541 VSS.n2644 VSS.n769 0.0950946
R5542 VSS.n1383 VSS.n1382 0.0950946
R5543 VSS.n1487 VSS.n1378 0.0950946
R5544 VSS.n1527 VSS.n1526 0.0950946
R5545 VSS.n1520 VSS.n1305 0.0950946
R5546 VSS.n1407 VSS.n1406 0.0950946
R5547 VSS.n1452 VSS.n1405 0.0950946
R5548 VSS.n1257 VSS.n1256 0.0950946
R5549 VSS.n1950 VSS.n1255 0.0950946
R5550 VSS.n2523 VSS.n2522 0.0950946
R5551 VSS.n2515 VSS.n2514 0.0950946
R5552 VSS.n1617 VSS.n1616 0.0950946
R5553 VSS.n2605 VSS.n832 0.0950946
R5554 VSS.n1690 VSS.n1562 0.0950946
R5555 VSS.n1684 VSS.n1565 0.0950946
R5556 VSS.n1725 VSS.n1724 0.0950946
R5557 VSS.n1547 VSS.n1546 0.0950946
R5558 VSS.n900 VSS.n866 0.0950946
R5559 VSS.n894 VSS.n869 0.0950946
R5560 VSS.n1651 VSS.n1590 0.0950946
R5561 VSS.n1645 VSS.n1593 0.0950946
R5562 VSS.n2021 VSS.n1230 0.0950946
R5563 VSS.n2015 VSS.n1987 0.0950946
R5564 VSS.n1909 VSS.n1908 0.0950946
R5565 VSS.n1982 VSS.n1237 0.0950946
R5566 VSS.n1835 VSS.n1296 0.0950946
R5567 VSS.n1735 VSS.n1734 0.0950946
R5568 VSS.n2535 VSS.n951 0.0950946
R5569 VSS.n980 VSS.n955 0.0950946
R5570 VSS.n1874 VSS.n1873 0.0950946
R5571 VSS.n1878 VSS.n1275 0.0950946
R5572 VSS.n1801 VSS.n1769 0.0950946
R5573 VSS.n1795 VSS.n1773 0.0950946
R5574 VSS.n1749 VSS.n1743 0.0950946
R5575 VSS.n1827 VSS.n1740 0.0950946
R5576 VSS.n2427 VSS.n2426 0.0950946
R5577 VSS.n2452 VSS.n2423 0.0950946
R5578 VSS.n2489 VSS.n2402 0.0950946
R5579 VSS.n2483 VSS.n2406 0.0950946
R5580 VSS.n2374 VSS.n2373 0.0950946
R5581 VSS.n2346 VSS.n1022 0.0950946
R5582 VSS.n3016 VSS.n266 0.0950946
R5583 VSS.n3005 VSS.n3002 0.0950946
R5584 VSS.n52 VSS 0.09425
R5585 VSS.n3142 VSS 0.09425
R5586 VSS VSS.n3307 0.09425
R5587 VSS.n3168 VSS.n3166 0.0934947
R5588 VSS.n2931 VSS.n2930 0.0916458
R5589 VSS.n647 VSS.n646 0.0916458
R5590 VSS.n2617 VSS.n2616 0.0916458
R5591 VSS.n864 VSS.n862 0.0916458
R5592 VSS.n2342 VSS.n1024 0.0916458
R5593 VSS.n2921 VSS.n570 0.0915625
R5594 VSS.n2091 VSS.n722 0.0915625
R5595 VSS.n2123 VSS.n741 0.0915625
R5596 VSS.n2149 VSS.n759 0.0915625
R5597 VSS.n2874 VSS.n2873 0.0915625
R5598 VSS.n2870 VSS.n567 0.0915625
R5599 VSS.n2378 VSS 0.0907344
R5600 VSS.n129 VSS 0.0906442
R5601 VSS.n134 VSS 0.0906442
R5602 VSS.n139 VSS 0.0906442
R5603 VSS.n144 VSS 0.0906442
R5604 VSS.n149 VSS 0.0906442
R5605 VSS.n154 VSS 0.0906442
R5606 VSS.n159 VSS 0.0906442
R5607 VSS.n164 VSS 0.0906442
R5608 VSS.n169 VSS 0.0906442
R5609 VSS.n2937 VSS.n523 0.0900105
R5610 VSS.n2814 VSS.n2813 0.0900105
R5611 VSS.n2302 VSS.n2298 0.0898892
R5612 VSS.n2303 VSS.n1049 0.0898892
R5613 VSS.n3434 VSS 0.0881354
R5614 VSS.n3165 VSS 0.0881354
R5615 VSS.n79 VSS 0.0881354
R5616 VSS.n2220 VSS.n1120 0.0864375
R5617 VSS.n2101 VSS.n2041 0.0864375
R5618 VSS.n2728 VSS.n725 0.0864375
R5619 VSS.n1588 VSS.n1584 0.0864375
R5620 VSS.n2026 VSS.n1226 0.0864375
R5621 VSS.n1064 VSS.n1063 0.0864375
R5622 VSS.n3468 VSS.n0 0.0853293
R5623 VSS.n2192 VSS.n2191 0.0838333
R5624 VSS.n1126 VSS.n1122 0.0838333
R5625 VSS.n2251 VSS.n1138 0.0838333
R5626 VSS.n2959 VSS.n2958 0.0838333
R5627 VSS.n543 VSS.n542 0.0838333
R5628 VSS.n2128 VSS.n1206 0.0838333
R5629 VSS.n2051 VSS.n2050 0.0838333
R5630 VSS.n2917 VSS.n572 0.0838333
R5631 VSS.n2912 VSS.n2906 0.0838333
R5632 VSS.n634 VSS.n633 0.0838333
R5633 VSS.n2699 VSS.n2698 0.0838333
R5634 VSS.n727 VSS.n719 0.0838333
R5635 VSS.n2774 VSS.n699 0.0838333
R5636 VSS.n2838 VSS.n677 0.0838333
R5637 VSS.n1525 VSS.n1524 0.0838333
R5638 VSS.n1492 VSS.n1376 0.0838333
R5639 VSS.n1402 VSS.n1399 0.0838333
R5640 VSS.n1451 VSS.n1410 0.0838333
R5641 VSS.n2649 VSS.n2648 0.0838333
R5642 VSS.n799 VSS.n795 0.0838333
R5643 VSS.n1691 VSS.n1561 0.0838333
R5644 VSS.n1595 VSS.n1594 0.0838333
R5645 VSS.n1614 VSS.n1613 0.0838333
R5646 VSS.n2604 VSS.n833 0.0838333
R5647 VSS.n2576 VSS.n849 0.0838333
R5648 VSS.n1872 VSS.n1871 0.0838333
R5649 VSS.n1903 VSS.n1900 0.0838333
R5650 VSS.n1949 VSS.n1260 0.0838333
R5651 VSS.n2568 VSS.n2567 0.0838333
R5652 VSS.n1989 VSS.n1988 0.0838333
R5653 VSS.n2490 VSS.n2401 0.0838333
R5654 VSS.n3011 VSS.n269 0.0838333
R5655 VSS.n1072 VSS.n1056 0.0838333
R5656 VSS.n1083 VSS.n1081 0.0838333
R5657 VSS.n2971 VSS.n500 0.0838333
R5658 VSS.n2312 VSS.n1038 0.0838333
R5659 VSS.n2347 VSS.n1027 0.0838333
R5660 VSS.n2611 VSS 0.0827875
R5661 VSS.n2529 VSS 0.0827875
R5662 VSS.n506 VSS 0.0827875
R5663 VSS.n2925 VSS 0.0827875
R5664 VSS.n2871 VSS 0.0827875
R5665 VSS.n761 VSS 0.0827875
R5666 VSS VSS.n880 0.082648
R5667 VSS.n1713 VSS 0.082648
R5668 VSS.n2430 VSS 0.0773229
R5669 VSS.n3054 VSS.n228 0.0766574
R5670 VSS.n3201 VSS.n181 0.0766574
R5671 VSS.n1167 VSS.n1165 0.0760208
R5672 VSS.n2129 VSS.n1203 0.0760208
R5673 VSS.n746 VSS.n744 0.0760208
R5674 VSS.n1303 VSS.n1301 0.0760208
R5675 VSS.n1692 VSS.n1557 0.0760208
R5676 VSS.n1282 VSS.n1280 0.0760208
R5677 VSS.n1803 VSS.n1766 0.0760208
R5678 VSS.n3017 VSS.n265 0.0760208
R5679 VSS.n2377 VSS.n1016 0.0747188
R5680 VSS.n3439 VSS.n3435 0.0721146
R5681 VSS.n101 VSS.n96 0.0721146
R5682 VSS.n3164 VSS.n210 0.0708554
R5683 VSS.n3458 VSS.n17 0.0708125
R5684 VSS.n3132 VSS.n3131 0.0708125
R5685 VSS.n3331 VSS.n111 0.0708125
R5686 VSS.n2159 VSS.n2156 0.0708125
R5687 VSS.n2288 VSS.n2287 0.0708125
R5688 VSS.n513 VSS.n511 0.0708125
R5689 VSS.n1186 VSS.n1184 0.0708125
R5690 VSS.n2096 VSS.n2044 0.0708125
R5691 VSS.n2880 VSS.n586 0.0708125
R5692 VSS.n2667 VSS.n2664 0.0708125
R5693 VSS.n2731 VSS.n716 0.0708125
R5694 VSS.n2800 VSS.n2795 0.0708125
R5695 VSS.n1330 VSS.n1329 0.0708125
R5696 VSS.n1493 VSS.n1375 0.0708125
R5697 VSS.n767 VSS.n765 0.0708125
R5698 VSS.n1539 VSS.n1537 0.0708125
R5699 VSS.n1652 VSS.n1589 0.0708125
R5700 VSS.n847 VSS.n846 0.0708125
R5701 VSS.n1730 VSS.n1293 0.0708125
R5702 VSS.n1907 VSS.n1906 0.0708125
R5703 VSS.n1756 VSS.n1754 0.0708125
R5704 VSS.n2022 VSS.n1229 0.0708125
R5705 VSS.n2491 VSS.n2400 0.0708125
R5706 VSS.n254 VSS.n252 0.0708125
R5707 VSS.n2313 VSS.n1045 0.0708125
R5708 VSS.n1141 VSS 0.0695104
R5709 VSS.n2767 VSS 0.0695104
R5710 VSS.n2771 VSS.n570 0.0692375
R5711 VSS.n2735 VSS.n722 0.0692375
R5712 VSS.n2703 VSS.n741 0.0692375
R5713 VSS.n2673 VSS.n759 0.0692375
R5714 VSS.n2873 VSS.n669 0.0692375
R5715 VSS.n2870 VSS.n2869 0.0692375
R5716 VSS.n1439 VSS.n1438 0.0685851
R5717 VSS.n2259 VSS.n2258 0.068325
R5718 VSS.n709 VSS.n704 0.068325
R5719 VSS.n2310 VSS.n1047 0.0680676
R5720 VSS.n1047 VSS.n1037 0.0680676
R5721 VSS.n251 VSS.n250 0.0680676
R5722 VSS.n251 VSS.n236 0.0680676
R5723 VSS.n2566 VSS.n928 0.0680676
R5724 VSS.n2566 VSS.n2565 0.0680676
R5725 VSS.n1071 VSS.n1069 0.0680676
R5726 VSS.n1071 VSS.n1070 0.0680676
R5727 VSS.n2575 VSS.n2574 0.0680676
R5728 VSS.n2574 VSS.n851 0.0680676
R5729 VSS.n1089 VSS.n1087 0.0680676
R5730 VSS.n1089 VSS.n1088 0.0680676
R5731 VSS.n2957 VSS.n512 0.0680676
R5732 VSS.n2957 VSS.n2956 0.0680676
R5733 VSS.n2280 VSS.n1121 0.0680676
R5734 VSS.n2282 VSS.n2280 0.0680676
R5735 VSS.n2190 VSS.n1166 0.0680676
R5736 VSS.n2190 VSS.n2189 0.0680676
R5737 VSS.n2158 VSS.n2154 0.0680676
R5738 VSS.n2158 VSS.n2157 0.0680676
R5739 VSS.n541 VSS.n539 0.0680676
R5740 VSS.n541 VSS.n540 0.0680676
R5741 VSS.n1144 VSS.n1135 0.0680676
R5742 VSS.n1144 VSS.n1136 0.0680676
R5743 VSS.n2126 VSS.n1208 0.0680676
R5744 VSS.n1210 VSS.n1208 0.0680676
R5745 VSS.n1189 VSS.n1183 0.0680676
R5746 VSS.n1191 VSS.n1189 0.0680676
R5747 VSS.n632 VSS.n607 0.0680676
R5748 VSS.n632 VSS.n608 0.0680676
R5749 VSS.n2877 VSS.n588 0.0680676
R5750 VSS.n590 VSS.n588 0.0680676
R5751 VSS.n2094 VSS.n2046 0.0680676
R5752 VSS.n2048 VSS.n2046 0.0680676
R5753 VSS.n2907 VSS.n573 0.0680676
R5754 VSS.n2909 VSS.n2907 0.0680676
R5755 VSS.n2697 VSS.n745 0.0680676
R5756 VSS.n2697 VSS.n2696 0.0680676
R5757 VSS.n2666 VSS.n2662 0.0680676
R5758 VSS.n2666 VSS.n2665 0.0680676
R5759 VSS.n2855 VSS.n675 0.0680676
R5760 VSS.n2857 VSS.n2855 0.0680676
R5761 VSS.n2806 VSS.n688 0.0680676
R5762 VSS.n2807 VSS.n2806 0.0680676
R5763 VSS.n729 VSS.n728 0.0680676
R5764 VSS.n728 VSS.n726 0.0680676
R5765 VSS.n707 VSS.n705 0.0680676
R5766 VSS.n707 VSS.n706 0.0680676
R5767 VSS.n1331 VSS.n1317 0.0680676
R5768 VSS.n1332 VSS.n1331 0.0680676
R5769 VSS.n798 VSS.n796 0.0680676
R5770 VSS.n798 VSS.n797 0.0680676
R5771 VSS.n2647 VSS.n766 0.0680676
R5772 VSS.n2647 VSS.n2646 0.0680676
R5773 VSS.n1491 VSS.n1377 0.0680676
R5774 VSS.n1491 VSS.n1490 0.0680676
R5775 VSS.n1523 VSS.n1302 0.0680676
R5776 VSS.n1523 VSS.n1522 0.0680676
R5777 VSS.n1456 VSS.n1404 0.0680676
R5778 VSS.n1456 VSS.n1455 0.0680676
R5779 VSS.n1954 VSS.n1254 0.0680676
R5780 VSS.n1954 VSS.n1953 0.0680676
R5781 VSS.n992 VSS.n987 0.0680676
R5782 VSS.n994 VSS.n992 0.0680676
R5783 VSS.n1621 VSS.n1619 0.0680676
R5784 VSS.n1621 VSS.n1620 0.0680676
R5785 VSS.n1689 VSS.n1563 0.0680676
R5786 VSS.n1564 VSS.n1563 0.0680676
R5787 VSS.n1542 VSS.n1536 0.0680676
R5788 VSS.n1544 VSS.n1542 0.0680676
R5789 VSS.n899 VSS.n867 0.0680676
R5790 VSS.n868 VSS.n867 0.0680676
R5791 VSS.n1650 VSS.n1591 0.0680676
R5792 VSS.n1592 VSS.n1591 0.0680676
R5793 VSS.n2020 VSS.n1231 0.0680676
R5794 VSS.n1986 VSS.n1231 0.0680676
R5795 VSS.n1902 VSS.n1899 0.0680676
R5796 VSS.n1902 VSS.n1901 0.0680676
R5797 VSS.n1731 VSS.n1729 0.0680676
R5798 VSS.n1732 VSS.n1731 0.0680676
R5799 VSS.n2534 VSS.n952 0.0680676
R5800 VSS.n954 VSS.n952 0.0680676
R5801 VSS.n1870 VSS.n1281 0.0680676
R5802 VSS.n1870 VSS.n1869 0.0680676
R5803 VSS.n1800 VSS.n1770 0.0680676
R5804 VSS.n1772 VSS.n1770 0.0680676
R5805 VSS.n1753 VSS.n1751 0.0680676
R5806 VSS.n1753 VSS.n1752 0.0680676
R5807 VSS.n2456 VSS.n2422 0.0680676
R5808 VSS.n2456 VSS.n2455 0.0680676
R5809 VSS.n2488 VSS.n2403 0.0680676
R5810 VSS.n2405 VSS.n2403 0.0680676
R5811 VSS.n1026 VSS.n1021 0.0680676
R5812 VSS.n1026 VSS.n1020 0.0680676
R5813 VSS.n3013 VSS.n3012 0.0680676
R5814 VSS.n3012 VSS.n268 0.0680676
R5815 VSS.n2521 VSS 0.0669062
R5816 VSS.n2200 VSS.n1159 0.0656042
R5817 VSS.n1146 VSS.n1145 0.0656042
R5818 VSS.n538 VSS.n534 0.0656042
R5819 VSS.n1214 VSS.n1213 0.0656042
R5820 VSS.n2913 VSS.n574 0.0656042
R5821 VSS.n631 VSS.n630 0.0656042
R5822 VSS.n2707 VSS.n738 0.0656042
R5823 VSS.n2762 VSS.n708 0.0656042
R5824 VSS.n2865 VSS.n2864 0.0656042
R5825 VSS.n2861 VSS.n2860 0.0656042
R5826 VSS.n1519 VSS.n1518 0.0656042
R5827 VSS.n1457 VSS.n1403 0.0656042
R5828 VSS.n800 VSS.n794 0.0656042
R5829 VSS.n822 VSS.n791 0.0656042
R5830 VSS.n1568 VSS.n1566 0.0656042
R5831 VSS.n1622 VSS.n1615 0.0656042
R5832 VSS.n901 VSS.n865 0.0656042
R5833 VSS.n893 VSS.n872 0.0656042
R5834 VSS.n1283 VSS.n1274 0.0656042
R5835 VSS.n1955 VSS.n1253 0.0656042
R5836 VSS.n2536 VSS.n950 0.0656042
R5837 VSS.n979 VSS.n958 0.0656042
R5838 VSS.n2517 VSS.n988 0.0656042
R5839 VSS.n2451 VSS.n2431 0.0656042
R5840 VSS.n3007 VSS.n270 0.0656042
R5841 VSS.n1090 VSS.n1084 0.0656042
R5842 VSS.n2372 VSS.n2371 0.0656042
R5843 VSS.n2368 VSS.n2367 0.0656042
R5844 VSS.n227 VSS 0.064875
R5845 VSS.n288 VSS 0.064875
R5846 VSS.n287 VSS 0.064875
R5847 VSS.n327 VSS 0.064875
R5848 VSS.n331 VSS 0.064875
R5849 VSS.n374 VSS 0.064875
R5850 VSS.n351 VSS 0.064875
R5851 VSS.n349 VSS 0.064875
R5852 VSS.n3240 VSS 0.064875
R5853 VSS.n3272 VSS 0.064875
R5854 VSS.n3221 VSS 0.064875
R5855 VSS.n3219 VSS 0.064875
R5856 VSS.n200 VSS 0.064875
R5857 VSS.n3200 VSS 0.064875
R5858 VSS.n3384 VSS 0.064875
R5859 VSS.n3274 VSS 0.064875
R5860 VSS.n2161 VSS 0.0643021
R5861 VSS.n2145 VSS 0.0643021
R5862 VSS.n2669 VSS 0.0643021
R5863 VSS.n1322 VSS 0.0643021
R5864 VSS.n1723 VSS 0.0643021
R5865 VSS.n1295 VSS 0.0643021
R5866 VSS VSS.n1910 0.0643021
R5867 VSS.n1748 VSS 0.0643021
R5868 VSS.n248 VSS 0.0643021
R5869 VSS.n3053 VSS.n3052 0.063797
R5870 VSS.n3068 VSS 0.063625
R5871 VSS.n3048 VSS.n233 0.0635047
R5872 VSS.n3066 VSS 0.063
R5873 VSS.n3432 VSS.n41 0.0616979
R5874 VSS.n3163 VSS.n211 0.0616979
R5875 VSS.n3379 VSS.n80 0.0616979
R5876 VSS.n59 VSS 0.0603958
R5877 VSS VSS.n3425 0.0603958
R5878 VSS.n3409 VSS 0.0603958
R5879 VSS.n3410 VSS 0.0603958
R5880 VSS VSS.n3416 0.0603958
R5881 VSS VSS.n36 0.0603958
R5882 VSS.n3443 VSS 0.0603958
R5883 VSS.n45 VSS 0.0603958
R5884 VSS.n5 VSS 0.0603958
R5885 VSS.n13 VSS 0.0603958
R5886 VSS.n14 VSS 0.0603958
R5887 VSS.n3458 VSS 0.0603958
R5888 VSS VSS.n3457 0.0603958
R5889 VSS VSS.n3456 0.0603958
R5890 VSS.n20 VSS 0.0603958
R5891 VSS.n3450 VSS 0.0603958
R5892 VSS VSS.n34 0.0603958
R5893 VSS.n3135 VSS 0.0603958
R5894 VSS.n3086 VSS 0.0603958
R5895 VSS.n3093 VSS 0.0603958
R5896 VSS VSS.n217 0.0603958
R5897 VSS.n3131 VSS 0.0603958
R5898 VSS.n3127 VSS 0.0603958
R5899 VSS VSS.n3126 0.0603958
R5900 VSS VSS.n3119 0.0603958
R5901 VSS VSS.n3102 0.0603958
R5902 VSS VSS.n3112 0.0603958
R5903 VSS.n3159 VSS 0.0603958
R5904 VSS.n3153 VSS 0.0603958
R5905 VSS.n3188 VSS 0.0603958
R5906 VSS VSS.n3187 0.0603958
R5907 VSS.n3181 VSS 0.0603958
R5908 VSS.n194 VSS 0.0603958
R5909 VSS VSS.n3172 0.0603958
R5910 VSS.n82 VSS 0.0603958
R5911 VSS VSS.n3372 0.0603958
R5912 VSS.n87 VSS 0.0603958
R5913 VSS.n88 VSS 0.0603958
R5914 VSS VSS.n3363 0.0603958
R5915 VSS.n3358 VSS 0.0603958
R5916 VSS VSS.n105 0.0603958
R5917 VSS.n3314 VSS 0.0603958
R5918 VSS.n3318 VSS 0.0603958
R5919 VSS.n3326 VSS 0.0603958
R5920 VSS.n3327 VSS 0.0603958
R5921 VSS VSS.n3331 0.0603958
R5922 VSS.n3332 VSS 0.0603958
R5923 VSS.n3333 VSS 0.0603958
R5924 VSS.n3338 VSS 0.0603958
R5925 VSS.n3339 VSS 0.0603958
R5926 VSS.n3351 VSS 0.0603958
R5927 VSS.n2174 VSS 0.0603958
R5928 VSS.n2183 VSS 0.0603958
R5929 VSS VSS.n2221 0.0603958
R5930 VSS VSS.n2220 0.0603958
R5931 VSS VSS.n2279 0.0603958
R5932 VSS VSS.n2234 0.0603958
R5933 VSS.n2231 VSS 0.0603958
R5934 VSS.n2953 VSS.n514 0.0603958
R5935 VSS.n2953 VSS.n2952 0.0603958
R5936 VSS.n559 VSS 0.0603958
R5937 VSS.n2140 VSS 0.0603958
R5938 VSS VSS.n2133 0.0603958
R5939 VSS.n2102 VSS 0.0603958
R5940 VSS.n2088 VSS.n2052 0.0603958
R5941 VSS.n2088 VSS.n2087 0.0603958
R5942 VSS VSS.n2079 0.0603958
R5943 VSS.n2887 VSS 0.0603958
R5944 VSS.n595 VSS.n594 0.0603958
R5945 VSS.n635 VSS 0.0603958
R5946 VSS.n624 VSS 0.0603958
R5947 VSS VSS.n611 0.0603958
R5948 VSS.n616 VSS 0.0603958
R5949 VSS.n2681 VSS 0.0603958
R5950 VSS.n2690 VSS 0.0603958
R5951 VSS.n2727 VSS 0.0603958
R5952 VSS.n2728 VSS 0.0603958
R5953 VSS VSS.n715 0.0603958
R5954 VSS.n2793 VSS 0.0603958
R5955 VSS.n2804 VSS.n689 0.0603958
R5956 VSS.n689 VSS.n685 0.0603958
R5957 VSS VSS.n683 0.0603958
R5958 VSS.n2825 VSS 0.0603958
R5959 VSS.n2833 VSS 0.0603958
R5960 VSS.n1338 VSS 0.0603958
R5961 VSS.n1342 VSS 0.0603958
R5962 VSS.n1350 VSS 0.0603958
R5963 VSS VSS.n1355 0.0603958
R5964 VSS.n1356 VSS 0.0603958
R5965 VSS VSS.n1512 0.0603958
R5966 VSS.n1499 VSS 0.0603958
R5967 VSS VSS.n1498 0.0603958
R5968 VSS VSS.n1386 0.0603958
R5969 VSS VSS.n1486 0.0603958
R5970 VSS VSS.n1411 0.0603958
R5971 VSS.n1414 VSS 0.0603958
R5972 VSS VSS.n1414 0.0603958
R5973 VSS.n1445 VSS 0.0603958
R5974 VSS VSS.n1444 0.0603958
R5975 VSS VSS.n1435 0.0603958
R5976 VSS VSS.n1434 0.0603958
R5977 VSS.n1426 VSS 0.0603958
R5978 VSS.n2643 VSS.n768 0.0603958
R5979 VSS.n2643 VSS.n2642 0.0603958
R5980 VSS.n821 VSS 0.0603958
R5981 VSS.n817 VSS 0.0603958
R5982 VSS VSS.n1712 0.0603958
R5983 VSS VSS.n1697 0.0603958
R5984 VSS.n1668 VSS 0.0603958
R5985 VSS.n1660 VSS 0.0603958
R5986 VSS VSS.n1659 0.0603958
R5987 VSS.n1644 VSS.n1596 0.0603958
R5988 VSS.n1644 VSS.n1643 0.0603958
R5989 VSS.n1640 VSS 0.0603958
R5990 VSS VSS.n1607 0.0603958
R5991 VSS.n1609 VSS 0.0603958
R5992 VSS VSS.n1626 0.0603958
R5993 VSS VSS.n837 0.0603958
R5994 VSS.n2597 VSS 0.0603958
R5995 VSS VSS.n2595 0.0603958
R5996 VSS.n2591 VSS 0.0603958
R5997 VSS.n2585 VSS.n2584 0.0603958
R5998 VSS.n2584 VSS.n850 0.0603958
R5999 VSS VSS.n921 0.0603958
R6000 VSS.n862 VSS 0.0603958
R6001 VSS.n881 VSS 0.0603958
R6002 VSS.n1847 VSS 0.0603958
R6003 VSS.n1849 VSS 0.0603958
R6004 VSS.n1857 VSS 0.0603958
R6005 VSS.n1860 VSS 0.0603958
R6006 VSS VSS.n1880 0.0603958
R6007 VSS.n1881 VSS 0.0603958
R6008 VSS VSS.n1269 0.0603958
R6009 VSS VSS.n1894 0.0603958
R6010 VSS.n1895 VSS 0.0603958
R6011 VSS.n1912 VSS 0.0603958
R6012 VSS VSS.n1911 0.0603958
R6013 VSS.n1981 VSS.n1238 0.0603958
R6014 VSS.n1981 VSS.n1980 0.0603958
R6015 VSS.n1975 VSS 0.0603958
R6016 VSS VSS.n1974 0.0603958
R6017 VSS.n1246 VSS 0.0603958
R6018 VSS VSS.n1965 0.0603958
R6019 VSS VSS.n1942 0.0603958
R6020 VSS VSS.n1932 0.0603958
R6021 VSS.n1929 VSS 0.0603958
R6022 VSS VSS.n1928 0.0603958
R6023 VSS.n929 VSS 0.0603958
R6024 VSS.n2562 VSS.n930 0.0603958
R6025 VSS.n2562 VSS.n2561 0.0603958
R6026 VSS.n935 VSS 0.0603958
R6027 VSS.n2546 VSS 0.0603958
R6028 VSS.n1821 VSS 0.0603958
R6029 VSS VSS.n1820 0.0603958
R6030 VSS.n1815 VSS 0.0603958
R6031 VSS VSS.n1807 0.0603958
R6032 VSS.n1777 VSS 0.0603958
R6033 VSS.n1787 VSS 0.0603958
R6034 VSS.n1785 VSS 0.0603958
R6035 VSS VSS.n1224 0.0603958
R6036 VSS.n2027 VSS 0.0603958
R6037 VSS.n2014 VSS.n1990 0.0603958
R6038 VSS.n2014 VSS.n2013 0.0603958
R6039 VSS.n2010 VSS 0.0603958
R6040 VSS.n2008 VSS 0.0603958
R6041 VSS.n2005 VSS 0.0603958
R6042 VSS VSS.n2004 0.0603958
R6043 VSS VSS.n1997 0.0603958
R6044 VSS VSS.n2511 0.0603958
R6045 VSS.n2502 VSS 0.0603958
R6046 VSS.n2500 VSS 0.0603958
R6047 VSS.n2396 VSS 0.0603958
R6048 VSS.n2496 VSS 0.0603958
R6049 VSS.n2408 VSS.n2407 0.0603958
R6050 VSS.n2409 VSS.n2408 0.0603958
R6051 VSS.n2471 VSS 0.0603958
R6052 VSS.n2469 VSS 0.0603958
R6053 VSS.n2466 VSS 0.0603958
R6054 VSS VSS.n2465 0.0603958
R6055 VSS.n2458 VSS 0.0603958
R6056 VSS.n2450 VSS 0.0603958
R6057 VSS.n2447 VSS 0.0603958
R6058 VSS VSS.n2446 0.0603958
R6059 VSS VSS.n2433 0.0603958
R6060 VSS.n2441 VSS 0.0603958
R6061 VSS VSS.n3033 0.0603958
R6062 VSS VSS.n3018 0.0603958
R6063 VSS.n1058 VSS 0.0603958
R6064 VSS.n1073 VSS 0.0603958
R6065 VSS.n1114 VSS.n1053 0.0603958
R6066 VSS.n1114 VSS.n1113 0.0603958
R6067 VSS.n1040 VSS 0.0603958
R6068 VSS.n1044 VSS 0.0603958
R6069 VSS.n2317 VSS.n2316 0.0603958
R6070 VSS.n2317 VSS.n1036 0.0603958
R6071 VSS.n2333 VSS 0.0603958
R6072 VSS.n2335 VSS 0.0603958
R6073 VSS VSS.n1029 0.0603958
R6074 VSS.n3432 VSS.n3431 0.0590938
R6075 VSS VSS.n3449 0.0590938
R6076 VSS.n3104 VSS 0.0590938
R6077 VSS.n3163 VSS.n3162 0.0590938
R6078 VSS.n3379 VSS.n3378 0.0590938
R6079 VSS.n3355 VSS 0.0590938
R6080 VSS.n2922 VSS.n504 0.0574875
R6081 VSS.n2292 VSS.n1118 0.0574875
R6082 VSS.n2196 VSS.n1163 0.0574875
R6083 VSS.n2166 VSS.n2151 0.0574875
R6084 VSS.n2963 VSS.n509 0.0574875
R6085 VSS.n2927 VSS.n2926 0.0574875
R6086 VSS.n2564 VSS.n926 0.0574697
R6087 VSS.n2573 VSS.n923 0.0574697
R6088 VSS.n2955 VSS.n510 0.0574697
R6089 VSS.n2281 VSS.n1119 0.0574697
R6090 VSS.n1164 VSS.n1161 0.0574697
R6091 VSS.n531 VSS.n529 0.0574697
R6092 VSS.n2255 VSS.n2254 0.0574697
R6093 VSS.n2125 VSS.n1209 0.0574697
R6094 VSS.n1190 VSS.n1181 0.0574697
R6095 VSS.n643 VSS.n642 0.0574697
R6096 VSS.n2876 VSS.n589 0.0574697
R6097 VSS.n2093 VSS.n2047 0.0574697
R6098 VSS.n2908 VSS.n571 0.0574697
R6099 VSS.n743 VSS.n740 0.0574697
R6100 VSS.n2660 VSS.n756 0.0574697
R6101 VSS.n2856 VSS.n673 0.0574697
R6102 VSS.n2808 VSS.n687 0.0574697
R6103 VSS.n724 VSS.n721 0.0574697
R6104 VSS.n703 VSS.n701 0.0574697
R6105 VSS.n789 VSS.n788 0.0574697
R6106 VSS.n2645 VSS.n764 0.0574697
R6107 VSS.n1489 VSS.n1379 0.0574697
R6108 VSS.n1521 VSS.n1300 0.0574697
R6109 VSS.n1454 VSS.n1409 0.0574697
R6110 VSS.n1952 VSS.n1259 0.0574697
R6111 VSS.n993 VSS.n985 0.0574697
R6112 VSS.n1618 VSS.n829 0.0574697
R6113 VSS.n2606 VSS.n831 0.0574697
R6114 VSS.n1688 VSS.n1686 0.0574697
R6115 VSS.n1543 VSS.n1534 0.0574697
R6116 VSS.n898 VSS.n896 0.0574697
R6117 VSS.n1649 VSS.n1647 0.0574697
R6118 VSS.n2019 VSS.n1232 0.0574697
R6119 VSS.n1898 VSS.n1235 0.0574697
R6120 VSS.n1983 VSS.n1236 0.0574697
R6121 VSS.n2533 VSS.n953 0.0574697
R6122 VSS.n1279 VSS.n1276 0.0574697
R6123 VSS.n1799 VSS.n1771 0.0574697
R6124 VSS.n1750 VSS.n1738 0.0574697
R6125 VSS.n1828 VSS.n1739 0.0574697
R6126 VSS.n2454 VSS.n2429 0.0574697
R6127 VSS.n2487 VSS.n2404 0.0574697
R6128 VSS.n232 VSS.n231 0.0574529
R6129 VSS VSS.n3399 0.0557885
R6130 VSS VSS.n3398 0.0557885
R6131 VSS VSS.n3397 0.0557885
R6132 VSS.n126 VSS 0.0557885
R6133 VSS.n128 VSS 0.0557885
R6134 VSS.n133 VSS 0.0557885
R6135 VSS.n138 VSS 0.0557885
R6136 VSS.n143 VSS 0.0557885
R6137 VSS.n148 VSS 0.0557885
R6138 VSS.n153 VSS 0.0557885
R6139 VSS.n158 VSS 0.0557885
R6140 VSS.n163 VSS 0.0557885
R6141 VSS.n168 VSS 0.0557885
R6142 VSS.n3293 VSS 0.0557885
R6143 VSS.n2188 VSS.n1159 0.0551875
R6144 VSS.n1145 VSS.n1143 0.0551875
R6145 VSS.n534 VSS.n527 0.0551875
R6146 VSS.n564 VSS.n563 0.0551875
R6147 VSS.n1213 VSS.n1212 0.0551875
R6148 VSS.n2916 VSS.n574 0.0551875
R6149 VSS.n630 VSS.n605 0.0551875
R6150 VSS.n639 VSS.n638 0.0551875
R6151 VSS.n2695 VSS.n738 0.0551875
R6152 VSS.n2766 VSS.n708 0.0551875
R6153 VSS.n2865 VSS.n676 0.0551875
R6154 VSS.n2860 VSS.n2854 0.0551875
R6155 VSS.n1458 VSS.n1457 0.0551875
R6156 VSS.n794 VSS.n786 0.0551875
R6157 VSS.n822 VSS.n821 0.0551875
R6158 VSS.n1569 VSS.n1568 0.0551875
R6159 VSS.n1623 VSS.n1622 0.0551875
R6160 VSS.n902 VSS.n901 0.0551875
R6161 VSS.n893 VSS.n892 0.0551875
R6162 VSS.n1868 VSS.n1283 0.0551875
R6163 VSS.n1956 VSS.n1955 0.0551875
R6164 VSS.n2537 VSS.n2536 0.0551875
R6165 VSS.n979 VSS.n978 0.0551875
R6166 VSS.n2520 VSS.n988 0.0551875
R6167 VSS.n2451 VSS.n2450 0.0551875
R6168 VSS.n3010 VSS.n270 0.0551875
R6169 VSS.n1091 VSS.n1090 0.0551875
R6170 VSS.n2372 VSS.n1025 0.0551875
R6171 VSS.n2367 VSS.n2366 0.0551875
R6172 VSS.n3381 VSS 0.0527529
R6173 VSS VSS.n1250 0.0525833
R6174 VSS.n1802 VSS 0.0525833
R6175 VSS.n3381 VSS.n3380 0.0519696
R6176 VSS.n3295 VSS 0.0518289
R6177 VSS.n17 VSS.n14 0.0499792
R6178 VSS.n3132 VSS.n217 0.0499792
R6179 VSS.n3327 VSS.n111 0.0499792
R6180 VSS.n2160 VSS.n2159 0.0499792
R6181 VSS.n2230 VSS.n511 0.0499792
R6182 VSS.n2144 VSS.n1184 0.0499792
R6183 VSS.n586 VSS.n584 0.0499792
R6184 VSS.n2668 VSS.n2667 0.0499792
R6185 VSS.n1330 VSS.n1318 0.0499792
R6186 VSS.n1427 VSS.n765 0.0499792
R6187 VSS.n1722 VSS.n1537 0.0499792
R6188 VSS.n1653 VSS.n1652 0.0499792
R6189 VSS.n2589 VSS.n846 0.0499792
R6190 VSS.n1730 VSS.n1294 0.0499792
R6191 VSS.n1907 VSS.n1897 0.0499792
R6192 VSS.n1754 VSS.n1742 0.0499792
R6193 VSS.n2023 VSS.n2022 0.0499792
R6194 VSS.n2400 VSS.n2398 0.0499792
R6195 VSS.n252 VSS.n241 0.0499792
R6196 VSS.n1045 VSS.n1044 0.0499792
R6197 VSS.n3442 VSS.n3435 0.0486771
R6198 VSS.n3171 VSS.n3166 0.0486771
R6199 VSS.n104 VSS.n96 0.0486771
R6200 VSS.n2155 VSS 0.047375
R6201 VSS.n1192 VSS 0.047375
R6202 VSS.n2663 VSS 0.047375
R6203 VSS.n1319 VSS 0.047375
R6204 VSS.n1545 VSS 0.047375
R6205 VSS.n1733 VSS 0.047375
R6206 VSS.n1755 VSS 0.047375
R6207 VSS.n253 VSS 0.047375
R6208 VSS.n3466 VSS 0.0460729
R6209 VSS VSS.n3134 0.0460729
R6210 VSS VSS.n3298 0.0460729
R6211 VSS.n2183 VSS.n1165 0.0447708
R6212 VSS.n2133 VSS.n1203 0.0447708
R6213 VSS.n2690 VSS.n744 0.0447708
R6214 VSS.n1357 VSS.n1301 0.0447708
R6215 VSS.n1696 VSS.n1557 0.0447708
R6216 VSS.n1862 VSS.n1280 0.0447708
R6217 VSS.n1806 VSS.n1766 0.0447708
R6218 VSS.n3018 VSS.n3017 0.0447708
R6219 VSS.n3470 VSS.n3469 0.0423452
R6220 VSS.n3471 VSS.n3470 0.0423452
R6221 VSS.n3472 VSS.n3471 0.0423452
R6222 VSS.n3473 VSS.n3472 0.0423452
R6223 VSS.n3474 VSS.n3473 0.0423452
R6224 VSS.n3475 VSS.n3474 0.0423452
R6225 VSS.n3476 VSS.n3475 0.0423452
R6226 VSS.n3477 VSS.n3476 0.0423452
R6227 VSS.n3478 VSS.n3477 0.0423452
R6228 VSS.n3479 VSS.n3478 0.0423452
R6229 VSS.n3480 VSS.n3479 0.0423452
R6230 VSS.n3481 VSS.n3480 0.0423452
R6231 VSS.n3482 VSS.n3481 0.0423452
R6232 VSS.n3483 VSS.n3482 0.0423452
R6233 VSS.n3484 VSS.n3483 0.0423452
R6234 VSS.n3485 VSS.n3484 0.0423452
R6235 VSS.n3486 VSS.n3485 0.0423452
R6236 VSS.n3487 VSS.n3486 0.0423452
R6237 VSS.n3488 VSS.n3487 0.0423452
R6238 VSS.n3489 VSS.n3488 0.0423452
R6239 VSS.n3490 VSS.n3489 0.0423452
R6240 VSS.n3491 VSS.n3490 0.0423452
R6241 VSS.n871 VSS 0.0421667
R6242 VSS.n957 VSS 0.0421667
R6243 VSS.n2516 VSS 0.0421667
R6244 VSS.n2513 VSS 0.0421667
R6245 VSS.n3051 VSS.n230 0.0416941
R6246 VSS.n2385 VSS.n2383 0.0414836
R6247 VSS.n2311 VSS.n2310 0.0410405
R6248 VSS.n2318 VSS.n1037 0.0410405
R6249 VSS.n250 VSS.n249 0.0410405
R6250 VSS.n238 VSS.n236 0.0410405
R6251 VSS.n2569 VSS.n928 0.0410405
R6252 VSS.n2565 VSS.n2563 0.0410405
R6253 VSS.n1069 VSS.n1067 0.0410405
R6254 VSS.n1070 VSS.n1052 0.0410405
R6255 VSS.n2577 VSS.n2575 0.0410405
R6256 VSS.n2583 VSS.n851 0.0410405
R6257 VSS.n1087 VSS.n1086 0.0410405
R6258 VSS.n1088 VSS.n501 0.0410405
R6259 VSS.n2960 VSS.n512 0.0410405
R6260 VSS.n2956 VSS.n2954 0.0410405
R6261 VSS.n2289 VSS.n1121 0.0410405
R6262 VSS.n2283 VSS.n2282 0.0410405
R6263 VSS.n2193 VSS.n1166 0.0410405
R6264 VSS.n2189 VSS.n1160 0.0410405
R6265 VSS.n2162 VSS.n2154 0.0410405
R6266 VSS.n2157 VSS.n1176 0.0410405
R6267 VSS.n539 VSS.n528 0.0410405
R6268 VSS.n540 VSS.n532 0.0410405
R6269 VSS.n1135 VSS.n1134 0.0410405
R6270 VSS.n1137 VSS.n1136 0.0410405
R6271 VSS.n2127 VSS.n2126 0.0410405
R6272 VSS.n1211 VSS.n1210 0.0410405
R6273 VSS.n2146 VSS.n1183 0.0410405
R6274 VSS.n1193 VSS.n1191 0.0410405
R6275 VSS.n607 VSS.n606 0.0410405
R6276 VSS.n609 VSS.n608 0.0410405
R6277 VSS.n2878 VSS.n2877 0.0410405
R6278 VSS.n591 VSS.n590 0.0410405
R6279 VSS.n2095 VSS.n2094 0.0410405
R6280 VSS.n2049 VSS.n2048 0.0410405
R6281 VSS.n2918 VSS.n573 0.0410405
R6282 VSS.n2911 VSS.n2909 0.0410405
R6283 VSS.n2700 VSS.n745 0.0410405
R6284 VSS.n2696 VSS.n739 0.0410405
R6285 VSS.n2670 VSS.n2662 0.0410405
R6286 VSS.n2665 VSS.n755 0.0410405
R6287 VSS.n2866 VSS.n675 0.0410405
R6288 VSS.n2858 VSS.n2857 0.0410405
R6289 VSS.n2798 VSS.n688 0.0410405
R6290 VSS.n2807 VSS.n686 0.0410405
R6291 VSS.n2732 VSS.n729 0.0410405
R6292 VSS.n726 VSS.n720 0.0410405
R6293 VSS.n2768 VSS.n705 0.0410405
R6294 VSS.n706 VSS.n700 0.0410405
R6295 VSS.n1323 VSS.n1317 0.0410405
R6296 VSS.n1332 VSS.n1315 0.0410405
R6297 VSS.n796 VSS.n787 0.0410405
R6298 VSS.n797 VSS.n790 0.0410405
R6299 VSS.n2650 VSS.n766 0.0410405
R6300 VSS.n2646 VSS.n2644 0.0410405
R6301 VSS.n1382 VSS.n1377 0.0410405
R6302 VSS.n1490 VSS.n1378 0.0410405
R6303 VSS.n1526 VSS.n1302 0.0410405
R6304 VSS.n1522 VSS.n1520 0.0410405
R6305 VSS.n1406 VSS.n1404 0.0410405
R6306 VSS.n1455 VSS.n1405 0.0410405
R6307 VSS.n1256 VSS.n1254 0.0410405
R6308 VSS.n1953 VSS.n1255 0.0410405
R6309 VSS.n2522 VSS.n987 0.0410405
R6310 VSS.n2515 VSS.n994 0.0410405
R6311 VSS.n1619 VSS.n1617 0.0410405
R6312 VSS.n1620 VSS.n832 0.0410405
R6313 VSS.n1690 VSS.n1689 0.0410405
R6314 VSS.n1565 VSS.n1564 0.0410405
R6315 VSS.n1724 VSS.n1536 0.0410405
R6316 VSS.n1546 VSS.n1544 0.0410405
R6317 VSS.n900 VSS.n899 0.0410405
R6318 VSS.n869 VSS.n868 0.0410405
R6319 VSS.n1651 VSS.n1650 0.0410405
R6320 VSS.n1593 VSS.n1592 0.0410405
R6321 VSS.n2021 VSS.n2020 0.0410405
R6322 VSS.n1987 VSS.n1986 0.0410405
R6323 VSS.n1908 VSS.n1899 0.0410405
R6324 VSS.n1901 VSS.n1237 0.0410405
R6325 VSS.n1729 VSS.n1296 0.0410405
R6326 VSS.n1734 VSS.n1732 0.0410405
R6327 VSS.n2535 VSS.n2534 0.0410405
R6328 VSS.n955 VSS.n954 0.0410405
R6329 VSS.n1873 VSS.n1281 0.0410405
R6330 VSS.n1869 VSS.n1275 0.0410405
R6331 VSS.n1801 VSS.n1800 0.0410405
R6332 VSS.n1773 VSS.n1772 0.0410405
R6333 VSS.n1751 VSS.n1749 0.0410405
R6334 VSS.n1752 VSS.n1740 0.0410405
R6335 VSS.n2426 VSS.n2422 0.0410405
R6336 VSS.n2455 VSS.n2423 0.0410405
R6337 VSS.n2489 VSS.n2488 0.0410405
R6338 VSS.n2406 VSS.n2405 0.0410405
R6339 VSS.n2373 VSS.n1021 0.0410405
R6340 VSS.n2346 VSS.n1020 0.0410405
R6341 VSS.n3013 VSS.n266 0.0410405
R6342 VSS.n3002 VSS.n268 0.0410405
R6343 VSS.n2301 VSS.n2299 0.0393869
R6344 VSS.n594 VSS 0.0382604
R6345 VSS.n2169 VSS 0.0369583
R6346 VSS.n1195 VSS 0.0369583
R6347 VSS.n592 VSS 0.0369583
R6348 VSS.n2676 VSS 0.0369583
R6349 VSS.n2805 VSS 0.0369583
R6350 VSS.n1336 VSS 0.0369583
R6351 VSS.n1548 VSS 0.0369583
R6352 VSS.n922 VSS 0.0369583
R6353 VSS VSS.n1291 0.0369583
R6354 VSS VSS.n932 0.0369583
R6355 VSS.n1826 VSS 0.0369583
R6356 VSS.n3042 VSS 0.0369583
R6357 VSS.n2378 VSS.n2377 0.0352656
R6358 VSS.n827 VSS.n702 0.0351625
R6359 VSS.n1385 VSS.n723 0.0351625
R6360 VSS.n1529 VSS.n742 0.0351625
R6361 VSS.n2659 VSS.n760 0.0351625
R6362 VSS.n2654 VSS.n2653 0.0351625
R6363 VSS.n2613 VSS.n672 0.0351625
R6364 VSS.n210 VSS 0.0346243
R6365 VSS.n3465 VSS 0.0343542
R6366 VSS VSS.n216 0.0343542
R6367 VSS VSS.n3317 0.0343542
R6368 VSS.n2161 VSS.n2160 0.0343542
R6369 VSS.n2218 VSS.n1120 0.0343542
R6370 VSS.n2145 VSS.n2144 0.0343542
R6371 VSS.n2097 VSS.n2041 0.0343542
R6372 VSS.n2669 VSS.n2668 0.0343542
R6373 VSS.n2730 VSS.n725 0.0343542
R6374 VSS.n1322 VSS.n1318 0.0343542
R6375 VSS.n1338 VSS 0.0343542
R6376 VSS.n1381 VSS.n1371 0.0343542
R6377 VSS.n1723 VSS.n1722 0.0343542
R6378 VSS.n1718 VSS 0.0343542
R6379 VSS.n1653 VSS.n1588 0.0343542
R6380 VSS.n1295 VSS.n1294 0.0343542
R6381 VSS.n1841 VSS 0.0343542
R6382 VSS.n1910 VSS.n1897 0.0343542
R6383 VSS.n1973 VSS 0.0343542
R6384 VSS.n1929 VSS 0.0343542
R6385 VSS.n1748 VSS.n1742 0.0343542
R6386 VSS.n2023 VSS.n1226 0.0343542
R6387 VSS.n248 VSS.n241 0.0343542
R6388 VSS.n1065 VSS.n1064 0.0343542
R6389 VSS.n1041 VSS 0.0343542
R6390 VSS.n2526 VSS.n830 0.0339875
R6391 VSS.n1985 VSS.n1984 0.0339875
R6392 VSS.n1876 VSS.n1278 0.0339875
R6393 VSS.n1832 VSS.n1831 0.0339875
R6394 VSS.n2572 VSS.n925 0.0339875
R6395 VSS.n2531 VSS.n2530 0.0339875
R6396 VSS VSS.n3409 0.0330521
R6397 VSS VSS.n13 0.0330521
R6398 VSS.n3093 VSS 0.0330521
R6399 VSS.n3188 VSS 0.0330521
R6400 VSS VSS.n87 0.0330521
R6401 VSS VSS.n3326 0.0330521
R6402 VSS.n2222 VSS 0.0330521
R6403 VSS.n2235 VSS 0.0330521
R6404 VSS VSS.n2040 0.0330521
R6405 VSS VSS.n583 0.0330521
R6406 VSS.n2724 VSS 0.0330521
R6407 VSS.n2789 VSS 0.0330521
R6408 VSS.n1519 VSS 0.0330521
R6409 VSS.n1499 VSS 0.0330521
R6410 VSS.n1435 VSS 0.0330521
R6411 VSS.n1660 VSS 0.0330521
R6412 VSS VSS.n1895 0.0330521
R6413 VSS.n1932 VSS 0.0330521
R6414 VSS VSS.n1224 0.0330521
R6415 VSS VSS.n2396 0.0330521
R6416 VSS.n2425 VSS 0.0330521
R6417 VSS VSS.n279 0.0330521
R6418 VSS VSS.n494 0.0330521
R6419 VSS VSS.n37 0.03175
R6420 VSS.n3173 VSS 0.03175
R6421 VSS.n106 VSS 0.03175
R6422 VSS.n2221 VSS 0.03175
R6423 VSS.n563 VSS 0.03175
R6424 VSS VSS.n2727 0.03175
R6425 VSS.n2833 VSS 0.03175
R6426 VSS VSS.n674 0.03175
R6427 VSS VSS.n1337 0.03175
R6428 VSS.n1445 VSS 0.03175
R6429 VSS.n1434 VSS 0.03175
R6430 VSS.n1912 VSS 0.03175
R6431 VSS.n1252 VSS 0.03175
R6432 VSS.n949 VSS 0.03175
R6433 VSS.n1774 VSS 0.03175
R6434 VSS VSS.n1775 0.03175
R6435 VSS.n2005 VSS 0.03175
R6436 VSS.n2512 VSS 0.03175
R6437 VSS.n2466 VSS 0.03175
R6438 VSS.n2447 VSS 0.03175
R6439 VSS.n2381 VSS.n1018 0.0308279
R6440 VSS.n3399 VSS 0.0305481
R6441 VSS.n3398 VSS 0.0305481
R6442 VSS.n3397 VSS 0.0305481
R6443 VSS VSS.n126 0.0305481
R6444 VSS VSS.n3293 0.0305481
R6445 VSS.n2524 VSS.n985 0.0292489
R6446 VSS.n993 VSS.n984 0.0292489
R6447 VSS.n1259 VSS.n1258 0.0292489
R6448 VSS.n1952 VSS.n1951 0.0292489
R6449 VSS.n1409 VSS.n1408 0.0292489
R6450 VSS.n1454 VSS.n1453 0.0292489
R6451 VSS.n2770 VSS.n703 0.0292489
R6452 VSS.n2772 VSS.n701 0.0292489
R6453 VSS.n2920 VSS.n571 0.0292489
R6454 VSS.n2908 VSS.n569 0.0292489
R6455 VSS.n2256 VSS.n2255 0.0292489
R6456 VSS.n2254 VSS.n2253 0.0292489
R6457 VSS.n831 VSS.n828 0.0292489
R6458 VSS.n1618 VSS.n828 0.0292489
R6459 VSS.n2019 VSS.n2018 0.0292489
R6460 VSS.n2016 VSS.n1232 0.0292489
R6461 VSS.n1649 VSS.n1648 0.0292489
R6462 VSS.n1647 VSS.n1646 0.0292489
R6463 VSS.n1384 VSS.n1379 0.0292489
R6464 VSS.n1489 VSS.n1488 0.0292489
R6465 VSS.n2734 VSS.n724 0.0292489
R6466 VSS.n2736 VSS.n721 0.0292489
R6467 VSS.n2093 VSS.n2092 0.0292489
R6468 VSS.n2090 VSS.n2047 0.0292489
R6469 VSS.n2291 VSS.n1119 0.0292489
R6470 VSS.n2281 VSS.n1117 0.0292489
R6471 VSS.n1236 VSS.n1234 0.0292489
R6472 VSS.n1898 VSS.n1234 0.0292489
R6473 VSS.n1799 VSS.n1798 0.0292489
R6474 VSS.n1796 VSS.n1771 0.0292489
R6475 VSS.n1875 VSS.n1279 0.0292489
R6476 VSS.n1877 VSS.n1276 0.0292489
R6477 VSS.n1688 VSS.n1687 0.0292489
R6478 VSS.n1686 VSS.n1685 0.0292489
R6479 VSS.n1528 VSS.n1300 0.0292489
R6480 VSS.n1521 VSS.n1299 0.0292489
R6481 VSS.n2702 VSS.n743 0.0292489
R6482 VSS.n2704 VSS.n740 0.0292489
R6483 VSS.n2125 VSS.n2124 0.0292489
R6484 VSS.n2122 VSS.n1209 0.0292489
R6485 VSS.n2195 VSS.n1164 0.0292489
R6486 VSS.n2197 VSS.n1161 0.0292489
R6487 VSS.n1726 VSS.n1534 0.0292489
R6488 VSS.n1543 VSS.n1533 0.0292489
R6489 VSS.n2672 VSS.n2660 0.0292489
R6490 VSS.n2674 VSS.n756 0.0292489
R6491 VSS.n2148 VSS.n1181 0.0292489
R6492 VSS.n1190 VSS.n1180 0.0292489
R6493 VSS.n1739 VSS.n1737 0.0292489
R6494 VSS.n1750 VSS.n1737 0.0292489
R6495 VSS.n2487 VSS.n2486 0.0292489
R6496 VSS.n2484 VSS.n2404 0.0292489
R6497 VSS.n2571 VSS.n926 0.0292489
R6498 VSS.n2564 VSS.n924 0.0292489
R6499 VSS.n2579 VSS.n2573 0.0292489
R6500 VSS.n2581 VSS.n923 0.0292489
R6501 VSS.n2652 VSS.n764 0.0292489
R6502 VSS.n2645 VSS.n762 0.0292489
R6503 VSS.n2796 VSS.n687 0.0292489
R6504 VSS.n2809 VSS.n2808 0.0292489
R6505 VSS.n2876 VSS.n2875 0.0292489
R6506 VSS.n668 VSS.n589 0.0292489
R6507 VSS.n2962 VSS.n510 0.0292489
R6508 VSS.n2955 VSS.n508 0.0292489
R6509 VSS.n2429 VSS.n2428 0.0292489
R6510 VSS.n2454 VSS.n2453 0.0292489
R6511 VSS.n2533 VSS.n2532 0.0292489
R6512 VSS.n981 VSS.n953 0.0292489
R6513 VSS.n898 VSS.n897 0.0292489
R6514 VSS.n896 VSS.n895 0.0292489
R6515 VSS.n2614 VSS.n788 0.0292489
R6516 VSS.n824 VSS.n789 0.0292489
R6517 VSS.n2868 VSS.n673 0.0292489
R6518 VSS.n2856 VSS.n671 0.0292489
R6519 VSS.n644 VSS.n643 0.0292489
R6520 VSS.n642 VSS.n641 0.0292489
R6521 VSS.n2928 VSS.n529 0.0292489
R6522 VSS.n566 VSS.n531 0.0292489
R6523 VSS.n2191 VSS.n2188 0.0291458
R6524 VSS.n1143 VSS.n1141 0.0291458
R6525 VSS.n2930 VSS.n527 0.0291458
R6526 VSS.n1212 VSS.n1206 0.0291458
R6527 VSS.n2917 VSS.n2916 0.0291458
R6528 VSS.n646 VSS.n605 0.0291458
R6529 VSS.n2698 VSS.n2695 0.0291458
R6530 VSS.n2767 VSS.n2766 0.0291458
R6531 VSS.n676 VSS.n674 0.0291458
R6532 VSS.n1524 VSS.n1304 0.0291458
R6533 VSS.n1458 VSS.n1402 0.0291458
R6534 VSS.n2616 VSS.n786 0.0291458
R6535 VSS.n1569 VSS.n1561 0.0291458
R6536 VSS.n1623 VSS.n1614 0.0291458
R6537 VSS.n902 VSS.n864 0.0291458
R6538 VSS.n1871 VSS.n1868 0.0291458
R6539 VSS.n1956 VSS.n1252 0.0291458
R6540 VSS.n2537 VSS.n949 0.0291458
R6541 VSS.n1775 VSS.n1774 0.0291458
R6542 VSS.n2521 VSS.n2520 0.0291458
R6543 VSS.n2424 VSS.n2418 0.0291458
R6544 VSS.n3011 VSS.n3010 0.0291458
R6545 VSS.n1091 VSS.n1083 0.0291458
R6546 VSS.n1025 VSS.n1024 0.0291458
R6547 VSS.n2288 VSS 0.0278438
R6548 VSS VSS.n2096 0.0278438
R6549 VSS.n2731 VSS 0.0278438
R6550 VSS.n1375 VSS 0.0278438
R6551 VSS VSS.n927 0.0278438
R6552 VSS.n1066 VSS 0.0278438
R6553 VSS.n1381 VSS 0.0265417
R6554 VSS.n1825 VSS 0.0252396
R6555 VSS.n1807 VSS 0.0252396
R6556 VSS.n1787 VSS 0.0252396
R6557 VSS.n2010 VSS 0.0252396
R6558 VSS.n2502 VSS 0.0252396
R6559 VSS.n2471 VSS 0.0252396
R6560 VSS.n2446 VSS 0.0252396
R6561 VSS VSS.n2333 0.0252396
R6562 VSS.n2376 VSS.n2375 0.024993
R6563 VSS.n2285 VSS.n1126 0.0239375
R6564 VSS.n2958 VSS.n514 0.0239375
R6565 VSS.n2952 VSS.n516 0.0239375
R6566 VSS.n2052 VSS.n2051 0.0239375
R6567 VSS.n593 VSS.n592 0.0239375
R6568 VSS.n666 VSS.n595 0.0239375
R6569 VSS.n2738 VSS.n719 0.0239375
R6570 VSS.n2805 VSS.n2804 0.0239375
R6571 VSS.n2811 VSS.n685 0.0239375
R6572 VSS.n1337 VSS.n1336 0.0239375
R6573 VSS.n1386 VSS.n1376 0.0239375
R6574 VSS.n2648 VSS.n768 0.0239375
R6575 VSS.n2642 VSS.n770 0.0239375
R6576 VSS.n1719 VSS.n1548 0.0239375
R6577 VSS.n1596 VSS.n1595 0.0239375
R6578 VSS.n1640 VSS 0.0239375
R6579 VSS.n2585 VSS.n849 0.0239375
R6580 VSS.n922 VSS.n850 0.0239375
R6581 VSS.n881 VSS 0.0239375
R6582 VSS.n1840 VSS.n1291 0.0239375
R6583 VSS VSS.n1860 0.0239375
R6584 VSS.n1900 VSS.n1238 0.0239375
R6585 VSS.n2567 VSS.n930 0.0239375
R6586 VSS.n2561 VSS.n932 0.0239375
R6587 VSS.n1826 VSS.n1825 0.0239375
R6588 VSS.n1776 VSS 0.0239375
R6589 VSS.n1990 VSS.n1989 0.0239375
R6590 VSS.n2407 VSS.n2401 0.0239375
R6591 VSS.n2482 VSS.n2409 0.0239375
R6592 VSS.n3042 VSS.n3041 0.0239375
R6593 VSS.n1056 VSS.n1053 0.0239375
R6594 VSS.n2316 VSS.n1038 0.0239375
R6595 VSS.n2320 VSS.n1036 0.0239375
R6596 VSS.n2968 VSS.n2967 0.0234125
R6597 VSS.n2294 VSS.n2293 0.0234125
R6598 VSS.n1162 VSS.n267 0.0234125
R6599 VSS.n1179 VSS.n237 0.0234125
R6600 VSS.n2964 VSS.n507 0.0234125
R6601 VSS.n1023 VSS.n530 0.0234125
R6602 VSS.n3431 VSS 0.0226354
R6603 VSS.n3426 VSS 0.0226354
R6604 VSS VSS.n62 0.0226354
R6605 VSS.n3417 VSS 0.0226354
R6606 VSS.n3412 VSS 0.0226354
R6607 VSS.n3438 VSS 0.0226354
R6608 VSS.n5 VSS 0.0226354
R6609 VSS VSS.n12 0.0226354
R6610 VSS.n3457 VSS 0.0226354
R6611 VSS VSS.n19 0.0226354
R6612 VSS.n35 VSS 0.0226354
R6613 VSS.n27 VSS 0.0226354
R6614 VSS.n3086 VSS 0.0226354
R6615 VSS VSS.n3092 0.0226354
R6616 VSS.n3127 VSS 0.0226354
R6617 VSS.n3120 VSS 0.0226354
R6618 VSS.n3113 VSS 0.0226354
R6619 VSS.n3162 VSS 0.0226354
R6620 VSS VSS.n3147 0.0226354
R6621 VSS.n3149 VSS 0.0226354
R6622 VSS VSS.n190 0.0226354
R6623 VSS VSS.n193 0.0226354
R6624 VSS.n3378 VSS 0.0226354
R6625 VSS.n3373 VSS 0.0226354
R6626 VSS VSS.n85 0.0226354
R6627 VSS.n3364 VSS 0.0226354
R6628 VSS VSS.n91 0.0226354
R6629 VSS.n100 VSS 0.0226354
R6630 VSS.n3318 VSS 0.0226354
R6631 VSS VSS.n3325 0.0226354
R6632 VSS VSS.n3332 0.0226354
R6633 VSS VSS.n3337 0.0226354
R6634 VSS.n3354 VSS 0.0226354
R6635 VSS.n3344 VSS 0.0226354
R6636 VSS VSS.n2216 0.0226354
R6637 VSS.n2218 VSS 0.0226354
R6638 VSS.n2285 VSS 0.0226354
R6639 VSS VSS.n1131 0.0226354
R6640 VSS.n2238 VSS 0.0226354
R6641 VSS.n2234 VSS 0.0226354
R6642 VSS.n2940 VSS 0.0226354
R6643 VSS.n544 VSS 0.0226354
R6644 VSS.n552 VSS 0.0226354
R6645 VSS.n2107 VSS 0.0226354
R6646 VSS.n2097 VSS 0.0226354
R6647 VSS.n2080 VSS 0.0226354
R6648 VSS VSS.n2062 0.0226354
R6649 VSS.n2905 VSS 0.0226354
R6650 VSS VSS.n580 0.0226354
R6651 VSS VSS.n593 0.0226354
R6652 VSS.n638 VSS 0.0226354
R6653 VSS.n616 VSS 0.0226354
R6654 VSS VSS.n2723 0.0226354
R6655 VSS VSS.n2730 0.0226354
R6656 VSS.n2738 VSS 0.0226354
R6657 VSS.n2757 VSS 0.0226354
R6658 VSS VSS.n2788 0.0226354
R6659 VSS VSS.n2793 0.0226354
R6660 VSS.n2826 VSS 0.0226354
R6661 VSS VSS.n2832 0.0226354
R6662 VSS.n2847 VSS 0.0226354
R6663 VSS VSS.n1349 0.0226354
R6664 VSS.n1350 VSS 0.0226354
R6665 VSS VSS.n1304 0.0226354
R6666 VSS.n1513 VSS 0.0226354
R6667 VSS VSS.n1367 0.0226354
R6668 VSS.n1497 VSS 0.0226354
R6669 VSS VSS.n1371 0.0226354
R6670 VSS.n1486 VSS 0.0226354
R6671 VSS.n1436 VSS 0.0226354
R6672 VSS VSS.n1426 0.0226354
R6673 VSS VSS.n778 0.0226354
R6674 VSS.n810 VSS 0.0226354
R6675 VSS.n1698 VSS 0.0226354
R6676 VSS VSS.n1576 0.0226354
R6677 VSS VSS.n1579 0.0226354
R6678 VSS.n1643 VSS 0.0226354
R6679 VSS VSS.n1609 0.0226354
R6680 VSS.n1627 VSS 0.0226354
R6681 VSS.n2595 VSS 0.0226354
R6682 VSS.n906 VSS 0.0226354
R6683 VSS VSS.n873 0.0226354
R6684 VSS VSS.n1847 0.0226354
R6685 VSS VSS.n1848 0.0226354
R6686 VSS.n1881 VSS 0.0226354
R6687 VSS.n1886 VSS 0.0226354
R6688 VSS.n1911 VSS 0.0226354
R6689 VSS.n1966 VSS 0.0226354
R6690 VSS.n1965 VSS 0.0226354
R6691 VSS.n1943 VSS 0.0226354
R6692 VSS.n1933 VSS 0.0226354
R6693 VSS.n1928 VSS 0.0226354
R6694 VSS.n1923 VSS 0.0226354
R6695 VSS VSS.n941 0.0226354
R6696 VSS VSS.n945 0.0226354
R6697 VSS VSS.n965 0.0226354
R6698 VSS.n1808 VSS 0.0226354
R6699 VSS.n2013 VSS 0.0226354
R6700 VSS.n2505 VSS 0.0226354
R6701 VSS VSS.n2410 0.0226354
R6702 VSS VSS.n2418 0.0226354
R6703 VSS.n2436 VSS 0.0226354
R6704 VSS.n3034 VSS 0.0226354
R6705 VSS.n3019 VSS 0.0226354
R6706 VSS.n2990 VSS 0.0226354
R6707 VSS VSS.n1065 0.0226354
R6708 VSS.n2983 VSS 0.0226354
R6709 VSS.n2330 VSS 0.0226354
R6710 VSS.n2360 VSS 0.0226354
R6711 VSS.n2352 VSS 0.0226354
R6712 VSS.n3294 VSS 0.0219286
R6713 VSS.n2303 VSS.n2302 0.0218125
R6714 VSS.n2812 VSS 0.0213333
R6715 VSS.n2597 VSS 0.0213333
R6716 VSS VSS.n128 0.0209327
R6717 VSS.n130 VSS 0.0209327
R6718 VSS VSS.n133 0.0209327
R6719 VSS.n135 VSS 0.0209327
R6720 VSS VSS.n138 0.0209327
R6721 VSS.n140 VSS 0.0209327
R6722 VSS VSS.n143 0.0209327
R6723 VSS.n145 VSS 0.0209327
R6724 VSS VSS.n148 0.0209327
R6725 VSS.n150 VSS 0.0209327
R6726 VSS VSS.n153 0.0209327
R6727 VSS.n155 VSS 0.0209327
R6728 VSS VSS.n158 0.0209327
R6729 VSS.n160 VSS 0.0209327
R6730 VSS VSS.n163 0.0209327
R6731 VSS.n165 VSS 0.0209327
R6732 VSS VSS.n168 0.0209327
R6733 VSS.n170 VSS 0.0209327
R6734 VSS VSS.n2153 0.0200312
R6735 VSS VSS.n1182 0.0200312
R6736 VSS VSS.n2661 0.0200312
R6737 VSS.n1327 VSS 0.0200312
R6738 VSS VSS.n1535 0.0200312
R6739 VSS.n1836 VSS 0.0200312
R6740 VSS VSS.n1747 0.0200312
R6741 VSS VSS.n1761 0.0200312
R6742 VSS VSS.n247 0.0200312
R6743 VSS.n2200 VSS.n2199 0.0187292
R6744 VSS.n1146 VSS.n1138 0.0187292
R6745 VSS.n2251 VSS.n2250 0.0187292
R6746 VSS.n542 VSS.n538 0.0187292
R6747 VSS.n544 VSS.n543 0.0187292
R6748 VSS.n2120 VSS.n1214 0.0187292
R6749 VSS.n2913 VSS.n2912 0.0187292
R6750 VSS.n2906 VSS.n2905 0.0187292
R6751 VSS.n633 VSS.n631 0.0187292
R6752 VSS.n635 VSS.n634 0.0187292
R6753 VSS.n2707 VSS.n2706 0.0187292
R6754 VSS.n2762 VSS.n699 0.0187292
R6755 VSS.n2775 VSS.n2774 0.0187292
R6756 VSS.n2864 VSS.n677 0.0187292
R6757 VSS.n2861 VSS.n2838 0.0187292
R6758 VSS.n1518 VSS.n1306 0.0187292
R6759 VSS.n1410 VSS.n1403 0.0187292
R6760 VSS.n1451 VSS.n1450 0.0187292
R6761 VSS.n800 VSS.n799 0.0187292
R6762 VSS.n795 VSS.n791 0.0187292
R6763 VSS.n1683 VSS.n1566 0.0187292
R6764 VSS.n1615 VSS.n833 0.0187292
R6765 VSS.n2604 VSS.n2603 0.0187292
R6766 VSS.n870 VSS.n865 0.0187292
R6767 VSS.n872 VSS.n871 0.0187292
R6768 VSS.n1879 VSS.n1274 0.0187292
R6769 VSS.n1260 VSS.n1253 0.0187292
R6770 VSS.n1949 VSS.n1948 0.0187292
R6771 VSS.n956 VSS.n950 0.0187292
R6772 VSS.n958 VSS.n957 0.0187292
R6773 VSS.n1794 VSS.n1777 0.0187292
R6774 VSS.n2517 VSS.n2516 0.0187292
R6775 VSS.n2513 VSS.n2512 0.0187292
R6776 VSS.n2458 VSS.n2457 0.0187292
R6777 VSS.n2431 VSS.n2430 0.0187292
R6778 VSS.n3007 VSS.n3006 0.0187292
R6779 VSS.n1084 VSS.n500 0.0187292
R6780 VSS.n2972 VSS.n2971 0.0187292
R6781 VSS.n2371 VSS.n1027 0.0187292
R6782 VSS.n2368 VSS.n2347 0.0187292
R6783 VSS.n2297 VSS.n2296 0.0183038
R6784 VSS.n2298 VSS.n2295 0.0182893
R6785 VSS VSS.n986 0.0174271
R6786 VSS.n472 VSS.n471 0.0158654
R6787 VSS.n3466 VSS.n3465 0.0148229
R6788 VSS.n3134 VSS.n216 0.0148229
R6789 VSS.n3317 VSS.n3298 0.0148229
R6790 VSS.n2258 VSS 0.0148229
R6791 VSS VSS.n704 0.0148229
R6792 VSS.n3047 VSS 0.0140546
R6793 VSS.n2156 VSS.n2155 0.0135208
R6794 VSS.n2287 VSS.n1122 0.0135208
R6795 VSS.n2959 VSS.n513 0.0135208
R6796 VSS.n1192 VSS.n1186 0.0135208
R6797 VSS.n2050 VSS.n2044 0.0135208
R6798 VSS.n2880 VSS.n2879 0.0135208
R6799 VSS.n2664 VSS.n2663 0.0135208
R6800 VSS.n727 VSS.n716 0.0135208
R6801 VSS.n2800 VSS.n2799 0.0135208
R6802 VSS.n1329 VSS.n1319 0.0135208
R6803 VSS.n1493 VSS.n1492 0.0135208
R6804 VSS.n2649 VSS.n767 0.0135208
R6805 VSS.n1545 VSS.n1539 0.0135208
R6806 VSS.n1594 VSS.n1589 0.0135208
R6807 VSS.n2576 VSS.n847 0.0135208
R6808 VSS.n1733 VSS.n1293 0.0135208
R6809 VSS.n1906 VSS.n1903 0.0135208
R6810 VSS.n2568 VSS.n929 0.0135208
R6811 VSS.n1756 VSS.n1755 0.0135208
R6812 VSS.n1988 VSS.n1229 0.0135208
R6813 VSS.n2491 VSS.n2490 0.0135208
R6814 VSS.n254 VSS.n253 0.0135208
R6815 VSS.n1073 VSS.n1072 0.0135208
R6816 VSS.n2313 VSS.n2312 0.0135208
R6817 VSS VSS.n927 0.0109167
R6818 VSS.n1066 VSS 0.0109167
R6819 VSS.n2879 VSS 0.00961458
R6820 VSS.n2799 VSS 0.00961458
R6821 VSS.n2152 VSS.n1177 0.00878194
R6822 VSS.n1333 VSS.n1316 0.00878194
R6823 VSS.n1728 VSS.n1298 0.00878194
R6824 VSS.n242 VSS.n235 0.00838554
R6825 VSS.n3045 VSS.n3044 0.00838554
R6826 VSS.n2192 VSS.n1167 0.0083125
R6827 VSS.n2129 VSS.n2128 0.0083125
R6828 VSS.n2065 VSS.n572 0.0083125
R6829 VSS.n2699 VSS.n746 0.0083125
R6830 VSS.n1525 VSS.n1303 0.0083125
R6831 VSS.n1462 VSS.n1399 0.0083125
R6832 VSS.n1692 VSS.n1691 0.0083125
R6833 VSS.n1626 VSS.n1613 0.0083125
R6834 VSS.n1872 VSS.n1282 0.0083125
R6835 VSS.n1959 VSS.n1250 0.0083125
R6836 VSS.n1803 VSS.n1802 0.0083125
R6837 VSS.n1997 VSS.n986 0.0083125
R6838 VSS.n269 VSS.n265 0.0083125
R6839 VSS.n1094 VSS.n1081 0.0083125
R6840 VSS.n2386 VSS.n2381 0.00808197
R6841 VSS.n3046 VSS.n235 0.00790157
R6842 VSS.n3046 VSS.n3045 0.00790157
R6843 VSS.n2525 VSS 0.00755
R6844 VSS.n2017 VSS 0.00755
R6845 VSS.n1797 VSS 0.00755
R6846 VSS.n1829 VSS 0.00755
R6847 VSS.n2485 VSS 0.00755
R6848 VSS.n982 VSS 0.00755
R6849 VSS.n3047 VSS.n3046 0.0070355
R6850 VSS.n2457 VSS 0.00701042
R6851 VSS.n1051 VSS.n1049 0.00653911
R6852 VSS.n3003 VSS.n234 0.00640857
R6853 VSS.n3015 VSS.n3014 0.00636298
R6854 VSS.n3004 VSS.n3003 0.00636298
R6855 VSS.n2304 VSS.n502 0.00631183
R6856 VSS.n1068 VSS.n1050 0.00624332
R6857 VSS.n1116 VSS.n1051 0.00624332
R6858 VSS.n1048 VSS.n503 0.00604629
R6859 VSS.n2969 VSS.n502 0.00604629
R6860 VSS.n2309 VSS.n2308 0.00579577
R6861 VSS.n564 VSS 0.00570833
R6862 VSS.n639 VSS 0.00570833
R6863 VSS VSS.n1776 0.00570833
R6864 VSS.n2425 VSS 0.00570833
R6865 VSS.n3014 VSS.n234 0.00533429
R6866 VSS.n2295 VSS.n2294 0.0052
R6867 VSS.n2296 VSS.n267 0.0052
R6868 VSS.n2299 VSS.n507 0.0052
R6869 VSS.n2300 VSS.n1023 0.0052
R6870 VSS.n2165 VSS.n2164 0.00513595
R6871 VSS.n1325 VSS.n1324 0.00513595
R6872 VSS.n1834 VSS.n1833 0.00513595
R6873 VSS.n1833 VSS.n1298 0.00513595
R6874 VSS.n1736 VSS.n1728 0.00513595
R6875 VSS.n1324 VSS.n1316 0.00513595
R6876 VSS.n1334 VSS.n1333 0.00513595
R6877 VSS.n2165 VSS.n2152 0.00513595
R6878 VSS.n2167 VSS.n1177 0.00513595
R6879 VSS.n1068 VSS.n1049 0.00496369
R6880 VSS.n2304 VSS.n1048 0.0047957
R6881 VSS.n52 VSS.n51 0.00440625
R6882 VSS.n3142 VSS.n3141 0.00440625
R6883 VSS.n3307 VSS.n3300 0.00440625
R6884 VSS.n2199 VSS 0.00440625
R6885 VSS.n2120 VSS 0.00440625
R6886 VSS.n2706 VSS 0.00440625
R6887 VSS VSS.n956 0.00440625
R6888 VSS.n2309 VSS.n2306 0.00364583
R6889 VSS.n2307 VSS.n1019 0.00364583
R6890 VSS.n2308 VSS.n2307 0.00364583
R6891 VSS.n2306 VSS.n2305 0.00364583
R6892 VSS VSS.n870 0.00310417
R6893 VSS.n37 VSS.n36 0.00180208
R6894 VSS.n3449 VSS.n35 0.00180208
R6895 VSS.n3113 VSS.n3104 0.00180208
R6896 VSS.n3173 VSS.n194 0.00180208
R6897 VSS.n3358 VSS.n106 0.00180208
R6898 VSS.n3355 VSS.n3354 0.00180208
R6899 VSS.n2386 VSS.n2385 0.00152459
R6900 VSS.n2608 VSS.n2607 0.0010875
R6901 VSS.n1380 VSS.n1233 0.0010875
R6902 VSS.n1530 VSS.n1277 0.0010875
R6903 VSS.n1727 VSS.n1532 0.0010875
R6904 VSS.n2580 VSS.n763 0.0010875
R6905 VSS.n2612 VSS.n825 0.0010875
R6906 VDPWR.n711 VDPWR.n707 8629.41
R6907 VDPWR.n711 VDPWR.n708 8629.41
R6908 VDPWR.n713 VDPWR.n707 8629.41
R6909 VDPWR.n713 VDPWR.n708 8629.41
R6910 VDPWR.n696 VDPWR.n692 8629.41
R6911 VDPWR.n696 VDPWR.n693 8629.41
R6912 VDPWR.n698 VDPWR.n692 8629.41
R6913 VDPWR.n698 VDPWR.n693 8629.41
R6914 VDPWR.n680 VDPWR.n676 8629.41
R6915 VDPWR.n680 VDPWR.n677 8629.41
R6916 VDPWR.n682 VDPWR.n676 8629.41
R6917 VDPWR.n682 VDPWR.n677 8629.41
R6918 VDPWR.n666 VDPWR.n660 8629.41
R6919 VDPWR.n664 VDPWR.n660 8629.41
R6920 VDPWR.n666 VDPWR.n662 8629.41
R6921 VDPWR.n664 VDPWR.n662 8629.41
R6922 VDPWR.n522 VDPWR.n518 8629.41
R6923 VDPWR.n522 VDPWR.n519 8629.41
R6924 VDPWR.n524 VDPWR.n518 8629.41
R6925 VDPWR.n524 VDPWR.n519 8629.41
R6926 VDPWR.n507 VDPWR.n503 8629.41
R6927 VDPWR.n507 VDPWR.n504 8629.41
R6928 VDPWR.n509 VDPWR.n503 8629.41
R6929 VDPWR.n509 VDPWR.n504 8629.41
R6930 VDPWR.n491 VDPWR.n487 8629.41
R6931 VDPWR.n491 VDPWR.n488 8629.41
R6932 VDPWR.n493 VDPWR.n487 8629.41
R6933 VDPWR.n493 VDPWR.n488 8629.41
R6934 VDPWR.n474 VDPWR.n470 8629.41
R6935 VDPWR.n474 VDPWR.n471 8629.41
R6936 VDPWR.n476 VDPWR.n470 8629.41
R6937 VDPWR.n476 VDPWR.n471 8629.41
R6938 VDPWR.n412 VDPWR.n406 8629.41
R6939 VDPWR.n412 VDPWR.n407 8629.41
R6940 VDPWR.n410 VDPWR.n407 8629.41
R6941 VDPWR.n410 VDPWR.n406 8629.41
R6942 VDPWR.n385 VDPWR.n379 8629.41
R6943 VDPWR.n382 VDPWR.n381 8629.41
R6944 VDPWR.n397 VDPWR.n391 8629.41
R6945 VDPWR.n394 VDPWR.n393 8629.41
R6946 VDPWR.n453 VDPWR.n449 8629.41
R6947 VDPWR.n453 VDPWR.n450 8629.41
R6948 VDPWR.n455 VDPWR.n449 8629.41
R6949 VDPWR.n455 VDPWR.n450 8629.41
R6950 VDPWR.n437 VDPWR.n433 8629.41
R6951 VDPWR.n437 VDPWR.n434 8629.41
R6952 VDPWR.n439 VDPWR.n433 8629.41
R6953 VDPWR.n439 VDPWR.n434 8629.41
R6954 VDPWR.n423 VDPWR.n417 8629.41
R6955 VDPWR.n421 VDPWR.n417 8629.41
R6956 VDPWR.n423 VDPWR.n419 8629.41
R6957 VDPWR.n421 VDPWR.n419 8629.41
R6958 VDPWR.n766 VDPWR.n762 8629.41
R6959 VDPWR.n766 VDPWR.n763 8629.41
R6960 VDPWR.n768 VDPWR.n762 8629.41
R6961 VDPWR.n768 VDPWR.n763 8629.41
R6962 VDPWR.n3160 VDPWR.n3154 8629.41
R6963 VDPWR.n3160 VDPWR.n3155 8629.41
R6964 VDPWR.n3158 VDPWR.n3155 8629.41
R6965 VDPWR.n3158 VDPWR.n3154 8629.41
R6966 VDPWR.n3144 VDPWR.n3138 8629.41
R6967 VDPWR.n3144 VDPWR.n3139 8629.41
R6968 VDPWR.n3142 VDPWR.n3139 8629.41
R6969 VDPWR.n3142 VDPWR.n3138 8629.41
R6970 VDPWR.n3125 VDPWR.n3121 8629.41
R6971 VDPWR.n3125 VDPWR.n3122 8629.41
R6972 VDPWR.n3127 VDPWR.n3121 8629.41
R6973 VDPWR.n3127 VDPWR.n3122 8629.41
R6974 VDPWR.n734 VDPWR.n731 5460
R6975 VDPWR.n736 VDPWR.n731 5460
R6976 VDPWR.n734 VDPWR.n732 5460
R6977 VDPWR.n736 VDPWR.n732 5460
R6978 VDPWR.n748 VDPWR.n742 4260
R6979 VDPWR.n746 VDPWR.n745 4260
R6980 VDPWR.t315 VDPWR.n711 2459.29
R6981 VDPWR.n713 VDPWR.t314 2459.29
R6982 VDPWR.t760 VDPWR.n696 2459.29
R6983 VDPWR.n698 VDPWR.t761 2459.29
R6984 VDPWR.t281 VDPWR.n680 2459.29
R6985 VDPWR.n682 VDPWR.t282 2459.29
R6986 VDPWR.t763 VDPWR.n660 2459.29
R6987 VDPWR.t762 VDPWR.n662 2459.29
R6988 VDPWR.t1036 VDPWR.n522 2459.29
R6989 VDPWR.n524 VDPWR.t1035 2459.29
R6990 VDPWR.t67 VDPWR.n507 2459.29
R6991 VDPWR.n509 VDPWR.t13 2459.29
R6992 VDPWR.t122 VDPWR.n491 2459.29
R6993 VDPWR.n493 VDPWR.t121 2459.29
R6994 VDPWR.t956 VDPWR.n474 2459.29
R6995 VDPWR.n476 VDPWR.t957 2459.29
R6996 VDPWR.t345 VDPWR.n410 2459.29
R6997 VDPWR.n412 VDPWR.t1037 2459.29
R6998 VDPWR.t68 VDPWR.n453 2459.29
R6999 VDPWR.n455 VDPWR.t69 2459.29
R7000 VDPWR.t120 VDPWR.n437 2459.29
R7001 VDPWR.n439 VDPWR.t123 2459.29
R7002 VDPWR.t958 VDPWR.n417 2459.29
R7003 VDPWR.t959 VDPWR.n419 2459.29
R7004 VDPWR.t1012 VDPWR.n766 2459.29
R7005 VDPWR.n768 VDPWR.t118 2459.29
R7006 VDPWR.t239 VDPWR.n3158 2459.29
R7007 VDPWR.n3160 VDPWR.t1093 2459.29
R7008 VDPWR.t49 VDPWR.n3142 2459.29
R7009 VDPWR.n3144 VDPWR.t50 2459.29
R7010 VDPWR.t1094 VDPWR.n3125 2459.29
R7011 VDPWR.n3127 VDPWR.t1095 2459.29
R7012 VDPWR.n712 VDPWR.t315 2298.92
R7013 VDPWR.t314 VDPWR.n712 2298.92
R7014 VDPWR.n697 VDPWR.t760 2298.92
R7015 VDPWR.t761 VDPWR.n697 2298.92
R7016 VDPWR.n681 VDPWR.t281 2298.92
R7017 VDPWR.t282 VDPWR.n681 2298.92
R7018 VDPWR.n665 VDPWR.t763 2298.92
R7019 VDPWR.n665 VDPWR.t762 2298.92
R7020 VDPWR.n523 VDPWR.t1036 2298.92
R7021 VDPWR.t1035 VDPWR.n523 2298.92
R7022 VDPWR.n508 VDPWR.t67 2298.92
R7023 VDPWR.t13 VDPWR.n508 2298.92
R7024 VDPWR.n492 VDPWR.t122 2298.92
R7025 VDPWR.t121 VDPWR.n492 2298.92
R7026 VDPWR.n475 VDPWR.t956 2298.92
R7027 VDPWR.t957 VDPWR.n475 2298.92
R7028 VDPWR.n411 VDPWR.t345 2298.92
R7029 VDPWR.t1037 VDPWR.n411 2298.92
R7030 VDPWR.n454 VDPWR.t68 2298.92
R7031 VDPWR.t69 VDPWR.n454 2298.92
R7032 VDPWR.n438 VDPWR.t120 2298.92
R7033 VDPWR.t123 VDPWR.n438 2298.92
R7034 VDPWR.n422 VDPWR.t958 2298.92
R7035 VDPWR.n422 VDPWR.t959 2298.92
R7036 VDPWR.n767 VDPWR.t1012 2298.92
R7037 VDPWR.t118 VDPWR.n767 2298.92
R7038 VDPWR.n3159 VDPWR.t239 2298.92
R7039 VDPWR.t1093 VDPWR.n3159 2298.92
R7040 VDPWR.n3143 VDPWR.t49 2298.92
R7041 VDPWR.t50 VDPWR.n3143 2298.92
R7042 VDPWR.n3126 VDPWR.t1094 2298.92
R7043 VDPWR.t1095 VDPWR.n3126 2298.92
R7044 VDPWR.n1367 VDPWR.n1349 2296.22
R7045 VDPWR.n1700 VDPWR.n1682 2296.22
R7046 VDPWR.n1623 VDPWR.n1622 2296.22
R7047 VDPWR.n2453 VDPWR.n2452 2291.62
R7048 VDPWR.n2452 VDPWR.n2442 1418.92
R7049 VDPWR.n1367 VDPWR.n1366 1408
R7050 VDPWR.n1700 VDPWR.n1699 1408
R7051 VDPWR.n1622 VDPWR.n1621 1408
R7052 VDPWR VDPWR.t565 975.178
R7053 VDPWR VDPWR.t465 975.178
R7054 VDPWR VDPWR.t459 975.178
R7055 VDPWR.n710 VDPWR.n709 920.471
R7056 VDPWR.n695 VDPWR.n694 920.471
R7057 VDPWR.n679 VDPWR.n678 920.471
R7058 VDPWR.n663 VDPWR.n659 920.471
R7059 VDPWR.n521 VDPWR.n520 920.471
R7060 VDPWR.n506 VDPWR.n505 920.471
R7061 VDPWR.n490 VDPWR.n489 920.471
R7062 VDPWR.n473 VDPWR.n472 920.471
R7063 VDPWR.n409 VDPWR.n408 920.471
R7064 VDPWR.n386 VDPWR.n380 920.471
R7065 VDPWR.n398 VDPWR.n392 920.471
R7066 VDPWR.n452 VDPWR.n451 920.471
R7067 VDPWR.n436 VDPWR.n435 920.471
R7068 VDPWR.n420 VDPWR.n416 920.471
R7069 VDPWR.n765 VDPWR.n764 920.471
R7070 VDPWR.n3157 VDPWR.n3156 920.471
R7071 VDPWR.n3141 VDPWR.n3140 920.471
R7072 VDPWR.n3124 VDPWR.n3123 920.471
R7073 VDPWR.n387 VDPWR.n386 917.46
R7074 VDPWR.n399 VDPWR.n398 917.46
R7075 VDPWR.n709 VDPWR.n705 914.447
R7076 VDPWR.n694 VDPWR.n689 914.447
R7077 VDPWR.n678 VDPWR.n673 914.447
R7078 VDPWR.n663 VDPWR.n658 914.447
R7079 VDPWR.n520 VDPWR.n516 914.447
R7080 VDPWR.n505 VDPWR.n500 914.447
R7081 VDPWR.n489 VDPWR.n484 914.447
R7082 VDPWR.n472 VDPWR.n468 914.447
R7083 VDPWR.n408 VDPWR.n404 914.447
R7084 VDPWR.n451 VDPWR.n446 914.447
R7085 VDPWR.n435 VDPWR.n430 914.447
R7086 VDPWR.n420 VDPWR.n415 914.447
R7087 VDPWR.n764 VDPWR.n760 914.447
R7088 VDPWR.n3156 VDPWR.n3151 914.447
R7089 VDPWR.n3140 VDPWR.n3135 914.447
R7090 VDPWR.n3123 VDPWR.n3119 914.447
R7091 VDPWR.t565 VDPWR 877.827
R7092 VDPWR.t465 VDPWR 877.827
R7093 VDPWR.t459 VDPWR 877.827
R7094 VDPWR.n2359 VDPWR.t389 843.261
R7095 VDPWR.n1871 VDPWR.t43 842.073
R7096 VDPWR.n3051 VDPWR.t1151 842.073
R7097 VDPWR.n1184 VDPWR.t349 832.876
R7098 VDPWR.n1826 VDPWR.t576 812.014
R7099 VDPWR.n2107 VDPWR.t493 811.918
R7100 VDPWR.n2172 VDPWR.t706 811.793
R7101 VDPWR.n2865 VDPWR.t309 808.141
R7102 VDPWR.n1239 VDPWR.t612 807.567
R7103 VDPWR.n2459 VDPWR.t512 807.548
R7104 VDPWR.n1796 VDPWR.t651 807.481
R7105 VDPWR.n1767 VDPWR.t753 807.481
R7106 VDPWR.n1761 VDPWR.t552 807.462
R7107 VDPWR.n1834 VDPWR.t454 806.484
R7108 VDPWR.n1327 VDPWR.t675 806.423
R7109 VDPWR.n1127 VDPWR.t547 806.423
R7110 VDPWR.n807 VDPWR.t266 804.845
R7111 VDPWR.n1528 VDPWR.t609 804.731
R7112 VDPWR.n1521 VDPWR.t608 804.731
R7113 VDPWR.n1528 VDPWR.t461 804.731
R7114 VDPWR.n1521 VDPWR.t460 804.731
R7115 VDPWR.n1520 VDPWR.t655 804.731
R7116 VDPWR.n1296 VDPWR.t654 804.731
R7117 VDPWR.n1482 VDPWR.t623 804.731
R7118 VDPWR.n1311 VDPWR.t622 804.731
R7119 VDPWR.n1482 VDPWR.t467 804.731
R7120 VDPWR.n1311 VDPWR.t466 804.731
R7121 VDPWR.n1312 VDPWR.t710 804.731
R7122 VDPWR.n1323 VDPWR.t709 804.731
R7123 VDPWR.n1312 VDPWR.t567 804.731
R7124 VDPWR.n1323 VDPWR.t566 804.731
R7125 VDPWR.n1326 VDPWR.t488 804.731
R7126 VDPWR.n1328 VDPWR.t621 804.731
R7127 VDPWR.n1405 VDPWR.t674 804.731
R7128 VDPWR.n1397 VDPWR.t620 804.731
R7129 VDPWR.n1339 VDPWR.t524 804.731
R7130 VDPWR.n1350 VDPWR.t523 804.731
R7131 VDPWR.n1353 VDPWR.t458 804.731
R7132 VDPWR.n1356 VDPWR.t647 804.731
R7133 VDPWR.n1360 VDPWR.t431 804.731
R7134 VDPWR.n1365 VDPWR.t634 804.731
R7135 VDPWR.n1540 VDPWR.t452 804.731
R7136 VDPWR.n1543 VDPWR.t649 804.731
R7137 VDPWR.n1213 VDPWR.t455 804.731
R7138 VDPWR.n1829 VDPWR.t745 804.731
R7139 VDPWR.n1798 VDPWR.t575 804.731
R7140 VDPWR.n1810 VDPWR.t652 804.731
R7141 VDPWR.n1769 VDPWR.t611 804.731
R7142 VDPWR.n1791 VDPWR.t754 804.731
R7143 VDPWR.n1260 VDPWR.t725 804.731
R7144 VDPWR.n1743 VDPWR.t470 804.731
R7145 VDPWR.n1735 VDPWR.t551 804.731
R7146 VDPWR.n1727 VDPWR.t469 804.731
R7147 VDPWR.n1275 VDPWR.t582 804.731
R7148 VDPWR.n1683 VDPWR.t581 804.731
R7149 VDPWR.n1686 VDPWR.t691 804.731
R7150 VDPWR.n1689 VDPWR.t538 804.731
R7151 VDPWR.n1693 VDPWR.t521 804.731
R7152 VDPWR.n1698 VDPWR.t703 804.731
R7153 VDPWR.n1201 VDPWR.t748 804.731
R7154 VDPWR.n1204 VDPWR.t615 804.731
R7155 VDPWR.n1208 VDPWR.t743 804.731
R7156 VDPWR.n1895 VDPWR.t604 804.731
R7157 VDPWR.n1602 VDPWR.t578 804.731
R7158 VDPWR.n1628 VDPWR.t560 804.731
R7159 VDPWR.n1644 VDPWR.t579 804.731
R7160 VDPWR.n2059 VDPWR.t561 804.731
R7161 VDPWR.n1639 VDPWR.t546 804.731
R7162 VDPWR.t448 VDPWR.n2048 804.731
R7163 VDPWR.n2047 VDPWR.t750 804.731
R7164 VDPWR.n1134 VDPWR.t665 804.731
R7165 VDPWR.n2027 VDPWR.t751 804.731
R7166 VDPWR.n1155 VDPWR.t666 804.731
R7167 VDPWR.n1153 VDPWR.t644 804.731
R7168 VDPWR.n1156 VDPWR.t659 804.731
R7169 VDPWR.n1177 VDPWR.t645 804.731
R7170 VDPWR.n1995 VDPWR.t660 804.731
R7171 VDPWR.n1606 VDPWR.t618 804.731
R7172 VDPWR.n1612 VDPWR.t695 804.731
R7173 VDPWR.n1615 VDPWR.t443 804.731
R7174 VDPWR.n1619 VDPWR.t535 804.731
R7175 VDPWR.t606 VDPWR.n1924 804.731
R7176 VDPWR.n1939 VDPWR.t515 804.731
R7177 VDPWR.n1942 VDPWR.t593 804.731
R7178 VDPWR.n2098 VDPWR.t527 804.731
R7179 VDPWR.n2101 VDPWR.t636 804.731
R7180 VDPWR.n2265 VDPWR.t591 804.731
R7181 VDPWR.n2284 VDPWR.t590 804.731
R7182 VDPWR.n1051 VDPWR.t632 804.731
R7183 VDPWR.n1029 VDPWR.t631 804.731
R7184 VDPWR.n2316 VDPWR.t738 804.731
R7185 VDPWR.n2207 VDPWR.t737 804.731
R7186 VDPWR.n2203 VDPWR.t434 804.731
R7187 VDPWR.n2185 VDPWR.t433 804.731
R7188 VDPWR.n1108 VDPWR.t563 804.731
R7189 VDPWR.n2166 VDPWR.t642 804.731
R7190 VDPWR.n2141 VDPWR.t705 804.731
R7191 VDPWR.n2136 VDPWR.t641 804.731
R7192 VDPWR.n2080 VDPWR.t494 804.731
R7193 VDPWR.n2094 VDPWR.t679 804.731
R7194 VDPWR.n1071 VDPWR.t585 804.731
R7195 VDPWR.n1074 VDPWR.t693 804.731
R7196 VDPWR.n2731 VDPWR.t626 804.731
R7197 VDPWR.n2734 VDPWR.t723 804.731
R7198 VDPWR.n2959 VDPWR.t689 804.731
R7199 VDPWR.n2940 VDPWR.t688 804.731
R7200 VDPWR.n939 VDPWR.t716 804.731
R7201 VDPWR.n2903 VDPWR.t715 804.731
R7202 VDPWR.t588 VDPWR.n2726 804.731
R7203 VDPWR.n2728 VDPWR.t572 804.731
R7204 VDPWR.n2743 VDPWR.t587 804.731
R7205 VDPWR.n932 VDPWR.t677 804.731
R7206 VDPWR.n2972 VDPWR.t446 804.731
R7207 VDPWR.n2552 VDPWR.t708 804.731
R7208 VDPWR.n2555 VDPWR.t491 804.731
R7209 VDPWR.n2559 VDPWR.t721 804.731
R7210 VDPWR.n2564 VDPWR.t500 804.731
R7211 VDPWR.n2597 VDPWR.t497 804.731
R7212 VDPWR.n891 VDPWR.t732 804.731
R7213 VDPWR.n2991 VDPWR.t428 804.731
R7214 VDPWR.n2999 VDPWR.t549 804.731
R7215 VDPWR.n819 VDPWR.t509 804.731
R7216 VDPWR.n2373 VDPWR.t476 804.731
R7217 VDPWR.n2376 VDPWR.t595 804.731
R7218 VDPWR.n2474 VDPWR.t734 804.731
R7219 VDPWR.n2450 VDPWR.t511 804.731
R7220 VDPWR.n834 VDPWR.t533 804.731
R7221 VDPWR.n838 VDPWR.t657 804.731
R7222 VDPWR.n1003 VDPWR.t1119 783.403
R7223 VDPWR.n2210 VDPWR.t419 779.372
R7224 VDPWR.n1065 VDPWR.t1082 779.372
R7225 VDPWR.t664 VDPWR.t749 772.086
R7226 VDPWR.t658 VDPWR.t643 772.086
R7227 VDPWR.t745 VDPWR.n1828 751.692
R7228 VDPWR.t725 VDPWR.n1259 751.692
R7229 VDPWR.t748 VDPWR.n1200 751.692
R7230 VDPWR.t615 VDPWR.n1203 751.692
R7231 VDPWR.n2049 VDPWR.t448 751.692
R7232 VDPWR.n1925 VDPWR.t606 751.692
R7233 VDPWR.t563 VDPWR.n1107 751.692
R7234 VDPWR.n2740 VDPWR.t588 751.692
R7235 VDPWR.t572 VDPWR.n2727 751.692
R7236 VDPWR.t587 VDPWR.n2742 751.692
R7237 VDPWR.t721 VDPWR.n2558 751.692
R7238 VDPWR.t500 VDPWR.n2563 751.692
R7239 VDPWR.t734 VDPWR.n2473 751.692
R7240 VDPWR.t488 VDPWR.n1325 725.173
R7241 VDPWR.t458 VDPWR.n1352 725.173
R7242 VDPWR.t647 VDPWR.n1355 725.173
R7243 VDPWR.t431 VDPWR.n1359 725.173
R7244 VDPWR.t634 VDPWR.n1364 725.173
R7245 VDPWR.t452 VDPWR.n1539 725.173
R7246 VDPWR.t649 VDPWR.n1542 725.173
R7247 VDPWR.t691 VDPWR.n1685 725.173
R7248 VDPWR.t538 VDPWR.n1688 725.173
R7249 VDPWR.t521 VDPWR.n1692 725.173
R7250 VDPWR.t703 VDPWR.n1697 725.173
R7251 VDPWR.t743 VDPWR.n1207 725.173
R7252 VDPWR.t604 VDPWR.n1894 725.173
R7253 VDPWR.t618 VDPWR.n1605 725.173
R7254 VDPWR.t695 VDPWR.n1611 725.173
R7255 VDPWR.t443 VDPWR.n1614 725.173
R7256 VDPWR.t535 VDPWR.n1618 725.173
R7257 VDPWR.t515 VDPWR.n1938 725.173
R7258 VDPWR.t593 VDPWR.n1941 725.173
R7259 VDPWR.t527 VDPWR.n2097 725.173
R7260 VDPWR.t636 VDPWR.n2100 725.173
R7261 VDPWR.t679 VDPWR.n2093 725.173
R7262 VDPWR.t585 VDPWR.n1070 725.173
R7263 VDPWR.t693 VDPWR.n1073 725.173
R7264 VDPWR.t626 VDPWR.n2730 725.173
R7265 VDPWR.t723 VDPWR.n2733 725.173
R7266 VDPWR.t677 VDPWR.n931 725.173
R7267 VDPWR.t446 VDPWR.n2971 725.173
R7268 VDPWR.t708 VDPWR.n2551 725.173
R7269 VDPWR.t491 VDPWR.n2554 725.173
R7270 VDPWR.t497 VDPWR.n2596 725.173
R7271 VDPWR.t732 VDPWR.n890 725.173
R7272 VDPWR.t428 VDPWR.n2990 725.173
R7273 VDPWR.t549 VDPWR.n2998 725.173
R7274 VDPWR.t509 VDPWR.n818 725.173
R7275 VDPWR.t476 VDPWR.n2372 725.173
R7276 VDPWR.t595 VDPWR.n2375 725.173
R7277 VDPWR.t533 VDPWR.n833 725.173
R7278 VDPWR.t657 VDPWR.n837 725.173
R7279 VDPWR.n2637 VDPWR.n2636 717.729
R7280 VDPWR.n2643 VDPWR.n2642 717.729
R7281 VDPWR.n1919 VDPWR.n1916 713.462
R7282 VDPWR.n571 VDPWR.t1024 675.542
R7283 VDPWR.n291 VDPWR.t107 675.542
R7284 VDPWR.n33 VDPWR.t927 675.542
R7285 VDPWR.n879 VDPWR.t915 671.408
R7286 VDPWR.n789 VDPWR.t871 671.408
R7287 VDPWR.n3091 VDPWR.t869 671.408
R7288 VDPWR.n560 VDPWR.t146 671.376
R7289 VDPWR.n280 VDPWR.t765 671.376
R7290 VDPWR.n22 VDPWR.t988 671.376
R7291 VDPWR.n2852 VDPWR.t365 669.655
R7292 VDPWR.n1872 VDPWR.t3 667.734
R7293 VDPWR.n1966 VDPWR.t997 667.734
R7294 VDPWR.n965 VDPWR.t380 667.734
R7295 VDPWR.n2714 VDPWR.t830 667.734
R7296 VDPWR.n2714 VDPWR.t1145 667.734
R7297 VDPWR.n3045 VDPWR.t205 667.734
R7298 VDPWR.n3040 VDPWR.t213 667.734
R7299 VDPWR.n2834 VDPWR.t1135 666.677
R7300 VDPWR.n2668 VDPWR.t1161 666.677
R7301 VDPWR.n2700 VDPWR.t12 666.677
R7302 VDPWR.n2700 VDPWR.t264 666.677
R7303 VDPWR.n3024 VDPWR.t251 666.677
R7304 VDPWR.n3019 VDPWR.t10 666.677
R7305 VDPWR.t504 VDPWR 666.343
R7306 VDPWR.t717 VDPWR 666.343
R7307 VDPWR VDPWR.t752 666.343
R7308 VDPWR VDPWR.t650 666.343
R7309 VDPWR.t477 VDPWR 666.343
R7310 VDPWR.t556 VDPWR 666.343
R7311 VDPWR VDPWR.t684 664.664
R7312 VDPWR.n2657 VDPWR.t35 664.37
R7313 VDPWR.n2909 VDPWR.t813 664.279
R7314 VDPWR.n2677 VDPWR.t382 664.279
R7315 VDPWR.n2684 VDPWR.t317 664.279
R7316 VDPWR.n2938 VDPWR.t978 663.024
R7317 VDPWR.n1841 VDPWR.t175 662.571
R7318 VDPWR.n1987 VDPWR.t919 662.571
R7319 VDPWR.n2793 VDPWR.t162 659.593
R7320 VDPWR.n2417 VDPWR.t834 659.593
R7321 VDPWR.n2434 VDPWR.t325 659.593
R7322 VDPWR.n980 VDPWR.n979 642.188
R7323 VDPWR.n251 VDPWR.t892 633.369
R7324 VDPWR VDPWR.t516 630.375
R7325 VDPWR VDPWR.t435 630.375
R7326 VDPWR VDPWR.t568 630.375
R7327 VDPWR.t673 VDPWR.t619 617.668
R7328 VDPWR.t550 VDPWR.t468 617.668
R7329 VDPWR.t545 VDPWR.t559 617.668
R7330 VDPWR.n814 VDPWR.n813 614.562
R7331 VDPWR.n2860 VDPWR.n2859 613.71
R7332 VDPWR.n1968 VDPWR.n1967 611.178
R7333 VDPWR.n2633 VDPWR.n2625 611.178
R7334 VDPWR.n2657 VDPWR.n2647 611.178
R7335 VDPWR.n2782 VDPWR.n2781 610.861
R7336 VDPWR.n2773 VDPWR.n2772 609.847
R7337 VDPWR.n1001 VDPWR.n1000 609.717
R7338 VDPWR.n1057 VDPWR.n1050 609.303
R7339 VDPWR.n2202 VDPWR.n2201 606.42
R7340 VDPWR.n2231 VDPWR.n2199 606.42
R7341 VDPWR.n2205 VDPWR.n2204 606.42
R7342 VDPWR.n1062 VDPWR.n1061 606.42
R7343 VDPWR.n2282 VDPWR.n1058 606.42
R7344 VDPWR.n998 VDPWR.n997 606.42
R7345 VDPWR.n2221 VDPWR.n2208 605.581
R7346 VDPWR.n2276 VDPWR.n1064 605.581
R7347 VDPWR.n2196 VDPWR.n2195 605.186
R7348 VDPWR.n2194 VDPWR.n1098 605.186
R7349 VDPWR.n1100 VDPWR.n1099 605.186
R7350 VDPWR.n1041 VDPWR.n1040 605.186
R7351 VDPWR.n1039 VDPWR.n1038 605.186
R7352 VDPWR.n2303 VDPWR.n1035 605.186
R7353 VDPWR.n2790 VDPWR.n996 605.186
R7354 VDPWR.n2794 VDPWR.n2792 605.186
R7355 VDPWR.n2814 VDPWR.n983 605.186
R7356 VDPWR.n1990 VDPWR.n1989 604.394
R7357 VDPWR.n2830 VDPWR.n2829 604.394
R7358 VDPWR.n2620 VDPWR.n2619 604.394
R7359 VDPWR.n2649 VDPWR.n2648 604.394
R7360 VDPWR.n2587 VDPWR.n2585 604.394
R7361 VDPWR.n2587 VDPWR.n2586 604.394
R7362 VDPWR.n916 VDPWR.n915 604.394
R7363 VDPWR.n2635 VDPWR.n2634 603.231
R7364 VDPWR.n2353 VDPWR.n2352 603.231
R7365 VDPWR.n1960 VDPWR.n1927 603.052
R7366 VDPWR.n630 VDPWR.n565 602.456
R7367 VDPWR.n651 VDPWR.n540 602.456
R7368 VDPWR.n350 VDPWR.n285 602.456
R7369 VDPWR.n371 VDPWR.n260 602.456
R7370 VDPWR.n2777 VDPWR.n2776 602.456
R7371 VDPWR.n92 VDPWR.n27 602.456
R7372 VDPWR.n113 VDPWR.n2 602.456
R7373 VDPWR.n1221 VDPWR.n1220 601.097
R7374 VDPWR.n937 VDPWR.n936 601.097
R7375 VDPWR.n3014 VDPWR.n919 601.097
R7376 VDPWR.n2890 VDPWR.n2887 599.159
R7377 VDPWR.n2791 VDPWR.n995 596.442
R7378 VDPWR.n2421 VDPWR.n2419 596.442
R7379 VDPWR.n2519 VDPWR.n2436 596.442
R7380 VDPWR.n2771 VDPWR.n2770 589.481
R7381 VDPWR.n2872 VDPWR.n961 588.318
R7382 VDPWR.n546 VDPWR.n545 585
R7383 VDPWR.n544 VDPWR.n543 585
R7384 VDPWR.n266 VDPWR.n265 585
R7385 VDPWR.n264 VDPWR.n263 585
R7386 VDPWR.n2836 VDPWR.n2835 585
R7387 VDPWR.n2874 VDPWR.n2873 585
R7388 VDPWR.n2769 VDPWR.n2768 585
R7389 VDPWR.n8 VDPWR.n7 585
R7390 VDPWR.n6 VDPWR.n5 585
R7391 VDPWR.n737 VDPWR.n730 582.4
R7392 VDPWR.n733 VDPWR.n730 582.4
R7393 VDPWR.t610 VDPWR 568.994
R7394 VDPWR.t574 VDPWR 568.994
R7395 VDPWR VDPWR.t447 568.994
R7396 VDPWR.t498 VDPWR.t489 540.46
R7397 VDPWR VDPWR.n250 535.705
R7398 VDPWR.n733 VDPWR.n729 531.923
R7399 VDPWR.n738 VDPWR.n737 531.427
R7400 VDPWR.t640 VDPWR 511.926
R7401 VDPWR VDPWR.t670 510.248
R7402 VDPWR.t1081 VDPWR.t696 496.82
R7403 VDPWR VDPWR.n1166 491.784
R7404 VDPWR.n409 VDPWR.n405 480.764
R7405 VDPWR.n3157 VDPWR.n3152 480.764
R7406 VDPWR.n3141 VDPWR.n3136 480.764
R7407 VDPWR.n710 VDPWR.n706 480.764
R7408 VDPWR.n695 VDPWR.n690 480.764
R7409 VDPWR.n679 VDPWR.n674 480.764
R7410 VDPWR.n667 VDPWR.n659 480.764
R7411 VDPWR.n521 VDPWR.n517 480.764
R7412 VDPWR.n506 VDPWR.n501 480.764
R7413 VDPWR.n490 VDPWR.n485 480.764
R7414 VDPWR.n473 VDPWR.n469 480.764
R7415 VDPWR.n380 VDPWR.n378 480.764
R7416 VDPWR.n392 VDPWR.n390 480.764
R7417 VDPWR.n452 VDPWR.n447 480.764
R7418 VDPWR.n436 VDPWR.n431 480.764
R7419 VDPWR.n424 VDPWR.n416 480.764
R7420 VDPWR.n765 VDPWR.n761 480.764
R7421 VDPWR.n3124 VDPWR.n3120 480.764
R7422 VDPWR VDPWR.t370 470.562
R7423 VDPWR VDPWR.t76 470.562
R7424 VDPWR VDPWR.t246 470.562
R7425 VDPWR VDPWR.t84 470.562
R7426 VDPWR VDPWR.t90 470.562
R7427 VDPWR VDPWR.t310 470.562
R7428 VDPWR VDPWR.t273 470.562
R7429 VDPWR VDPWR.t279 470.562
R7430 VDPWR.t429 VDPWR.t456 463.252
R7431 VDPWR.t519 VDPWR.t536 463.252
R7432 VDPWR.t616 VDPWR.t441 463.252
R7433 VDPWR.t678 VDPWR.t525 463.252
R7434 VDPWR.t704 VDPWR.t640 463.252
R7435 VDPWR.t687 VDPWR.t462 463.252
R7436 VDPWR VDPWR.t699 458.724
R7437 VDPWR.t516 VDPWR 458.724
R7438 VDPWR VDPWR.t596 458.724
R7439 VDPWR.t435 VDPWR 458.724
R7440 VDPWR VDPWR.t711 458.724
R7441 VDPWR.t568 VDPWR 458.724
R7442 VDPWR.t998 VDPWR.t128 458.216
R7443 VDPWR.n749 VDPWR.n741 454.401
R7444 VDPWR.n743 VDPWR.n741 454.401
R7445 VDPWR.n743 VDPWR.n740 448.736
R7446 VDPWR.n750 VDPWR.n749 448.288
R7447 VDPWR.n178 VDPWR 435.082
R7448 VDPWR.n621 VDPWR.t943 420.25
R7449 VDPWR.n341 VDPWR.t1096 420.25
R7450 VDPWR.t904 VDPWR.n176 420.25
R7451 VDPWR.n83 VDPWR.t949 420.25
R7452 VDPWR.t653 VDPWR 414.577
R7453 VDPWR VDPWR.t492 414.577
R7454 VDPWR VDPWR.t704 414.577
R7455 VDPWR.t462 VDPWR 414.577
R7456 VDPWR.t670 VDPWR 414.577
R7457 VDPWR.n857 VDPWR.t473 390.875
R7458 VDPWR.n1257 VDPWR.t726 389.526
R7459 VDPWR.n2471 VDPWR.t735 389.361
R7460 VDPWR.n1222 VDPWR.t746 388.721
R7461 VDPWR.n320 VDPWR.t437 388.656
R7462 VDPWR.n1350 VDPWR.t505 388.656
R7463 VDPWR.n1391 VDPWR.t506 388.656
R7464 VDPWR.n1503 VDPWR.t685 388.656
R7465 VDPWR.n1292 VDPWR.t686 388.656
R7466 VDPWR.n1683 VDPWR.t718 388.656
R7467 VDPWR.n1721 VDPWR.t719 388.656
R7468 VDPWR.n1133 VDPWR.t449 388.656
R7469 VDPWR.n1602 VDPWR.t478 388.656
R7470 VDPWR.n1627 VDPWR.t479 388.656
R7471 VDPWR.n2090 VDPWR.t557 388.656
R7472 VDPWR.n2082 VDPWR.t558 388.656
R7473 VDPWR.n2179 VDPWR.t564 388.656
R7474 VDPWR.n2628 VDPWR.t484 388.656
R7475 VDPWR.n884 VDPWR.t485 388.656
R7476 VDPWR.n830 VDPWR.t544 388.656
R7477 VDPWR.n596 VDPWR.t517 388.656
R7478 VDPWR.n600 VDPWR.t518 388.656
R7479 VDPWR.n588 VDPWR.t700 388.656
R7480 VDPWR.n624 VDPWR.t701 388.656
R7481 VDPWR.n574 VDPWR.t668 388.656
R7482 VDPWR.n583 VDPWR.t669 388.656
R7483 VDPWR.n548 VDPWR.t682 388.656
R7484 VDPWR.n553 VDPWR.t683 388.656
R7485 VDPWR.n316 VDPWR.t436 388.656
R7486 VDPWR.n308 VDPWR.t597 388.656
R7487 VDPWR.n344 VDPWR.t598 388.656
R7488 VDPWR.n294 VDPWR.t600 388.656
R7489 VDPWR.n303 VDPWR.t601 388.656
R7490 VDPWR.n268 VDPWR.t540 388.656
R7491 VDPWR.n273 VDPWR.t541 388.656
R7492 VDPWR.n1179 VDPWR.t740 388.656
R7493 VDPWR.n1995 VDPWR.t741 388.656
R7494 VDPWR.n1928 VDPWR.t607 388.656
R7495 VDPWR.n2211 VDPWR.t728 388.656
R7496 VDPWR.n1019 VDPWR.t729 388.656
R7497 VDPWR.n1066 VDPWR.t697 388.656
R7498 VDPWR.n2265 VDPWR.t698 388.656
R7499 VDPWR.n2884 VDPWR.t502 388.656
R7500 VDPWR.n2889 VDPWR.t503 388.656
R7501 VDPWR.n2762 VDPWR.t573 388.656
R7502 VDPWR.n2952 VDPWR.t463 388.656
R7503 VDPWR.n2959 VDPWR.t464 388.656
R7504 VDPWR.n917 VDPWR.t554 388.656
R7505 VDPWR.n2987 VDPWR.t555 388.656
R7506 VDPWR.n2411 VDPWR.t638 388.656
R7507 VDPWR.n2420 VDPWR.t639 388.656
R7508 VDPWR.n2398 VDPWR.t439 388.656
R7509 VDPWR.n2357 VDPWR.t440 388.656
R7510 VDPWR.n2525 VDPWR.t481 388.656
R7511 VDPWR.n2437 VDPWR.t482 388.656
R7512 VDPWR.n2450 VDPWR.t671 388.656
R7513 VDPWR.n2485 VDPWR.t672 388.656
R7514 VDPWR.n792 VDPWR.t628 388.656
R7515 VDPWR.n798 VDPWR.t629 388.656
R7516 VDPWR.n864 VDPWR.t472 388.656
R7517 VDPWR.n58 VDPWR.t569 388.656
R7518 VDPWR.n62 VDPWR.t570 388.656
R7519 VDPWR.n50 VDPWR.t712 388.656
R7520 VDPWR.n86 VDPWR.t713 388.656
R7521 VDPWR.n36 VDPWR.t529 388.656
R7522 VDPWR.n45 VDPWR.t530 388.656
R7523 VDPWR.n10 VDPWR.t662 388.656
R7524 VDPWR.n15 VDPWR.t663 388.656
R7525 VDPWR.n1199 VDPWR.t747 387.682
R7526 VDPWR.n1202 VDPWR.t614 387.682
R7527 VDPWR.n2557 VDPWR.t720 387.682
R7528 VDPWR.n2562 VDPWR.t499 387.682
R7529 VDPWR.n1167 VDPWR.t739 386.043
R7530 VDPWR.n820 VDPWR.t543 385.026
R7531 VDPWR.n2091 VDPWR.t680 383.42
R7532 VDPWR VDPWR.t837 381.007
R7533 VDPWR.n1324 VDPWR.t487 380.193
R7534 VDPWR.n1351 VDPWR.t457 380.193
R7535 VDPWR.n1354 VDPWR.t646 380.193
R7536 VDPWR.n1358 VDPWR.t430 380.193
R7537 VDPWR.n1363 VDPWR.t633 380.193
R7538 VDPWR.n1538 VDPWR.t451 380.193
R7539 VDPWR.n1541 VDPWR.t648 380.193
R7540 VDPWR.n1684 VDPWR.t690 380.193
R7541 VDPWR.n1687 VDPWR.t537 380.193
R7542 VDPWR.n1691 VDPWR.t520 380.193
R7543 VDPWR.n1696 VDPWR.t702 380.193
R7544 VDPWR.n1206 VDPWR.t742 380.193
R7545 VDPWR.n1893 VDPWR.t603 380.193
R7546 VDPWR.n1604 VDPWR.t617 380.193
R7547 VDPWR.n1610 VDPWR.t694 380.193
R7548 VDPWR.n1613 VDPWR.t442 380.193
R7549 VDPWR.n1617 VDPWR.t534 380.193
R7550 VDPWR.n1937 VDPWR.t514 380.193
R7551 VDPWR.n1940 VDPWR.t592 380.193
R7552 VDPWR.n2096 VDPWR.t526 380.193
R7553 VDPWR.n2099 VDPWR.t635 380.193
R7554 VDPWR.n1069 VDPWR.t584 380.193
R7555 VDPWR.n1072 VDPWR.t692 380.193
R7556 VDPWR.n2729 VDPWR.t625 380.193
R7557 VDPWR.n2732 VDPWR.t722 380.193
R7558 VDPWR.n930 VDPWR.t676 380.193
R7559 VDPWR.n2970 VDPWR.t445 380.193
R7560 VDPWR.n2550 VDPWR.t707 380.193
R7561 VDPWR.n2553 VDPWR.t490 380.193
R7562 VDPWR.n2595 VDPWR.t496 380.193
R7563 VDPWR.n889 VDPWR.t731 380.193
R7564 VDPWR.n2989 VDPWR.t427 380.193
R7565 VDPWR.n2997 VDPWR.t548 380.193
R7566 VDPWR.n817 VDPWR.t508 380.193
R7567 VDPWR.n2371 VDPWR.t475 380.193
R7568 VDPWR.n2374 VDPWR.t594 380.193
R7569 VDPWR.n832 VDPWR.t532 380.193
R7570 VDPWR.n836 VDPWR.t656 380.193
R7571 VDPWR.n716 VDPWR.n706 379.2
R7572 VDPWR.n700 VDPWR.n690 379.2
R7573 VDPWR.n684 VDPWR.n674 379.2
R7574 VDPWR.n668 VDPWR.n667 379.2
R7575 VDPWR.n527 VDPWR.n517 379.2
R7576 VDPWR.n511 VDPWR.n501 379.2
R7577 VDPWR.n495 VDPWR.n485 379.2
R7578 VDPWR.n479 VDPWR.n469 379.2
R7579 VDPWR.n463 VDPWR.n405 379.2
R7580 VDPWR.n388 VDPWR.n378 379.2
R7581 VDPWR.n400 VDPWR.n390 379.2
R7582 VDPWR.n457 VDPWR.n447 379.2
R7583 VDPWR.n441 VDPWR.n431 379.2
R7584 VDPWR.n425 VDPWR.n424 379.2
R7585 VDPWR.n3168 VDPWR.n761 379.2
R7586 VDPWR.n3162 VDPWR.n3152 379.2
R7587 VDPWR.n3146 VDPWR.n3136 379.2
R7588 VDPWR.n3130 VDPWR.n3120 379.2
R7589 VDPWR VDPWR.t116 369.938
R7590 VDPWR VDPWR.t853 369.938
R7591 VDPWR VDPWR.t1045 369.938
R7592 VDPWR VDPWR.t237 369.938
R7593 VDPWR.t172 VDPWR 369.938
R7594 VDPWR.t182 VDPWR 369.938
R7595 VDPWR.t888 VDPWR 369.938
R7596 VDPWR.t884 VDPWR 369.938
R7597 VDPWR.t291 VDPWR 369.938
R7598 VDPWR.t842 VDPWR 369.938
R7599 VDPWR.t840 VDPWR 369.938
R7600 VDPWR.t898 VDPWR 369.938
R7601 VDPWR VDPWR.t1021 369.938
R7602 VDPWR VDPWR.t59 369.938
R7603 VDPWR VDPWR.t613 360.866
R7604 VDPWR.t619 VDPWR 357.51
R7605 VDPWR.t468 VDPWR 357.51
R7606 VDPWR.t559 VDPWR 357.51
R7607 VDPWR.t586 VDPWR 355.83
R7608 VDPWR.t157 VDPWR.t812 352.474
R7609 VDPWR.t829 VDPWR.t320 352.474
R7610 VDPWR.n141 VDPWR.t859 348.849
R7611 VDPWR.n2828 VDPWR.t774 340.212
R7612 VDPWR VDPWR.t474 337.368
R7613 VDPWR.n2177 VDPWR.t255 336.524
R7614 VDPWR.n1028 VDPWR.t1157 336.524
R7615 VDPWR.n2687 VDPWR.n2603 334.247
R7616 VDPWR VDPWR.t624 334.012
R7617 VDPWR.n1922 VDPWR.n1921 333.99
R7618 VDPWR.n1875 VDPWR.n1874 333.348
R7619 VDPWR.n953 VDPWR.n952 333.348
R7620 VDPWR.n2547 VDPWR.n2546 333.348
R7621 VDPWR.n894 VDPWR.n893 333.348
R7622 VDPWR.n2866 VDPWR.n964 333.346
R7623 VDPWR.n2608 VDPWR.n2607 333.346
R7624 VDPWR.n2547 VDPWR.n2545 333.346
R7625 VDPWR.n897 VDPWR.n896 333.346
R7626 VDPWR.n2386 VDPWR.n2366 328.036
R7627 VDPWR.n1403 VDPWR.t1192 328.005
R7628 VDPWR.n1733 VDPWR.t1286 328.005
R7629 VDPWR.n1630 VDPWR.t1208 328.005
R7630 VDPWR.n2470 VDPWR.n2461 326.202
R7631 VDPWR.n3052 VDPWR.n887 325.639
R7632 VDPWR.n1876 VDPWR.n1873 324.74
R7633 VDPWR.n577 VDPWR.n570 322.329
R7634 VDPWR.n555 VDPWR.n551 322.329
R7635 VDPWR.n297 VDPWR.n290 322.329
R7636 VDPWR.n275 VDPWR.n271 322.329
R7637 VDPWR.n2627 VDPWR.n2626 322.329
R7638 VDPWR.n796 VDPWR.n795 322.329
R7639 VDPWR.n39 VDPWR.n32 322.329
R7640 VDPWR.n17 VDPWR.n13 322.329
R7641 VDPWR.t269 VDPWR.t214 322.262
R7642 VDPWR.n1031 VDPWR.t1216 321.911
R7643 VDPWR.n140 VDPWR.n139 320.976
R7644 VDPWR.n1848 VDPWR.n1847 320.976
R7645 VDPWR.n2916 VDPWR.n2915 320.976
R7646 VDPWR.n2676 VDPWR.n2609 320.976
R7647 VDPWR.n2707 VDPWR.n2582 320.976
R7648 VDPWR.n900 VDPWR.n899 320.976
R7649 VDPWR.n1918 VDPWR.n1917 320.976
R7650 VDPWR.n2853 VDPWR.n2851 320.976
R7651 VDPWR.n2669 VDPWR.n2612 320.976
R7652 VDPWR.n2707 VDPWR.n2581 320.976
R7653 VDPWR.n3026 VDPWR.n913 320.976
R7654 VDPWR.t147 VDPWR.t11 315.548
R7655 VDPWR.t167 VDPWR.t388 315.548
R7656 VDPWR.n2816 VDPWR.n2815 315.089
R7657 VDPWR.n2824 VDPWR.n2823 314.447
R7658 VDPWR.t379 VDPWR.t308 313.87
R7659 VDPWR.n1982 VDPWR.n1981 312.829
R7660 VDPWR.n2406 VDPWR.n2355 312.053
R7661 VDPWR.n2386 VDPWR.n2368 312.053
R7662 VDPWR.n2381 VDPWR.n2370 312.053
R7663 VDPWR.n2513 VDPWR.n2441 312.053
R7664 VDPWR.n2824 VDPWR.n2822 312.051
R7665 VDPWR.n2179 VDPWR.n2178 311.151
R7666 VDPWR.n2310 VDPWR.n1030 311.151
R7667 VDPWR.n2186 VDPWR.n1102 310.904
R7668 VDPWR.n1034 VDPWR.n1033 310.904
R7669 VDPWR.n2514 VDPWR.n2438 310.5
R7670 VDPWR.t522 VDPWR.t504 308.834
R7671 VDPWR.n1430 VDPWR.t486 308.834
R7672 VDPWR.t580 VDPWR.t717 308.834
R7673 VDPWR.t752 VDPWR.t610 308.834
R7674 VDPWR.t650 VDPWR.t574 308.834
R7675 VDPWR.t577 VDPWR.t477 308.834
R7676 VDPWR.t736 VDPWR.t727 308.834
R7677 VDPWR.t571 VDPWR.t586 308.834
R7678 VDPWR.n826 VDPWR.n825 308.755
R7679 VDPWR.n800 VDPWR.n799 308.755
R7680 VDPWR.n2463 VDPWR.n2462 308.755
R7681 VDPWR.n2480 VDPWR.n2458 308.755
R7682 VDPWR.n2531 VDPWR.n2347 308.755
R7683 VDPWR VDPWR.n821 308.755
R7684 VDPWR.n1519 VDPWR.n1291 308.755
R7685 VDPWR.n2761 VDPWR.n1005 308.755
R7686 VDPWR.n2784 VDPWR.n2783 307.204
R7687 VDPWR.n2431 VDPWR.n2348 307.204
R7688 VDPWR.n1440 VDPWR.t1252 306.735
R7689 VDPWR.n1440 VDPWR.t1281 306.735
R7690 VDPWR.n1309 VDPWR.t1168 306.735
R7691 VDPWR.n1309 VDPWR.t1191 306.735
R7692 VDPWR.n1343 VDPWR.t1272 306.735
R7693 VDPWR.n1411 VDPWR.t1213 306.735
R7694 VDPWR.n1506 VDPWR.t1222 306.735
R7695 VDPWR.n1524 VDPWR.t1170 306.735
R7696 VDPWR.n1524 VDPWR.t1195 306.735
R7697 VDPWR.n1279 VDPWR.t1246 306.735
R7698 VDPWR.n1741 VDPWR.t1260 306.735
R7699 VDPWR.n1776 VDPWR.t1235 306.735
R7700 VDPWR.n1770 VDPWR.t1175 306.735
R7701 VDPWR.n1804 VDPWR.t1177 306.735
R7702 VDPWR.n1237 VDPWR.t1223 306.735
R7703 VDPWR.n1835 VDPWR.t1219 306.735
R7704 VDPWR.n1158 VDPWR.t1174 306.735
R7705 VDPWR.n1154 VDPWR.t1184 306.735
R7706 VDPWR.n1150 VDPWR.t1172 306.735
R7707 VDPWR.n1132 VDPWR.t1271 306.735
R7708 VDPWR.n1633 VDPWR.t1224 306.735
R7709 VDPWR.n1625 VDPWR.t1210 306.735
R7710 VDPWR.n2117 VDPWR.t1238 306.735
R7711 VDPWR.n2079 VDPWR.t1209 306.735
R7712 VDPWR.n2077 VDPWR.t1279 306.735
R7713 VDPWR.n2192 VDPWR.t1283 306.735
R7714 VDPWR.n2209 VDPWR.t1173 306.735
R7715 VDPWR.n1063 VDPWR.t1230 306.735
R7716 VDPWR.n950 VDPWR.t1178 306.735
R7717 VDPWR.n2945 VDPWR.t1187 306.735
R7718 VDPWR.n2456 VDPWR.t1264 306.735
R7719 VDPWR.t418 VDPWR 290.372
R7720 VDPWR VDPWR.t450 280.3
R7721 VDPWR VDPWR.t602 280.3
R7722 VDPWR.t994 VDPWR 280.3
R7723 VDPWR VDPWR.t513 280.3
R7724 VDPWR VDPWR.t583 280.3
R7725 VDPWR VDPWR.t444 280.3
R7726 VDPWR VDPWR.t426 280.3
R7727 VDPWR VDPWR.t531 280.3
R7728 VDPWR.t790 VDPWR.t220 278.623
R7729 VDPWR.n147 VDPWR.n146 272.274
R7730 VDPWR.n147 VDPWR.n134 272.274
R7731 VDPWR.n176 VDPWR.n134 272.274
R7732 VDPWR.t47 VDPWR 261.837
R7733 VDPWR VDPWR.t522 260.159
R7734 VDPWR VDPWR.t673 260.159
R7735 VDPWR VDPWR.t580 260.159
R7736 VDPWR VDPWR.t550 260.159
R7737 VDPWR.t724 VDPWR 260.159
R7738 VDPWR.t744 VDPWR 260.159
R7739 VDPWR.t613 VDPWR 260.159
R7740 VDPWR VDPWR.t577 260.159
R7741 VDPWR VDPWR.t545 260.159
R7742 VDPWR.t739 VDPWR 260.159
R7743 VDPWR.t727 VDPWR 260.159
R7744 VDPWR.t696 VDPWR 260.159
R7745 VDPWR VDPWR.t498 260.159
R7746 VDPWR VDPWR.t438 260.159
R7747 VDPWR.t922 VDPWR 260.159
R7748 VDPWR.t63 VDPWR 260.159
R7749 VDPWR.t38 VDPWR 260.159
R7750 VDPWR.n634 VDPWR.n632 259.697
R7751 VDPWR.n354 VDPWR.n352 259.697
R7752 VDPWR.n96 VDPWR.n94 259.697
R7753 VDPWR.n610 VDPWR.t854 255.905
R7754 VDPWR.n615 VDPWR.t117 255.905
R7755 VDPWR.n591 VDPWR.t944 255.905
R7756 VDPWR.n631 VDPWR.t970 255.905
R7757 VDPWR.n539 VDPWR.t187 255.905
R7758 VDPWR.n330 VDPWR.t238 255.905
R7759 VDPWR.n335 VDPWR.t1046 255.905
R7760 VDPWR.n311 VDPWR.t1097 255.905
R7761 VDPWR.n351 VDPWR.t850 255.905
R7762 VDPWR.n259 VDPWR.t177 255.905
R7763 VDPWR.n183 VDPWR.t899 255.905
R7764 VDPWR.n188 VDPWR.t841 255.905
R7765 VDPWR.n193 VDPWR.t843 255.905
R7766 VDPWR.n198 VDPWR.t292 255.905
R7767 VDPWR.n129 VDPWR.t885 255.905
R7768 VDPWR.n159 VDPWR.t889 255.905
R7769 VDPWR.n164 VDPWR.t183 255.905
R7770 VDPWR.n169 VDPWR.t173 255.905
R7771 VDPWR.n135 VDPWR.t905 255.905
R7772 VDPWR.n72 VDPWR.t60 255.905
R7773 VDPWR.n77 VDPWR.t1022 255.905
R7774 VDPWR.n53 VDPWR.t950 255.905
R7775 VDPWR.n93 VDPWR.t1138 255.905
R7776 VDPWR.n1 VDPWR.t881 255.905
R7777 VDPWR.n246 VDPWR.t371 255.904
R7778 VDPWR.n123 VDPWR.t77 255.904
R7779 VDPWR.n124 VDPWR.t247 255.904
R7780 VDPWR.n125 VDPWR.t85 255.904
R7781 VDPWR.n126 VDPWR.t91 255.904
R7782 VDPWR.n204 VDPWR.t311 255.904
R7783 VDPWR.n205 VDPWR.t274 255.904
R7784 VDPWR.n206 VDPWR.t280 255.904
R7785 VDPWR.n119 VDPWR.t893 255.904
R7786 VDPWR.n581 VDPWR.t982 254.475
R7787 VDPWR.n301 VDPWR.t1009 254.475
R7788 VDPWR.n43 VDPWR.t211 254.475
R7789 VDPWR.n606 VDPWR.t58 252.95
R7790 VDPWR.n611 VDPWR.t115 252.95
R7791 VDPWR.n616 VDPWR.t953 252.95
R7792 VDPWR.n650 VDPWR.t185 252.95
R7793 VDPWR.n645 VDPWR.t1163 252.95
R7794 VDPWR.n326 VDPWR.t234 252.95
R7795 VDPWR.n331 VDPWR.t815 252.95
R7796 VDPWR.n336 VDPWR.t1099 252.95
R7797 VDPWR.n370 VDPWR.t179 252.95
R7798 VDPWR.n365 VDPWR.t73 252.95
R7799 VDPWR.n179 VDPWR.t897 252.95
R7800 VDPWR.n184 VDPWR.t839 252.95
R7801 VDPWR.n189 VDPWR.t845 252.95
R7802 VDPWR.n194 VDPWR.t290 252.95
R7803 VDPWR.n199 VDPWR.t883 252.95
R7804 VDPWR.n155 VDPWR.t887 252.95
R7805 VDPWR.n160 VDPWR.t181 252.95
R7806 VDPWR.n165 VDPWR.t171 252.95
R7807 VDPWR.n170 VDPWR.t903 252.95
R7808 VDPWR.n68 VDPWR.t1032 252.95
R7809 VDPWR.n73 VDPWR.t929 252.95
R7810 VDPWR.n78 VDPWR.t947 252.95
R7811 VDPWR.n112 VDPWR.t879 252.95
R7812 VDPWR.n107 VDPWR.t305 252.95
R7813 VDPWR.n120 VDPWR.t369 252.948
R7814 VDPWR.n245 VDPWR.t75 252.948
R7815 VDPWR.n240 VDPWR.t245 252.948
R7816 VDPWR.n235 VDPWR.t87 252.948
R7817 VDPWR.n230 VDPWR.t89 252.948
R7818 VDPWR.n225 VDPWR.t313 252.948
R7819 VDPWR.n220 VDPWR.t276 252.948
R7820 VDPWR.n215 VDPWR.t278 252.948
R7821 VDPWR.n210 VDPWR.t895 252.948
R7822 VDPWR.n630 VDPWR.t980 251.516
R7823 VDPWR.n350 VDPWR.t1011 251.516
R7824 VDPWR.n92 VDPWR.t209 251.516
R7825 VDPWR.n541 VDPWR.t1165 250.724
R7826 VDPWR.n261 VDPWR.t71 250.724
R7827 VDPWR.n3 VDPWR.t307 250.724
R7828 VDPWR.n144 VDPWR.t241 249.363
R7829 VDPWR.t943 VDPWR.t952 248.599
R7830 VDPWR.t116 VDPWR.t114 248.599
R7831 VDPWR.t853 VDPWR.t57 248.599
R7832 VDPWR.t1096 VDPWR.t1098 248.599
R7833 VDPWR.t1045 VDPWR.t814 248.599
R7834 VDPWR.t237 VDPWR.t233 248.599
R7835 VDPWR.t370 VDPWR.t368 248.599
R7836 VDPWR.t76 VDPWR.t74 248.599
R7837 VDPWR.t246 VDPWR.t244 248.599
R7838 VDPWR.t84 VDPWR.t86 248.599
R7839 VDPWR.t90 VDPWR.t88 248.599
R7840 VDPWR.t310 VDPWR.t312 248.599
R7841 VDPWR.t273 VDPWR.t275 248.599
R7842 VDPWR.t279 VDPWR.t277 248.599
R7843 VDPWR.t892 VDPWR.t894 248.599
R7844 VDPWR.t860 VDPWR.t858 248.599
R7845 VDPWR.t242 VDPWR.t860 248.599
R7846 VDPWR.t240 VDPWR.t242 248.599
R7847 VDPWR.t902 VDPWR.t904 248.599
R7848 VDPWR.t170 VDPWR.t172 248.599
R7849 VDPWR.t180 VDPWR.t182 248.599
R7850 VDPWR.t886 VDPWR.t888 248.599
R7851 VDPWR.t882 VDPWR.t884 248.599
R7852 VDPWR.t289 VDPWR.t291 248.599
R7853 VDPWR.t844 VDPWR.t842 248.599
R7854 VDPWR.t838 VDPWR.t840 248.599
R7855 VDPWR.t896 VDPWR.t898 248.599
R7856 VDPWR.t949 VDPWR.t946 248.599
R7857 VDPWR.t1021 VDPWR.t928 248.599
R7858 VDPWR.t59 VDPWR.t1031 248.599
R7859 VDPWR.n633 VDPWR.t972 248.219
R7860 VDPWR.n353 VDPWR.t852 248.219
R7861 VDPWR.n95 VDPWR.t1137 248.219
R7862 VDPWR.n2093 VDPWR.t1188 246.71
R7863 VDPWR.n1325 VDPWR.t1244 245.667
R7864 VDPWR.n1352 VDPWR.t1258 245.667
R7865 VDPWR.n1355 VDPWR.t1225 245.667
R7866 VDPWR.n1359 VDPWR.t1262 245.667
R7867 VDPWR.n1364 VDPWR.t1233 245.667
R7868 VDPWR.n1539 VDPWR.t1257 245.667
R7869 VDPWR.n1542 VDPWR.t1226 245.667
R7870 VDPWR.n1685 VDPWR.t1221 245.667
R7871 VDPWR.n1688 VDPWR.t1266 245.667
R7872 VDPWR.n1692 VDPWR.t1227 245.667
R7873 VDPWR.n1697 VDPWR.t1197 245.667
R7874 VDPWR.n1207 VDPWR.t1220 245.667
R7875 VDPWR.n1894 VDPWR.t1242 245.667
R7876 VDPWR.n1605 VDPWR.t1186 245.667
R7877 VDPWR.n1611 VDPWR.t1169 245.667
R7878 VDPWR.n1614 VDPWR.t1251 245.667
R7879 VDPWR.n1618 VDPWR.t1229 245.667
R7880 VDPWR.n1938 VDPWR.t1232 245.667
R7881 VDPWR.n1941 VDPWR.t1203 245.667
R7882 VDPWR.n2097 VDPWR.t1254 245.667
R7883 VDPWR.n2100 VDPWR.t1183 245.667
R7884 VDPWR.n1070 VDPWR.t1234 245.667
R7885 VDPWR.n1073 VDPWR.t1167 245.667
R7886 VDPWR.n2730 VDPWR.t1218 245.667
R7887 VDPWR.n2733 VDPWR.t1277 245.667
R7888 VDPWR.n931 VDPWR.t1190 245.667
R7889 VDPWR.n2971 VDPWR.t1253 245.667
R7890 VDPWR.n2551 VDPWR.t1179 245.667
R7891 VDPWR.n2554 VDPWR.t1278 245.667
R7892 VDPWR.n2596 VDPWR.t1267 245.667
R7893 VDPWR.n890 VDPWR.t1180 245.667
R7894 VDPWR.n2990 VDPWR.t1285 245.667
R7895 VDPWR.n2998 VDPWR.t1256 245.667
R7896 VDPWR.n818 VDPWR.t1265 245.667
R7897 VDPWR.n2372 VDPWR.t1274 245.667
R7898 VDPWR.n2375 VDPWR.t1211 245.667
R7899 VDPWR.n833 VDPWR.t1248 245.667
R7900 VDPWR.n837 VDPWR.t1185 245.667
R7901 VDPWR.n962 VDPWR.t796 245.064
R7902 VDPWR.n1182 VDPWR.t103 243.512
R7903 VDPWR.n797 VDPWR.t129 241.767
R7904 VDPWR.n2946 VDPWR.t873 240.215
R7905 VDPWR.n2987 VDPWR.t877 240.214
R7906 VDPWR.n1828 VDPWR.t1181 235.319
R7907 VDPWR.n2432 VDPWR.t7 234.982
R7908 VDPWR VDPWR.t872 233.304
R7909 VDPWR.t733 VDPWR.t846 231.625
R7910 VDPWR.t795 VDPWR.t14 229.947
R7911 VDPWR.n146 VDPWR 224.923
R7912 VDPWR.n2405 VDPWR.n2356 223.868
R7913 VDPWR.t831 VDPWR 223.233
R7914 VDPWR.t318 VDPWR 223.233
R7915 VDPWR.n621 VDPWR 221.964
R7916 VDPWR.n341 VDPWR 221.964
R7917 VDPWR.n83 VDPWR 221.964
R7918 VDPWR.t168 VDPWR.t26 221.555
R7919 VDPWR.t920 VDPWR.t1053 221.555
R7920 VDPWR.t200 VDPWR.t198 221.555
R7921 VDPWR.n2633 VDPWR.n2623 221.314
R7922 VDPWR.n1259 VDPWR.t1189 215.827
R7923 VDPWR.n2473 VDPWR.t1280 215.827
R7924 VDPWR VDPWR.t153 213.163
R7925 VDPWR VDPWR.t974 213.163
R7926 VDPWR.n1200 VDPWR.t1166 213.148
R7927 VDPWR.n1203 VDPWR.t1237 213.148
R7928 VDPWR.n2558 VDPWR.t1176 213.148
R7929 VDPWR.n2563 VDPWR.t1276 213.148
R7930 VDPWR.n581 VDPWR.n578 213.119
R7931 VDPWR.n301 VDPWR.n298 213.119
R7932 VDPWR.n43 VDPWR.n40 213.119
R7933 VDPWR.n622 VDPWR.n621 213.119
R7934 VDPWR.n641 VDPWR.n640 213.119
R7935 VDPWR.n342 VDPWR.n341 213.119
R7936 VDPWR.n361 VDPWR.n360 213.119
R7937 VDPWR.n176 VDPWR.n175 213.119
R7938 VDPWR.n136 VDPWR.n134 213.119
R7939 VDPWR.n148 VDPWR.n147 213.119
R7940 VDPWR.n146 VDPWR.n145 213.119
R7941 VDPWR.n2811 VDPWR.n954 213.119
R7942 VDPWR.n3053 VDPWR.n886 213.119
R7943 VDPWR.n3096 VDPWR.n791 213.119
R7944 VDPWR.n84 VDPWR.n83 213.119
R7945 VDPWR.n103 VDPWR.n102 213.119
R7946 VDPWR.n533 VDPWR.t942 212.081
R7947 VDPWR.n534 VDPWR.t951 212.081
R7948 VDPWR.n3173 VDPWR.t948 212.081
R7949 VDPWR.n3174 VDPWR.t945 212.081
R7950 VDPWR.n1106 VDPWR.t1240 211.263
R7951 VDPWR.n598 VDPWR.t1205 210.964
R7952 VDPWR.n589 VDPWR.t1261 210.964
R7953 VDPWR.n575 VDPWR.t1214 210.964
R7954 VDPWR.n550 VDPWR.t1207 210.964
R7955 VDPWR.n318 VDPWR.t1263 210.964
R7956 VDPWR.n309 VDPWR.t1201 210.964
R7957 VDPWR.n295 VDPWR.t1200 210.964
R7958 VDPWR.n270 VDPWR.t1228 210.964
R7959 VDPWR.n1181 VDPWR.t1275 210.964
R7960 VDPWR.n1018 VDPWR.t1273 210.964
R7961 VDPWR.n1068 VDPWR.t1284 210.964
R7962 VDPWR.n2885 VDPWR.t1236 210.964
R7963 VDPWR.n878 VDPWR.t1270 210.964
R7964 VDPWR.n2399 VDPWR.t1269 210.964
R7965 VDPWR.n60 VDPWR.t1215 210.964
R7966 VDPWR.n51 VDPWR.t1282 210.964
R7967 VDPWR.n37 VDPWR.t1268 210.964
R7968 VDPWR.n12 VDPWR.t1217 210.964
R7969 VDPWR.n1431 VDPWR.n1430 209.368
R7970 VDPWR.n1825 VDPWR.n1223 209.368
R7971 VDPWR.n1760 VDPWR.n1262 209.368
R7972 VDPWR.n2001 VDPWR.n1167 209.368
R7973 VDPWR.n1166 VDPWR.n1126 209.368
R7974 VDPWR.n2317 VDPWR.n1024 209.368
R7975 VDPWR.n1110 VDPWR.n1109 209.368
R7976 VDPWR.n2813 VDPWR.n2812 209.368
R7977 VDPWR.n2686 VDPWR.n2685 209.368
R7978 VDPWR.t267 VDPWR 206.45
R7979 VDPWR VDPWR.t744 203.093
R7980 VDPWR.t447 VDPWR 203.093
R7981 VDPWR.t749 VDPWR 203.093
R7982 VDPWR.t643 VDPWR 203.093
R7983 VDPWR VDPWR.t471 203.093
R7984 VDPWR VDPWR.t918 201.413
R7985 VDPWR VDPWR.t992 199.736
R7986 VDPWR VDPWR.t194 199.736
R7987 VDPWR.t952 VDPWR 198.287
R7988 VDPWR.t114 VDPWR 198.287
R7989 VDPWR.t57 VDPWR 198.287
R7990 VDPWR.t1098 VDPWR 198.287
R7991 VDPWR.t814 VDPWR 198.287
R7992 VDPWR.t233 VDPWR 198.287
R7993 VDPWR VDPWR.t902 198.287
R7994 VDPWR VDPWR.t170 198.287
R7995 VDPWR VDPWR.t180 198.287
R7996 VDPWR VDPWR.t886 198.287
R7997 VDPWR VDPWR.t882 198.287
R7998 VDPWR VDPWR.t289 198.287
R7999 VDPWR VDPWR.t844 198.287
R8000 VDPWR VDPWR.t838 198.287
R8001 VDPWR VDPWR.t896 198.287
R8002 VDPWR.t946 VDPWR 198.287
R8003 VDPWR.t928 VDPWR 198.287
R8004 VDPWR.t1031 VDPWR 198.287
R8005 VDPWR.t1150 VDPWR.t202 198.058
R8006 VDPWR.n2051 VDPWR.n2050 197.508
R8007 VDPWR.t25 VDPWR.t2 191.344
R8008 VDPWR.t812 VDPWR.t803 191.344
R8009 VDPWR.t152 VDPWR.t829 191.344
R8010 VDPWR.t1146 VDPWR.t248 189.665
R8011 VDPWR VDPWR.t240 189.409
R8012 VDPWR.n2811 VDPWR 184.63
R8013 VDPWR.n791 VDPWR 184.63
R8014 VDPWR.n643 VDPWR.n642 183.673
R8015 VDPWR.n363 VDPWR.n362 183.673
R8016 VDPWR.n105 VDPWR.n104 183.673
R8017 VDPWR.n535 VDPWR.n534 183.441
R8018 VDPWR.n3175 VDPWR.n3174 183.441
R8019 VDPWR VDPWR.t4 182.952
R8020 VDPWR VDPWR.n641 182.952
R8021 VDPWR.t287 VDPWR 182.952
R8022 VDPWR VDPWR.t302 182.952
R8023 VDPWR VDPWR.n361 182.952
R8024 VDPWR.t285 VDPWR 182.952
R8025 VDPWR VDPWR.t429 182.952
R8026 VDPWR.t486 VDPWR 182.952
R8027 VDPWR.t450 VDPWR 182.952
R8028 VDPWR VDPWR.t519 182.952
R8029 VDPWR.n1223 VDPWR 182.952
R8030 VDPWR.t602 VDPWR 182.952
R8031 VDPWR VDPWR.t616 182.952
R8032 VDPWR.t513 VDPWR 182.952
R8033 VDPWR.t583 VDPWR 182.952
R8034 VDPWR.t444 VDPWR 182.952
R8035 VDPWR.t426 VDPWR 182.952
R8036 VDPWR.t507 VDPWR 182.952
R8037 VDPWR.t531 VDPWR 182.952
R8038 VDPWR VDPWR.t206 182.952
R8039 VDPWR VDPWR.n103 182.952
R8040 VDPWR.t260 VDPWR 182.952
R8041 VDPWR.t1132 VDPWR.t354 181.273
R8042 VDPWR.n1429 VDPWR 179.595
R8043 VDPWR.n1262 VDPWR 179.595
R8044 VDPWR.n1109 VDPWR 179.595
R8045 VDPWR.n1024 VDPWR 179.595
R8046 VDPWR.n2432 VDPWR 179.595
R8047 VDPWR.t356 VDPWR.t1040 174.559
R8048 VDPWR.t227 VDPWR.t799 174.559
R8049 VDPWR.t165 VDPWR.t168 172.881
R8050 VDPWR.t1053 VDPWR.t155 172.881
R8051 VDPWR.t149 VDPWR.t200 172.881
R8052 VDPWR.t1000 VDPWR.t80 172.881
R8053 VDPWR.t914 VDPWR 169.524
R8054 VDPWR.t1040 VDPWR.t833 167.845
R8055 VDPWR.t163 VDPWR.t453 164.488
R8056 VDPWR.t366 VDPWR.t1148 162.81
R8057 VDPWR.t862 VDPWR.t293 162.81
R8058 VDPWR.t250 VDPWR.t973 161.131
R8059 VDPWR.t912 VDPWR.t352 161.131
R8060 VDPWR.n545 VDPWR.n544 159.476
R8061 VDPWR.n265 VDPWR.n264 159.476
R8062 VDPWR.n2873 VDPWR.n2872 159.476
R8063 VDPWR.n2770 VDPWR.n2769 159.476
R8064 VDPWR.n7 VDPWR.n6 159.476
R8065 VDPWR.t24 VDPWR.t165 159.452
R8066 VDPWR.t827 VDPWR.t983 159.452
R8067 VDPWR.t190 VDPWR.t986 159.452
R8068 VDPWR.t155 VDPWR.t804 159.452
R8069 VDPWR.t198 VDPWR.t150 159.452
R8070 VDPWR.t151 VDPWR.t149 159.452
R8071 VDPWR.t142 VDPWR.t283 159.452
R8072 VDPWR.t962 VDPWR.t542 157.774
R8073 VDPWR.n632 VDPWR.t925 157.014
R8074 VDPWR.n352 VDPWR.t105 157.014
R8075 VDPWR.n94 VDPWR.t931 157.014
R8076 VDPWR.t1164 VDPWR.t910 154.417
R8077 VDPWR.t70 VDPWR.t1089 154.417
R8078 VDPWR.t684 VDPWR.t653 154.417
R8079 VDPWR.t346 VDPWR.t134 154.417
R8080 VDPWR.t492 VDPWR.t556 154.417
R8081 VDPWR.t973 VDPWR.t334 154.417
R8082 VDPWR.t306 VDPWR.t55 154.417
R8083 VDPWR VDPWR.t126 152.739
R8084 VDPWR.t453 VDPWR.t174 151.06
R8085 VDPWR.t501 VDPWR.t1141 151.06
R8086 VDPWR.t324 VDPWR.t480 151.06
R8087 VDPWR.t1002 VDPWR.t94 149.382
R8088 VDPWR.t932 VDPWR.t47 149.382
R8089 VDPWR.t30 VDPWR.t924 147.703
R8090 VDPWR.t848 VDPWR.t104 147.703
R8091 VDPWR.t1087 VDPWR.t40 147.703
R8092 VDPWR.t954 VDPWR.t900 147.703
R8093 VDPWR.t194 VDPWR.t22 147.703
R8094 VDPWR.t7 VDPWR.t801 147.703
R8095 VDPWR.t223 VDPWR.t922 147.703
R8096 VDPWR.t159 VDPWR.t63 147.703
R8097 VDPWR.t757 VDPWR.t962 147.703
R8098 VDPWR.t938 VDPWR.t78 147.703
R8099 VDPWR.t960 VDPWR.t930 147.703
R8100 VDPWR.t759 VDPWR.t932 144.346
R8101 VDPWR.t254 VDPWR.t1019 144.346
R8102 VDPWR.t258 VDPWR.t256 144.346
R8103 VDPWR.t256 VDPWR.t416 144.346
R8104 VDPWR.t416 VDPWR.t410 144.346
R8105 VDPWR.t410 VDPWR.t420 144.346
R8106 VDPWR.t420 VDPWR.t424 144.346
R8107 VDPWR.t424 VDPWR.t396 144.346
R8108 VDPWR.t400 VDPWR.t422 144.346
R8109 VDPWR.t422 VDPWR.t394 144.346
R8110 VDPWR.t398 VDPWR.t402 144.346
R8111 VDPWR.t402 VDPWR.t412 144.346
R8112 VDPWR.t406 VDPWR.t408 144.346
R8113 VDPWR.t408 VDPWR.t404 144.346
R8114 VDPWR.t404 VDPWR.t414 144.346
R8115 VDPWR.t414 VDPWR.t418 144.346
R8116 VDPWR.t1156 VDPWR.t1152 144.346
R8117 VDPWR.t1152 VDPWR.t779 144.346
R8118 VDPWR.t779 VDPWR.t1154 144.346
R8119 VDPWR.t1154 VDPWR.t1061 144.346
R8120 VDPWR.t1061 VDPWR.t1067 144.346
R8121 VDPWR.t1071 VDPWR.t1075 144.346
R8122 VDPWR.t1075 VDPWR.t1065 144.346
R8123 VDPWR.t1065 VDPWR.t1069 144.346
R8124 VDPWR.t1069 VDPWR.t1073 144.346
R8125 VDPWR.t1073 VDPWR.t1063 144.346
R8126 VDPWR.t1079 VDPWR.t1085 144.346
R8127 VDPWR.t1085 VDPWR.t1057 144.346
R8128 VDPWR.t1057 VDPWR.t1059 144.346
R8129 VDPWR.t1059 VDPWR.t1083 144.346
R8130 VDPWR.t1083 VDPWR.t1055 144.346
R8131 VDPWR.t1055 VDPWR.t1077 144.346
R8132 VDPWR.t1112 VDPWR.t1118 144.346
R8133 VDPWR.t1122 VDPWR.t1130 144.346
R8134 VDPWR.t1116 VDPWR.t1126 144.346
R8135 VDPWR.t1106 VDPWR.t1108 144.346
R8136 VDPWR.t775 VDPWR.t773 144.346
R8137 VDPWR.t799 VDPWR.t297 144.346
R8138 VDPWR.t174 VDPWR.t24 142.668
R8139 VDPWR.t394 VDPWR.t398 142.668
R8140 VDPWR.t1124 VDPWR.t1120 142.668
R8141 VDPWR.t804 VDPWR.t977 142.668
R8142 VDPWR.t11 VDPWR.t151 142.668
R8143 VDPWR.t1160 VDPWR.t1000 142.668
R8144 VDPWR.t1033 VDPWR.t1023 140.989
R8145 VDPWR.t924 VDPWR.t971 140.989
R8146 VDPWR.t184 VDPWR.t186 140.989
R8147 VDPWR.t1162 VDPWR.t1164 140.989
R8148 VDPWR.t145 VDPWR.t328 140.989
R8149 VDPWR.t1091 VDPWR.t106 140.989
R8150 VDPWR.t104 VDPWR.t851 140.989
R8151 VDPWR.t178 VDPWR.t176 140.989
R8152 VDPWR.t72 VDPWR.t70 140.989
R8153 VDPWR.t764 VDPWR.t61 140.989
R8154 VDPWR.t825 VDPWR.t163 140.989
R8155 VDPWR.t42 VDPWR.t936 140.989
R8156 VDPWR.t992 VDPWR.t994 140.989
R8157 VDPWR.t810 VDPWR.t157 140.989
R8158 VDPWR.t803 VDPWR.t156 140.989
R8159 VDPWR.t153 VDPWR.t390 140.989
R8160 VDPWR.t320 VDPWR.t831 140.989
R8161 VDPWR.t150 VDPWR.t152 140.989
R8162 VDPWR.t783 VDPWR.t147 140.989
R8163 VDPWR.t80 VDPWR.t322 140.989
R8164 VDPWR.t1029 VDPWR.t221 140.989
R8165 VDPWR.t771 VDPWR.t326 140.989
R8166 VDPWR.t337 VDPWR.t336 140.989
R8167 VDPWR.t974 VDPWR.t392 140.989
R8168 VDPWR.t96 VDPWR.t387 140.989
R8169 VDPWR.t805 VDPWR.t96 140.989
R8170 VDPWR.t868 VDPWR.t916 140.989
R8171 VDPWR.t908 VDPWR.t926 140.989
R8172 VDPWR.t930 VDPWR.t1136 140.989
R8173 VDPWR.t878 VDPWR.t880 140.989
R8174 VDPWR.t304 VDPWR.t306 140.989
R8175 VDPWR.t987 VDPWR.t792 140.989
R8176 VDPWR.n533 VDPWR.t1193 139.78
R8177 VDPWR.n534 VDPWR.t1202 139.78
R8178 VDPWR.n3173 VDPWR.t1206 139.78
R8179 VDPWR.n3174 VDPWR.t1212 139.78
R8180 VDPWR.t1148 VDPWR.t1134 139.311
R8181 VDPWR.t936 VDPWR.t906 137.633
R8182 VDPWR.t940 VDPWR.t0 137.633
R8183 VDPWR.n632 VDPWR.t29 137.079
R8184 VDPWR.n352 VDPWR.t111 137.079
R8185 VDPWR.n94 VDPWR.t1039 137.079
R8186 VDPWR.t348 VDPWR.t133 135.954
R8187 VDPWR.t781 VDPWR.t331 135.954
R8188 VDPWR.t92 VDPWR.t231 135.954
R8189 VDPWR.t81 VDPWR.t797 135.954
R8190 VDPWR.t294 VDPWR.t1015 135.954
R8191 VDPWR.t876 VDPWR 135.954
R8192 VDPWR.n2835 VDPWR.t93 135.268
R8193 VDPWR.t300 VDPWR.t1049 134.276
R8194 VDPWR.t336 VDPWR.t212 130.919
R8195 VDPWR.t338 VDPWR.t890 130.919
R8196 VDPWR.n934 VDPWR.t1247 129.344
R8197 VDPWR.n3015 VDPWR.t1250 129.344
R8198 VDPWR.n863 VDPWR.t1259 129.344
R8199 VDPWR.n2524 VDPWR.t1255 129.344
R8200 VDPWR.n2351 VDPWR.t1194 129.344
R8201 VDPWR VDPWR.t166 129.24
R8202 VDPWR.n2453 VDPWR.t1182 127.695
R8203 VDPWR.t866 VDPWR.t1114 127.562
R8204 VDPWR.n2685 VDPWR.t316 127.562
R8205 VDPWR.t350 VDPWR.t358 127.562
R8206 VDPWR VDPWR.t1132 127.562
R8207 VDPWR.n578 VDPWR 125.883
R8208 VDPWR.n642 VDPWR 125.883
R8209 VDPWR.n298 VDPWR 125.883
R8210 VDPWR.n362 VDPWR 125.883
R8211 VDPWR.t456 VDPWR 125.883
R8212 VDPWR.n1430 VDPWR 125.883
R8213 VDPWR VDPWR.n1429 125.883
R8214 VDPWR.t536 VDPWR 125.883
R8215 VDPWR.n1262 VDPWR 125.883
R8216 VDPWR VDPWR.n1223 125.883
R8217 VDPWR.t441 VDPWR 125.883
R8218 VDPWR.n1166 VDPWR 125.883
R8219 VDPWR.n1167 VDPWR 125.883
R8220 VDPWR.t525 VDPWR 125.883
R8221 VDPWR.n1109 VDPWR 125.883
R8222 VDPWR VDPWR.n1024 125.883
R8223 VDPWR.t624 VDPWR 125.883
R8224 VDPWR.t828 VDPWR.t362 125.883
R8225 VDPWR VDPWR.n2811 125.883
R8226 VDPWR.t489 VDPWR 125.883
R8227 VDPWR.n2685 VDPWR 125.883
R8228 VDPWR.t283 VDPWR.t381 125.883
R8229 VDPWR.t755 VDPWR.t98 125.883
R8230 VDPWR VDPWR.n886 125.883
R8231 VDPWR.t474 VDPWR 125.883
R8232 VDPWR VDPWR.n791 125.883
R8233 VDPWR.n40 VDPWR 125.883
R8234 VDPWR.n104 VDPWR 125.883
R8235 VDPWR.n2741 VDPWR.t1231 124.953
R8236 VDPWR.t968 VDPWR.t1112 124.206
R8237 VDPWR.t316 VDPWR.t383 124.206
R8238 VDPWR.t32 VDPWR.t1025 124.206
R8239 VDPWR.t46 VDPWR 122.526
R8240 VDPWR.t1128 VDPWR.t360 122.526
R8241 VDPWR.t1102 VDPWR.t1042 122.526
R8242 VDPWR.n2812 VDPWR.t1106 122.526
R8243 VDPWR.t53 VDPWR.t1143 122.526
R8244 VDPWR.t589 VDPWR.t1081 120.849
R8245 VDPWR.t299 VDPWR.t364 120.849
R8246 VDPWR.t872 VDPWR.t1044 120.849
R8247 VDPWR.t967 VDPWR.t876 120.849
R8248 VDPWR.n823 VDPWR.t1245 120.76
R8249 VDPWR.n2727 VDPWR.t1204 119.007
R8250 VDPWR.n1925 VDPWR.t1196 118.853
R8251 VDPWR.n2835 VDPWR.t1048 118.549
R8252 VDPWR.t202 VDPWR.t991 117.492
R8253 VDPWR.n2783 VDPWR.t361 117.451
R8254 VDPWR.n2348 VDPWR.t1052 117.451
R8255 VDPWR.n2438 VDPWR.t298 117.451
R8256 VDPWR.n1505 VDPWR.t1171 117.294
R8257 VDPWR.n2116 VDPWR.t1243 117.294
R8258 VDPWR.n3090 VDPWR.t1198 117.294
R8259 VDPWR.n2461 VDPWR.t127 116.343
R8260 VDPWR.n570 VDPWR.t1034 116.341
R8261 VDPWR.n551 VDPWR.t329 116.341
R8262 VDPWR.n290 VDPWR.t1092 116.341
R8263 VDPWR.n271 VDPWR.t62 116.341
R8264 VDPWR.n2626 VDPWR.t355 116.341
R8265 VDPWR.n795 VDPWR.t917 116.341
R8266 VDPWR.n32 VDPWR.t909 116.341
R8267 VDPWR.n13 VDPWR.t793 116.341
R8268 VDPWR.t1027 VDPWR 115.814
R8269 VDPWR.n2859 VDPWR.t363 114.918
R8270 VDPWR.n813 VDPWR.t1147 114.918
R8271 VDPWR.n1349 VDPWR.t1239 114.546
R8272 VDPWR.n1682 VDPWR.t1199 114.546
R8273 VDPWR.n1623 VDPWR.t1241 114.546
R8274 VDPWR.t102 VDPWR.t136 114.135
R8275 VDPWR.t1120 VDPWR.t262 114.135
R8276 VDPWR.n1847 VDPWR.t169 113.98
R8277 VDPWR.n1917 VDPWR.t1003 113.98
R8278 VDPWR.n2851 VDPWR.t232 113.98
R8279 VDPWR.n2915 VDPWR.t1054 113.98
R8280 VDPWR.n2612 VDPWR.t1001 113.98
R8281 VDPWR.n2609 VDPWR.t376 113.98
R8282 VDPWR.n2582 VDPWR.t201 113.98
R8283 VDPWR.n2581 VDPWR.t794 113.98
R8284 VDPWR.n913 VDPWR.t891 113.98
R8285 VDPWR.n899 VDPWR.t865 113.98
R8286 VDPWR.t1023 VDPWR 112.457
R8287 VDPWR.t971 VDPWR 112.457
R8288 VDPWR VDPWR.t145 112.457
R8289 VDPWR.t106 VDPWR 112.457
R8290 VDPWR.t851 VDPWR 112.457
R8291 VDPWR VDPWR.t764 112.457
R8292 VDPWR VDPWR.t868 112.457
R8293 VDPWR.t926 VDPWR 112.457
R8294 VDPWR.t1136 VDPWR 112.457
R8295 VDPWR VDPWR.t987 112.457
R8296 VDPWR.t1004 VDPWR 110.778
R8297 VDPWR.t1019 VDPWR 110.778
R8298 VDPWR.t204 VDPWR.t36 110.778
R8299 VDPWR VDPWR.t964 109.1
R8300 VDPWR VDPWR.t188 109.1
R8301 VDPWR.t40 VDPWR 109.1
R8302 VDPWR VDPWR.t954 109.1
R8303 VDPWR VDPWR.t385 109.1
R8304 VDPWR.t1141 VDPWR 109.1
R8305 VDPWR.t100 VDPWR 109.1
R8306 VDPWR.t192 VDPWR 109.1
R8307 VDPWR VDPWR.t140 109.1
R8308 VDPWR VDPWR.t807 109.1
R8309 VDPWR.t51 VDPWR 109.1
R8310 VDPWR.t248 VDPWR 109.1
R8311 VDPWR.t78 VDPWR 109.1
R8312 VDPWR VDPWR.t216 109.1
R8313 VDPWR.t6 VDPWR 107.421
R8314 VDPWR.t934 VDPWR.t996 107.421
R8315 VDPWR.t1044 VDPWR 107.421
R8316 VDPWR.t553 VDPWR 107.421
R8317 VDPWR.n1429 VDPWR.n1297 106.561
R8318 VDPWR.n2433 VDPWR.n2432 106.559
R8319 VDPWR.n717 VDPWR.n705 105.788
R8320 VDPWR.n701 VDPWR.n689 105.788
R8321 VDPWR.n685 VDPWR.n673 105.788
R8322 VDPWR.n669 VDPWR.n658 105.788
R8323 VDPWR.n528 VDPWR.n516 105.788
R8324 VDPWR.n512 VDPWR.n500 105.788
R8325 VDPWR.n496 VDPWR.n484 105.788
R8326 VDPWR.n480 VDPWR.n468 105.788
R8327 VDPWR.n464 VDPWR.n404 105.788
R8328 VDPWR.n458 VDPWR.n446 105.788
R8329 VDPWR.n442 VDPWR.n430 105.788
R8330 VDPWR.n426 VDPWR.n415 105.788
R8331 VDPWR.n3169 VDPWR.n760 105.788
R8332 VDPWR.n3163 VDPWR.n3151 105.788
R8333 VDPWR.n3147 VDPWR.n3135 105.788
R8334 VDPWR.n3131 VDPWR.n3119 105.788
R8335 VDPWR VDPWR.t664 105.743
R8336 VDPWR VDPWR.t658 105.743
R8337 VDPWR VDPWR.t571 105.743
R8338 VDPWR.t510 VDPWR 105.743
R8339 VDPWR.t265 VDPWR.t38 105.743
R8340 VDPWR.t667 VDPWR.t1033 104.064
R8341 VDPWR.t328 VDPWR.t681 104.064
R8342 VDPWR.t599 VDPWR.t1091 104.064
R8343 VDPWR.t61 VDPWR.t539 104.064
R8344 VDPWR.t1104 VDPWR 104.064
R8345 VDPWR.t1158 VDPWR 104.064
R8346 VDPWR VDPWR.t835 104.064
R8347 VDPWR.t916 VDPWR.t627 104.064
R8348 VDPWR.t528 VDPWR.t908 104.064
R8349 VDPWR.t792 VDPWR.t661 104.064
R8350 VDPWR.t855 VDPWR 102.385
R8351 VDPWR.t235 VDPWR 102.385
R8352 VDPWR.t377 VDPWR.t795 102.385
R8353 VDPWR.t977 VDPWR 102.385
R8354 VDPWR.t34 VDPWR 102.385
R8355 VDPWR.t542 VDPWR 102.385
R8356 VDPWR.t130 VDPWR 102.385
R8357 VDPWR.n2050 VDPWR.n2049 101.591
R8358 VDPWR VDPWR.t20 100.707
R8359 VDPWR.t981 VDPWR 99.0288
R8360 VDPWR.t1008 VDPWR 99.0288
R8361 VDPWR.t630 VDPWR.t1071 99.0288
R8362 VDPWR.t14 VDPWR 99.0288
R8363 VDPWR VDPWR.t768 99.0288
R8364 VDPWR.t210 VDPWR 99.0288
R8365 VDPWR.t368 VDPWR 97.6641
R8366 VDPWR.t74 VDPWR 97.6641
R8367 VDPWR.t244 VDPWR 97.6641
R8368 VDPWR.t86 VDPWR 97.6641
R8369 VDPWR.t88 VDPWR 97.6641
R8370 VDPWR.t312 VDPWR 97.6641
R8371 VDPWR.t275 VDPWR 97.6641
R8372 VDPWR.t277 VDPWR 97.6641
R8373 VDPWR.t894 VDPWR 97.6641
R8374 VDPWR.t1047 VDPWR.t827 97.3503
R8375 VDPWR.n565 VDPWR.t31 96.1553
R8376 VDPWR.n540 VDPWR.t19 96.1553
R8377 VDPWR.n285 VDPWR.t849 96.1553
R8378 VDPWR.n260 VDPWR.t990 96.1553
R8379 VDPWR.n979 VDPWR.t1149 96.1553
R8380 VDPWR.n2887 VDPWR.t23 96.1553
R8381 VDPWR.n2776 VDPWR.t867 96.1553
R8382 VDPWR.n27 VDPWR.t961 96.1553
R8383 VDPWR.n2 VDPWR.t197 96.1553
R8384 VDPWR.t381 VDPWR.t375 95.6719
R8385 VDPWR.t375 VDPWR.t817 95.6719
R8386 VDPWR.t83 VDPWR.t766 95.6719
R8387 VDPWR.n1916 VDPWR.t45 93.81
R8388 VDPWR.n2636 VDPWR.t756 93.81
R8389 VDPWR.n2642 VDPWR.t798 93.81
R8390 VDPWR.n746 VDPWR.n741 92.5005
R8391 VDPWR.n742 VDPWR.n740 92.5005
R8392 VDPWR VDPWR.t18 92.315
R8393 VDPWR VDPWR.t989 92.315
R8394 VDPWR.t1100 VDPWR.t225 92.315
R8395 VDPWR VDPWR.t196 92.315
R8396 VDPWR.t166 VDPWR.t857 90.6365
R8397 VDPWR.t483 VDPWR.t914 90.6365
R8398 VDPWR.t976 VDPWR.t333 90.6365
R8399 VDPWR.t271 VDPWR.t338 90.6365
R8400 VDPWR.n744 VDPWR.n742 89.0328
R8401 VDPWR.n747 VDPWR.n746 89.0328
R8402 VDPWR.t412 VDPWR 88.9581
R8403 VDPWR.t65 VDPWR.t44 87.2797
R8404 VDPWR.t124 VDPWR.t870 87.2797
R8405 VDPWR VDPWR.t966 87.2797
R8406 VDPWR.n544 VDPWR.t911 86.7743
R8407 VDPWR.n264 VDPWR.t1090 86.7743
R8408 VDPWR.n2872 VDPWR.t195 86.7743
R8409 VDPWR.n2770 VDPWR.t969 86.7743
R8410 VDPWR.n995 VDPWR.t1043 86.7743
R8411 VDPWR.n995 VDPWR.t226 86.7743
R8412 VDPWR.n2419 VDPWR.t1041 86.7743
R8413 VDPWR.n2419 VDPWR.t357 86.7743
R8414 VDPWR.n2436 VDPWR.t228 86.7743
R8415 VDPWR.n2436 VDPWR.t800 86.7743
R8416 VDPWR.n6 VDPWR.t56 86.7743
R8417 VDPWR VDPWR.t1079 85.6012
R8418 VDPWR.t837 VDPWR 85.6012
R8419 VDPWR.n578 VDPWR.t981 83.9228
R8420 VDPWR.n298 VDPWR.t1008 83.9228
R8421 VDPWR.t135 VDPWR.t1017 83.9228
R8422 VDPWR.t132 VDPWR.t934 83.9228
R8423 VDPWR.t768 VDPWR.t495 83.9228
R8424 VDPWR.n40 VDPWR.t210 83.9228
R8425 VDPWR.t773 VDPWR 82.2443
R8426 VDPWR.t864 VDPWR.t976 82.2443
R8427 VDPWR.n641 VDPWR.t28 80.5659
R8428 VDPWR.n361 VDPWR.t110 80.5659
R8429 VDPWR.t777 VDPWR 80.5659
R8430 VDPWR.t156 VDPWR.t714 80.5659
R8431 VDPWR.t390 VDPWR 80.5659
R8432 VDPWR VDPWR.t783 80.5659
R8433 VDPWR.t785 VDPWR 80.5659
R8434 VDPWR.t36 VDPWR.t337 80.5659
R8435 VDPWR.t392 VDPWR 80.5659
R8436 VDPWR.n103 VDPWR.t1038 80.5659
R8437 VDPWR.t364 VDPWR.t190 78.8874
R8438 VDPWR.t714 VDPWR.t920 78.8874
R8439 VDPWR.t138 VDPWR.t1160 78.8874
R8440 VDPWR VDPWR.t1051 78.8874
R8441 VDPWR.t297 VDPWR 78.8874
R8442 VDPWR.t4 VDPWR.t667 77.209
R8443 VDPWR.t681 VDPWR.t287 77.209
R8444 VDPWR.t302 VDPWR.t599 77.209
R8445 VDPWR.t539 VDPWR.t285 77.209
R8446 VDPWR.t817 VDPWR.t143 77.209
R8447 VDPWR.t627 VDPWR.t998 77.209
R8448 VDPWR.t471 VDPWR.t507 77.209
R8449 VDPWR.t206 VDPWR.t528 77.209
R8450 VDPWR.t661 VDPWR.t260 77.209
R8451 VDPWR.t396 VDPWR.t432 75.5305
R8452 VDPWR.t161 VDPWR.t1100 75.5305
R8453 VDPWR VDPWR.t912 75.5305
R8454 VDPWR.t1051 VDPWR 75.5305
R8455 VDPWR.t339 VDPWR.n734 75.1466
R8456 VDPWR.n736 VDPWR.t343 75.1466
R8457 VDPWR.t2 VDPWR.t42 73.8521
R8458 VDPWR.t767 VDPWR.t1139 73.8521
R8459 VDPWR.t326 VDPWR.t730 73.8521
R8460 VDPWR.t9 VDPWR 73.8521
R8461 VDPWR.t94 VDPWR.t65 72.1736
R8462 VDPWR.t44 VDPWR.t135 72.1736
R8463 VDPWR.t1108 VDPWR 72.1736
R8464 VDPWR VDPWR.t777 72.1736
R8465 VDPWR.n745 VDPWR.n744 70.6952
R8466 VDPWR.n748 VDPWR.n747 70.6952
R8467 VDPWR.t432 VDPWR.t400 68.8168
R8468 VDPWR.t1110 VDPWR.t161 68.8168
R8469 VDPWR.t333 VDPWR.t271 68.8168
R8470 VDPWR VDPWR.t356 68.8168
R8471 VDPWR VDPWR.t810 67.1383
R8472 VDPWR.t383 VDPWR.t767 67.1383
R8473 VDPWR.t1139 VDPWR.t142 67.1383
R8474 VDPWR.t730 VDPWR.t1027 67.1383
R8475 VDPWR.t966 VDPWR 67.1383
R8476 VDPWR.n545 VDPWR.t965 66.8398
R8477 VDPWR.n265 VDPWR.t189 66.8398
R8478 VDPWR.n2873 VDPWR.t15 66.8398
R8479 VDPWR.n2769 VDPWR.t268 66.8398
R8480 VDPWR.n7 VDPWR.t217 66.8398
R8481 VDPWR.t362 VDPWR.t379 65.4599
R8482 VDPWR VDPWR.t771 65.4599
R8483 VDPWR.t387 VDPWR 65.4599
R8484 VDPWR.n387 VDPWR.n379 64.4072
R8485 VDPWR.n399 VDPWR.n391 64.4072
R8486 VDPWR.t1006 VDPWR.t828 63.7814
R8487 VDPWR.t143 VDPWR.t83 63.7814
R8488 VDPWR.t766 VDPWR.t138 63.7814
R8489 VDPWR.n700 VDPWR.n699 63.3551
R8490 VDPWR.n684 VDPWR.n683 63.3551
R8491 VDPWR.n511 VDPWR.n510 63.3551
R8492 VDPWR.n495 VDPWR.n494 63.3551
R8493 VDPWR.n457 VDPWR.n456 63.3551
R8494 VDPWR.n441 VDPWR.n440 63.3551
R8495 VDPWR.n3162 VDPWR.n3161 63.3551
R8496 VDPWR.n3146 VDPWR.n3145 63.3551
R8497 VDPWR.n565 VDPWR.t856 63.3219
R8498 VDPWR.n540 VDPWR.t789 63.3219
R8499 VDPWR.n285 VDPWR.t236 63.3219
R8500 VDPWR.n260 VDPWR.t109 63.3219
R8501 VDPWR.n1967 VDPWR.t1018 63.3219
R8502 VDPWR.n1967 VDPWR.t935 63.3219
R8503 VDPWR.n2887 VDPWR.t1142 63.3219
R8504 VDPWR.n2776 VDPWR.t386 63.3219
R8505 VDPWR.n2625 VDPWR.t351 63.3219
R8506 VDPWR.n2625 VDPWR.t101 63.3219
R8507 VDPWR.n2647 VDPWR.t1030 63.3219
R8508 VDPWR.n2647 VDPWR.t222 63.3219
R8509 VDPWR.n27 VDPWR.t131 63.3219
R8510 VDPWR.n2 VDPWR.t113 63.3219
R8511 VDPWR.n716 VDPWR.n715 62.2257
R8512 VDPWR.n527 VDPWR.n526 62.2257
R8513 VDPWR.n463 VDPWR.n462 62.2257
R8514 VDPWR.n3168 VDPWR.n3167 62.2257
R8515 VDPWR VDPWR.t30 62.103
R8516 VDPWR VDPWR.t848 62.103
R8517 VDPWR.t816 VDPWR 62.103
R8518 VDPWR VDPWR.t960 62.103
R8519 VDPWR.n711 VDPWR.n710 61.6672
R8520 VDPWR.n714 VDPWR.n713 61.6672
R8521 VDPWR.n696 VDPWR.n695 61.6672
R8522 VDPWR.n699 VDPWR.n698 61.6672
R8523 VDPWR.n680 VDPWR.n679 61.6672
R8524 VDPWR.n683 VDPWR.n682 61.6672
R8525 VDPWR.n660 VDPWR.n659 61.6672
R8526 VDPWR.n662 VDPWR.n661 61.6672
R8527 VDPWR.n522 VDPWR.n521 61.6672
R8528 VDPWR.n525 VDPWR.n524 61.6672
R8529 VDPWR.n507 VDPWR.n506 61.6672
R8530 VDPWR.n510 VDPWR.n509 61.6672
R8531 VDPWR.n491 VDPWR.n490 61.6672
R8532 VDPWR.n494 VDPWR.n493 61.6672
R8533 VDPWR.n474 VDPWR.n473 61.6672
R8534 VDPWR.n477 VDPWR.n476 61.6672
R8535 VDPWR.n410 VDPWR.n409 61.6672
R8536 VDPWR.n413 VDPWR.n412 61.6672
R8537 VDPWR.n381 VDPWR.n380 61.6672
R8538 VDPWR.n393 VDPWR.n392 61.6672
R8539 VDPWR.n453 VDPWR.n452 61.6672
R8540 VDPWR.n456 VDPWR.n455 61.6672
R8541 VDPWR.n437 VDPWR.n436 61.6672
R8542 VDPWR.n440 VDPWR.n439 61.6672
R8543 VDPWR.n417 VDPWR.n416 61.6672
R8544 VDPWR.n419 VDPWR.n418 61.6672
R8545 VDPWR.n766 VDPWR.n765 61.6672
R8546 VDPWR.n769 VDPWR.n768 61.6672
R8547 VDPWR.n3158 VDPWR.n3157 61.6672
R8548 VDPWR.n3161 VDPWR.n3160 61.6672
R8549 VDPWR.n3142 VDPWR.n3141 61.6672
R8550 VDPWR.n3145 VDPWR.n3144 61.6672
R8551 VDPWR.n3125 VDPWR.n3124 61.6672
R8552 VDPWR.n3128 VDPWR.n3127 61.6672
R8553 VDPWR.n668 VDPWR.n657 61.4728
R8554 VDPWR.n479 VDPWR.n478 61.4728
R8555 VDPWR.n425 VDPWR.n414 61.4728
R8556 VDPWR.n3130 VDPWR.n3129 61.4728
R8557 VDPWR.n534 VDPWR.n533 61.346
R8558 VDPWR.n3174 VDPWR.n3173 61.346
R8559 VDPWR.n383 VDPWR.n379 60.9564
R8560 VDPWR.n384 VDPWR.n381 60.9564
R8561 VDPWR.n395 VDPWR.n391 60.9564
R8562 VDPWR.n396 VDPWR.n393 60.9564
R8563 VDPWR.t870 VDPWR.t51 60.4245
R8564 VDPWR.t293 VDPWR.t864 58.7461
R8565 VDPWR VDPWR.t1002 57.0676
R8566 VDPWR.t1017 VDPWR.t132 57.0676
R8567 VDPWR.t1063 VDPWR 57.0676
R8568 VDPWR.t495 VDPWR.t318 57.0676
R8569 VDPWR.t910 VDPWR 55.3892
R8570 VDPWR.t1089 VDPWR 55.3892
R8571 VDPWR VDPWR.t406 55.3892
R8572 VDPWR.t55 VDPWR 55.3892
R8573 VDPWR VDPWR.t1156 53.7107
R8574 VDPWR.t788 VDPWR 52.0323
R8575 VDPWR.t108 VDPWR 52.0323
R8576 VDPWR VDPWR.t1087 52.0323
R8577 VDPWR VDPWR.t825 52.0323
R8578 VDPWR VDPWR.t1013 52.0323
R8579 VDPWR VDPWR.t736 52.0323
R8580 VDPWR.t900 VDPWR 52.0323
R8581 VDPWR.t225 VDPWR.t1102 52.0323
R8582 VDPWR VDPWR.t16 52.0323
R8583 VDPWR VDPWR.t1158 52.0323
R8584 VDPWR VDPWR.t1006 52.0323
R8585 VDPWR VDPWR.t34 52.0323
R8586 VDPWR VDPWR.t1029 52.0323
R8587 VDPWR.t835 VDPWR 52.0323
R8588 VDPWR.t20 VDPWR 52.0323
R8589 VDPWR.t295 VDPWR 52.0323
R8590 VDPWR.t801 VDPWR 52.0323
R8591 VDPWR VDPWR.t324 52.0323
R8592 VDPWR VDPWR.t159 52.0323
R8593 VDPWR VDPWR.t124 52.0323
R8594 VDPWR VDPWR.t874 52.0323
R8595 VDPWR VDPWR.t757 52.0323
R8596 VDPWR VDPWR.t938 52.0323
R8597 VDPWR.t112 VDPWR 52.0323
R8598 VDPWR.n2050 VDPWR.t1249 50.5057
R8599 VDPWR.t857 VDPWR.t25 50.3539
R8600 VDPWR VDPWR.t687 50.3539
R8601 VDPWR.t354 VDPWR.t483 50.3539
R8602 VDPWR VDPWR.t967 50.3539
R8603 VDPWR VDPWR.t724 48.6754
R8604 VDPWR VDPWR.t605 48.6754
R8605 VDPWR VDPWR.t562 48.6754
R8606 VDPWR VDPWR.t553 48.6754
R8607 VDPWR.t637 VDPWR 48.6754
R8608 VDPWR VDPWR.t510 48.6754
R8609 VDPWR VDPWR.t733 48.6754
R8610 VDPWR.n2051 VDPWR.n1130 46.0805
R8611 VDPWR VDPWR.t28 45.3185
R8612 VDPWR VDPWR.t110 45.3185
R8613 VDPWR.t1067 VDPWR.t630 45.3185
R8614 VDPWR.t1134 VDPWR.t1047 45.3185
R8615 VDPWR VDPWR.t790 45.3185
R8616 VDPWR VDPWR.t229 45.3185
R8617 VDPWR VDPWR.t1038 45.3185
R8618 VDPWR VDPWR.t192 43.6401
R8619 VDPWR.t140 VDPWR 43.6401
R8620 VDPWR.n2783 VDPWR.t263 42.3555
R8621 VDPWR.n2348 VDPWR.t374 42.3555
R8622 VDPWR.n2438 VDPWR.t230 42.3555
R8623 VDPWR VDPWR.t979 41.9616
R8624 VDPWR VDPWR.t1010 41.9616
R8625 VDPWR.t874 VDPWR.t265 41.9616
R8626 VDPWR VDPWR.t208 41.9616
R8627 VDPWR.n1220 VDPWR.t826 41.5552
R8628 VDPWR.n1220 VDPWR.t164 41.5552
R8629 VDPWR.n1989 VDPWR.t1014 41.5552
R8630 VDPWR.n1989 VDPWR.t137 41.5552
R8631 VDPWR.n2829 VDPWR.t1159 41.5552
R8632 VDPWR.n2829 VDPWR.t985 41.5552
R8633 VDPWR.n936 VDPWR.t154 41.5552
R8634 VDPWR.n936 VDPWR.t391 41.5552
R8635 VDPWR.n2619 VDPWR.t82 41.5552
R8636 VDPWR.n2619 VDPWR.t786 41.5552
R8637 VDPWR.n2648 VDPWR.t144 41.5552
R8638 VDPWR.n2648 VDPWR.t323 41.5552
R8639 VDPWR.n2585 VDPWR.t770 41.5552
R8640 VDPWR.n2585 VDPWR.t787 41.5552
R8641 VDPWR.n2586 VDPWR.t148 41.5552
R8642 VDPWR.n2586 VDPWR.t784 41.5552
R8643 VDPWR.n915 VDPWR.t335 41.5552
R8644 VDPWR.n915 VDPWR.t1016 41.5552
R8645 VDPWR.n919 VDPWR.t975 41.5552
R8646 VDPWR.n919 VDPWR.t393 41.5552
R8647 VDPWR.t821 VDPWR.t339 40.7512
R8648 VDPWR.t218 VDPWR.t821 40.7512
R8649 VDPWR.t252 VDPWR.t218 40.7512
R8650 VDPWR.t823 VDPWR.t341 40.7512
R8651 VDPWR.t819 VDPWR.t823 40.7512
R8652 VDPWR.t343 VDPWR.t819 40.7512
R8653 VDPWR VDPWR.t1110 40.2832
R8654 VDPWR.t308 VDPWR.t53 38.6047
R8655 VDPWR.n385 VDPWR.n384 38.5759
R8656 VDPWR.n383 VDPWR.n382 38.5759
R8657 VDPWR.n397 VDPWR.n396 38.5759
R8658 VDPWR.n395 VDPWR.n394 38.5759
R8659 VDPWR VDPWR.t984 36.9263
R8660 VDPWR.t983 VDPWR.t92 36.9263
R8661 VDPWR.t220 VDPWR.t32 36.9263
R8662 VDPWR.n1981 VDPWR.t347 36.4455
R8663 VDPWR.n1291 VDPWR.t1088 36.1587
R8664 VDPWR.n1291 VDPWR.t41 36.1587
R8665 VDPWR.n1005 VDPWR.t901 36.1587
R8666 VDPWR.n1005 VDPWR.t955 36.1587
R8667 VDPWR.n2822 VDPWR.t17 36.1587
R8668 VDPWR.n2822 VDPWR.t332 36.1587
R8669 VDPWR.n825 VDPWR.t939 36.1587
R8670 VDPWR.n825 VDPWR.t79 36.1587
R8671 VDPWR.n799 VDPWR.t875 36.1587
R8672 VDPWR.n799 VDPWR.t39 36.1587
R8673 VDPWR.n2462 VDPWR.t125 36.1587
R8674 VDPWR.n2462 VDPWR.t52 36.1587
R8675 VDPWR.n2458 VDPWR.t160 36.1587
R8676 VDPWR.n2458 VDPWR.t64 36.1587
R8677 VDPWR.n2347 VDPWR.t802 36.1587
R8678 VDPWR.n2347 VDPWR.t8 36.1587
R8679 VDPWR.n2355 VDPWR.t296 36.1587
R8680 VDPWR.n2355 VDPWR.t301 36.1587
R8681 VDPWR.n2368 VDPWR.t97 36.1587
R8682 VDPWR.n2368 VDPWR.t808 36.1587
R8683 VDPWR.n2370 VDPWR.t836 36.1587
R8684 VDPWR.n2370 VDPWR.t141 36.1587
R8685 VDPWR.n2441 VDPWR.t224 36.1587
R8686 VDPWR.n2441 VDPWR.t923 36.1587
R8687 VDPWR.n821 VDPWR.t758 36.1587
R8688 VDPWR.n821 VDPWR.t963 36.1587
R8689 VDPWR.n1847 VDPWR.t27 35.4605
R8690 VDPWR.n1917 VDPWR.t66 35.4605
R8691 VDPWR.n2851 VDPWR.t191 35.4605
R8692 VDPWR.n2915 VDPWR.t921 35.4605
R8693 VDPWR.n2612 VDPWR.t139 35.4605
R8694 VDPWR.n2609 VDPWR.t284 35.4605
R8695 VDPWR.n2582 VDPWR.t199 35.4605
R8696 VDPWR.n2581 VDPWR.t818 35.4605
R8697 VDPWR.n913 VDPWR.t272 35.4605
R8698 VDPWR.n899 VDPWR.t863 35.4605
R8699 VDPWR.t1025 VDPWR.t755 35.2479
R8700 VDPWR.n1969 VDPWR.n1920 34.6358
R8701 VDPWR.n2531 VDPWR.n2530 34.6358
R8702 VDPWR.n2469 VDPWR.n2463 34.6358
R8703 VDPWR.n3079 VDPWR.n800 34.6358
R8704 VDPWR.n1866 VDPWR.n1211 34.6358
R8705 VDPWR.n1870 VDPWR.n1211 34.6358
R8706 VDPWR.n1881 VDPWR.n1209 34.6358
R8707 VDPWR.n1882 VDPWR.n1881 34.6358
R8708 VDPWR.n1969 VDPWR.n1968 34.6358
R8709 VDPWR.n1980 VDPWR.n1186 34.6358
R8710 VDPWR.n2854 VDPWR.n2850 34.6358
R8711 VDPWR.n2858 VDPWR.n967 34.6358
R8712 VDPWR.n2868 VDPWR.n2867 34.6358
R8713 VDPWR.n2641 VDPWR.n2621 34.6358
R8714 VDPWR.n2679 VDPWR.n2678 34.6358
R8715 VDPWR.n2675 VDPWR.n2610 34.6358
R8716 VDPWR.n2671 VDPWR.n2610 34.6358
R8717 VDPWR.n2671 VDPWR.n2670 34.6358
R8718 VDPWR.n2683 VDPWR.n2605 34.6358
R8719 VDPWR.n2567 VDPWR.n2566 34.6358
R8720 VDPWR.n2713 VDPWR.n2712 34.6358
R8721 VDPWR.n2712 VDPWR.n2579 34.6358
R8722 VDPWR.n2708 VDPWR.n2579 34.6358
R8723 VDPWR.n2706 VDPWR.n2705 34.6358
R8724 VDPWR.n2705 VDPWR.n2583 34.6358
R8725 VDPWR.n2701 VDPWR.n2583 34.6358
R8726 VDPWR.n3050 VDPWR.n892 34.6358
R8727 VDPWR.n912 VDPWR.n911 34.6358
R8728 VDPWR.n3027 VDPWR.n912 34.6358
R8729 VDPWR.n2385 VDPWR.n2369 34.6358
R8730 VDPWR.n2512 VDPWR.n2442 34.6358
R8731 VDPWR.n812 VDPWR.n808 34.6358
R8732 VDPWR.n2623 VDPWR.t359 34.4755
R8733 VDPWR.n2356 VDPWR.t1050 34.4755
R8734 VDPWR.n2789 VDPWR.n2788 33.6462
R8735 VDPWR.n2796 VDPWR.n2795 33.6462
R8736 VDPWR.n2813 VDPWR.n984 33.6462
R8737 VDPWR VDPWR.t258 33.5694
R8738 VDPWR.t128 VDPWR 33.5694
R8739 VDPWR.n2859 VDPWR.t1007 33.4905
R8740 VDPWR.n2623 VDPWR.t193 33.4905
R8741 VDPWR.n2356 VDPWR.t21 33.4905
R8742 VDPWR.n813 VDPWR.t249 33.4905
R8743 VDPWR.n979 VDPWR.t367 32.7439
R8744 VDPWR.n388 VDPWR.n387 32.5881
R8745 VDPWR.n400 VDPWR.n399 32.5881
R8746 VDPWR.n2634 VDPWR.t1026 32.5055
R8747 VDPWR.n2634 VDPWR.t99 32.5055
R8748 VDPWR.n2352 VDPWR.t353 32.5055
R8749 VDPWR.n2352 VDPWR.t913 32.5055
R8750 VDPWR.n1983 VDPWR.n1184 32.377
R8751 VDPWR.n2850 VDPWR.n969 32.2581
R8752 VDPWR.n1988 VDPWR.n1987 32.0005
R8753 VDPWR.t1126 VDPWR 31.891
R8754 VDPWR.n752 VDPWR.t373 31.6605
R8755 VDPWR.n2679 VDPWR.n2608 31.624
R8756 VDPWR.n2578 VDPWR.n2547 31.624
R8757 VDPWR.n3046 VDPWR.n894 31.624
R8758 VDPWR.n3041 VDPWR.n897 31.624
R8759 VDPWR.n143 VDPWR.n140 30.8711
R8760 VDPWR.n1876 VDPWR.n1875 30.8711
R8761 VDPWR.n2866 VDPWR.n2865 30.8711
R8762 VDPWR.n2817 VDPWR.n2816 30.7205
R8763 VDPWR.n1927 VDPWR.t48 30.5355
R8764 VDPWR.n1877 VDPWR.n1872 30.4946
R8765 VDPWR.n2714 VDPWR.n2578 30.4946
R8766 VDPWR.n3046 VDPWR.n3045 30.4946
R8767 VDPWR.n3041 VDPWR.n3040 30.4946
R8768 VDPWR.t26 VDPWR 30.2125
R8769 VDPWR VDPWR.t678 30.2125
R8770 VDPWR.t1118 VDPWR.t267 30.2125
R8771 VDPWR.t262 VDPWR.t1116 30.2125
R8772 VDPWR.t98 VDPWR.t350 30.2125
R8773 VDPWR.t214 VDPWR.t204 30.2125
R8774 VDPWR.n2431 VDPWR.n2430 29.3652
R8775 VDPWR.n2785 VDPWR.n2782 29.2576
R8776 VDPWR.n2875 VDPWR.n2871 29.1064
R8777 VDPWR.n723 VDPWR.t340 28.6596
R8778 VDPWR.n725 VDPWR.t344 28.6583
R8779 VDPWR.n642 VDPWR 28.5341
R8780 VDPWR.n362 VDPWR 28.5341
R8781 VDPWR.n886 VDPWR 28.5341
R8782 VDPWR.t212 VDPWR.t862 28.5341
R8783 VDPWR.t846 VDPWR 28.5341
R8784 VDPWR.n104 VDPWR 28.5341
R8785 VDPWR.n2626 VDPWR.t1133 28.4453
R8786 VDPWR.n570 VDPWR.t5 28.4453
R8787 VDPWR.n551 VDPWR.t288 28.4453
R8788 VDPWR.n290 VDPWR.t303 28.4453
R8789 VDPWR.n271 VDPWR.t286 28.4453
R8790 VDPWR.n795 VDPWR.t999 28.4453
R8791 VDPWR.n32 VDPWR.t207 28.4453
R8792 VDPWR.n13 VDPWR.t261 28.4453
R8793 VDPWR.n2461 VDPWR.t847 28.4433
R8794 VDPWR.n1981 VDPWR.t1005 27.5805
R8795 VDPWR.n1927 VDPWR.t933 27.5805
R8796 VDPWR.n1050 VDPWR.t1064 27.5805
R8797 VDPWR.n2178 VDPWR.t1020 27.5805
R8798 VDPWR.n2178 VDPWR.t259 27.5805
R8799 VDPWR.n2201 VDPWR.t403 27.5805
R8800 VDPWR.n2201 VDPWR.t413 27.5805
R8801 VDPWR.n2199 VDPWR.t395 27.5805
R8802 VDPWR.n2195 VDPWR.t401 27.5805
R8803 VDPWR.n2195 VDPWR.t423 27.5805
R8804 VDPWR.n1098 VDPWR.t425 27.5805
R8805 VDPWR.n1098 VDPWR.t397 27.5805
R8806 VDPWR.n1099 VDPWR.t411 27.5805
R8807 VDPWR.n1099 VDPWR.t421 27.5805
R8808 VDPWR.n1102 VDPWR.t257 27.5805
R8809 VDPWR.n1102 VDPWR.t417 27.5805
R8810 VDPWR.n2208 VDPWR.t405 27.5805
R8811 VDPWR.n2208 VDPWR.t415 27.5805
R8812 VDPWR.n2204 VDPWR.t407 27.5805
R8813 VDPWR.n2204 VDPWR.t409 27.5805
R8814 VDPWR.n1030 VDPWR.t1153 27.5805
R8815 VDPWR.n1030 VDPWR.t780 27.5805
R8816 VDPWR.n1040 VDPWR.t1070 27.5805
R8817 VDPWR.n1040 VDPWR.t1074 27.5805
R8818 VDPWR.n1038 VDPWR.t1076 27.5805
R8819 VDPWR.n1038 VDPWR.t1066 27.5805
R8820 VDPWR.n1035 VDPWR.t1068 27.5805
R8821 VDPWR.n1035 VDPWR.t1072 27.5805
R8822 VDPWR.n1033 VDPWR.t1155 27.5805
R8823 VDPWR.n1033 VDPWR.t1062 27.5805
R8824 VDPWR.n1064 VDPWR.t1056 27.5805
R8825 VDPWR.n1064 VDPWR.t1078 27.5805
R8826 VDPWR.n1061 VDPWR.t1060 27.5805
R8827 VDPWR.n1061 VDPWR.t1084 27.5805
R8828 VDPWR.n1058 VDPWR.t1086 27.5805
R8829 VDPWR.n1058 VDPWR.t1058 27.5805
R8830 VDPWR.n2823 VDPWR.t782 27.5805
R8831 VDPWR.n2823 VDPWR.t776 27.5805
R8832 VDPWR.n2815 VDPWR.t1109 27.5805
R8833 VDPWR.n2815 VDPWR.t778 27.5805
R8834 VDPWR.n2772 VDPWR.t1113 27.5805
R8835 VDPWR.n2772 VDPWR.t1115 27.5805
R8836 VDPWR.n1000 VDPWR.t1131 27.5805
R8837 VDPWR.n1000 VDPWR.t1123 27.5805
R8838 VDPWR.n2781 VDPWR.t1127 27.5805
R8839 VDPWR.n2781 VDPWR.t1117 27.5805
R8840 VDPWR.n997 VDPWR.t1125 27.5805
R8841 VDPWR.n996 VDPWR.t1129 27.5805
R8842 VDPWR.n996 VDPWR.t1103 27.5805
R8843 VDPWR.n2792 VDPWR.t1101 27.5805
R8844 VDPWR.n2792 VDPWR.t1111 27.5805
R8845 VDPWR.n983 VDPWR.t1105 27.5805
R8846 VDPWR.n983 VDPWR.t1107 27.5805
R8847 VDPWR.n2837 VDPWR.n2834 27.4829
R8848 VDPWR.n2860 VDPWR.n2858 27.4829
R8849 VDPWR.n2635 VDPWR.n2633 27.4829
R8850 VDPWR.n2701 VDPWR.n2700 27.4829
R8851 VDPWR.n3025 VDPWR.n3024 27.4829
R8852 VDPWR.n1499 VDPWR.n1498 27.0566
R8853 VDPWR.n2904 VDPWR.n2902 27.0566
R8854 VDPWR.n1916 VDPWR.t95 26.9729
R8855 VDPWR.n2636 VDPWR.t33 26.9729
R8856 VDPWR.n2642 VDPWR.t791 26.9729
R8857 VDPWR.t1013 VDPWR.t102 26.8556
R8858 VDPWR.n1866 VDPWR.n1865 26.7859
R8859 VDPWR.n645 VDPWR.n644 26.7299
R8860 VDPWR.n365 VDPWR.n364 26.7299
R8861 VDPWR.n107 VDPWR.n106 26.7299
R8862 VDPWR.n2684 VDPWR.n2683 26.7299
R8863 VDPWR.n139 VDPWR.t861 26.5955
R8864 VDPWR.n139 VDPWR.t243 26.5955
R8865 VDPWR.n1873 VDPWR.t937 26.5955
R8866 VDPWR.n1873 VDPWR.t941 26.5955
R8867 VDPWR.n1874 VDPWR.t907 26.5955
R8868 VDPWR.n1874 VDPWR.t1 26.5955
R8869 VDPWR.n1921 VDPWR.t993 26.5955
R8870 VDPWR.n1921 VDPWR.t995 26.5955
R8871 VDPWR.n1050 VDPWR.t1080 26.5955
R8872 VDPWR.n2199 VDPWR.t399 26.5955
R8873 VDPWR.n964 VDPWR.t54 26.5955
R8874 VDPWR.n964 VDPWR.t378 26.5955
R8875 VDPWR.n997 VDPWR.t1121 26.5955
R8876 VDPWR.n952 VDPWR.t811 26.5955
R8877 VDPWR.n952 VDPWR.t158 26.5955
R8878 VDPWR.n2607 VDPWR.t384 26.5955
R8879 VDPWR.n2607 VDPWR.t1140 26.5955
R8880 VDPWR.n2546 VDPWR.t1144 26.5955
R8881 VDPWR.n2546 VDPWR.t330 26.5955
R8882 VDPWR.n2545 VDPWR.t832 26.5955
R8883 VDPWR.n2545 VDPWR.t321 26.5955
R8884 VDPWR.n2603 VDPWR.t319 26.5955
R8885 VDPWR.n2603 VDPWR.t769 26.5955
R8886 VDPWR.n887 VDPWR.t327 26.5955
R8887 VDPWR.n887 VDPWR.t1028 26.5955
R8888 VDPWR.n893 VDPWR.t203 26.5955
R8889 VDPWR.n893 VDPWR.t270 26.5955
R8890 VDPWR.n896 VDPWR.t215 26.5955
R8891 VDPWR.n896 VDPWR.t37 26.5955
R8892 VDPWR.n2366 VDPWR.t809 26.5955
R8893 VDPWR.n2366 VDPWR.t806 26.5955
R8894 VDPWR.n856 VDPWR.n820 26.3341
R8895 VDPWR.n144 VDPWR.n143 25.977
R8896 VDPWR.n644 VDPWR.n643 25.6953
R8897 VDPWR.n364 VDPWR.n363 25.6953
R8898 VDPWR.n106 VDPWR.n105 25.6953
R8899 VDPWR.n610 VDPWR.n594 25.224
R8900 VDPWR.n606 VDPWR.n594 25.224
R8901 VDPWR.n615 VDPWR.n593 25.224
R8902 VDPWR.n611 VDPWR.n593 25.224
R8903 VDPWR.n617 VDPWR.n591 25.224
R8904 VDPWR.n617 VDPWR.n616 25.224
R8905 VDPWR.n635 VDPWR.n631 25.224
R8906 VDPWR.n330 VDPWR.n314 25.224
R8907 VDPWR.n326 VDPWR.n314 25.224
R8908 VDPWR.n335 VDPWR.n313 25.224
R8909 VDPWR.n331 VDPWR.n313 25.224
R8910 VDPWR.n337 VDPWR.n311 25.224
R8911 VDPWR.n337 VDPWR.n336 25.224
R8912 VDPWR.n355 VDPWR.n351 25.224
R8913 VDPWR.n247 VDPWR.n120 25.224
R8914 VDPWR.n247 VDPWR.n246 25.224
R8915 VDPWR.n245 VDPWR.n244 25.224
R8916 VDPWR.n244 VDPWR.n123 25.224
R8917 VDPWR.n240 VDPWR.n239 25.224
R8918 VDPWR.n239 VDPWR.n124 25.224
R8919 VDPWR.n235 VDPWR.n234 25.224
R8920 VDPWR.n234 VDPWR.n125 25.224
R8921 VDPWR.n230 VDPWR.n229 25.224
R8922 VDPWR.n229 VDPWR.n126 25.224
R8923 VDPWR.n225 VDPWR.n224 25.224
R8924 VDPWR.n224 VDPWR.n204 25.224
R8925 VDPWR.n220 VDPWR.n219 25.224
R8926 VDPWR.n219 VDPWR.n205 25.224
R8927 VDPWR.n215 VDPWR.n214 25.224
R8928 VDPWR.n214 VDPWR.n206 25.224
R8929 VDPWR.n210 VDPWR.n209 25.224
R8930 VDPWR.n209 VDPWR.n119 25.224
R8931 VDPWR.n183 VDPWR.n133 25.224
R8932 VDPWR.n179 VDPWR.n133 25.224
R8933 VDPWR.n188 VDPWR.n132 25.224
R8934 VDPWR.n184 VDPWR.n132 25.224
R8935 VDPWR.n193 VDPWR.n131 25.224
R8936 VDPWR.n189 VDPWR.n131 25.224
R8937 VDPWR.n198 VDPWR.n130 25.224
R8938 VDPWR.n194 VDPWR.n130 25.224
R8939 VDPWR.n200 VDPWR.n129 25.224
R8940 VDPWR.n200 VDPWR.n199 25.224
R8941 VDPWR.n159 VDPWR.n154 25.224
R8942 VDPWR.n155 VDPWR.n154 25.224
R8943 VDPWR.n164 VDPWR.n153 25.224
R8944 VDPWR.n160 VDPWR.n153 25.224
R8945 VDPWR.n169 VDPWR.n152 25.224
R8946 VDPWR.n165 VDPWR.n152 25.224
R8947 VDPWR.n171 VDPWR.n135 25.224
R8948 VDPWR.n171 VDPWR.n170 25.224
R8949 VDPWR.n72 VDPWR.n56 25.224
R8950 VDPWR.n68 VDPWR.n56 25.224
R8951 VDPWR.n77 VDPWR.n55 25.224
R8952 VDPWR.n73 VDPWR.n55 25.224
R8953 VDPWR.n79 VDPWR.n53 25.224
R8954 VDPWR.n79 VDPWR.n78 25.224
R8955 VDPWR.n97 VDPWR.n93 25.224
R8956 VDPWR.n2632 VDPWR.n2629 25.1912
R8957 VDPWR.n2430 VDPWR.n2349 25.1912
R8958 VDPWR.n2412 VDPWR.n2410 25.1912
R8959 VDPWR.n3080 VDPWR.n3079 25.1912
R8960 VDPWR.t986 VDPWR 25.1772
R8961 VDPWR VDPWR.t1150 25.1772
R8962 VDPWR.t388 VDPWR 25.1772
R8963 VDPWR.n725 VDPWR.n724 25.0224
R8964 VDPWR.n727 VDPWR.n726 25.0224
R8965 VDPWR.n723 VDPWR.n722 25.0224
R8966 VDPWR.n1107 VDPWR.n1106 24.0557
R8967 VDPWR.n2687 VDPWR.n2686 23.7181
R8968 VDPWR.n581 VDPWR.n564 23.7181
R8969 VDPWR.n640 VDPWR.n562 23.7181
R8970 VDPWR.n301 VDPWR.n284 23.7181
R8971 VDPWR.n360 VDPWR.n282 23.7181
R8972 VDPWR.n1498 VDPWR.n1297 23.7181
R8973 VDPWR.n1882 VDPWR.n1205 23.7181
R8974 VDPWR.n2738 VDPWR.n2735 23.7181
R8975 VDPWR.n2744 VDPWR.n2738 23.7181
R8976 VDPWR.n2902 VDPWR.n954 23.7181
R8977 VDPWR.n2633 VDPWR.n2632 23.7181
R8978 VDPWR.n2657 VDPWR.n2656 23.7181
R8979 VDPWR.n2567 VDPWR.n2565 23.7181
R8980 VDPWR.n2687 VDPWR.n2594 23.7181
R8981 VDPWR.n2530 VDPWR.n2433 23.7181
R8982 VDPWR.n2380 VDPWR.n2377 23.7181
R8983 VDPWR.n3097 VDPWR.n3096 23.7181
R8984 VDPWR.n43 VDPWR.n26 23.7181
R8985 VDPWR.n102 VDPWR.n24 23.7181
R8986 VDPWR.t1077 VDPWR.t589 23.4987
R8987 VDPWR.t991 VDPWR.t269 23.4987
R8988 VDPWR.t352 VDPWR.t300 23.4987
R8989 VDPWR.n808 VDPWR.n807 22.9652
R8990 VDPWR.n1990 VDPWR.n1988 22.9652
R8991 VDPWR.n2657 VDPWR.n2620 22.9652
R8992 VDPWR.n2649 VDPWR.n2613 22.9652
R8993 VDPWR.n2699 VDPWR.n2587 22.9652
R8994 VDPWR.n3023 VDPWR.n916 22.9652
R8995 VDPWR.n2817 VDPWR.n2814 22.6748
R8996 VDPWR.n2828 VDPWR.n981 22.5887
R8997 VDPWR.n2643 VDPWR.n2641 22.5887
R8998 VDPWR.n2637 VDPWR.n2621 22.5887
R8999 VDPWR.n2774 VDPWR.n1001 22.3091
R9000 VDPWR.n1982 VDPWR.n1980 22.2123
R9001 VDPWR.n1983 VDPWR.n1982 22.2123
R9002 VDPWR.n2824 VDPWR.n2821 22.2123
R9003 VDPWR.n2824 VDPWR.n981 22.2123
R9004 VDPWR.n2387 VDPWR.n2386 22.2123
R9005 VDPWR.n2381 VDPWR.n2369 22.2123
R9006 VDPWR.n2386 VDPWR.n2385 22.2123
R9007 VDPWR.n2381 VDPWR.n2380 22.2123
R9008 VDPWR.n2513 VDPWR.n2512 22.2123
R9009 VDPWR.n2668 VDPWR.n2613 21.8358
R9010 VDPWR.n2700 VDPWR.n2699 21.8358
R9011 VDPWR.n3024 VDPWR.n3023 21.8358
R9012 VDPWR.t360 VDPWR.t1124 21.8203
R9013 VDPWR.t1042 VDPWR.t1128 21.8203
R9014 VDPWR.n2812 VDPWR.t1104 21.8203
R9015 VDPWR.t231 VDPWR.t299 21.8203
R9016 VDPWR.n630 VDPWR.n564 21.4593
R9017 VDPWR.n350 VDPWR.n284 21.4593
R9018 VDPWR.n2656 VDPWR.n2649 21.4593
R9019 VDPWR.n2594 VDPWR.n2587 21.4593
R9020 VDPWR.n92 VDPWR.n26 21.4593
R9021 VDPWR.n2763 VDPWR.n1003 21.05
R9022 VDPWR.n2106 VDPWR.n2091 20.912
R9023 VDPWR.n2780 VDPWR.n1001 20.8462
R9024 VDPWR.n857 VDPWR.n856 20.4852
R9025 VDPWR.n2774 VDPWR.n2773 20.4805
R9026 VDPWR.n735 VDPWR.t252 20.3758
R9027 VDPWR.t341 VDPWR.n735 20.3758
R9028 VDPWR.n611 VDPWR.n610 20.3299
R9029 VDPWR.n616 VDPWR.n615 20.3299
R9030 VDPWR.n331 VDPWR.n330 20.3299
R9031 VDPWR.n336 VDPWR.n335 20.3299
R9032 VDPWR.n246 VDPWR.n245 20.3299
R9033 VDPWR.n240 VDPWR.n123 20.3299
R9034 VDPWR.n235 VDPWR.n124 20.3299
R9035 VDPWR.n230 VDPWR.n125 20.3299
R9036 VDPWR.n225 VDPWR.n126 20.3299
R9037 VDPWR.n220 VDPWR.n204 20.3299
R9038 VDPWR.n215 VDPWR.n205 20.3299
R9039 VDPWR.n210 VDPWR.n206 20.3299
R9040 VDPWR.n184 VDPWR.n183 20.3299
R9041 VDPWR.n189 VDPWR.n188 20.3299
R9042 VDPWR.n194 VDPWR.n193 20.3299
R9043 VDPWR.n199 VDPWR.n198 20.3299
R9044 VDPWR.n155 VDPWR.n129 20.3299
R9045 VDPWR.n160 VDPWR.n159 20.3299
R9046 VDPWR.n165 VDPWR.n164 20.3299
R9047 VDPWR.n170 VDPWR.n169 20.3299
R9048 VDPWR.n73 VDPWR.n72 20.3299
R9049 VDPWR.n78 VDPWR.n77 20.3299
R9050 VDPWR.t18 VDPWR.t184 20.1418
R9051 VDPWR.t989 VDPWR.t178 20.1418
R9052 VDPWR.t1114 VDPWR.t968 20.1418
R9053 VDPWR.t221 VDPWR.t81 20.1418
R9054 VDPWR.t196 VDPWR.t878 20.1418
R9055 VDPWR.n2782 VDPWR.n2780 20.1148
R9056 VDPWR.n2053 VDPWR.n1130 20.0749
R9057 VDPWR.n2463 VDPWR.n789 19.9534
R9058 VDPWR.n2742 VDPWR.n2741 19.9237
R9059 VDPWR.n650 VDPWR.n649 19.8181
R9060 VDPWR.n370 VDPWR.n369 19.8181
R9061 VDPWR.n112 VDPWR.n111 19.8181
R9062 VDPWR.n2784 VDPWR.n998 19.7491
R9063 VDPWR.n2790 VDPWR.n2789 19.7491
R9064 VDPWR.n646 VDPWR.n645 19.6946
R9065 VDPWR.n366 VDPWR.n365 19.6946
R9066 VDPWR.n108 VDPWR.n107 19.6946
R9067 VDPWR.n1966 VDPWR.n1922 19.577
R9068 VDPWR.n2315 VDPWR.n1026 19.2067
R9069 VDPWR.n2226 VDPWR.n2225 18.7808
R9070 VDPWR.n1829 VDPWR.n1827 18.7591
R9071 VDPWR.t1143 VDPWR.t377 18.4634
R9072 VDPWR.t322 VDPWR.t816 18.4634
R9073 VDPWR.n1918 VDPWR.n1186 18.4476
R9074 VDPWR.n2854 VDPWR.n2853 18.4476
R9075 VDPWR.n2676 VDPWR.n2675 18.4476
R9076 VDPWR.n2707 VDPWR.n2706 18.4476
R9077 VDPWR.n911 VDPWR.n900 18.4476
R9078 VDPWR.n3026 VDPWR.n3025 18.4476
R9079 VDPWR.n2821 VDPWR.n982 18.0711
R9080 VDPWR.n2405 VDPWR.n2404 18.0382
R9081 VDPWR.n1576 VDPWR.n1575 17.9678
R9082 VDPWR VDPWR.n2359 17.6841
R9083 VDPWR.n2184 VDPWR.n1103 17.612
R9084 VDPWR.n622 VDPWR.n591 17.3181
R9085 VDPWR.n634 VDPWR.n633 17.3181
R9086 VDPWR.n640 VDPWR.n539 17.3181
R9087 VDPWR.n342 VDPWR.n311 17.3181
R9088 VDPWR.n354 VDPWR.n353 17.3181
R9089 VDPWR.n360 VDPWR.n259 17.3181
R9090 VDPWR.n251 VDPWR.n119 17.3181
R9091 VDPWR.n175 VDPWR.n135 17.3181
R9092 VDPWR.n84 VDPWR.n53 17.3181
R9093 VDPWR.n96 VDPWR.n95 17.3181
R9094 VDPWR.n102 VDPWR.n1 17.3181
R9095 VDPWR.n606 VDPWR.n605 17.2853
R9096 VDPWR.n326 VDPWR.n325 17.2853
R9097 VDPWR.n68 VDPWR.n67 17.2853
R9098 VDPWR.n3052 VDPWR.n3051 16.9417
R9099 VDPWR.n2410 VDPWR.n2353 16.9417
R9100 VDPWR.t1130 VDPWR.t866 16.785
R9101 VDPWR.t438 VDPWR.t167 16.785
R9102 VDPWR.t480 VDPWR.t227 16.785
R9103 VDPWR.n1830 VDPWR.n1829 16.7729
R9104 VDPWR.n2173 VDPWR.n1108 16.7729
R9105 VDPWR.n1466 VDPWR.n1465 16.6847
R9106 VDPWR.n2939 VDPWR.n2938 16.5825
R9107 VDPWR.n631 VDPWR.n630 16.5652
R9108 VDPWR.n635 VDPWR.n634 16.5652
R9109 VDPWR.n351 VDPWR.n350 16.5652
R9110 VDPWR.n355 VDPWR.n354 16.5652
R9111 VDPWR.n93 VDPWR.n92 16.5652
R9112 VDPWR.n97 VDPWR.n96 16.5652
R9113 VDPWR.n2794 VDPWR.n2793 16.4576
R9114 VDPWR.n2670 VDPWR.n2669 16.1887
R9115 VDPWR.n2708 VDPWR.n2707 16.1887
R9116 VDPWR.n3039 VDPWR.n900 16.1887
R9117 VDPWR.n3027 VDPWR.n3026 16.1887
R9118 VDPWR.n250 VDPWR.n120 15.8123
R9119 VDPWR.n179 VDPWR.n178 15.8123
R9120 VDPWR.n732 VDPWR.n730 15.4172
R9121 VDPWR.n735 VDPWR.n732 15.4172
R9122 VDPWR.n731 VDPWR.n729 15.4172
R9123 VDPWR.n735 VDPWR.n731 15.4172
R9124 VDPWR.n2795 VDPWR.n2794 15.3605
R9125 VDPWR.n1107 VDPWR.n1105 15.2281
R9126 VDPWR.n1827 VDPWR.n1222 15.101
R9127 VDPWR.n2861 VDPWR.n965 15.0593
R9128 VDPWR.n2714 VDPWR.n2713 15.0593
R9129 VDPWR.n3045 VDPWR.n3044 15.0593
R9130 VDPWR.n3040 VDPWR.n3039 15.0593
R9131 VDPWR.n2406 VDPWR.n2353 15.0593
R9132 VDPWR.n2514 VDPWR.n2513 15.0593
R9133 VDPWR.n1435 VDPWR.n1434 14.9
R9134 VDPWR.n3097 VDPWR.n789 14.6829
R9135 VDPWR.n1994 VDPWR.n1182 14.6484
R9136 VDPWR.n644 VDPWR.n560 14.6078
R9137 VDPWR.n364 VDPWR.n280 14.6078
R9138 VDPWR.n106 VDPWR.n22 14.6078
R9139 VDPWR.n1481 VDPWR.n1297 14.5851
R9140 VDPWR.n1549 VDPWR.n1537 14.5851
R9141 VDPWR.n2853 VDPWR.n2852 14.3064
R9142 VDPWR.n2643 VDPWR.n2620 14.3064
R9143 VDPWR.n3019 VDPWR.n916 14.3064
R9144 VDPWR.n623 VDPWR.n622 14.2735
R9145 VDPWR.n582 VDPWR.n581 14.2735
R9146 VDPWR.n343 VDPWR.n342 14.2735
R9147 VDPWR.n302 VDPWR.n301 14.2735
R9148 VDPWR.n1948 VDPWR.n1936 14.2735
R9149 VDPWR.n2888 VDPWR.n954 14.2735
R9150 VDPWR.n3053 VDPWR.n885 14.2735
R9151 VDPWR.n3000 VDPWR.n2988 14.2735
R9152 VDPWR.n2526 VDPWR.n2433 14.2735
R9153 VDPWR.n3096 VDPWR.n3095 14.2735
R9154 VDPWR.n843 VDPWR.n831 14.2735
R9155 VDPWR.n85 VDPWR.n84 14.2735
R9156 VDPWR.n44 VDPWR.n43 14.2735
R9157 VDPWR.n1919 VDPWR.n1918 13.9299
R9158 VDPWR.n2264 VDPWR.n1075 13.8955
R9159 VDPWR.n2973 VDPWR.n929 13.8955
R9160 VDPWR.n651 VDPWR.n650 13.5534
R9161 VDPWR.n371 VDPWR.n370 13.5534
R9162 VDPWR.n113 VDPWR.n112 13.5534
R9163 VDPWR VDPWR.n571 13.4732
R9164 VDPWR VDPWR.n291 13.4732
R9165 VDPWR VDPWR.n33 13.4732
R9166 VDPWR.t984 VDPWR.t366 13.4281
R9167 VDPWR.t22 VDPWR.t501 13.4281
R9168 VDPWR.t358 VDPWR.t100 13.4281
R9169 VDPWR.t1049 VDPWR.t295 13.4281
R9170 VDPWR VDPWR.t1146 13.4281
R9171 VDPWR.n2767 VDPWR.n1003 12.9181
R9172 VDPWR.n175 VDPWR.n136 12.8005
R9173 VDPWR.n148 VDPWR.n136 12.8005
R9174 VDPWR.n148 VDPWR.n145 12.8005
R9175 VDPWR.n145 VDPWR.n144 12.8005
R9176 VDPWR.n1366 VDPWR.n1357 12.8005
R9177 VDPWR.n1699 VDPWR.n1690 12.8005
R9178 VDPWR.n1896 VDPWR.n1205 12.8005
R9179 VDPWR.n1621 VDPWR.n1620 12.8005
R9180 VDPWR.n2102 VDPWR.n2095 12.8005
R9181 VDPWR.n2565 VDPWR.n2556 12.8005
R9182 VDPWR.n3053 VDPWR.n3052 12.8005
R9183 VDPWR.n2837 VDPWR.n2836 12.3976
R9184 VDPWR.n3019 VDPWR.n3018 12.3912
R9185 VDPWR.n651 VDPWR.n539 12.0476
R9186 VDPWR.n371 VDPWR.n259 12.0476
R9187 VDPWR.n113 VDPWR.n1 12.0476
R9188 VDPWR.t16 VDPWR.t781 11.7496
R9189 VDPWR.t890 VDPWR.t250 11.7496
R9190 VDPWR.n814 VDPWR.n812 11.6993
R9191 VDPWR.n807 VDPWR.n800 11.6711
R9192 VDPWR.n587 VDPWR.n586 11.4366
R9193 VDPWR.n307 VDPWR.n306 11.4366
R9194 VDPWR.n49 VDPWR.n48 11.4366
R9195 VDPWR VDPWR.n535 11.4331
R9196 VDPWR VDPWR.n3175 11.4331
R9197 VDPWR.n389 VDPWR.n388 11.3235
R9198 VDPWR.n401 VDPWR.n400 11.3235
R9199 VDPWR.n2830 VDPWR.n2828 11.2946
R9200 VDPWR.n2669 VDPWR.n2668 11.2946
R9201 VDPWR.n643 VDPWR.n561 11.2937
R9202 VDPWR.n363 VDPWR.n281 11.2937
R9203 VDPWR.n105 VDPWR.n23 11.2937
R9204 VDPWR.n628 VDPWR.n627 11.2737
R9205 VDPWR.n348 VDPWR.n347 11.2737
R9206 VDPWR.n90 VDPWR.n89 11.2737
R9207 VDPWR.n2814 VDPWR.n2813 10.9719
R9208 VDPWR.n141 VDPWR.n140 10.9345
R9209 VDPWR.n2861 VDPWR.n2860 10.9181
R9210 VDPWR.n2052 VDPWR.n2051 10.912
R9211 VDPWR.n2744 VDPWR.n2743 10.5744
R9212 VDPWR.n2406 VDPWR.n2405 10.5417
R9213 VDPWR.n560 VDPWR.n559 10.1786
R9214 VDPWR.n280 VDPWR.n279 10.1786
R9215 VDPWR.n22 VDPWR.n21 10.1786
R9216 VDPWR.n2834 VDPWR.n980 10.1652
R9217 VDPWR.t979 VDPWR.t855 10.0712
R9218 VDPWR.t1010 VDPWR.t235 10.0712
R9219 VDPWR.t605 VDPWR.t759 10.0712
R9220 VDPWR.t208 VDPWR.t130 10.0712
R9221 VDPWR.n2107 VDPWR.n2106 9.8812
R9222 VDPWR.n2830 VDPWR.n980 9.78874
R9223 VDPWR.n2637 VDPWR.n2635 9.78874
R9224 VDPWR.n1519 VDPWR.n1518 9.73273
R9225 VDPWR.n1762 VDPWR.n1760 9.73273
R9226 VDPWR.n1840 VDPWR.n1839 9.73273
R9227 VDPWR.n1842 VDPWR.n1218 9.73273
R9228 VDPWR.n1846 VDPWR.n1218 9.73273
R9229 VDPWR.n1850 VDPWR.n1846 9.73273
R9230 VDPWR.n1850 VDPWR.n1849 9.73273
R9231 VDPWR.n2171 VDPWR.n1110 9.73273
R9232 VDPWR.n2216 VDPWR.n2215 9.73273
R9233 VDPWR.n2309 VDPWR.n2308 9.73273
R9234 VDPWR.n2908 VDPWR.n2907 9.73273
R9235 VDPWR.n2914 VDPWR.n2913 9.73273
R9236 VDPWR.n2917 VDPWR.n2914 9.73273
R9237 VDPWR.n2921 VDPWR.n948 9.73273
R9238 VDPWR.n2922 VDPWR.n2921 9.73273
R9239 VDPWR.n2923 VDPWR.n2922 9.73273
R9240 VDPWR.n2947 VDPWR.n2944 9.73273
R9241 VDPWR.n2951 VDPWR.n935 9.73273
R9242 VDPWR.n2480 VDPWR.n2479 9.73273
R9243 VDPWR.n2479 VDPWR.n2478 9.73273
R9244 VDPWR.n2220 VDPWR.n2219 9.71972
R9245 VDPWR.n2275 VDPWR.n2274 9.71972
R9246 VDPWR.n2173 VDPWR.n2172 9.71084
R9247 VDPWR.n2188 VDPWR.n2187 9.65296
R9248 VDPWR.n2243 VDPWR.n2242 9.65296
R9249 VDPWR.n2233 VDPWR.n2232 9.65296
R9250 VDPWR.n2230 VDPWR.n2200 9.65296
R9251 VDPWR.n2305 VDPWR.n2304 9.65296
R9252 VDPWR.n2302 VDPWR.n1036 9.65296
R9253 VDPWR.n2298 VDPWR.n2297 9.65296
R9254 VDPWR.n2281 VDPWR.n1059 9.65296
R9255 VDPWR.n600 VDPWR.n599 9.60526
R9256 VDPWR.n588 VDPWR.n587 9.60526
R9257 VDPWR.n553 VDPWR.n552 9.60526
R9258 VDPWR.n320 VDPWR.n319 9.60526
R9259 VDPWR.n308 VDPWR.n307 9.60526
R9260 VDPWR.n273 VDPWR.n272 9.60526
R9261 VDPWR.n62 VDPWR.n61 9.60526
R9262 VDPWR.n50 VDPWR.n49 9.60526
R9263 VDPWR.n15 VDPWR.n14 9.60526
R9264 VDPWR.n2742 VDPWR.n2739 9.6005
R9265 VDPWR.n2782 VDPWR.n999 9.56172
R9266 VDPWR.n2944 VDPWR.n937 9.52116
R9267 VDPWR.n1830 VDPWR.n1826 9.49016
R9268 VDPWR.n2285 VDPWR.n1057 9.35121
R9269 VDPWR.n250 VDPWR 9.30627
R9270 VDPWR.n590 VDPWR.n566 9.3005
R9271 VDPWR.n626 VDPWR.n625 9.3005
R9272 VDPWR.n623 VDPWR.n567 9.3005
R9273 VDPWR.n622 VDPWR.n620 9.3005
R9274 VDPWR.n619 VDPWR.n591 9.3005
R9275 VDPWR.n618 VDPWR.n617 9.3005
R9276 VDPWR.n616 VDPWR.n592 9.3005
R9277 VDPWR.n615 VDPWR.n614 9.3005
R9278 VDPWR.n613 VDPWR.n593 9.3005
R9279 VDPWR.n612 VDPWR.n611 9.3005
R9280 VDPWR.n610 VDPWR.n609 9.3005
R9281 VDPWR.n608 VDPWR.n594 9.3005
R9282 VDPWR.n607 VDPWR.n606 9.3005
R9283 VDPWR.n605 VDPWR.n604 9.3005
R9284 VDPWR.n603 VDPWR.n602 9.3005
R9285 VDPWR.n601 VDPWR.n597 9.3005
R9286 VDPWR.n573 VDPWR.n572 9.3005
R9287 VDPWR.n576 VDPWR.n568 9.3005
R9288 VDPWR.n585 VDPWR.n584 9.3005
R9289 VDPWR.n582 VDPWR.n569 9.3005
R9290 VDPWR.n581 VDPWR.n580 9.3005
R9291 VDPWR.n579 VDPWR.n564 9.3005
R9292 VDPWR.n630 VDPWR.n629 9.3005
R9293 VDPWR.n631 VDPWR.n563 9.3005
R9294 VDPWR.n636 VDPWR.n635 9.3005
R9295 VDPWR.n637 VDPWR.n562 9.3005
R9296 VDPWR.n640 VDPWR.n639 9.3005
R9297 VDPWR.n638 VDPWR.n539 9.3005
R9298 VDPWR.n652 VDPWR.n651 9.3005
R9299 VDPWR.n650 VDPWR.n538 9.3005
R9300 VDPWR.n649 VDPWR.n648 9.3005
R9301 VDPWR.n647 VDPWR.n646 9.3005
R9302 VDPWR.n645 VDPWR.n542 9.3005
R9303 VDPWR.n644 VDPWR.n547 9.3005
R9304 VDPWR.n559 VDPWR.n558 9.3005
R9305 VDPWR.n557 VDPWR.n556 9.3005
R9306 VDPWR.n554 VDPWR.n549 9.3005
R9307 VDPWR.n310 VDPWR.n286 9.3005
R9308 VDPWR.n346 VDPWR.n345 9.3005
R9309 VDPWR.n343 VDPWR.n287 9.3005
R9310 VDPWR.n342 VDPWR.n340 9.3005
R9311 VDPWR.n339 VDPWR.n311 9.3005
R9312 VDPWR.n338 VDPWR.n337 9.3005
R9313 VDPWR.n336 VDPWR.n312 9.3005
R9314 VDPWR.n335 VDPWR.n334 9.3005
R9315 VDPWR.n333 VDPWR.n313 9.3005
R9316 VDPWR.n332 VDPWR.n331 9.3005
R9317 VDPWR.n330 VDPWR.n329 9.3005
R9318 VDPWR.n328 VDPWR.n314 9.3005
R9319 VDPWR.n327 VDPWR.n326 9.3005
R9320 VDPWR.n325 VDPWR.n324 9.3005
R9321 VDPWR.n323 VDPWR.n322 9.3005
R9322 VDPWR.n321 VDPWR.n317 9.3005
R9323 VDPWR.n293 VDPWR.n292 9.3005
R9324 VDPWR.n296 VDPWR.n288 9.3005
R9325 VDPWR.n305 VDPWR.n304 9.3005
R9326 VDPWR.n302 VDPWR.n289 9.3005
R9327 VDPWR.n301 VDPWR.n300 9.3005
R9328 VDPWR.n299 VDPWR.n284 9.3005
R9329 VDPWR.n350 VDPWR.n349 9.3005
R9330 VDPWR.n351 VDPWR.n283 9.3005
R9331 VDPWR.n356 VDPWR.n355 9.3005
R9332 VDPWR.n357 VDPWR.n282 9.3005
R9333 VDPWR.n360 VDPWR.n359 9.3005
R9334 VDPWR.n358 VDPWR.n259 9.3005
R9335 VDPWR.n372 VDPWR.n371 9.3005
R9336 VDPWR.n370 VDPWR.n258 9.3005
R9337 VDPWR.n369 VDPWR.n368 9.3005
R9338 VDPWR.n367 VDPWR.n366 9.3005
R9339 VDPWR.n365 VDPWR.n262 9.3005
R9340 VDPWR.n364 VDPWR.n267 9.3005
R9341 VDPWR.n279 VDPWR.n278 9.3005
R9342 VDPWR.n277 VDPWR.n276 9.3005
R9343 VDPWR.n274 VDPWR.n269 9.3005
R9344 VDPWR.n143 VDPWR.n142 9.3005
R9345 VDPWR.n144 VDPWR.n138 9.3005
R9346 VDPWR.n145 VDPWR.n137 9.3005
R9347 VDPWR.n149 VDPWR.n148 9.3005
R9348 VDPWR.n150 VDPWR.n136 9.3005
R9349 VDPWR.n175 VDPWR.n174 9.3005
R9350 VDPWR.n173 VDPWR.n135 9.3005
R9351 VDPWR.n172 VDPWR.n171 9.3005
R9352 VDPWR.n170 VDPWR.n151 9.3005
R9353 VDPWR.n169 VDPWR.n168 9.3005
R9354 VDPWR.n167 VDPWR.n152 9.3005
R9355 VDPWR.n166 VDPWR.n165 9.3005
R9356 VDPWR.n164 VDPWR.n163 9.3005
R9357 VDPWR.n162 VDPWR.n153 9.3005
R9358 VDPWR.n161 VDPWR.n160 9.3005
R9359 VDPWR.n159 VDPWR.n158 9.3005
R9360 VDPWR.n157 VDPWR.n154 9.3005
R9361 VDPWR.n156 VDPWR.n155 9.3005
R9362 VDPWR.n129 VDPWR.n127 9.3005
R9363 VDPWR.n201 VDPWR.n200 9.3005
R9364 VDPWR.n199 VDPWR.n128 9.3005
R9365 VDPWR.n198 VDPWR.n197 9.3005
R9366 VDPWR.n196 VDPWR.n130 9.3005
R9367 VDPWR.n195 VDPWR.n194 9.3005
R9368 VDPWR.n193 VDPWR.n192 9.3005
R9369 VDPWR.n191 VDPWR.n131 9.3005
R9370 VDPWR.n190 VDPWR.n189 9.3005
R9371 VDPWR.n188 VDPWR.n187 9.3005
R9372 VDPWR.n186 VDPWR.n132 9.3005
R9373 VDPWR.n185 VDPWR.n184 9.3005
R9374 VDPWR.n183 VDPWR.n182 9.3005
R9375 VDPWR.n181 VDPWR.n133 9.3005
R9376 VDPWR.n180 VDPWR.n179 9.3005
R9377 VDPWR.n178 VDPWR.n177 9.3005
R9378 VDPWR.n252 VDPWR.n251 9.3005
R9379 VDPWR.n249 VDPWR.n120 9.3005
R9380 VDPWR.n248 VDPWR.n247 9.3005
R9381 VDPWR.n246 VDPWR.n121 9.3005
R9382 VDPWR.n245 VDPWR.n122 9.3005
R9383 VDPWR.n244 VDPWR.n243 9.3005
R9384 VDPWR.n242 VDPWR.n123 9.3005
R9385 VDPWR.n241 VDPWR.n240 9.3005
R9386 VDPWR.n239 VDPWR.n238 9.3005
R9387 VDPWR.n237 VDPWR.n124 9.3005
R9388 VDPWR.n236 VDPWR.n235 9.3005
R9389 VDPWR.n234 VDPWR.n233 9.3005
R9390 VDPWR.n232 VDPWR.n125 9.3005
R9391 VDPWR.n231 VDPWR.n230 9.3005
R9392 VDPWR.n229 VDPWR.n228 9.3005
R9393 VDPWR.n227 VDPWR.n126 9.3005
R9394 VDPWR.n226 VDPWR.n225 9.3005
R9395 VDPWR.n224 VDPWR.n223 9.3005
R9396 VDPWR.n222 VDPWR.n204 9.3005
R9397 VDPWR.n221 VDPWR.n220 9.3005
R9398 VDPWR.n219 VDPWR.n218 9.3005
R9399 VDPWR.n217 VDPWR.n205 9.3005
R9400 VDPWR.n216 VDPWR.n215 9.3005
R9401 VDPWR.n214 VDPWR.n213 9.3005
R9402 VDPWR.n212 VDPWR.n206 9.3005
R9403 VDPWR.n211 VDPWR.n210 9.3005
R9404 VDPWR.n209 VDPWR.n208 9.3005
R9405 VDPWR.n207 VDPWR.n119 9.3005
R9406 VDPWR.n1549 VDPWR.n1548 9.3005
R9407 VDPWR.n1550 VDPWR.n1549 9.3005
R9408 VDPWR.n1549 VDPWR.n1535 9.3005
R9409 VDPWR.n1369 VDPWR.n1368 9.3005
R9410 VDPWR.n1376 VDPWR.n1375 9.3005
R9411 VDPWR.n1378 VDPWR.n1348 9.3005
R9412 VDPWR.n1380 VDPWR.n1379 9.3005
R9413 VDPWR.n1389 VDPWR.n1388 9.3005
R9414 VDPWR.n1390 VDPWR.n1342 9.3005
R9415 VDPWR.n1393 VDPWR.n1392 9.3005
R9416 VDPWR.n1394 VDPWR.n1341 9.3005
R9417 VDPWR.n1396 VDPWR.n1395 9.3005
R9418 VDPWR.n1398 VDPWR.n1340 9.3005
R9419 VDPWR.n1400 VDPWR.n1399 9.3005
R9420 VDPWR.n1402 VDPWR.n1401 9.3005
R9421 VDPWR.n1404 VDPWR.n1338 9.3005
R9422 VDPWR.n1407 VDPWR.n1406 9.3005
R9423 VDPWR.n1408 VDPWR.n1337 9.3005
R9424 VDPWR.n1410 VDPWR.n1409 9.3005
R9425 VDPWR.n1412 VDPWR.n1335 9.3005
R9426 VDPWR.n1415 VDPWR.n1414 9.3005
R9427 VDPWR.n1413 VDPWR.n1329 9.3005
R9428 VDPWR.n1428 VDPWR.n1427 9.3005
R9429 VDPWR.n1432 VDPWR.n1431 9.3005
R9430 VDPWR.n1436 VDPWR.n1435 9.3005
R9431 VDPWR.n1438 VDPWR.n1437 9.3005
R9432 VDPWR.n1439 VDPWR.n1322 9.3005
R9433 VDPWR.n1442 VDPWR.n1441 9.3005
R9434 VDPWR.n1443 VDPWR.n1321 9.3005
R9435 VDPWR.n1445 VDPWR.n1444 9.3005
R9436 VDPWR.n1447 VDPWR.n1446 9.3005
R9437 VDPWR.n1451 VDPWR.n1314 9.3005
R9438 VDPWR.n1461 VDPWR.n1460 9.3005
R9439 VDPWR.n1462 VDPWR.n1313 9.3005
R9440 VDPWR.n1464 VDPWR.n1463 9.3005
R9441 VDPWR.n1465 VDPWR 9.3005
R9442 VDPWR.n1467 VDPWR.n1466 9.3005
R9443 VDPWR.n1469 VDPWR.n1468 9.3005
R9444 VDPWR.n1470 VDPWR.n1310 9.3005
R9445 VDPWR.n1472 VDPWR.n1471 9.3005
R9446 VDPWR.n1474 VDPWR.n1473 9.3005
R9447 VDPWR.n1475 VDPWR.n1308 9.3005
R9448 VDPWR.n1477 VDPWR.n1476 9.3005
R9449 VDPWR.n1478 VDPWR.n1307 9.3005
R9450 VDPWR.n1480 VDPWR.n1479 9.3005
R9451 VDPWR.n1487 VDPWR.n1486 9.3005
R9452 VDPWR.n1485 VDPWR.n1484 9.3005
R9453 VDPWR.n1481 VDPWR.n1298 9.3005
R9454 VDPWR.n1496 VDPWR.n1297 9.3005
R9455 VDPWR.n1498 VDPWR.n1497 9.3005
R9456 VDPWR.n1500 VDPWR.n1499 9.3005
R9457 VDPWR.n1502 VDPWR.n1501 9.3005
R9458 VDPWR.n1504 VDPWR.n1295 9.3005
R9459 VDPWR.n1508 VDPWR.n1507 9.3005
R9460 VDPWR.n1509 VDPWR.n1294 9.3005
R9461 VDPWR.n1511 VDPWR.n1510 9.3005
R9462 VDPWR.n1512 VDPWR.n1293 9.3005
R9463 VDPWR.n1514 VDPWR.n1513 9.3005
R9464 VDPWR.n1516 VDPWR.n1515 9.3005
R9465 VDPWR.n1518 VDPWR.n1517 9.3005
R9466 VDPWR.n1519 VDPWR.n1289 9.3005
R9467 VDPWR.n1577 VDPWR.n1576 9.3005
R9468 VDPWR.n1575 VDPWR.n1574 9.3005
R9469 VDPWR.n1573 VDPWR.n1572 9.3005
R9470 VDPWR.n1571 VDPWR.n1523 9.3005
R9471 VDPWR.n1570 VDPWR.n1569 9.3005
R9472 VDPWR.n1568 VDPWR.n1567 9.3005
R9473 VDPWR.n1566 VDPWR.n1525 9.3005
R9474 VDPWR.n1565 VDPWR.n1564 9.3005
R9475 VDPWR.n1563 VDPWR.n1526 9.3005
R9476 VDPWR.n1562 VDPWR.n1561 9.3005
R9477 VDPWR.n1560 VDPWR.n1527 9.3005
R9478 VDPWR.n1559 VDPWR.n1558 9.3005
R9479 VDPWR.n1537 VDPWR.n1529 9.3005
R9480 VDPWR.n1897 VDPWR.n1896 9.3005
R9481 VDPWR.n1896 VDPWR.n1198 9.3005
R9482 VDPWR.n1896 VDPWR.n1892 9.3005
R9483 VDPWR.n1702 VDPWR.n1701 9.3005
R9484 VDPWR.n1704 VDPWR.n1703 9.3005
R9485 VDPWR.n1709 VDPWR.n1708 9.3005
R9486 VDPWR.n1707 VDPWR.n1706 9.3005
R9487 VDPWR.n1719 VDPWR.n1718 9.3005
R9488 VDPWR.n1720 VDPWR.n1278 9.3005
R9489 VDPWR.n1723 VDPWR.n1722 9.3005
R9490 VDPWR.n1724 VDPWR.n1277 9.3005
R9491 VDPWR.n1726 VDPWR.n1725 9.3005
R9492 VDPWR.n1728 VDPWR.n1276 9.3005
R9493 VDPWR.n1730 VDPWR.n1729 9.3005
R9494 VDPWR.n1732 VDPWR.n1731 9.3005
R9495 VDPWR.n1734 VDPWR.n1274 9.3005
R9496 VDPWR.n1737 VDPWR.n1736 9.3005
R9497 VDPWR.n1738 VDPWR.n1273 9.3005
R9498 VDPWR.n1740 VDPWR.n1739 9.3005
R9499 VDPWR.n1742 VDPWR.n1271 9.3005
R9500 VDPWR.n1746 VDPWR.n1745 9.3005
R9501 VDPWR.n1744 VDPWR.n1264 9.3005
R9502 VDPWR.n1758 VDPWR.n1263 9.3005
R9503 VDPWR.n1760 VDPWR.n1759 9.3005
R9504 VDPWR.n1763 VDPWR.n1762 9.3005
R9505 VDPWR.n1768 VDPWR.n1256 9.3005
R9506 VDPWR.n1772 VDPWR.n1771 9.3005
R9507 VDPWR.n1773 VDPWR.n1255 9.3005
R9508 VDPWR.n1775 VDPWR.n1774 9.3005
R9509 VDPWR.n1777 VDPWR.n1250 9.3005
R9510 VDPWR.n1779 VDPWR.n1778 9.3005
R9511 VDPWR.n1242 VDPWR.n1241 9.3005
R9512 VDPWR.n1789 VDPWR.n1788 9.3005
R9513 VDPWR.n1790 VDPWR.n1240 9.3005
R9514 VDPWR.n1793 VDPWR.n1792 9.3005
R9515 VDPWR.n1797 VDPWR.n1238 9.3005
R9516 VDPWR.n1800 VDPWR.n1799 9.3005
R9517 VDPWR.n1802 VDPWR.n1801 9.3005
R9518 VDPWR.n1803 VDPWR.n1236 9.3005
R9519 VDPWR.n1806 VDPWR.n1805 9.3005
R9520 VDPWR.n1807 VDPWR.n1235 9.3005
R9521 VDPWR.n1809 VDPWR.n1808 9.3005
R9522 VDPWR.n1815 VDPWR.n1814 9.3005
R9523 VDPWR.n1813 VDPWR.n1812 9.3005
R9524 VDPWR.n1225 VDPWR.n1224 9.3005
R9525 VDPWR.n1825 VDPWR.n1824 9.3005
R9526 VDPWR.n1831 VDPWR.n1830 9.3005
R9527 VDPWR.n1837 VDPWR.n1836 9.3005
R9528 VDPWR.n1839 VDPWR.n1838 9.3005
R9529 VDPWR.n1840 VDPWR.n1219 9.3005
R9530 VDPWR.n1843 VDPWR.n1842 9.3005
R9531 VDPWR.n1844 VDPWR.n1218 9.3005
R9532 VDPWR.n1846 VDPWR.n1845 9.3005
R9533 VDPWR.n1851 VDPWR.n1850 9.3005
R9534 VDPWR.n1849 VDPWR.n1214 9.3005
R9535 VDPWR.n1865 VDPWR.n1864 9.3005
R9536 VDPWR.n1867 VDPWR.n1866 9.3005
R9537 VDPWR.n1868 VDPWR.n1211 9.3005
R9538 VDPWR.n1870 VDPWR.n1869 9.3005
R9539 VDPWR.n1872 VDPWR.n1210 9.3005
R9540 VDPWR.n1878 VDPWR.n1877 9.3005
R9541 VDPWR.n1879 VDPWR.n1209 9.3005
R9542 VDPWR.n1881 VDPWR.n1880 9.3005
R9543 VDPWR.n1883 VDPWR.n1882 9.3005
R9544 VDPWR.n1885 VDPWR.n1205 9.3005
R9545 VDPWR.n1948 VDPWR.n1947 9.3005
R9546 VDPWR.n1949 VDPWR.n1948 9.3005
R9547 VDPWR.n1948 VDPWR.n1934 9.3005
R9548 VDPWR.n1608 VDPWR.n1603 9.3005
R9549 VDPWR.n1607 VDPWR.n1601 9.3005
R9550 VDPWR.n1667 VDPWR.n1666 9.3005
R9551 VDPWR.n1665 VDPWR.n1664 9.3005
R9552 VDPWR.n1656 VDPWR.n1655 9.3005
R9553 VDPWR.n1654 VDPWR.n1626 9.3005
R9554 VDPWR.n1653 VDPWR.n1652 9.3005
R9555 VDPWR.n1651 VDPWR.n1650 9.3005
R9556 VDPWR.n1649 VDPWR.n1648 9.3005
R9557 VDPWR.n1647 VDPWR.n1646 9.3005
R9558 VDPWR.n1645 VDPWR.n1629 9.3005
R9559 VDPWR.n1643 VDPWR.n1642 9.3005
R9560 VDPWR.n1641 VDPWR.n1640 9.3005
R9561 VDPWR.n1638 VDPWR.n1631 9.3005
R9562 VDPWR.n1637 VDPWR.n1636 9.3005
R9563 VDPWR.n1635 VDPWR.n1634 9.3005
R9564 VDPWR.n1632 VDPWR.n1121 9.3005
R9565 VDPWR.n1125 VDPWR.n1122 9.3005
R9566 VDPWR.n2061 VDPWR.n2060 9.3005
R9567 VDPWR.n2058 VDPWR.n2057 9.3005
R9568 VDPWR.n2056 VDPWR.n1126 9.3005
R9569 VDPWR.n2054 VDPWR.n2053 9.3005
R9570 VDPWR.n2046 VDPWR.n1129 9.3005
R9571 VDPWR.n2045 VDPWR.n2044 9.3005
R9572 VDPWR.n2043 VDPWR.n1131 9.3005
R9573 VDPWR.n2042 VDPWR.n2041 9.3005
R9574 VDPWR.n2040 VDPWR.n2039 9.3005
R9575 VDPWR.n1142 VDPWR.n1135 9.3005
R9576 VDPWR.n1148 VDPWR.n1147 9.3005
R9577 VDPWR.n1149 VDPWR.n1140 9.3005
R9578 VDPWR.n2030 VDPWR.n2029 9.3005
R9579 VDPWR.n2028 VDPWR.n1141 9.3005
R9580 VDPWR.n2026 VDPWR.n2025 9.3005
R9581 VDPWR.n2024 VDPWR.n1151 9.3005
R9582 VDPWR.n2023 VDPWR.n2022 9.3005
R9583 VDPWR.n2021 VDPWR.n1152 9.3005
R9584 VDPWR.n2020 VDPWR.n2019 9.3005
R9585 VDPWR.n2018 VDPWR.n2017 9.3005
R9586 VDPWR.n2016 VDPWR.n2015 9.3005
R9587 VDPWR.n2014 VDPWR.n2013 9.3005
R9588 VDPWR.n2012 VDPWR.n1157 9.3005
R9589 VDPWR.n2011 VDPWR.n2010 9.3005
R9590 VDPWR.n1169 VDPWR.n1168 9.3005
R9591 VDPWR.n1176 VDPWR.n1175 9.3005
R9592 VDPWR.n1178 VDPWR.n1165 9.3005
R9593 VDPWR.n2002 VDPWR.n2001 9.3005
R9594 VDPWR.n2000 VDPWR.n1999 9.3005
R9595 VDPWR.n1998 VDPWR.n1997 9.3005
R9596 VDPWR.n1996 VDPWR.n1180 9.3005
R9597 VDPWR.n1994 VDPWR.n1993 9.3005
R9598 VDPWR.n1992 VDPWR.n1182 9.3005
R9599 VDPWR.n1991 VDPWR.n1990 9.3005
R9600 VDPWR.n1988 VDPWR.n1183 9.3005
R9601 VDPWR.n1986 VDPWR.n1985 9.3005
R9602 VDPWR.n1984 VDPWR.n1983 9.3005
R9603 VDPWR.n1982 VDPWR.n1185 9.3005
R9604 VDPWR.n1980 VDPWR 9.3005
R9605 VDPWR.n1912 VDPWR.n1186 9.3005
R9606 VDPWR.n1920 VDPWR.n1914 9.3005
R9607 VDPWR.n1970 VDPWR.n1969 9.3005
R9608 VDPWR.n1966 VDPWR.n1965 9.3005
R9609 VDPWR.n1963 VDPWR.n1922 9.3005
R9610 VDPWR.n1962 VDPWR.n1961 9.3005
R9611 VDPWR.n1959 VDPWR.n1923 9.3005
R9612 VDPWR.n1958 VDPWR.n1957 9.3005
R9613 VDPWR.n1936 VDPWR.n1929 9.3005
R9614 VDPWR.n1086 VDPWR.n1075 9.3005
R9615 VDPWR.n1084 VDPWR.n1075 9.3005
R9616 VDPWR.n1077 VDPWR.n1075 9.3005
R9617 VDPWR.n2106 VDPWR.n2105 9.3005
R9618 VDPWR.n2109 VDPWR.n2108 9.3005
R9619 VDPWR.n2115 VDPWR.n2114 9.3005
R9620 VDPWR.n2119 VDPWR.n2118 9.3005
R9621 VDPWR.n2120 VDPWR.n2084 9.3005
R9622 VDPWR.n2129 VDPWR.n2128 9.3005
R9623 VDPWR.n2130 VDPWR.n2083 9.3005
R9624 VDPWR.n2132 VDPWR.n2131 9.3005
R9625 VDPWR.n2134 VDPWR.n2133 9.3005
R9626 VDPWR.n2135 VDPWR.n2081 9.3005
R9627 VDPWR.n2138 VDPWR.n2137 9.3005
R9628 VDPWR.n2140 VDPWR.n2139 9.3005
R9629 VDPWR.n2143 VDPWR.n2142 9.3005
R9630 VDPWR.n2145 VDPWR.n2144 9.3005
R9631 VDPWR.n2146 VDPWR.n2078 9.3005
R9632 VDPWR.n2148 VDPWR.n2147 9.3005
R9633 VDPWR.n2150 VDPWR.n2149 9.3005
R9634 VDPWR.n2152 VDPWR.n2151 9.3005
R9635 VDPWR.n1113 VDPWR.n1112 9.3005
R9636 VDPWR.n2165 VDPWR.n2164 9.3005
R9637 VDPWR.n2168 VDPWR.n2167 9.3005
R9638 VDPWR.n2169 VDPWR.n1110 9.3005
R9639 VDPWR.n2171 VDPWR.n2170 9.3005
R9640 VDPWR.n2174 VDPWR.n2173 9.3005
R9641 VDPWR.n2176 VDPWR.n2175 9.3005
R9642 VDPWR.n2181 VDPWR.n2180 9.3005
R9643 VDPWR.n2182 VDPWR.n1103 9.3005
R9644 VDPWR.n2184 VDPWR.n2183 9.3005
R9645 VDPWR.n2187 VDPWR.n1101 9.3005
R9646 VDPWR.n2189 VDPWR.n2188 9.3005
R9647 VDPWR.n2191 VDPWR.n2190 9.3005
R9648 VDPWR.n2193 VDPWR.n1096 9.3005
R9649 VDPWR.n2244 VDPWR.n2243 9.3005
R9650 VDPWR.n2242 VDPWR.n2241 9.3005
R9651 VDPWR.n2234 VDPWR.n2233 9.3005
R9652 VDPWR.n2232 VDPWR.n2198 9.3005
R9653 VDPWR.n2230 VDPWR.n2229 9.3005
R9654 VDPWR.n2228 VDPWR.n2200 9.3005
R9655 VDPWR.n2227 VDPWR.n2226 9.3005
R9656 VDPWR.n2225 VDPWR.n2224 9.3005
R9657 VDPWR.n2223 VDPWR.n2222 9.3005
R9658 VDPWR.n2220 VDPWR.n2206 9.3005
R9659 VDPWR.n2219 VDPWR.n2218 9.3005
R9660 VDPWR.n2217 VDPWR.n2216 9.3005
R9661 VDPWR.n2215 VDPWR.n2214 9.3005
R9662 VDPWR.n2213 VDPWR.n2212 9.3005
R9663 VDPWR.n2326 VDPWR.n2325 9.3005
R9664 VDPWR.n2324 VDPWR.n2323 9.3005
R9665 VDPWR.n1025 VDPWR.n1020 9.3005
R9666 VDPWR.n2318 VDPWR.n2317 9.3005
R9667 VDPWR.n2315 VDPWR.n2314 9.3005
R9668 VDPWR.n2313 VDPWR.n1026 9.3005
R9669 VDPWR.n2312 VDPWR.n2311 9.3005
R9670 VDPWR.n2309 VDPWR.n1027 9.3005
R9671 VDPWR.n2308 VDPWR.n2307 9.3005
R9672 VDPWR.n2306 VDPWR.n2305 9.3005
R9673 VDPWR.n2304 VDPWR.n1032 9.3005
R9674 VDPWR.n2302 VDPWR.n2301 9.3005
R9675 VDPWR.n2300 VDPWR.n1036 9.3005
R9676 VDPWR.n2299 VDPWR.n2298 9.3005
R9677 VDPWR.n2297 VDPWR.n2296 9.3005
R9678 VDPWR.n1053 VDPWR.n1052 9.3005
R9679 VDPWR.n1056 VDPWR.n1055 9.3005
R9680 VDPWR.n2286 VDPWR.n2285 9.3005
R9681 VDPWR.n2283 VDPWR.n1049 9.3005
R9682 VDPWR.n2281 VDPWR.n2280 9.3005
R9683 VDPWR.n2279 VDPWR.n1059 9.3005
R9684 VDPWR.n2278 VDPWR.n2277 9.3005
R9685 VDPWR.n2275 VDPWR.n1060 9.3005
R9686 VDPWR.n2274 VDPWR.n2273 9.3005
R9687 VDPWR.n2272 VDPWR.n2271 9.3005
R9688 VDPWR.n2270 VDPWR.n2269 9.3005
R9689 VDPWR.n2268 VDPWR.n2267 9.3005
R9690 VDPWR.n2266 VDPWR.n1067 9.3005
R9691 VDPWR.n2264 VDPWR.n2263 9.3005
R9692 VDPWR.n2974 VDPWR.n2973 9.3005
R9693 VDPWR.n2973 VDPWR.n928 9.3005
R9694 VDPWR.n2973 VDPWR.n2969 9.3005
R9695 VDPWR.n2738 VDPWR.n2737 9.3005
R9696 VDPWR.n2745 VDPWR.n2744 9.3005
R9697 VDPWR.n2750 VDPWR.n2749 9.3005
R9698 VDPWR.n2749 VDPWR.n2748 9.3005
R9699 VDPWR.n2760 VDPWR.n2759 9.3005
R9700 VDPWR.n2761 VDPWR.n1004 9.3005
R9701 VDPWR.n2764 VDPWR.n2763 9.3005
R9702 VDPWR.n2765 VDPWR.n1003 9.3005
R9703 VDPWR.n2767 VDPWR.n2766 9.3005
R9704 VDPWR.n2771 VDPWR.n1002 9.3005
R9705 VDPWR.n2775 VDPWR.n2774 9.3005
R9706 VDPWR.n2778 VDPWR.n2777 9.3005
R9707 VDPWR.n2780 VDPWR.n2779 9.3005
R9708 VDPWR.n2786 VDPWR.n2785 9.3005
R9709 VDPWR.n2788 VDPWR.n2787 9.3005
R9710 VDPWR.n2789 VDPWR.n993 9.3005
R9711 VDPWR.n2797 VDPWR.n2796 9.3005
R9712 VDPWR.n2795 VDPWR.n985 9.3005
R9713 VDPWR.n2809 VDPWR.n984 9.3005
R9714 VDPWR.n2813 VDPWR.n2810 9.3005
R9715 VDPWR.n2818 VDPWR.n2817 9.3005
R9716 VDPWR.n2819 VDPWR.n982 9.3005
R9717 VDPWR.n2821 VDPWR.n2820 9.3005
R9718 VDPWR.n2825 VDPWR.n2824 9.3005
R9719 VDPWR.n2826 VDPWR.n981 9.3005
R9720 VDPWR.n2828 VDPWR.n2827 9.3005
R9721 VDPWR.n2831 VDPWR.n2830 9.3005
R9722 VDPWR.n2832 VDPWR.n980 9.3005
R9723 VDPWR.n2834 VDPWR.n2833 9.3005
R9724 VDPWR.n2838 VDPWR.n2837 9.3005
R9725 VDPWR.n2839 VDPWR.n969 9.3005
R9726 VDPWR.n2850 VDPWR.n2849 9.3005
R9727 VDPWR.n2855 VDPWR.n2854 9.3005
R9728 VDPWR.n2856 VDPWR.n967 9.3005
R9729 VDPWR.n2858 VDPWR.n2857 9.3005
R9730 VDPWR.n2860 VDPWR.n966 9.3005
R9731 VDPWR.n2862 VDPWR.n2861 9.3005
R9732 VDPWR.n2863 VDPWR.n965 9.3005
R9733 VDPWR.n2865 VDPWR.n2864 9.3005
R9734 VDPWR.n2867 VDPWR.n963 9.3005
R9735 VDPWR.n2869 VDPWR.n2868 9.3005
R9736 VDPWR.n2871 VDPWR.n2870 9.3005
R9737 VDPWR.n2876 VDPWR.n2875 9.3005
R9738 VDPWR.n2883 VDPWR.n2882 9.3005
R9739 VDPWR.n2886 VDPWR.n959 9.3005
R9740 VDPWR.n2892 VDPWR.n2891 9.3005
R9741 VDPWR.n2888 VDPWR.n955 9.3005
R9742 VDPWR.n2900 VDPWR.n954 9.3005
R9743 VDPWR.n2902 VDPWR.n2901 9.3005
R9744 VDPWR.n2905 VDPWR.n2904 9.3005
R9745 VDPWR.n2907 VDPWR.n2906 9.3005
R9746 VDPWR.n2908 VDPWR.n951 9.3005
R9747 VDPWR.n2911 VDPWR.n2910 9.3005
R9748 VDPWR.n2913 VDPWR.n2912 9.3005
R9749 VDPWR.n2914 VDPWR.n949 9.3005
R9750 VDPWR.n2918 VDPWR.n2917 9.3005
R9751 VDPWR.n2919 VDPWR.n948 9.3005
R9752 VDPWR.n2921 VDPWR.n2920 9.3005
R9753 VDPWR.n2922 VDPWR.n947 9.3005
R9754 VDPWR.n2924 VDPWR.n2923 9.3005
R9755 VDPWR.n2937 VDPWR.n2936 9.3005
R9756 VDPWR.n2939 VDPWR.n938 9.3005
R9757 VDPWR.n2942 VDPWR.n2941 9.3005
R9758 VDPWR.n2944 VDPWR.n2943 9.3005
R9759 VDPWR.n2948 VDPWR.n2947 9.3005
R9760 VDPWR.n2949 VDPWR.n935 9.3005
R9761 VDPWR.n2951 VDPWR.n2950 9.3005
R9762 VDPWR.n2954 VDPWR.n2953 9.3005
R9763 VDPWR.n2955 VDPWR.n934 9.3005
R9764 VDPWR.n2957 VDPWR.n2956 9.3005
R9765 VDPWR.n2958 VDPWR.n933 9.3005
R9766 VDPWR.n2961 VDPWR.n2960 9.3005
R9767 VDPWR.n2962 VDPWR.n929 9.3005
R9768 VDPWR.n3001 VDPWR.n3000 9.3005
R9769 VDPWR.n3000 VDPWR.n2996 9.3005
R9770 VDPWR.n3000 VDPWR.n2993 9.3005
R9771 VDPWR.n2568 VDPWR.n2567 9.3005
R9772 VDPWR.n2566 VDPWR.n2548 9.3005
R9773 VDPWR.n2578 VDPWR.n2577 9.3005
R9774 VDPWR.n2715 VDPWR.n2714 9.3005
R9775 VDPWR.n2713 VDPWR.n2544 9.3005
R9776 VDPWR.n2712 VDPWR.n2711 9.3005
R9777 VDPWR.n2710 VDPWR.n2579 9.3005
R9778 VDPWR.n2709 VDPWR.n2708 9.3005
R9779 VDPWR.n2706 VDPWR.n2580 9.3005
R9780 VDPWR.n2705 VDPWR.n2704 9.3005
R9781 VDPWR.n2703 VDPWR.n2583 9.3005
R9782 VDPWR.n2702 VDPWR.n2701 9.3005
R9783 VDPWR.n2700 VDPWR.n2584 9.3005
R9784 VDPWR.n2699 VDPWR.n2698 9.3005
R9785 VDPWR.n2697 VDPWR.n2587 9.3005
R9786 VDPWR.n2594 VDPWR.n2588 9.3005
R9787 VDPWR.n2687 VDPWR.n2602 9.3005
R9788 VDPWR.n2687 VDPWR.n2593 9.3005
R9789 VDPWR.n2688 VDPWR.n2687 9.3005
R9790 VDPWR.n2686 VDPWR.n2604 9.3005
R9791 VDPWR.n2683 VDPWR.n2682 9.3005
R9792 VDPWR.n2681 VDPWR.n2605 9.3005
R9793 VDPWR.n2680 VDPWR.n2679 9.3005
R9794 VDPWR.n2678 VDPWR.n2606 9.3005
R9795 VDPWR.n2675 VDPWR.n2674 9.3005
R9796 VDPWR.n2673 VDPWR.n2610 9.3005
R9797 VDPWR.n2672 VDPWR.n2671 9.3005
R9798 VDPWR.n2670 VDPWR.n2611 9.3005
R9799 VDPWR.n2668 VDPWR.n2667 9.3005
R9800 VDPWR.n2614 VDPWR.n2613 9.3005
R9801 VDPWR.n2651 VDPWR.n2649 9.3005
R9802 VDPWR.n2656 VDPWR.n2655 9.3005
R9803 VDPWR.n2658 VDPWR.n2657 9.3005
R9804 VDPWR.n2657 VDPWR.n2646 9.3005
R9805 VDPWR.n2645 VDPWR.n2620 9.3005
R9806 VDPWR.n2644 VDPWR.n2643 9.3005
R9807 VDPWR.n2641 VDPWR.n2640 9.3005
R9808 VDPWR.n2639 VDPWR.n2621 9.3005
R9809 VDPWR.n2638 VDPWR.n2637 9.3005
R9810 VDPWR.n2635 VDPWR.n2622 9.3005
R9811 VDPWR.n2632 VDPWR.n2631 9.3005
R9812 VDPWR.n2630 VDPWR.n2629 9.3005
R9813 VDPWR.n3062 VDPWR.n3061 9.3005
R9814 VDPWR.n3060 VDPWR.n3059 9.3005
R9815 VDPWR.n885 VDPWR.n880 9.3005
R9816 VDPWR.n3054 VDPWR.n3053 9.3005
R9817 VDPWR.n3050 VDPWR.n3049 9.3005
R9818 VDPWR.n3048 VDPWR.n892 9.3005
R9819 VDPWR.n3047 VDPWR.n3046 9.3005
R9820 VDPWR.n3045 VDPWR.n895 9.3005
R9821 VDPWR.n3044 VDPWR.n3043 9.3005
R9822 VDPWR.n3042 VDPWR.n3041 9.3005
R9823 VDPWR.n3040 VDPWR.n898 9.3005
R9824 VDPWR.n3039 VDPWR.n3038 9.3005
R9825 VDPWR.n911 VDPWR.n910 9.3005
R9826 VDPWR.n912 VDPWR.n907 9.3005
R9827 VDPWR.n3028 VDPWR.n3027 9.3005
R9828 VDPWR.n3025 VDPWR.n908 9.3005
R9829 VDPWR.n3024 VDPWR.n914 9.3005
R9830 VDPWR.n3023 VDPWR.n3022 9.3005
R9831 VDPWR.n3021 VDPWR.n916 9.3005
R9832 VDPWR.n3020 VDPWR.n3019 9.3005
R9833 VDPWR.n3018 VDPWR.n3017 9.3005
R9834 VDPWR.n3016 VDPWR.n3015 9.3005
R9835 VDPWR.n3013 VDPWR.n918 9.3005
R9836 VDPWR.n3012 VDPWR.n3011 9.3005
R9837 VDPWR.n3010 VDPWR.n920 9.3005
R9838 VDPWR.n2988 VDPWR.n921 9.3005
R9839 VDPWR.n843 VDPWR.n842 9.3005
R9840 VDPWR.n843 VDPWR.n835 9.3005
R9841 VDPWR.n844 VDPWR.n843 9.3005
R9842 VDPWR.n2380 VDPWR.n2379 9.3005
R9843 VDPWR.n2382 VDPWR.n2381 9.3005
R9844 VDPWR.n2383 VDPWR.n2369 9.3005
R9845 VDPWR.n2385 VDPWR.n2384 9.3005
R9846 VDPWR.n2386 VDPWR.n2367 9.3005
R9847 VDPWR.n2388 VDPWR.n2387 9.3005
R9848 VDPWR.n2397 VDPWR.n2396 9.3005
R9849 VDPWR.n2400 VDPWR.n2358 9.3005
R9850 VDPWR.n2402 VDPWR.n2401 9.3005
R9851 VDPWR.n2404 VDPWR.n2403 9.3005
R9852 VDPWR.n2405 VDPWR.n2354 9.3005
R9853 VDPWR.n2407 VDPWR.n2406 9.3005
R9854 VDPWR.n2408 VDPWR.n2353 9.3005
R9855 VDPWR.n2410 VDPWR.n2409 9.3005
R9856 VDPWR.n2413 VDPWR.n2412 9.3005
R9857 VDPWR.n2414 VDPWR.n2351 9.3005
R9858 VDPWR.n2416 VDPWR.n2415 9.3005
R9859 VDPWR.n2418 VDPWR.n2350 9.3005
R9860 VDPWR.n2423 VDPWR.n2422 9.3005
R9861 VDPWR.n2425 VDPWR.n2349 9.3005
R9862 VDPWR.n2430 VDPWR.n2429 9.3005
R9863 VDPWR.n2532 VDPWR.n2531 9.3005
R9864 VDPWR.n2530 VDPWR.n2529 9.3005
R9865 VDPWR.n2528 VDPWR.n2433 9.3005
R9866 VDPWR.n2527 VDPWR.n2526 9.3005
R9867 VDPWR.n2524 VDPWR.n2523 9.3005
R9868 VDPWR.n2522 VDPWR.n2521 9.3005
R9869 VDPWR.n2520 VDPWR.n2435 9.3005
R9870 VDPWR.n2518 VDPWR.n2517 9.3005
R9871 VDPWR.n2516 VDPWR.n2515 9.3005
R9872 VDPWR.n2514 VDPWR.n2439 9.3005
R9873 VDPWR.n2513 VDPWR.n2440 9.3005
R9874 VDPWR.n2512 VDPWR.n2511 9.3005
R9875 VDPWR.n2443 VDPWR.n2442 9.3005
R9876 VDPWR.n2451 VDPWR.n2448 9.3005
R9877 VDPWR.n2493 VDPWR.n2492 9.3005
R9878 VDPWR.n2490 VDPWR.n2489 9.3005
R9879 VDPWR.n2488 VDPWR.n2454 9.3005
R9880 VDPWR.n2487 VDPWR.n2486 9.3005
R9881 VDPWR.n2484 VDPWR.n2455 9.3005
R9882 VDPWR.n2483 VDPWR.n2482 9.3005
R9883 VDPWR.n2481 VDPWR.n2480 9.3005
R9884 VDPWR.n2479 VDPWR.n2457 9.3005
R9885 VDPWR.n2478 VDPWR.n2477 9.3005
R9886 VDPWR.n2469 VDPWR.n2468 9.3005
R9887 VDPWR.n2463 VDPWR.n787 9.3005
R9888 VDPWR.n3098 VDPWR.n3097 9.3005
R9889 VDPWR.n3096 VDPWR.n790 9.3005
R9890 VDPWR.n3095 VDPWR.n3094 9.3005
R9891 VDPWR.n3093 VDPWR.n3092 9.3005
R9892 VDPWR.n3089 VDPWR.n3088 9.3005
R9893 VDPWR.n3087 VDPWR.n793 9.3005
R9894 VDPWR.n3086 VDPWR.n3085 9.3005
R9895 VDPWR.n3084 VDPWR.n794 9.3005
R9896 VDPWR.n3083 VDPWR.n3082 9.3005
R9897 VDPWR.n3081 VDPWR.n3080 9.3005
R9898 VDPWR.n3079 VDPWR.n3078 9.3005
R9899 VDPWR.n3077 VDPWR.n800 9.3005
R9900 VDPWR.n808 VDPWR.n801 9.3005
R9901 VDPWR.n812 VDPWR.n811 9.3005
R9902 VDPWR.n866 VDPWR.n865 9.3005
R9903 VDPWR.n863 VDPWR.n862 9.3005
R9904 VDPWR.n861 VDPWR.n815 9.3005
R9905 VDPWR.n860 VDPWR.n859 9.3005
R9906 VDPWR.n858 VDPWR.n816 9.3005
R9907 VDPWR.n856 VDPWR.n855 9.3005
R9908 VDPWR.n853 VDPWR.n852 9.3005
R9909 VDPWR.n851 VDPWR.n850 9.3005
R9910 VDPWR.n849 VDPWR.n826 9.3005
R9911 VDPWR.n831 VDPWR.n827 9.3005
R9912 VDPWR.n52 VDPWR.n28 9.3005
R9913 VDPWR.n88 VDPWR.n87 9.3005
R9914 VDPWR.n85 VDPWR.n29 9.3005
R9915 VDPWR.n84 VDPWR.n82 9.3005
R9916 VDPWR.n81 VDPWR.n53 9.3005
R9917 VDPWR.n80 VDPWR.n79 9.3005
R9918 VDPWR.n78 VDPWR.n54 9.3005
R9919 VDPWR.n77 VDPWR.n76 9.3005
R9920 VDPWR.n75 VDPWR.n55 9.3005
R9921 VDPWR.n74 VDPWR.n73 9.3005
R9922 VDPWR.n72 VDPWR.n71 9.3005
R9923 VDPWR.n70 VDPWR.n56 9.3005
R9924 VDPWR.n69 VDPWR.n68 9.3005
R9925 VDPWR.n67 VDPWR.n66 9.3005
R9926 VDPWR.n65 VDPWR.n64 9.3005
R9927 VDPWR.n63 VDPWR.n59 9.3005
R9928 VDPWR.n35 VDPWR.n34 9.3005
R9929 VDPWR.n38 VDPWR.n30 9.3005
R9930 VDPWR.n47 VDPWR.n46 9.3005
R9931 VDPWR.n44 VDPWR.n31 9.3005
R9932 VDPWR.n43 VDPWR.n42 9.3005
R9933 VDPWR.n41 VDPWR.n26 9.3005
R9934 VDPWR.n92 VDPWR.n91 9.3005
R9935 VDPWR.n93 VDPWR.n25 9.3005
R9936 VDPWR.n98 VDPWR.n97 9.3005
R9937 VDPWR.n99 VDPWR.n24 9.3005
R9938 VDPWR.n102 VDPWR.n101 9.3005
R9939 VDPWR.n100 VDPWR.n1 9.3005
R9940 VDPWR.n114 VDPWR.n113 9.3005
R9941 VDPWR.n112 VDPWR.n0 9.3005
R9942 VDPWR.n111 VDPWR.n110 9.3005
R9943 VDPWR.n109 VDPWR.n108 9.3005
R9944 VDPWR.n107 VDPWR.n4 9.3005
R9945 VDPWR.n106 VDPWR.n9 9.3005
R9946 VDPWR.n21 VDPWR.n20 9.3005
R9947 VDPWR.n19 VDPWR.n18 9.3005
R9948 VDPWR.n16 VDPWR.n11 9.3005
R9949 VDPWR.n1520 VDPWR.n1519 9.09802
R9950 VDPWR.n2317 VDPWR.n2316 9.09802
R9951 VDPWR.n2311 VDPWR.n1029 9.09802
R9952 VDPWR.n2311 VDPWR.n2310 9.09802
R9953 VDPWR.n2923 VDPWR.n939 9.09802
R9954 VDPWR.n2941 VDPWR.n2940 9.09802
R9955 VDPWR.n2222 VDPWR.n2207 9.02345
R9956 VDPWR.n1052 VDPWR.n1051 9.02345
R9957 VDPWR.n2284 VDPWR.n2283 9.02345
R9958 VDPWR.n1841 VDPWR.n1840 8.99224
R9959 VDPWR.n823 VDPWR.n820 8.9761
R9960 VDPWR.n2907 VDPWR.n953 8.88645
R9961 VDPWR.n2788 VDPWR.n998 8.77764
R9962 VDPWR.n2222 VDPWR.n2221 8.60378
R9963 VDPWR.n2277 VDPWR.n2276 8.60378
R9964 VDPWR.n1431 VDPWR.n1428 8.44958
R9965 VDPWR.n1760 VDPWR.n1263 8.44958
R9966 VDPWR.n1825 VDPWR.n1224 8.44958
R9967 VDPWR.n2001 VDPWR.n1178 8.44958
R9968 VDPWR.n2058 VDPWR.n1126 8.44958
R9969 VDPWR.n2167 VDPWR.n1110 8.44958
R9970 VDPWR.t331 VDPWR.t775 8.39273
R9971 VDPWR.n2282 VDPWR.n2281 8.28902
R9972 VDPWR.n1872 VDPWR.n1871 8.28285
R9973 VDPWR.n2677 VDPWR.n2676 8.28285
R9974 VDPWR.n671 VDPWR.n657 8.23557
R9975 VDPWR.n428 VDPWR.n414 8.23557
R9976 VDPWR.n2791 VDPWR.n2790 8.04621
R9977 VDPWR.n2274 VDPWR.n1065 8.04017
R9978 VDPWR.n1766 VDPWR.n1257 7.98741
R9979 VDPWR.n2480 VDPWR 7.93438
R9980 VDPWR.n2678 VDPWR.n2677 7.90638
R9981 VDPWR.n2686 VDPWR.n2684 7.90638
R9982 VDPWR.n1518 VDPWR.n1516 7.75995
R9983 VDPWR.n2001 VDPWR.n2000 7.75995
R9984 VDPWR.n2215 VDPWR.n2212 7.75995
R9985 VDPWR.n2317 VDPWR.n1025 7.75995
R9986 VDPWR.n2271 VDPWR.n2270 7.75995
R9987 VDPWR.n2953 VDPWR.n2951 7.75995
R9988 VDPWR.n2484 VDPWR.n2483 7.75995
R9989 VDPWR.n2203 VDPWR.n2202 7.65952
R9990 VDPWR.n718 VDPWR.n717 7.54407
R9991 VDPWR.n702 VDPWR.n701 7.54407
R9992 VDPWR.n686 VDPWR.n685 7.54407
R9993 VDPWR.n670 VDPWR.n669 7.54407
R9994 VDPWR.n529 VDPWR.n528 7.54407
R9995 VDPWR.n513 VDPWR.n512 7.54407
R9996 VDPWR.n497 VDPWR.n496 7.54407
R9997 VDPWR.n481 VDPWR.n480 7.54407
R9998 VDPWR.n459 VDPWR.n458 7.54407
R9999 VDPWR.n443 VDPWR.n442 7.54407
R10000 VDPWR.n427 VDPWR.n426 7.54407
R10001 VDPWR.n3170 VDPWR.n3169 7.54407
R10002 VDPWR.n3132 VDPWR.n3131 7.54407
R10003 VDPWR.n465 VDPWR.n464 7.54307
R10004 VDPWR.n3164 VDPWR.n3163 7.54307
R10005 VDPWR.n3148 VDPWR.n3147 7.54307
R10006 VDPWR.n2910 VDPWR.n2909 7.51124
R10007 VDPWR.n2515 VDPWR.n2514 7.49704
R10008 VDPWR.n1108 VDPWR.n1105 7.28326
R10009 VDPWR.n1106 VDPWR.n1104 7.23528
R10010 VDPWR.n2017 VDPWR.n2016 7.21067
R10011 VDPWR.n2026 VDPWR.n1151 7.21067
R10012 VDPWR.n2142 VDPWR.n2140 7.21067
R10013 VDPWR.n2186 VDPWR.n2185 7.17134
R10014 VDPWR.n1502 VDPWR.n1296 7.12524
R10015 VDPWR.n537 VDPWR.n532 7.10511
R10016 VDPWR.n2231 VDPWR.n2230 7.03001
R10017 VDPWR.n546 VDPWR.n543 6.8005
R10018 VDPWR.n266 VDPWR.n263 6.8005
R10019 VDPWR.n8 VDPWR.n5 6.8005
R10020 VDPWR.n1871 VDPWR.n1870 6.77697
R10021 VDPWR.n1990 VDPWR.n1182 6.77697
R10022 VDPWR.n3051 VDPWR.n3050 6.77697
R10023 VDPWR.n858 VDPWR.n857 6.73838
R10024 VDPWR.t136 VDPWR.t6 6.71428
R10025 VDPWR.t918 VDPWR.t348 6.71428
R10026 VDPWR.t1015 VDPWR.t9 6.71428
R10027 VDPWR.t807 VDPWR.t805 6.71428
R10028 VDPWR.t229 VDPWR.t223 6.71428
R10029 VDPWR.n1431 VDPWR.n1327 6.66496
R10030 VDPWR.n1762 VDPWR.n1761 6.66496
R10031 VDPWR.n1826 VDPWR.n1825 6.66496
R10032 VDPWR.n1836 VDPWR.n1834 6.66496
R10033 VDPWR.n1127 VDPWR.n1126 6.66496
R10034 VDPWR.n2172 VDPWR.n2171 6.66496
R10035 VDPWR.n2478 VDPWR.n2459 6.66496
R10036 VDPWR.n1396 VDPWR.n1341 6.52104
R10037 VDPWR.n1726 VDPWR.n1277 6.52104
R10038 VDPWR.n2135 VDPWR.n2134 6.52104
R10039 VDPWR.n2041 VDPWR.n2040 6.52104
R10040 VDPWR.n1650 VDPWR.n1649 6.52104
R10041 VDPWR.n2188 VDPWR.n1100 6.50542
R10042 VDPWR.n2304 VDPWR.n2303 6.50542
R10043 VDPWR.n1261 VDPWR.n1260 6.48583
R10044 VDPWR.n2475 VDPWR.n2474 6.48583
R10045 VDPWR.n2471 VDPWR.n2470 6.46951
R10046 VDPWR.n2865 VDPWR.n965 6.4005
R10047 VDPWR.n2387 VDPWR 6.4005
R10048 VDPWR.n2470 VDPWR.n2469 6.4005
R10049 VDPWR.n749 VDPWR.n748 6.37981
R10050 VDPWR.n745 VDPWR.n743 6.37981
R10051 VDPWR.n737 VDPWR.n736 6.37981
R10052 VDPWR.n734 VDPWR.n733 6.37981
R10053 VDPWR.n2771 VDPWR.n2768 6.3005
R10054 VDPWR.n720 VDPWR.n656 6.18087
R10055 VDPWR.n3177 VDPWR.n3172 6.12434
R10056 VDPWR.n714 VDPWR.n705 6.02403
R10057 VDPWR.n661 VDPWR.n658 6.02403
R10058 VDPWR.n525 VDPWR.n516 6.02403
R10059 VDPWR.n477 VDPWR.n468 6.02403
R10060 VDPWR.n413 VDPWR.n404 6.02403
R10061 VDPWR.n418 VDPWR.n415 6.02403
R10062 VDPWR.n769 VDPWR.n760 6.02403
R10063 VDPWR.n3128 VDPWR.n3119 6.02403
R10064 VDPWR.n2741 VDPWR.n2740 5.97436
R10065 VDPWR.n1259 VDPWR.n1258 5.8885
R10066 VDPWR.n2473 VDPWR.n2472 5.8885
R10067 VDPWR.n2796 VDPWR.n2791 5.85193
R10068 VDPWR.n3177 VDPWR.n3176 5.75618
R10069 VDPWR.n2233 VDPWR.n2196 5.66607
R10070 VDPWR.n1052 VDPWR.n1041 5.66607
R10071 VDPWR.n1439 VDPWR.n1438 5.66204
R10072 VDPWR.n1441 VDPWR.n1439 5.66204
R10073 VDPWR.n1445 VDPWR.n1321 5.66204
R10074 VDPWR.n1446 VDPWR.n1445 5.66204
R10075 VDPWR.n1446 VDPWR.n1314 5.66204
R10076 VDPWR.n1461 VDPWR.n1314 5.66204
R10077 VDPWR.n1462 VDPWR.n1461 5.66204
R10078 VDPWR.n1463 VDPWR.n1462 5.66204
R10079 VDPWR.n1470 VDPWR.n1469 5.66204
R10080 VDPWR.n1471 VDPWR.n1470 5.66204
R10081 VDPWR.n1475 VDPWR.n1474 5.66204
R10082 VDPWR.n1476 VDPWR.n1475 5.66204
R10083 VDPWR.n1476 VDPWR.n1307 5.66204
R10084 VDPWR.n1480 VDPWR.n1307 5.66204
R10085 VDPWR.n1486 VDPWR.n1480 5.66204
R10086 VDPWR.n1486 VDPWR.n1485 5.66204
R10087 VDPWR.n1399 VDPWR.n1398 5.66204
R10088 VDPWR.n1406 VDPWR.n1337 5.66204
R10089 VDPWR.n1410 VDPWR.n1337 5.66204
R10090 VDPWR.n1414 VDPWR.n1412 5.66204
R10091 VDPWR.n1414 VDPWR.n1413 5.66204
R10092 VDPWR.n1572 VDPWR.n1571 5.66204
R10093 VDPWR.n1571 VDPWR.n1570 5.66204
R10094 VDPWR.n1567 VDPWR.n1566 5.66204
R10095 VDPWR.n1566 VDPWR.n1565 5.66204
R10096 VDPWR.n1565 VDPWR.n1526 5.66204
R10097 VDPWR.n1561 VDPWR.n1526 5.66204
R10098 VDPWR.n1561 VDPWR.n1560 5.66204
R10099 VDPWR.n1560 VDPWR.n1559 5.66204
R10100 VDPWR.n1729 VDPWR.n1728 5.66204
R10101 VDPWR.n1736 VDPWR.n1273 5.66204
R10102 VDPWR.n1740 VDPWR.n1273 5.66204
R10103 VDPWR.n1745 VDPWR.n1742 5.66204
R10104 VDPWR.n1745 VDPWR.n1744 5.66204
R10105 VDPWR.n1775 VDPWR.n1255 5.66204
R10106 VDPWR.n1778 VDPWR.n1777 5.66204
R10107 VDPWR.n1778 VDPWR.n1241 5.66204
R10108 VDPWR.n1789 VDPWR.n1241 5.66204
R10109 VDPWR.n1790 VDPWR.n1789 5.66204
R10110 VDPWR.n1803 VDPWR.n1802 5.66204
R10111 VDPWR.n1805 VDPWR.n1235 5.66204
R10112 VDPWR.n1809 VDPWR.n1235 5.66204
R10113 VDPWR.n1814 VDPWR.n1809 5.66204
R10114 VDPWR.n1814 VDPWR.n1813 5.66204
R10115 VDPWR.n2013 VDPWR.n2012 5.66204
R10116 VDPWR.n2012 VDPWR.n2011 5.66204
R10117 VDPWR.n1176 VDPWR.n1168 5.66204
R10118 VDPWR.n2022 VDPWR.n2021 5.66204
R10119 VDPWR.n2021 VDPWR.n2020 5.66204
R10120 VDPWR.n1148 VDPWR.n1142 5.66204
R10121 VDPWR.n1149 VDPWR.n1148 5.66204
R10122 VDPWR.n2029 VDPWR.n2028 5.66204
R10123 VDPWR.n1638 VDPWR.n1637 5.66204
R10124 VDPWR.n1637 VDPWR.n1634 5.66204
R10125 VDPWR.n1632 VDPWR.n1125 5.66204
R10126 VDPWR.n2060 VDPWR.n1125 5.66204
R10127 VDPWR.n1646 VDPWR.n1645 5.66204
R10128 VDPWR.n2146 VDPWR.n2145 5.66204
R10129 VDPWR.n2147 VDPWR.n2146 5.66204
R10130 VDPWR.n2151 VDPWR.n2150 5.66204
R10131 VDPWR.n2151 VDPWR.n1112 5.66204
R10132 VDPWR.n2165 VDPWR.n1112 5.66204
R10133 VDPWR.n535 VDPWR 5.6325
R10134 VDPWR.n3175 VDPWR 5.6325
R10135 VDPWR.n1792 VDPWR.n1239 5.48759
R10136 VDPWR.n1768 VDPWR.n1767 5.42606
R10137 VDPWR.n1797 VDPWR.n1796 5.42606
R10138 VDPWR.n1833 VDPWR.n1222 5.3712
R10139 VDPWR.n1438 VDPWR.n1323 5.29281
R10140 VDPWR.n1463 VDPWR.n1312 5.29281
R10141 VDPWR.n1469 VDPWR.n1311 5.29281
R10142 VDPWR.n1485 VDPWR.n1482 5.29281
R10143 VDPWR.n1398 VDPWR.n1397 5.29281
R10144 VDPWR.n1399 VDPWR.n1339 5.29281
R10145 VDPWR.n1406 VDPWR.n1405 5.29281
R10146 VDPWR.n1413 VDPWR.n1328 5.29281
R10147 VDPWR.n1572 VDPWR.n1521 5.29281
R10148 VDPWR.n1559 VDPWR.n1528 5.29281
R10149 VDPWR.n1728 VDPWR.n1727 5.29281
R10150 VDPWR.n1729 VDPWR.n1275 5.29281
R10151 VDPWR.n1736 VDPWR.n1735 5.29281
R10152 VDPWR.n1744 VDPWR.n1743 5.29281
R10153 VDPWR.n1771 VDPWR.n1769 5.29281
R10154 VDPWR.n1791 VDPWR.n1790 5.29281
R10155 VDPWR.n1799 VDPWR.n1798 5.29281
R10156 VDPWR.n1813 VDPWR.n1810 5.29281
R10157 VDPWR.n2013 VDPWR.n1156 5.29281
R10158 VDPWR.n1177 VDPWR.n1176 5.29281
R10159 VDPWR.n2022 VDPWR.n1153 5.29281
R10160 VDPWR.n1142 VDPWR.n1134 5.29281
R10161 VDPWR.n2028 VDPWR.n2027 5.29281
R10162 VDPWR.n1639 VDPWR.n1638 5.29281
R10163 VDPWR.n2060 VDPWR.n2059 5.29281
R10164 VDPWR.n1646 VDPWR.n1628 5.29281
R10165 VDPWR.n1645 VDPWR.n1644 5.29281
R10166 VDPWR.n2137 VDPWR.n2136 5.29281
R10167 VDPWR.n2137 VDPWR.n2080 5.29281
R10168 VDPWR.n2166 VDPWR.n2165 5.29281
R10169 VDPWR.n2871 VDPWR.n962 5.27109
R10170 VDPWR.n2531 VDPWR.n2431 5.27109
R10171 VDPWR.n2095 VDPWR.n2094 5.25888
R10172 VDPWR.n2194 VDPWR.n2193 5.2464
R10173 VDPWR.n1039 VDPWR.n1036 5.2464
R10174 VDPWR.n1836 VDPWR.n1835 5.18397
R10175 VDPWR.n1849 VDPWR.n1848 5.18397
R10176 VDPWR.n2219 VDPWR.n2209 5.18397
R10177 VDPWR.n2910 VDPWR.n950 5.18397
R10178 VDPWR.n2916 VDPWR.n948 5.18397
R10179 VDPWR.n717 VDPWR.n716 5.18145
R10180 VDPWR.n701 VDPWR.n700 5.18145
R10181 VDPWR.n685 VDPWR.n684 5.18145
R10182 VDPWR.n669 VDPWR.n668 5.18145
R10183 VDPWR.n528 VDPWR.n527 5.18145
R10184 VDPWR.n512 VDPWR.n511 5.18145
R10185 VDPWR.n496 VDPWR.n495 5.18145
R10186 VDPWR.n480 VDPWR.n479 5.18145
R10187 VDPWR.n464 VDPWR.n463 5.18145
R10188 VDPWR.n458 VDPWR.n457 5.18145
R10189 VDPWR.n442 VDPWR.n441 5.18145
R10190 VDPWR.n426 VDPWR.n425 5.18145
R10191 VDPWR.n3169 VDPWR.n3168 5.18145
R10192 VDPWR.n3163 VDPWR.n3162 5.18145
R10193 VDPWR.n3147 VDPWR.n3146 5.18145
R10194 VDPWR.n3131 VDPWR.n3130 5.18145
R10195 VDPWR.n2192 VDPWR.n2191 5.14148
R10196 VDPWR.n2785 VDPWR.n2784 5.1205
R10197 VDPWR.n2308 VDPWR.n1031 5.103
R10198 VDPWR.n1063 VDPWR.n1062 5.03657
R10199 VDPWR.t133 VDPWR.t346 5.03584
R10200 VDPWR.t134 VDPWR.t1004 5.03584
R10201 VDPWR.t562 VDPWR.t254 5.03584
R10202 VDPWR.t797 VDPWR.t785 5.03584
R10203 VDPWR.t334 VDPWR.t294 5.03584
R10204 VDPWR.n824 VDPWR.n822 4.98336
R10205 VDPWR.n2874 VDPWR.n961 4.9005
R10206 VDPWR.n699 VDPWR.n691 4.89462
R10207 VDPWR.n675 VDPWR.n673 4.89462
R10208 VDPWR.n510 VDPWR.n502 4.89462
R10209 VDPWR.n486 VDPWR.n484 4.89462
R10210 VDPWR.n456 VDPWR.n448 4.89462
R10211 VDPWR.n432 VDPWR.n430 4.89462
R10212 VDPWR.n3161 VDPWR.n3153 4.89462
R10213 VDPWR.n3137 VDPWR.n3135 4.89462
R10214 VDPWR.n3133 VDPWR.n3118 4.72727
R10215 VDPWR.n2108 VDPWR.n2107 4.69218
R10216 VDPWR.n602 VDPWR.n601 4.67352
R10217 VDPWR.n625 VDPWR.n590 4.67352
R10218 VDPWR.n322 VDPWR.n321 4.67352
R10219 VDPWR.n345 VDPWR.n310 4.67352
R10220 VDPWR.n1959 VDPWR.n1958 4.67352
R10221 VDPWR.n2891 VDPWR.n2886 4.67352
R10222 VDPWR.n2761 VDPWR.n2760 4.67352
R10223 VDPWR.n3061 VDPWR.n3060 4.67352
R10224 VDPWR.n3013 VDPWR.n3012 4.67352
R10225 VDPWR.n3012 VDPWR.n920 4.67352
R10226 VDPWR.n2416 VDPWR.n2351 4.67352
R10227 VDPWR.n2422 VDPWR.n2418 4.67352
R10228 VDPWR.n2401 VDPWR.n2400 4.67352
R10229 VDPWR.n2521 VDPWR.n2520 4.67352
R10230 VDPWR.n3089 VDPWR.n793 4.67352
R10231 VDPWR.n3085 VDPWR.n3084 4.67352
R10232 VDPWR.n3084 VDPWR.n3083 4.67352
R10233 VDPWR.n863 VDPWR.n815 4.67352
R10234 VDPWR.n859 VDPWR.n815 4.67352
R10235 VDPWR.n859 VDPWR.n858 4.67352
R10236 VDPWR.n852 VDPWR.n851 4.67352
R10237 VDPWR.n851 VDPWR.n826 4.67352
R10238 VDPWR.n64 VDPWR.n63 4.67352
R10239 VDPWR.n87 VDPWR.n52 4.67352
R10240 VDPWR.n751 VDPWR.n750 4.6505
R10241 VDPWR.n1968 VDPWR.n1915 4.62124
R10242 VDPWR.n2633 VDPWR.n2624 4.62124
R10243 VDPWR.n1764 VDPWR.n1261 4.62124
R10244 VDPWR.n1766 VDPWR.n1765 4.62124
R10245 VDPWR.n1795 VDPWR.n1794 4.62124
R10246 VDPWR.n2104 VDPWR.n2095 4.62124
R10247 VDPWR.n2476 VDPWR.n2475 4.62124
R10248 VDPWR.n2470 VDPWR.n2460 4.62124
R10249 VDPWR.n2743 VDPWR.n2739 4.5918
R10250 VDPWR.n1961 VDPWR.n1960 4.57193
R10251 VDPWR.n3014 VDPWR.n3013 4.57193
R10252 VDPWR.n2913 VDPWR.n950 4.54926
R10253 VDPWR.n2917 VDPWR.n2916 4.54926
R10254 VDPWR.n2946 VDPWR.n2945 4.54926
R10255 VDPWR.n2945 VDPWR.n935 4.54926
R10256 VDPWR.n2180 VDPWR.n2177 4.52113
R10257 VDPWR.n2868 VDPWR.n962 4.51815
R10258 VDPWR.n2696 VDPWR.n2695 4.51401
R10259 VDPWR.n2690 VDPWR.n2689 4.51401
R10260 VDPWR.n2666 VDPWR.n2665 4.51401
R10261 VDPWR.n2660 VDPWR.n2659 4.51401
R10262 VDPWR.n2510 VDPWR.n2509 4.51401
R10263 VDPWR.n2449 VDPWR.n2446 4.51401
R10264 VDPWR.n1490 VDPWR.n1302 4.51401
R10265 VDPWR.n1495 VDPWR.n1494 4.51401
R10266 VDPWR.n1454 VDPWR.n1319 4.51401
R10267 VDPWR.n1459 VDPWR.n1458 4.51401
R10268 VDPWR.n1421 VDPWR.n1333 4.51401
R10269 VDPWR.n1426 VDPWR.n1425 4.51401
R10270 VDPWR.n1374 VDPWR.n1373 4.51401
R10271 VDPWR.n1387 VDPWR.n1386 4.51401
R10272 VDPWR.n1557 VDPWR.n1556 4.51401
R10273 VDPWR.n1547 VDPWR.n1546 4.51401
R10274 VDPWR.n1586 VDPWR.n1287 4.51401
R10275 VDPWR.n1522 VDPWR.n1290 4.51401
R10276 VDPWR.n1818 VDPWR.n1230 4.51401
R10277 VDPWR.n1823 VDPWR.n1822 4.51401
R10278 VDPWR.n1782 VDPWR.n1248 4.51401
R10279 VDPWR.n1787 VDPWR.n1786 4.51401
R10280 VDPWR.n1752 VDPWR.n1269 4.51401
R10281 VDPWR.n1757 VDPWR.n1756 4.51401
R10282 VDPWR.n1712 VDPWR.n1677 4.51401
R10283 VDPWR.n1717 VDPWR.n1716 4.51401
R10284 VDPWR.n1887 VDPWR.n1886 4.51401
R10285 VDPWR.n1898 VDPWR.n1195 4.51401
R10286 VDPWR.n1856 VDPWR.n1217 4.51401
R10287 VDPWR.n1861 VDPWR.n1212 4.51401
R10288 VDPWR.n2009 VDPWR.n2008 4.51401
R10289 VDPWR.n2004 VDPWR.n2003 4.51401
R10290 VDPWR.n2038 VDPWR.n2037 4.51401
R10291 VDPWR.n2032 VDPWR.n2031 4.51401
R10292 VDPWR.n2070 VDPWR.n1119 4.51401
R10293 VDPWR.n1124 VDPWR.n1123 4.51401
R10294 VDPWR.n1670 VDPWR.n1598 4.51401
R10295 VDPWR.n1661 VDPWR.n1657 4.51401
R10296 VDPWR.n1956 VDPWR.n1955 4.51401
R10297 VDPWR.n1946 VDPWR.n1945 4.51401
R10298 VDPWR.n1188 VDPWR.n1187 4.51401
R10299 VDPWR.n1972 VDPWR.n1971 4.51401
R10300 VDPWR.n2329 VDPWR.n1015 4.51401
R10301 VDPWR.n2320 VDPWR.n2319 4.51401
R10302 VDPWR.n2247 VDPWR.n1094 4.51401
R10303 VDPWR.n2240 VDPWR.n2239 4.51401
R10304 VDPWR.n2157 VDPWR.n2075 4.51401
R10305 VDPWR.n2161 VDPWR.n1111 4.51401
R10306 VDPWR.n2113 VDPWR.n2112 4.51401
R10307 VDPWR.n2127 VDPWR.n2126 4.51401
R10308 VDPWR.n1078 VDPWR.n1076 4.51401
R10309 VDPWR.n1088 VDPWR.n1087 4.51401
R10310 VDPWR.n1043 VDPWR.n1037 4.51401
R10311 VDPWR.n2288 VDPWR.n2287 4.51401
R10312 VDPWR.n2881 VDPWR.n2880 4.51401
R10313 VDPWR.n2899 VDPWR.n2898 4.51401
R10314 VDPWR.n2842 VDPWR.n976 4.51401
R10315 VDPWR.n2846 VDPWR.n968 4.51401
R10316 VDPWR.n2803 VDPWR.n991 4.51401
R10317 VDPWR.n2808 VDPWR.n2807 4.51401
R10318 VDPWR.n2753 VDPWR.n2721 4.51401
R10319 VDPWR.n2758 VDPWR.n2757 4.51401
R10320 VDPWR.n2964 VDPWR.n2963 4.51401
R10321 VDPWR.n2975 VDPWR.n925 4.51401
R10322 VDPWR.n2930 VDPWR.n945 4.51401
R10323 VDPWR.n2935 VDPWR.n2934 4.51401
R10324 VDPWR.n903 VDPWR.n901 4.51401
R10325 VDPWR.n3030 VDPWR.n3029 4.51401
R10326 VDPWR.n3065 VDPWR.n875 4.51401
R10327 VDPWR.n3056 VDPWR.n3055 4.51401
R10328 VDPWR.n2464 VDPWR.n785 4.51401
R10329 VDPWR.n788 VDPWR.n784 4.51401
R10330 VDPWR.n2569 VDPWR.n2549 4.51401
R10331 VDPWR.n2717 VDPWR.n2716 4.51401
R10332 VDPWR.n3009 VDPWR.n3008 4.51401
R10333 VDPWR.n3003 VDPWR.n3002 4.51401
R10334 VDPWR.n2424 VDPWR.n2344 4.51401
R10335 VDPWR.n2346 VDPWR.n2342 4.51401
R10336 VDPWR.n2391 VDPWR.n2365 4.51401
R10337 VDPWR.n2393 VDPWR.n2361 4.51401
R10338 VDPWR.n848 VDPWR.n847 4.51401
R10339 VDPWR.n841 VDPWR.n772 4.51401
R10340 VDPWR.n3076 VDPWR.n3075 4.51401
R10341 VDPWR.n806 VDPWR.n804 4.51401
R10342 VDPWR.n2193 VDPWR.n2192 4.51198
R10343 VDPWR.n2277 VDPWR.n1063 4.51198
R10344 VDPWR.n537 VDPWR.n536 4.5005
R10345 VDPWR.n1534 VDPWR.n1530 4.5005
R10346 VDPWR.n1552 VDPWR.n1551 4.5005
R10347 VDPWR.n1544 VDPWR.n1536 4.5005
R10348 VDPWR.n1371 VDPWR.n1370 4.5005
R10349 VDPWR.n1382 VDPWR.n1381 4.5005
R10350 VDPWR.n1345 VDPWR.n1344 4.5005
R10351 VDPWR.n1420 VDPWR.n1419 4.5005
R10352 VDPWR.n1418 VDPWR.n1417 4.5005
R10353 VDPWR.n1336 VDPWR.n1330 4.5005
R10354 VDPWR.n1453 VDPWR.n1452 4.5005
R10355 VDPWR.n1450 VDPWR.n1449 4.5005
R10356 VDPWR.n1316 VDPWR.n1315 4.5005
R10357 VDPWR.n1489 VDPWR.n1488 4.5005
R10358 VDPWR.n1306 VDPWR.n1305 4.5005
R10359 VDPWR.n1483 VDPWR.n1299 4.5005
R10360 VDPWR.n1585 VDPWR.n1584 4.5005
R10361 VDPWR.n1583 VDPWR.n1582 4.5005
R10362 VDPWR.n1579 VDPWR.n1578 4.5005
R10363 VDPWR.n1890 VDPWR.n1889 4.5005
R10364 VDPWR.n1891 VDPWR.n1197 4.5005
R10365 VDPWR.n1900 VDPWR.n1899 4.5005
R10366 VDPWR.n1711 VDPWR.n1710 4.5005
R10367 VDPWR.n1681 VDPWR.n1680 4.5005
R10368 VDPWR.n1281 VDPWR.n1280 4.5005
R10369 VDPWR.n1751 VDPWR.n1750 4.5005
R10370 VDPWR.n1749 VDPWR.n1748 4.5005
R10371 VDPWR.n1272 VDPWR.n1265 4.5005
R10372 VDPWR.n1781 VDPWR.n1780 4.5005
R10373 VDPWR.n1254 VDPWR.n1253 4.5005
R10374 VDPWR.n1251 VDPWR.n1243 4.5005
R10375 VDPWR.n1817 VDPWR.n1816 4.5005
R10376 VDPWR.n1234 VDPWR.n1233 4.5005
R10377 VDPWR.n1811 VDPWR.n1226 4.5005
R10378 VDPWR.n1855 VDPWR.n1854 4.5005
R10379 VDPWR.n1853 VDPWR.n1852 4.5005
R10380 VDPWR.n1863 VDPWR.n1862 4.5005
R10381 VDPWR.n1933 VDPWR.n1930 4.5005
R10382 VDPWR.n1951 VDPWR.n1950 4.5005
R10383 VDPWR.n1943 VDPWR.n1935 4.5005
R10384 VDPWR.n1669 VDPWR.n1668 4.5005
R10385 VDPWR.n1658 VDPWR.n1600 4.5005
R10386 VDPWR.n1663 VDPWR.n1662 4.5005
R10387 VDPWR.n2069 VDPWR.n2068 4.5005
R10388 VDPWR.n2067 VDPWR.n2066 4.5005
R10389 VDPWR.n2063 VDPWR.n2062 4.5005
R10390 VDPWR.n1143 VDPWR.n1136 4.5005
R10391 VDPWR.n1146 VDPWR.n1145 4.5005
R10392 VDPWR.n1144 VDPWR.n1139 4.5005
R10393 VDPWR.n1160 VDPWR.n1159 4.5005
R10394 VDPWR.n1173 VDPWR.n1172 4.5005
R10395 VDPWR.n1174 VDPWR.n1164 4.5005
R10396 VDPWR.n1979 VDPWR.n1978 4.5005
R10397 VDPWR.n1911 VDPWR.n1189 4.5005
R10398 VDPWR.n1913 VDPWR.n1910 4.5005
R10399 VDPWR.n2262 VDPWR.n2261 4.5005
R10400 VDPWR.n1083 VDPWR.n1079 4.5005
R10401 VDPWR.n1085 VDPWR.n1082 4.5005
R10402 VDPWR.n2110 VDPWR.n2089 4.5005
R10403 VDPWR.n2122 VDPWR.n2121 4.5005
R10404 VDPWR.n2086 VDPWR.n2085 4.5005
R10405 VDPWR.n2156 VDPWR.n2155 4.5005
R10406 VDPWR.n2154 VDPWR.n2153 4.5005
R10407 VDPWR.n2163 VDPWR.n2162 4.5005
R10408 VDPWR.n2246 VDPWR.n2245 4.5005
R10409 VDPWR.n2235 VDPWR.n1097 4.5005
R10410 VDPWR.n2238 VDPWR.n2197 4.5005
R10411 VDPWR.n2328 VDPWR.n2327 4.5005
R10412 VDPWR.n1021 VDPWR.n1017 4.5005
R10413 VDPWR.n2322 VDPWR.n2321 4.5005
R10414 VDPWR.n2295 VDPWR.n2294 4.5005
R10415 VDPWR.n1044 VDPWR.n1042 4.5005
R10416 VDPWR.n1054 VDPWR.n1048 4.5005
R10417 VDPWR.n2967 VDPWR.n2966 4.5005
R10418 VDPWR.n2968 VDPWR.n927 4.5005
R10419 VDPWR.n2977 VDPWR.n2976 4.5005
R10420 VDPWR.n2752 VDPWR.n2751 4.5005
R10421 VDPWR.n2725 VDPWR.n2724 4.5005
R10422 VDPWR.n2747 VDPWR.n1007 4.5005
R10423 VDPWR.n2802 VDPWR.n2801 4.5005
R10424 VDPWR.n2800 VDPWR.n2799 4.5005
R10425 VDPWR.n994 VDPWR.n986 4.5005
R10426 VDPWR.n2841 VDPWR.n2840 4.5005
R10427 VDPWR.n977 VDPWR.n970 4.5005
R10428 VDPWR.n2848 VDPWR.n2847 4.5005
R10429 VDPWR.n2878 VDPWR.n2877 4.5005
R10430 VDPWR.n2894 VDPWR.n2893 4.5005
R10431 VDPWR.n960 VDPWR.n956 4.5005
R10432 VDPWR.n2929 VDPWR.n2928 4.5005
R10433 VDPWR.n2927 VDPWR.n2926 4.5005
R10434 VDPWR.n941 VDPWR.n940 4.5005
R10435 VDPWR.n2571 VDPWR.n2570 4.5005
R10436 VDPWR.n2576 VDPWR.n2575 4.5005
R10437 VDPWR.n2543 VDPWR.n2542 4.5005
R10438 VDPWR.n2598 VDPWR.n2589 4.5005
R10439 VDPWR.n2600 VDPWR.n2599 4.5005
R10440 VDPWR.n2601 VDPWR.n2592 4.5005
R10441 VDPWR.n2650 VDPWR.n2615 4.5005
R10442 VDPWR.n2653 VDPWR.n2652 4.5005
R10443 VDPWR.n2654 VDPWR.n2618 4.5005
R10444 VDPWR.n3064 VDPWR.n3063 4.5005
R10445 VDPWR.n881 VDPWR.n877 4.5005
R10446 VDPWR.n3058 VDPWR.n3057 4.5005
R10447 VDPWR.n3037 VDPWR.n3036 4.5005
R10448 VDPWR.n904 VDPWR.n902 4.5005
R10449 VDPWR.n909 VDPWR.n906 4.5005
R10450 VDPWR.n2992 VDPWR.n922 4.5005
R10451 VDPWR.n2995 VDPWR.n2994 4.5005
R10452 VDPWR.n2986 VDPWR.n2985 4.5005
R10453 VDPWR.n846 VDPWR.n845 4.5005
R10454 VDPWR.n829 VDPWR.n828 4.5005
R10455 VDPWR.n840 VDPWR.n839 4.5005
R10456 VDPWR.n2390 VDPWR.n2389 4.5005
R10457 VDPWR.n2363 VDPWR.n2360 4.5005
R10458 VDPWR.n2395 VDPWR.n2394 4.5005
R10459 VDPWR.n2427 VDPWR.n2426 4.5005
R10460 VDPWR.n2428 VDPWR.n2345 4.5005
R10461 VDPWR.n2534 VDPWR.n2533 4.5005
R10462 VDPWR.n2447 VDPWR.n2444 4.5005
R10463 VDPWR.n2497 VDPWR.n2496 4.5005
R10464 VDPWR.n2495 VDPWR.n2494 4.5005
R10465 VDPWR.n2466 VDPWR.n2465 4.5005
R10466 VDPWR.n2467 VDPWR.n786 4.5005
R10467 VDPWR.n3100 VDPWR.n3099 4.5005
R10468 VDPWR.n809 VDPWR.n802 4.5005
R10469 VDPWR.n810 VDPWR.n805 4.5005
R10470 VDPWR.n868 VDPWR.n867 4.5005
R10471 VDPWR.n2048 VDPWR.n1130 4.49637
R10472 VDPWR.n2243 VDPWR.n2194 4.40706
R10473 VDPWR.n2298 VDPWR.n1039 4.40706
R10474 VDPWR.n759 VDPWR.n758 4.38372
R10475 VDPWR.n601 VDPWR.n600 4.36875
R10476 VDPWR.n625 VDPWR.n624 4.36875
R10477 VDPWR.n584 VDPWR.n583 4.36875
R10478 VDPWR.n554 VDPWR.n553 4.36875
R10479 VDPWR.n321 VDPWR.n320 4.36875
R10480 VDPWR.n345 VDPWR.n344 4.36875
R10481 VDPWR.n304 VDPWR.n303 4.36875
R10482 VDPWR.n274 VDPWR.n273 4.36875
R10483 VDPWR.n1958 VDPWR.n1928 4.36875
R10484 VDPWR.n2180 VDPWR.n2179 4.36875
R10485 VDPWR.n2762 VDPWR.n2761 4.36875
R10486 VDPWR.n3015 VDPWR.n917 4.36875
R10487 VDPWR.n2987 VDPWR.n920 4.36875
R10488 VDPWR.n2411 VDPWR.n2351 4.36875
R10489 VDPWR.n2418 VDPWR.n2417 4.36875
R10490 VDPWR.n2401 VDPWR.n2357 4.36875
R10491 VDPWR.n2525 VDPWR.n2524 4.36875
R10492 VDPWR.n2521 VDPWR.n2434 4.36875
R10493 VDPWR.n2518 VDPWR.n2437 4.36875
R10494 VDPWR.n3092 VDPWR.n792 4.36875
R10495 VDPWR.n864 VDPWR.n863 4.36875
R10496 VDPWR.n830 VDPWR.n826 4.36875
R10497 VDPWR.n63 VDPWR.n62 4.36875
R10498 VDPWR.n87 VDPWR.n86 4.36875
R10499 VDPWR.n46 VDPWR.n45 4.36875
R10500 VDPWR.n16 VDPWR.n15 4.36875
R10501 VDPWR.n2405 VDPWR 4.3525
R10502 VDPWR.n1835 VDPWR.n1221 4.33769
R10503 VDPWR.n2093 VDPWR.n2092 4.29023
R10504 VDPWR.n2890 VDPWR.n2889 4.26717
R10505 VDPWR.n1968 VDPWR.n1966 4.14168
R10506 VDPWR.n3172 VDPWR.n3171 4.06613
R10507 VDPWR.n720 VDPWR.n719 4.05291
R10508 VDPWR.n1434 VDPWR.n1326 4.02033
R10509 VDPWR.n1357 VDPWR.n1353 4.02033
R10510 VDPWR.n1357 VDPWR.n1356 4.02033
R10511 VDPWR.n1366 VDPWR.n1360 4.02033
R10512 VDPWR.n1366 VDPWR.n1365 4.02033
R10513 VDPWR.n1549 VDPWR.n1540 4.02033
R10514 VDPWR.n1549 VDPWR.n1543 4.02033
R10515 VDPWR.n1690 VDPWR.n1686 4.02033
R10516 VDPWR.n1690 VDPWR.n1689 4.02033
R10517 VDPWR.n1699 VDPWR.n1693 4.02033
R10518 VDPWR.n1699 VDPWR.n1698 4.02033
R10519 VDPWR.n1896 VDPWR.n1208 4.02033
R10520 VDPWR.n1896 VDPWR.n1895 4.02033
R10521 VDPWR.n2048 VDPWR.n1128 4.02033
R10522 VDPWR.n1621 VDPWR.n1606 4.02033
R10523 VDPWR.n1621 VDPWR.n1612 4.02033
R10524 VDPWR.n1620 VDPWR.n1615 4.02033
R10525 VDPWR.n1620 VDPWR.n1619 4.02033
R10526 VDPWR.n1948 VDPWR.n1939 4.02033
R10527 VDPWR.n1948 VDPWR.n1942 4.02033
R10528 VDPWR.n2102 VDPWR.n2098 4.02033
R10529 VDPWR.n2102 VDPWR.n2101 4.02033
R10530 VDPWR.n1075 VDPWR.n1071 4.02033
R10531 VDPWR.n1075 VDPWR.n1074 4.02033
R10532 VDPWR.n2735 VDPWR.n2731 4.02033
R10533 VDPWR.n2735 VDPWR.n2734 4.02033
R10534 VDPWR.n2973 VDPWR.n932 4.02033
R10535 VDPWR.n2973 VDPWR.n2972 4.02033
R10536 VDPWR.n2556 VDPWR.n2552 4.02033
R10537 VDPWR.n2556 VDPWR.n2555 4.02033
R10538 VDPWR.n2687 VDPWR.n2597 4.02033
R10539 VDPWR.n3052 VDPWR.n891 4.02033
R10540 VDPWR.n3000 VDPWR.n2991 4.02033
R10541 VDPWR.n3000 VDPWR.n2999 4.02033
R10542 VDPWR.n2377 VDPWR.n2373 4.02033
R10543 VDPWR.n2377 VDPWR.n2376 4.02033
R10544 VDPWR.n843 VDPWR.n834 4.02033
R10545 VDPWR.n843 VDPWR.n838 4.02033
R10546 VDPWR.n2242 VDPWR.n2196 3.98739
R10547 VDPWR.n2297 VDPWR.n1041 3.98739
R10548 VDPWR.n1848 VDPWR.n1213 3.91455
R10549 VDPWR.n2519 VDPWR.n2518 3.86082
R10550 VDPWR.n1767 VDPWR.n1766 3.78037
R10551 VDPWR.n1796 VDPWR.n1795 3.78037
R10552 VDPWR.n1761 VDPWR.n1261 3.75517
R10553 VDPWR.n1828 VDPWR.n1827 3.75222
R10554 VDPWR.n1795 VDPWR.n1239 3.69446
R10555 VDPWR.n2475 VDPWR.n2459 3.66983
R10556 VDPWR.n724 VDPWR.t824 3.61217
R10557 VDPWR.n724 VDPWR.t820 3.61217
R10558 VDPWR.n726 VDPWR.t253 3.61217
R10559 VDPWR.n726 VDPWR.t342 3.61217
R10560 VDPWR.n722 VDPWR.t822 3.61217
R10561 VDPWR.n722 VDPWR.t219 3.61217
R10562 VDPWR.n2421 VDPWR.n2420 3.55606
R10563 VDPWR.n2092 VDPWR.n2091 3.53179
R10564 VDPWR.n2836 VDPWR.n969 3.4812
R10565 VDPWR.n1379 VDPWR.n1378 3.47425
R10566 VDPWR.n1390 VDPWR.n1389 3.47425
R10567 VDPWR.n1392 VDPWR.n1390 3.47425
R10568 VDPWR.n1511 VDPWR.n1294 3.47425
R10569 VDPWR.n1512 VDPWR.n1511 3.47425
R10570 VDPWR.n1513 VDPWR.n1512 3.47425
R10571 VDPWR.n1708 VDPWR.n1707 3.47425
R10572 VDPWR.n1720 VDPWR.n1719 3.47425
R10573 VDPWR.n1722 VDPWR.n1720 3.47425
R10574 VDPWR.n1997 VDPWR.n1996 3.47425
R10575 VDPWR.n2046 VDPWR.n2045 3.47425
R10576 VDPWR.n2045 VDPWR.n1131 3.47425
R10577 VDPWR.n1666 VDPWR.n1665 3.47425
R10578 VDPWR.n1655 VDPWR.n1654 3.47425
R10579 VDPWR.n1654 VDPWR.n1653 3.47425
R10580 VDPWR.n2129 VDPWR.n2084 3.47425
R10581 VDPWR.n2130 VDPWR.n2129 3.47425
R10582 VDPWR.n2131 VDPWR.n2130 3.47425
R10583 VDPWR.n2325 VDPWR.n2324 3.47425
R10584 VDPWR.n2267 VDPWR.n2266 3.47425
R10585 VDPWR.n2957 VDPWR.n934 3.47425
R10586 VDPWR.n2958 VDPWR.n2957 3.47425
R10587 VDPWR.n2960 VDPWR.n2958 3.47425
R10588 VDPWR.n2490 VDPWR.n2454 3.47425
R10589 VDPWR.n3178 VDPWR.n3177 3.44037
R10590 VDPWR.n2691 VDPWR.n2690 3.43925
R10591 VDPWR.n2695 VDPWR.n2694 3.43925
R10592 VDPWR.n2661 VDPWR.n2660 3.43925
R10593 VDPWR.n2665 VDPWR.n2664 3.43925
R10594 VDPWR.n1494 VDPWR.n1493 3.43925
R10595 VDPWR.n1491 VDPWR.n1490 3.43925
R10596 VDPWR.n1458 VDPWR.n1457 3.43925
R10597 VDPWR.n1455 VDPWR.n1454 3.43925
R10598 VDPWR.n1425 VDPWR.n1424 3.43925
R10599 VDPWR.n1422 VDPWR.n1421 3.43925
R10600 VDPWR.n1386 VDPWR.n1385 3.43925
R10601 VDPWR.n1373 VDPWR.n1372 3.43925
R10602 VDPWR.n1546 VDPWR.n1545 3.43925
R10603 VDPWR.n1556 VDPWR.n1555 3.43925
R10604 VDPWR.n1290 VDPWR.n1285 3.43925
R10605 VDPWR.n1587 VDPWR.n1586 3.43925
R10606 VDPWR.n1822 VDPWR.n1821 3.43925
R10607 VDPWR.n1819 VDPWR.n1818 3.43925
R10608 VDPWR.n1786 VDPWR.n1785 3.43925
R10609 VDPWR.n1783 VDPWR.n1782 3.43925
R10610 VDPWR.n1756 VDPWR.n1755 3.43925
R10611 VDPWR.n1753 VDPWR.n1752 3.43925
R10612 VDPWR.n1716 VDPWR.n1715 3.43925
R10613 VDPWR.n1713 VDPWR.n1712 3.43925
R10614 VDPWR.n1903 VDPWR.n1195 3.43925
R10615 VDPWR.n1887 VDPWR.n1194 3.43925
R10616 VDPWR.n1861 VDPWR.n1860 3.43925
R10617 VDPWR.n1857 VDPWR.n1856 3.43925
R10618 VDPWR.n2005 VDPWR.n2004 3.43925
R10619 VDPWR.n2008 VDPWR.n2007 3.43925
R10620 VDPWR.n2033 VDPWR.n2032 3.43925
R10621 VDPWR.n2037 VDPWR.n2036 3.43925
R10622 VDPWR.n1123 VDPWR.n1117 3.43925
R10623 VDPWR.n2071 VDPWR.n2070 3.43925
R10624 VDPWR.n1661 VDPWR.n1595 3.43925
R10625 VDPWR.n1671 VDPWR.n1670 3.43925
R10626 VDPWR.n1945 VDPWR.n1944 3.43925
R10627 VDPWR.n1955 VDPWR.n1954 3.43925
R10628 VDPWR.n1973 VDPWR.n1972 3.43925
R10629 VDPWR.n1975 VDPWR.n1188 3.43925
R10630 VDPWR.n2320 VDPWR.n1013 3.43925
R10631 VDPWR.n2330 VDPWR.n2329 3.43925
R10632 VDPWR.n2239 VDPWR.n1092 3.43925
R10633 VDPWR.n2248 VDPWR.n2247 3.43925
R10634 VDPWR.n2161 VDPWR.n2160 3.43925
R10635 VDPWR.n2158 VDPWR.n2157 3.43925
R10636 VDPWR.n2126 VDPWR.n2125 3.43925
R10637 VDPWR.n2112 VDPWR.n2111 3.43925
R10638 VDPWR.n2257 VDPWR.n1088 3.43925
R10639 VDPWR.n1080 VDPWR.n1078 3.43925
R10640 VDPWR.n2289 VDPWR.n2288 3.43925
R10641 VDPWR.n2291 VDPWR.n1043 3.43925
R10642 VDPWR.n2898 VDPWR.n2897 3.43925
R10643 VDPWR.n2880 VDPWR.n2879 3.43925
R10644 VDPWR.n2846 VDPWR.n2845 3.43925
R10645 VDPWR.n2843 VDPWR.n2842 3.43925
R10646 VDPWR.n2807 VDPWR.n2806 3.43925
R10647 VDPWR.n2804 VDPWR.n2803 3.43925
R10648 VDPWR.n2757 VDPWR.n2756 3.43925
R10649 VDPWR.n2754 VDPWR.n2753 3.43925
R10650 VDPWR.n2980 VDPWR.n925 3.43925
R10651 VDPWR.n2964 VDPWR.n924 3.43925
R10652 VDPWR.n2934 VDPWR.n2933 3.43925
R10653 VDPWR.n2931 VDPWR.n2930 3.43925
R10654 VDPWR.n3031 VDPWR.n3030 3.43925
R10655 VDPWR.n3033 VDPWR.n903 3.43925
R10656 VDPWR.n3056 VDPWR.n873 3.43925
R10657 VDPWR.n3066 VDPWR.n3065 3.43925
R10658 VDPWR.n3004 VDPWR.n3003 3.43925
R10659 VDPWR.n3008 VDPWR.n3007 3.43925
R10660 VDPWR.n2491 VDPWR.n2490 3.43649
R10661 VDPWR.n656 VDPWR.n655 3.4105
R10662 VDPWR.n2693 VDPWR.n2590 3.4105
R10663 VDPWR.n2692 VDPWR.n2591 3.4105
R10664 VDPWR.n2663 VDPWR.n2616 3.4105
R10665 VDPWR.n2662 VDPWR.n2617 3.4105
R10666 VDPWR.n1303 VDPWR.n1301 3.4105
R10667 VDPWR.n1304 VDPWR.n1300 3.4105
R10668 VDPWR.n1320 VDPWR.n1318 3.4105
R10669 VDPWR.n1448 VDPWR.n1317 3.4105
R10670 VDPWR.n1334 VDPWR.n1332 3.4105
R10671 VDPWR.n1416 VDPWR.n1331 3.4105
R10672 VDPWR.n1347 VDPWR.n1346 3.4105
R10673 VDPWR.n1384 VDPWR.n1383 3.4105
R10674 VDPWR.n1554 VDPWR.n1553 3.4105
R10675 VDPWR.n1533 VDPWR.n1532 3.4105
R10676 VDPWR.n1288 VDPWR.n1286 3.4105
R10677 VDPWR.n1581 VDPWR.n1580 3.4105
R10678 VDPWR.n1231 VDPWR.n1229 3.4105
R10679 VDPWR.n1232 VDPWR.n1227 3.4105
R10680 VDPWR.n1249 VDPWR.n1247 3.4105
R10681 VDPWR.n1252 VDPWR.n1244 3.4105
R10682 VDPWR.n1270 VDPWR.n1268 3.4105
R10683 VDPWR.n1747 VDPWR.n1266 3.4105
R10684 VDPWR.n1678 VDPWR.n1676 3.4105
R10685 VDPWR.n1679 VDPWR.n1282 3.4105
R10686 VDPWR.n1888 VDPWR.n1196 3.4105
R10687 VDPWR.n1902 VDPWR.n1901 3.4105
R10688 VDPWR.n1858 VDPWR.n1216 3.4105
R10689 VDPWR.n1859 VDPWR.n1215 3.4105
R10690 VDPWR.n1170 VDPWR.n1161 3.4105
R10691 VDPWR.n1171 VDPWR.n1163 3.4105
R10692 VDPWR.n2035 VDPWR.n1137 3.4105
R10693 VDPWR.n2034 VDPWR.n1138 3.4105
R10694 VDPWR.n1120 VDPWR.n1118 3.4105
R10695 VDPWR.n2065 VDPWR.n2064 3.4105
R10696 VDPWR.n1599 VDPWR.n1597 3.4105
R10697 VDPWR.n1660 VDPWR.n1659 3.4105
R10698 VDPWR.n1953 VDPWR.n1952 3.4105
R10699 VDPWR.n1932 VDPWR.n1931 3.4105
R10700 VDPWR.n1977 VDPWR.n1976 3.4105
R10701 VDPWR.n1909 VDPWR.n1190 3.4105
R10702 VDPWR.n1016 VDPWR.n1014 3.4105
R10703 VDPWR.n1023 VDPWR.n1022 3.4105
R10704 VDPWR.n1095 VDPWR.n1093 3.4105
R10705 VDPWR.n2237 VDPWR.n2236 3.4105
R10706 VDPWR.n2076 VDPWR.n2074 3.4105
R10707 VDPWR.n1115 VDPWR.n1114 3.4105
R10708 VDPWR.n2088 VDPWR.n2087 3.4105
R10709 VDPWR.n2124 VDPWR.n2123 3.4105
R10710 VDPWR.n2260 VDPWR.n2259 3.4105
R10711 VDPWR.n2258 VDPWR.n1081 3.4105
R10712 VDPWR.n2293 VDPWR.n2292 3.4105
R10713 VDPWR.n1047 VDPWR.n1045 3.4105
R10714 VDPWR.n958 VDPWR.n957 3.4105
R10715 VDPWR.n2896 VDPWR.n2895 3.4105
R10716 VDPWR.n978 VDPWR.n975 3.4105
R10717 VDPWR.n972 VDPWR.n971 3.4105
R10718 VDPWR.n992 VDPWR.n990 3.4105
R10719 VDPWR.n2798 VDPWR.n987 3.4105
R10720 VDPWR.n2722 VDPWR.n2720 3.4105
R10721 VDPWR.n2723 VDPWR.n1008 3.4105
R10722 VDPWR.n2965 VDPWR.n926 3.4105
R10723 VDPWR.n2979 VDPWR.n2978 3.4105
R10724 VDPWR.n946 VDPWR.n944 3.4105
R10725 VDPWR.n2925 VDPWR.n942 3.4105
R10726 VDPWR.n3035 VDPWR.n3034 3.4105
R10727 VDPWR.n3032 VDPWR.n905 3.4105
R10728 VDPWR.n876 VDPWR.n874 3.4105
R10729 VDPWR.n883 VDPWR.n882 3.4105
R10730 VDPWR.n3102 VDPWR.n784 3.4105
R10731 VDPWR.n3102 VDPWR.n785 3.4105
R10732 VDPWR.n3102 VDPWR.n783 3.4105
R10733 VDPWR.n3102 VDPWR.n3101 3.4105
R10734 VDPWR.n2508 VDPWR.n2446 3.4105
R10735 VDPWR.n2509 VDPWR.n2508 3.4105
R10736 VDPWR.n2508 VDPWR.n2498 3.4105
R10737 VDPWR.n2508 VDPWR.n2445 3.4105
R10738 VDPWR.n2719 VDPWR.n2718 3.4105
R10739 VDPWR.n2719 VDPWR.n2338 3.4105
R10740 VDPWR.n2718 VDPWR.n2717 3.4105
R10741 VDPWR.n2549 VDPWR.n2338 3.4105
R10742 VDPWR.n2573 VDPWR.n2572 3.4105
R10743 VDPWR.n2574 VDPWR.n2541 3.4105
R10744 VDPWR.n3006 VDPWR.n2983 3.4105
R10745 VDPWR.n3005 VDPWR.n2984 3.4105
R10746 VDPWR.n2536 VDPWR.n2342 3.4105
R10747 VDPWR.n2536 VDPWR.n2344 3.4105
R10748 VDPWR.n2536 VDPWR.n2341 3.4105
R10749 VDPWR.n2536 VDPWR.n2535 3.4105
R10750 VDPWR.n2393 VDPWR.n2392 3.4105
R10751 VDPWR.n2392 VDPWR.n2391 3.4105
R10752 VDPWR.n2392 VDPWR.n2364 3.4105
R10753 VDPWR.n2392 VDPWR.n2362 3.4105
R10754 VDPWR.n3074 VDPWR.n804 3.4105
R10755 VDPWR.n3075 VDPWR.n3074 3.4105
R10756 VDPWR.n3074 VDPWR.n803 3.4105
R10757 VDPWR.n3074 VDPWR.n869 3.4105
R10758 VDPWR.n3113 VDPWR.n771 3.4105
R10759 VDPWR.n847 VDPWR.n771 3.4105
R10760 VDPWR.n3114 VDPWR.n773 3.4105
R10761 VDPWR.n3114 VDPWR.n774 3.4105
R10762 VDPWR.n3114 VDPWR.n772 3.4105
R10763 VDPWR.t186 VDPWR.t788 3.35739
R10764 VDPWR.t964 VDPWR.t1162 3.35739
R10765 VDPWR.t176 VDPWR.t108 3.35739
R10766 VDPWR.t188 VDPWR.t72 3.35739
R10767 VDPWR.t906 VDPWR.t940 3.35739
R10768 VDPWR.t0 VDPWR.t46 3.35739
R10769 VDPWR.t385 VDPWR.t1122 3.35739
R10770 VDPWR.t833 VDPWR.t637 3.35739
R10771 VDPWR.t880 VDPWR.t112 3.35739
R10772 VDPWR.t216 VDPWR.t304 3.35739
R10773 VDPWR.n1376 VDPWR.n1350 3.2477
R10774 VDPWR.n1392 VDPWR.n1391 3.2477
R10775 VDPWR.n1504 VDPWR.n1503 3.2477
R10776 VDPWR.n1513 VDPWR.n1292 3.2477
R10777 VDPWR.n1704 VDPWR.n1683 3.2477
R10778 VDPWR.n1722 VDPWR.n1721 3.2477
R10779 VDPWR.n1996 VDPWR.n1995 3.2477
R10780 VDPWR.n2047 VDPWR.n2046 3.2477
R10781 VDPWR.n1602 VDPWR.n1601 3.2477
R10782 VDPWR.n1653 VDPWR.n1627 3.2477
R10783 VDPWR.n2115 VDPWR.n2090 3.2477
R10784 VDPWR.n2131 VDPWR.n2082 3.2477
R10785 VDPWR.n2324 VDPWR.n1019 3.2477
R10786 VDPWR.n2266 VDPWR.n2265 3.2477
R10787 VDPWR.n2952 VDPWR.n934 3.2477
R10788 VDPWR.n2960 VDPWR.n2959 3.2477
R10789 VDPWR.n2492 VDPWR.n2450 3.2477
R10790 VDPWR.n2486 VDPWR.n2485 3.2477
R10791 VDPWR.n478 VDPWR.n467 3.24308
R10792 VDPWR.n3129 VDPWR.n3118 3.24308
R10793 VDPWR.n691 VDPWR.n688 3.23917
R10794 VDPWR.n502 VDPWR.n499 3.23917
R10795 VDPWR.n448 VDPWR.n445 3.23917
R10796 VDPWR.n3153 VDPWR.n3150 3.23917
R10797 VDPWR.n675 VDPWR.n672 3.23136
R10798 VDPWR.n486 VDPWR.n483 3.23136
R10799 VDPWR.n432 VDPWR.n429 3.23136
R10800 VDPWR.n3137 VDPWR.n3134 3.23136
R10801 VDPWR.n462 VDPWR.n461 3.22655
R10802 VDPWR.n715 VDPWR.n704 3.22655
R10803 VDPWR.n526 VDPWR.n515 3.22655
R10804 VDPWR.n3167 VDPWR.n3166 3.22655
R10805 VDPWR.n2760 VDPWR.n1006 3.2005
R10806 VDPWR.n1258 VDPWR.n1257 3.151
R10807 VDPWR.n2191 VDPWR.n1100 3.14804
R10808 VDPWR.n2303 VDPWR.n2302 3.14804
R10809 VDPWR.n859 VDPWR.n819 3.12116
R10810 VDPWR.n1361 VDPWR.n1357 3.05586
R10811 VDPWR.n1694 VDPWR.n1690 3.05586
R10812 VDPWR.n1620 VDPWR.n1616 3.05586
R10813 VDPWR.n2103 VDPWR.n2102 3.05586
R10814 VDPWR.n2736 VDPWR.n2735 3.05586
R10815 VDPWR.n2560 VDPWR.n2556 3.05586
R10816 VDPWR.n2378 VDPWR.n2377 3.05586
R10817 VDPWR.n1366 VDPWR.n1362 3.04861
R10818 VDPWR.n1699 VDPWR.n1695 3.04861
R10819 VDPWR.n1884 VDPWR.n1205 3.04861
R10820 VDPWR.n1621 VDPWR.n1609 3.04861
R10821 VDPWR.n3052 VDPWR.n888 3.04861
R10822 VDPWR.n1434 VDPWR.n1433 3.04861
R10823 VDPWR.n1833 VDPWR.n1832 3.04861
R10824 VDPWR.n2055 VDPWR.n1128 3.04861
R10825 VDPWR.n1964 VDPWR.n1922 3.04861
R10826 VDPWR.n2749 VDPWR.n2746 3.04861
R10827 VDPWR.n854 VDPWR.n822 3.04861
R10828 VDPWR.n1441 VDPWR.n1440 3.01588
R10829 VDPWR.n1471 VDPWR.n1309 3.01588
R10830 VDPWR.n1411 VDPWR.n1410 3.01588
R10831 VDPWR.n1570 VDPWR.n1524 3.01588
R10832 VDPWR.n1741 VDPWR.n1740 3.01588
R10833 VDPWR.n1771 VDPWR.n1770 3.01588
R10834 VDPWR.n1776 VDPWR.n1775 3.01588
R10835 VDPWR.n1799 VDPWR.n1237 3.01588
R10836 VDPWR.n1804 VDPWR.n1803 3.01588
R10837 VDPWR.n2011 VDPWR.n1158 3.01588
R10838 VDPWR.n2020 VDPWR.n1154 3.01588
R10839 VDPWR.n1150 VDPWR.n1149 3.01588
R10840 VDPWR.n1634 VDPWR.n1633 3.01588
R10841 VDPWR.n2147 VDPWR.n2077 3.01588
R10842 VDPWR.n1875 VDPWR.n1209 3.01226
R10843 VDPWR.n2867 VDPWR.n2866 3.01226
R10844 VDPWR.n2608 VDPWR.n2605 3.01226
R10845 VDPWR.n2566 VDPWR.n2547 3.01226
R10846 VDPWR.n894 VDPWR.n892 3.01226
R10847 VDPWR.n3044 VDPWR.n897 3.01226
R10848 VDPWR.n1961 VDPWR.n1926 2.99733
R10849 VDPWR.n852 VDPWR.n824 2.99733
R10850 VDPWR.n1205 VDPWR.n1201 2.91308
R10851 VDPWR.n1205 VDPWR.n1204 2.91308
R10852 VDPWR.n2565 VDPWR.n2559 2.91308
R10853 VDPWR.n2565 VDPWR.n2564 2.91308
R10854 VDPWR.n1924 VDPWR.n1922 2.87861
R10855 VDPWR.n2210 VDPWR.n2209 2.8567
R10856 VDPWR.n709 VDPWR.n708 2.84665
R10857 VDPWR.n712 VDPWR.n708 2.84665
R10858 VDPWR.n707 VDPWR.n706 2.84665
R10859 VDPWR.n712 VDPWR.n707 2.84665
R10860 VDPWR.n694 VDPWR.n693 2.84665
R10861 VDPWR.n697 VDPWR.n693 2.84665
R10862 VDPWR.n692 VDPWR.n690 2.84665
R10863 VDPWR.n697 VDPWR.n692 2.84665
R10864 VDPWR.n678 VDPWR.n677 2.84665
R10865 VDPWR.n681 VDPWR.n677 2.84665
R10866 VDPWR.n676 VDPWR.n674 2.84665
R10867 VDPWR.n681 VDPWR.n676 2.84665
R10868 VDPWR.n664 VDPWR.n663 2.84665
R10869 VDPWR.n665 VDPWR.n664 2.84665
R10870 VDPWR.n667 VDPWR.n666 2.84665
R10871 VDPWR.n666 VDPWR.n665 2.84665
R10872 VDPWR.n520 VDPWR.n519 2.84665
R10873 VDPWR.n523 VDPWR.n519 2.84665
R10874 VDPWR.n518 VDPWR.n517 2.84665
R10875 VDPWR.n523 VDPWR.n518 2.84665
R10876 VDPWR.n505 VDPWR.n504 2.84665
R10877 VDPWR.n508 VDPWR.n504 2.84665
R10878 VDPWR.n503 VDPWR.n501 2.84665
R10879 VDPWR.n508 VDPWR.n503 2.84665
R10880 VDPWR.n489 VDPWR.n488 2.84665
R10881 VDPWR.n492 VDPWR.n488 2.84665
R10882 VDPWR.n487 VDPWR.n485 2.84665
R10883 VDPWR.n492 VDPWR.n487 2.84665
R10884 VDPWR.n472 VDPWR.n471 2.84665
R10885 VDPWR.n475 VDPWR.n471 2.84665
R10886 VDPWR.n470 VDPWR.n469 2.84665
R10887 VDPWR.n475 VDPWR.n470 2.84665
R10888 VDPWR.n406 VDPWR.n405 2.84665
R10889 VDPWR.n411 VDPWR.n406 2.84665
R10890 VDPWR.n408 VDPWR.n407 2.84665
R10891 VDPWR.n411 VDPWR.n407 2.84665
R10892 VDPWR.n386 VDPWR.n385 2.84665
R10893 VDPWR.n382 VDPWR.n378 2.84665
R10894 VDPWR.n398 VDPWR.n397 2.84665
R10895 VDPWR.n394 VDPWR.n390 2.84665
R10896 VDPWR.n451 VDPWR.n450 2.84665
R10897 VDPWR.n454 VDPWR.n450 2.84665
R10898 VDPWR.n449 VDPWR.n447 2.84665
R10899 VDPWR.n454 VDPWR.n449 2.84665
R10900 VDPWR.n435 VDPWR.n434 2.84665
R10901 VDPWR.n438 VDPWR.n434 2.84665
R10902 VDPWR.n433 VDPWR.n431 2.84665
R10903 VDPWR.n438 VDPWR.n433 2.84665
R10904 VDPWR.n421 VDPWR.n420 2.84665
R10905 VDPWR.n422 VDPWR.n421 2.84665
R10906 VDPWR.n424 VDPWR.n423 2.84665
R10907 VDPWR.n423 VDPWR.n422 2.84665
R10908 VDPWR.n764 VDPWR.n763 2.84665
R10909 VDPWR.n767 VDPWR.n763 2.84665
R10910 VDPWR.n762 VDPWR.n761 2.84665
R10911 VDPWR.n767 VDPWR.n762 2.84665
R10912 VDPWR.n3154 VDPWR.n3152 2.84665
R10913 VDPWR.n3159 VDPWR.n3154 2.84665
R10914 VDPWR.n3156 VDPWR.n3155 2.84665
R10915 VDPWR.n3159 VDPWR.n3155 2.84665
R10916 VDPWR.n3138 VDPWR.n3136 2.84665
R10917 VDPWR.n3143 VDPWR.n3138 2.84665
R10918 VDPWR.n3140 VDPWR.n3139 2.84665
R10919 VDPWR.n3143 VDPWR.n3139 2.84665
R10920 VDPWR.n3123 VDPWR.n3122 2.84665
R10921 VDPWR.n3126 VDPWR.n3122 2.84665
R10922 VDPWR.n3121 VDPWR.n3120 2.84665
R10923 VDPWR.n3126 VDPWR.n3121 2.84665
R10924 VDPWR.n1260 VDPWR.n1258 2.8165
R10925 VDPWR.n2474 VDPWR.n2472 2.8165
R10926 VDPWR.n1377 VDPWR.n1349 2.6965
R10927 VDPWR.n1705 VDPWR.n1682 2.6965
R10928 VDPWR.n1624 VDPWR.n1623 2.6965
R10929 VDPWR.n3060 VDPWR.n879 2.69256
R10930 VDPWR.n1440 VDPWR.n1321 2.64665
R10931 VDPWR.n1474 VDPWR.n1309 2.64665
R10932 VDPWR.n1412 VDPWR.n1411 2.64665
R10933 VDPWR.n1567 VDPWR.n1524 2.64665
R10934 VDPWR.n1742 VDPWR.n1741 2.64665
R10935 VDPWR.n1770 VDPWR.n1255 2.64665
R10936 VDPWR.n1777 VDPWR.n1776 2.64665
R10937 VDPWR.n1802 VDPWR.n1237 2.64665
R10938 VDPWR.n1805 VDPWR.n1804 2.64665
R10939 VDPWR.n1168 VDPWR.n1158 2.64665
R10940 VDPWR.n2029 VDPWR.n1150 2.64665
R10941 VDPWR.n1633 VDPWR.n1632 2.64665
R10942 VDPWR.n2141 VDPWR.n2079 2.64665
R10943 VDPWR.n2145 VDPWR.n2079 2.64665
R10944 VDPWR.n2150 VDPWR.n2077 2.64665
R10945 VDPWR.n1987 VDPWR.n1986 2.63579
R10946 VDPWR.n1326 VDPWR.n1324 2.63539
R10947 VDPWR.n1353 VDPWR.n1351 2.63539
R10948 VDPWR.n1356 VDPWR.n1354 2.63539
R10949 VDPWR.n1360 VDPWR.n1358 2.63539
R10950 VDPWR.n1365 VDPWR.n1363 2.63539
R10951 VDPWR.n1540 VDPWR.n1538 2.63539
R10952 VDPWR.n1543 VDPWR.n1541 2.63539
R10953 VDPWR.n1686 VDPWR.n1684 2.63539
R10954 VDPWR.n1689 VDPWR.n1687 2.63539
R10955 VDPWR.n1693 VDPWR.n1691 2.63539
R10956 VDPWR.n1698 VDPWR.n1696 2.63539
R10957 VDPWR.n1208 VDPWR.n1206 2.63539
R10958 VDPWR.n1895 VDPWR.n1893 2.63539
R10959 VDPWR.n1606 VDPWR.n1604 2.63539
R10960 VDPWR.n1612 VDPWR.n1610 2.63539
R10961 VDPWR.n1615 VDPWR.n1613 2.63539
R10962 VDPWR.n1619 VDPWR.n1617 2.63539
R10963 VDPWR.n1939 VDPWR.n1937 2.63539
R10964 VDPWR.n1942 VDPWR.n1940 2.63539
R10965 VDPWR.n2098 VDPWR.n2096 2.63539
R10966 VDPWR.n2101 VDPWR.n2099 2.63539
R10967 VDPWR.n1071 VDPWR.n1069 2.63539
R10968 VDPWR.n1074 VDPWR.n1072 2.63539
R10969 VDPWR.n2731 VDPWR.n2729 2.63539
R10970 VDPWR.n2734 VDPWR.n2732 2.63539
R10971 VDPWR.n932 VDPWR.n930 2.63539
R10972 VDPWR.n2972 VDPWR.n2970 2.63539
R10973 VDPWR.n2552 VDPWR.n2550 2.63539
R10974 VDPWR.n2555 VDPWR.n2553 2.63539
R10975 VDPWR.n2597 VDPWR.n2595 2.63539
R10976 VDPWR.n891 VDPWR.n889 2.63539
R10977 VDPWR.n2991 VDPWR.n2989 2.63539
R10978 VDPWR.n2999 VDPWR.n2997 2.63539
R10979 VDPWR.n819 VDPWR.n817 2.63539
R10980 VDPWR.n2373 VDPWR.n2371 2.63539
R10981 VDPWR.n2376 VDPWR.n2374 2.63539
R10982 VDPWR.n834 VDPWR.n832 2.63539
R10983 VDPWR.n838 VDPWR.n836 2.63539
R10984 VDPWR.n2232 VDPWR.n2231 2.62345
R10985 VDPWR.n1926 VDPWR.n1925 2.61352
R10986 VDPWR.n1034 VDPWR.n1031 2.56175
R10987 VDPWR.n577 VDPWR.n576 2.54018
R10988 VDPWR.n556 VDPWR.n555 2.54018
R10989 VDPWR.n297 VDPWR.n296 2.54018
R10990 VDPWR.n276 VDPWR.n275 2.54018
R10991 VDPWR.n796 VDPWR.n793 2.54018
R10992 VDPWR.n39 VDPWR.n38 2.54018
R10993 VDPWR.n18 VDPWR.n17 2.54018
R10994 VDPWR.n3083 VDPWR.n797 2.3878
R10995 VDPWR.n824 VDPWR.n823 2.37764
R10996 VDPWR.n1325 VDPWR.n1324 2.37495
R10997 VDPWR.n1355 VDPWR.n1354 2.37495
R10998 VDPWR.n1352 VDPWR.n1351 2.37495
R10999 VDPWR.n1364 VDPWR.n1363 2.37495
R11000 VDPWR.n1359 VDPWR.n1358 2.37495
R11001 VDPWR.n1542 VDPWR.n1541 2.37495
R11002 VDPWR.n1539 VDPWR.n1538 2.37495
R11003 VDPWR.n1688 VDPWR.n1687 2.37495
R11004 VDPWR.n1685 VDPWR.n1684 2.37495
R11005 VDPWR.n1697 VDPWR.n1696 2.37495
R11006 VDPWR.n1692 VDPWR.n1691 2.37495
R11007 VDPWR.n1894 VDPWR.n1893 2.37495
R11008 VDPWR.n1207 VDPWR.n1206 2.37495
R11009 VDPWR.n1611 VDPWR.n1610 2.37495
R11010 VDPWR.n1605 VDPWR.n1604 2.37495
R11011 VDPWR.n1618 VDPWR.n1617 2.37495
R11012 VDPWR.n1614 VDPWR.n1613 2.37495
R11013 VDPWR.n1941 VDPWR.n1940 2.37495
R11014 VDPWR.n1938 VDPWR.n1937 2.37495
R11015 VDPWR.n2100 VDPWR.n2099 2.37495
R11016 VDPWR.n2097 VDPWR.n2096 2.37495
R11017 VDPWR.n1073 VDPWR.n1072 2.37495
R11018 VDPWR.n1070 VDPWR.n1069 2.37495
R11019 VDPWR.n2733 VDPWR.n2732 2.37495
R11020 VDPWR.n2730 VDPWR.n2729 2.37495
R11021 VDPWR.n2971 VDPWR.n2970 2.37495
R11022 VDPWR.n931 VDPWR.n930 2.37495
R11023 VDPWR.n2554 VDPWR.n2553 2.37495
R11024 VDPWR.n2551 VDPWR.n2550 2.37495
R11025 VDPWR.n2596 VDPWR.n2595 2.37495
R11026 VDPWR.n890 VDPWR.n889 2.37495
R11027 VDPWR.n2998 VDPWR.n2997 2.37495
R11028 VDPWR.n2990 VDPWR.n2989 2.37495
R11029 VDPWR.n818 VDPWR.n817 2.37495
R11030 VDPWR.n2375 VDPWR.n2374 2.37495
R11031 VDPWR.n2372 VDPWR.n2371 2.37495
R11032 VDPWR.n837 VDPWR.n836 2.37495
R11033 VDPWR.n833 VDPWR.n832 2.37495
R11034 VDPWR.n602 VDPWR.n598 2.33701
R11035 VDPWR.n590 VDPWR.n589 2.33701
R11036 VDPWR.n576 VDPWR.n575 2.33701
R11037 VDPWR.n556 VDPWR.n550 2.33701
R11038 VDPWR.n322 VDPWR.n318 2.33701
R11039 VDPWR.n310 VDPWR.n309 2.33701
R11040 VDPWR.n296 VDPWR.n295 2.33701
R11041 VDPWR.n276 VDPWR.n270 2.33701
R11042 VDPWR.n1105 VDPWR.n1104 2.33701
R11043 VDPWR.n2886 VDPWR.n2885 2.33701
R11044 VDPWR.n3061 VDPWR.n878 2.33701
R11045 VDPWR.n2400 VDPWR.n2399 2.33701
R11046 VDPWR.n64 VDPWR.n60 2.33701
R11047 VDPWR.n52 VDPWR.n51 2.33701
R11048 VDPWR.n38 VDPWR.n37 2.33701
R11049 VDPWR.n18 VDPWR.n12 2.33701
R11050 VDPWR.n1434 VDPWR.n1327 2.32777
R11051 VDPWR.n1128 VDPWR.n1127 2.32777
R11052 VDPWR.n1834 VDPWR.n1833 2.28432
R11053 VDPWR.n2749 VDPWR.n2726 2.28407
R11054 VDPWR.n2749 VDPWR.n2728 2.28407
R11055 VDPWR.n2094 VDPWR.n2092 2.28374
R11056 VDPWR.n1155 VDPWR.n1154 2.27742
R11057 VDPWR.n1920 VDPWR.n1919 2.25932
R11058 VDPWR.n1986 VDPWR.n1184 2.25932
R11059 VDPWR.n2565 VDPWR.n2561 2.25293
R11060 VDPWR.n3090 VDPWR.n3089 2.23542
R11061 VDPWR.n2909 VDPWR.n2908 2.22199
R11062 VDPWR.n3118 VDPWR.n3117 2.16151
R11063 VDPWR.n402 VDPWR.n401 2.13883
R11064 VDPWR.n483 VDPWR.n482 2.13544
R11065 VDPWR.n584 VDPWR.n577 2.13383
R11066 VDPWR.n555 VDPWR.n554 2.13383
R11067 VDPWR.n304 VDPWR.n297 2.13383
R11068 VDPWR.n275 VDPWR.n274 2.13383
R11069 VDPWR.n3085 VDPWR.n796 2.13383
R11070 VDPWR.n46 VDPWR.n39 2.13383
R11071 VDPWR.n17 VDPWR.n16 2.13383
R11072 VDPWR.n1057 VDPWR.n1056 2.0932
R11073 VDPWR.n2740 VDPWR.n2739 2.07374
R11074 VDPWR.n2727 VDPWR.n1006 2.07374
R11075 VDPWR.n598 VDPWR.n596 2.03225
R11076 VDPWR.n589 VDPWR.n588 2.03225
R11077 VDPWR.n575 VDPWR.n574 2.03225
R11078 VDPWR.n550 VDPWR.n548 2.03225
R11079 VDPWR.n318 VDPWR.n316 2.03225
R11080 VDPWR.n309 VDPWR.n308 2.03225
R11081 VDPWR.n295 VDPWR.n294 2.03225
R11082 VDPWR.n270 VDPWR.n268 2.03225
R11083 VDPWR.n2885 VDPWR.n2884 2.03225
R11084 VDPWR.n2399 VDPWR.n2398 2.03225
R11085 VDPWR.n60 VDPWR.n58 2.03225
R11086 VDPWR.n51 VDPWR.n50 2.03225
R11087 VDPWR.n37 VDPWR.n36 2.03225
R11088 VDPWR.n12 VDPWR.n10 2.03225
R11089 VDPWR.n1201 VDPWR.n1199 2.01703
R11090 VDPWR.n1204 VDPWR.n1202 2.01703
R11091 VDPWR.n2559 VDPWR.n2557 2.01703
R11092 VDPWR.n2564 VDPWR.n2562 2.01703
R11093 VDPWR.n3092 VDPWR.n3091 1.98145
R11094 VDPWR.n798 VDPWR.n797 1.98145
R11095 VDPWR.n482 VDPWR.n467 1.95379
R11096 VDPWR.n2187 VDPWR.n2186 1.88902
R11097 VDPWR.n2305 VDPWR.n1034 1.88902
R11098 VDPWR.n1203 VDPWR.n1202 1.88416
R11099 VDPWR.n1200 VDPWR.n1199 1.88416
R11100 VDPWR.n2563 VDPWR.n2562 1.88416
R11101 VDPWR.n2558 VDPWR.n2557 1.88416
R11102 VDPWR.n1643 VDPWR.n1630 1.88325
R11103 VDPWR.n1403 VDPWR.n1402 1.88295
R11104 VDPWR.n1733 VDPWR.n1732 1.88295
R11105 VDPWR.n661 VDPWR.n657 1.88285
R11106 VDPWR.n478 VDPWR.n477 1.88285
R11107 VDPWR.n418 VDPWR.n414 1.88285
R11108 VDPWR.n3129 VDPWR.n3128 1.88285
R11109 VDPWR.n2852 VDPWR.n967 1.88285
R11110 VDPWR.n1377 VDPWR.n1376 1.85065
R11111 VDPWR.n1379 VDPWR.n1343 1.85065
R11112 VDPWR.n1507 VDPWR.n1506 1.85065
R11113 VDPWR.n1705 VDPWR.n1704 1.85065
R11114 VDPWR.n1707 VDPWR.n1279 1.85065
R11115 VDPWR.n1132 VDPWR.n1131 1.85065
R11116 VDPWR.n1624 VDPWR.n1601 1.85065
R11117 VDPWR.n1665 VDPWR.n1625 1.85065
R11118 VDPWR.n2118 VDPWR.n2117 1.85065
R11119 VDPWR.n2456 VDPWR.n2454 1.85065
R11120 VDPWR.n2793 VDPWR.n984 1.82907
R11121 VDPWR.n2628 VDPWR.n2627 1.82907
R11122 VDPWR.n1505 VDPWR.n1504 1.81289
R11123 VDPWR.n2116 VDPWR.n2115 1.81289
R11124 VDPWR.n2483 VDPWR 1.79885
R11125 VDPWR.n654 VDPWR.n653 1.753
R11126 VDPWR.n374 VDPWR.n373 1.753
R11127 VDPWR.n116 VDPWR.n115 1.753
R11128 VDPWR.n1997 VDPWR.n1181 1.73737
R11129 VDPWR.n2325 VDPWR.n1018 1.73737
R11130 VDPWR.n2267 VDPWR.n1068 1.73737
R11131 VDPWR.n2216 VDPWR.n2210 1.69306
R11132 VDPWR.n2271 VDPWR.n1065 1.69306
R11133 VDPWR.n3031 VDPWR.n870 1.69188
R11134 VDPWR.n3033 VDPWR.n870 1.69188
R11135 VDPWR.n2933 VDPWR.n2932 1.69188
R11136 VDPWR.n2932 VDPWR.n2931 1.69188
R11137 VDPWR.n2290 VDPWR.n2289 1.69188
R11138 VDPWR.n2291 VDPWR.n2290 1.69188
R11139 VDPWR.n1974 VDPWR.n1973 1.69188
R11140 VDPWR.n1975 VDPWR.n1974 1.69188
R11141 VDPWR.n1860 VDPWR.n1191 1.69188
R11142 VDPWR.n1857 VDPWR.n1191 1.69188
R11143 VDPWR.n1588 VDPWR.n1285 1.69188
R11144 VDPWR.n1588 VDPWR.n1587 1.69188
R11145 VDPWR.n3067 VDPWR.n873 1.69188
R11146 VDPWR.n3067 VDPWR.n3066 1.69188
R11147 VDPWR.n2897 VDPWR.n872 1.69188
R11148 VDPWR.n2879 VDPWR.n872 1.69188
R11149 VDPWR.n2331 VDPWR.n1013 1.69188
R11150 VDPWR.n2331 VDPWR.n2330 1.69188
R11151 VDPWR.n2006 VDPWR.n2005 1.69188
R11152 VDPWR.n2007 VDPWR.n2006 1.69188
R11153 VDPWR.n1821 VDPWR.n1820 1.69188
R11154 VDPWR.n1820 VDPWR.n1819 1.69188
R11155 VDPWR.n1493 VDPWR.n1492 1.69188
R11156 VDPWR.n1492 VDPWR.n1491 1.69188
R11157 VDPWR.n2661 VDPWR.n974 1.69188
R11158 VDPWR.n2664 VDPWR.n974 1.69188
R11159 VDPWR.n2845 VDPWR.n2844 1.69188
R11160 VDPWR.n2844 VDPWR.n2843 1.69188
R11161 VDPWR.n2249 VDPWR.n1092 1.69188
R11162 VDPWR.n2249 VDPWR.n2248 1.69188
R11163 VDPWR.n2033 VDPWR.n1091 1.69188
R11164 VDPWR.n2036 VDPWR.n1091 1.69188
R11165 VDPWR.n1785 VDPWR.n1784 1.69188
R11166 VDPWR.n1784 VDPWR.n1783 1.69188
R11167 VDPWR.n1457 VDPWR.n1456 1.69188
R11168 VDPWR.n1456 VDPWR.n1455 1.69188
R11169 VDPWR.n2756 VDPWR.n2755 1.69188
R11170 VDPWR.n2755 VDPWR.n2754 1.69188
R11171 VDPWR.n2125 VDPWR.n1009 1.69188
R11172 VDPWR.n2111 VDPWR.n1009 1.69188
R11173 VDPWR.n1672 VDPWR.n1595 1.69188
R11174 VDPWR.n1672 VDPWR.n1671 1.69188
R11175 VDPWR.n1715 VDPWR.n1714 1.69188
R11176 VDPWR.n1714 VDPWR.n1713 1.69188
R11177 VDPWR.n1385 VDPWR.n1283 1.69188
R11178 VDPWR.n1372 VDPWR.n1283 1.69188
R11179 VDPWR.n2719 VDPWR.n2337 1.69188
R11180 VDPWR.n3007 VDPWR.n2982 1.69188
R11181 VDPWR.n3004 VDPWR.n2982 1.69188
R11182 VDPWR.n2981 VDPWR.n924 1.69188
R11183 VDPWR.n2981 VDPWR.n2980 1.69188
R11184 VDPWR.n2256 VDPWR.n1080 1.69188
R11185 VDPWR.n2257 VDPWR.n2256 1.69188
R11186 VDPWR.n1954 VDPWR.n1089 1.69188
R11187 VDPWR.n1944 VDPWR.n1089 1.69188
R11188 VDPWR.n1904 VDPWR.n1194 1.69188
R11189 VDPWR.n1904 VDPWR.n1903 1.69188
R11190 VDPWR.n1555 VDPWR.n1531 1.69188
R11191 VDPWR.n1545 VDPWR.n1531 1.69188
R11192 VDPWR.n2691 VDPWR.n989 1.69188
R11193 VDPWR.n2694 VDPWR.n989 1.69188
R11194 VDPWR.n2806 VDPWR.n2805 1.69188
R11195 VDPWR.n2805 VDPWR.n2804 1.69188
R11196 VDPWR.n2160 VDPWR.n2159 1.69188
R11197 VDPWR.n2159 VDPWR.n2158 1.69188
R11198 VDPWR.n2072 VDPWR.n1117 1.69188
R11199 VDPWR.n2072 VDPWR.n2071 1.69188
R11200 VDPWR.n1755 VDPWR.n1754 1.69188
R11201 VDPWR.n1754 VDPWR.n1753 1.69188
R11202 VDPWR.n1424 VDPWR.n1423 1.69188
R11203 VDPWR.n1423 VDPWR.n1422 1.69188
R11204 VDPWR.t996 VDPWR 1.67895
R11205 VDPWR.t126 VDPWR 1.67895
R11206 VDPWR.n884 VDPWR.n879 1.67669
R11207 VDPWR.n1507 VDPWR.n1505 1.66186
R11208 VDPWR.n2118 VDPWR.n2116 1.66186
R11209 VDPWR.n2491 VDPWR.n2453 1.64857
R11210 VDPWR.n1378 VDPWR.n1377 1.6241
R11211 VDPWR.n1389 VDPWR.n1343 1.6241
R11212 VDPWR.n1506 VDPWR.n1294 1.6241
R11213 VDPWR.n1708 VDPWR.n1705 1.6241
R11214 VDPWR.n1719 VDPWR.n1279 1.6241
R11215 VDPWR.n1666 VDPWR.n1624 1.6241
R11216 VDPWR.n1655 VDPWR.n1625 1.6241
R11217 VDPWR.n2117 VDPWR.n2084 1.6241
R11218 VDPWR.n2486 VDPWR.n2456 1.6241
R11219 VDPWR.n1404 VDPWR.n1403 1.62167
R11220 VDPWR.n1734 VDPWR.n1733 1.62167
R11221 VDPWR.n1640 VDPWR.n1630 1.62136
R11222 VDPWR.n3172 VDPWR.n117 1.59405
R11223 VDPWR.n754 VDPWR.n753 1.57294
R11224 VDPWR.n747 VDPWR.t372 1.53603
R11225 VDPWR.n744 VDPWR.t372 1.53603
R11226 VDPWR.n531 VDPWR.n530 1.51493
R11227 VDPWR.n1181 VDPWR.n1179 1.51082
R11228 VDPWR.n2211 VDPWR.n1018 1.51082
R11229 VDPWR.n1068 VDPWR.n1066 1.51082
R11230 VDPWR.n758 VDPWR 1.48239
R11231 VDPWR.n573 VDPWR.n571 1.46504
R11232 VDPWR.n293 VDPWR.n291 1.46504
R11233 VDPWR.n35 VDPWR.n33 1.46504
R11234 VDPWR.n532 VDPWR.n253 1.42384
R11235 VDPWR.n646 VDPWR.n546 1.4005
R11236 VDPWR.n366 VDPWR.n266 1.4005
R11237 VDPWR.n2875 VDPWR.n2874 1.4005
R11238 VDPWR.n2768 VDPWR.n2767 1.4005
R11239 VDPWR.n108 VDPWR.n8 1.4005
R11240 VDPWR.n1133 VDPWR.n1132 1.39755
R11241 VDPWR.n2202 VDPWR.n2200 1.36443
R11242 VDPWR.n2283 VDPWR.n2282 1.36443
R11243 VDPWR.n758 VDPWR.n757 1.34339
R11244 VDPWR.n2883 VDPWR.n961 1.3232
R11245 VDPWR.n402 VDPWR.n389 1.28133
R11246 VDPWR.n1926 VDPWR.n1924 1.2502
R11247 VDPWR.n257 VDPWR.n256 1.16828
R11248 VDPWR.n3133 VDPWR.n3132 1.16528
R11249 VDPWR.n755 VDPWR.n118 1.15151
R11250 VDPWR.n703 VDPWR.n702 1.143
R11251 VDPWR.n687 VDPWR.n686 1.143
R11252 VDPWR.n514 VDPWR.n513 1.143
R11253 VDPWR.n498 VDPWR.n497 1.143
R11254 VDPWR.n460 VDPWR.n459 1.143
R11255 VDPWR.n444 VDPWR.n443 1.143
R11256 VDPWR.n3165 VDPWR.n3164 1.143
R11257 VDPWR.n3149 VDPWR.n3148 1.143
R11258 VDPWR.n719 VDPWR.n718 1.13925
R11259 VDPWR.n530 VDPWR.n529 1.13925
R11260 VDPWR.n466 VDPWR.n465 1.13925
R11261 VDPWR.n3171 VDPWR.n3170 1.13925
R11262 VDPWR.n3114 VDPWR.n3113 1.13717
R11263 VDPWR.n671 VDPWR.n670 1.13675
R11264 VDPWR.n482 VDPWR.n481 1.13675
R11265 VDPWR.n428 VDPWR.n427 1.13675
R11266 VDPWR.n715 VDPWR.n714 1.12991
R11267 VDPWR.n691 VDPWR.n689 1.12991
R11268 VDPWR.n683 VDPWR.n675 1.12991
R11269 VDPWR.n526 VDPWR.n525 1.12991
R11270 VDPWR.n502 VDPWR.n500 1.12991
R11271 VDPWR.n494 VDPWR.n486 1.12991
R11272 VDPWR.n462 VDPWR.n413 1.12991
R11273 VDPWR.n448 VDPWR.n446 1.12991
R11274 VDPWR.n440 VDPWR.n432 1.12991
R11275 VDPWR.n3167 VDPWR.n769 1.12991
R11276 VDPWR.n3153 VDPWR.n3151 1.12991
R11277 VDPWR.n3145 VDPWR.n3137 1.12991
R11278 VDPWR.n2472 VDPWR.n2471 1.11173
R11279 VDPWR.n2397 VDPWR.n2359 1.08324
R11280 VDPWR.n721 VDPWR.n720 1.06914
R11281 VDPWR.n595 VDPWR 1.06099
R11282 VDPWR.n315 VDPWR 1.06099
R11283 VDPWR.n57 VDPWR 1.06099
R11284 VDPWR.n1368 VDPWR.n1367 1.05773
R11285 VDPWR.n1701 VDPWR.n1700 1.05773
R11286 VDPWR.n1622 VDPWR.n1603 1.05773
R11287 VDPWR.n2452 VDPWR.n2451 1.05773
R11288 VDPWR.n2221 VDPWR.n2220 1.04968
R11289 VDPWR.n2276 VDPWR.n2275 1.04968
R11290 VDPWR.n2739 VDPWR.n2726 0.992049
R11291 VDPWR.n2728 VDPWR.n1006 0.992049
R11292 VDPWR.n3117 VDPWR.n117 0.973454
R11293 VDPWR.n2049 VDPWR.n1130 0.899674
R11294 VDPWR VDPWR.n118 0.891339
R11295 VDPWR.n756 VDPWR.n755 0.884173
R11296 VDPWR.n2176 VDPWR.n1104 0.863992
R11297 VDPWR.n376 VDPWR.n375 0.853
R11298 VDPWR.n3102 VDPWR.n782 0.853
R11299 VDPWR.n2508 VDPWR.n2507 0.853
R11300 VDPWR.n2537 VDPWR.n2536 0.853
R11301 VDPWR.n2392 VDPWR.n2339 0.853
R11302 VDPWR.n3074 VDPWR.n3073 0.853
R11303 VDPWR.n688 VDPWR.n687 0.849559
R11304 VDPWR.n445 VDPWR.n444 0.849559
R11305 VDPWR.n499 VDPWR.n498 0.849559
R11306 VDPWR.n531 VDPWR.n377 0.843267
R11307 VDPWR.n2422 VDPWR.n2421 0.813198
R11308 VDPWR.n2520 VDPWR.n2519 0.813198
R11309 VDPWR.n532 VDPWR.n531 0.810458
R11310 VDPWR VDPWR.n3116 0.778686
R11311 VDPWR.n822 VDPWR 0.777643
R11312 VDPWR.n739 VDPWR.n738 0.7755
R11313 VDPWR.n672 VDPWR.n671 0.770881
R11314 VDPWR.n429 VDPWR.n428 0.770881
R11315 VDPWR.n403 VDPWR.n402 0.767167
R11316 VDPWR.n375 VDPWR.n374 0.763912
R11317 VDPWR.n633 VDPWR.n562 0.753441
R11318 VDPWR.n353 VDPWR.n282 0.753441
R11319 VDPWR.n1877 VDPWR.n1876 0.753441
R11320 VDPWR.n95 VDPWR.n24 0.753441
R11321 VDPWR.n1842 VDPWR.n1841 0.740996
R11322 VDPWR.n461 VDPWR.n460 0.73614
R11323 VDPWR.n704 VDPWR.n703 0.717512
R11324 VDPWR.n515 VDPWR.n514 0.717512
R11325 VDPWR.n2938 VDPWR.n2937 0.706789
R11326 VDPWR.n758 VDPWR.n118 0.70421
R11327 VDPWR.n255 VDPWR 0.659186
R11328 VDPWR.n865 VDPWR.n814 0.65125
R11329 VDPWR.n1499 VDPWR.n1296 0.635211
R11330 VDPWR.n1576 VDPWR.n1520 0.635211
R11331 VDPWR.n1865 VDPWR.n1213 0.635211
R11332 VDPWR.n2185 VDPWR.n2184 0.635211
R11333 VDPWR.n2316 VDPWR.n2315 0.635211
R11334 VDPWR.n2310 VDPWR.n2309 0.635211
R11335 VDPWR.n2904 VDPWR.n2903 0.635211
R11336 VDPWR.n2937 VDPWR.n939 0.635211
R11337 VDPWR.n2940 VDPWR.n2939 0.635211
R11338 VDPWR.n2947 VDPWR.n2946 0.635211
R11339 VDPWR.n2226 VDPWR.n2203 0.630008
R11340 VDPWR.n1056 VDPWR.n1051 0.630008
R11341 VDPWR.n2285 VDPWR.n2284 0.630008
R11342 VDPWR.n656 VDPWR.n537 0.624567
R11343 VDPWR.n543 VDPWR.n541 0.6005
R11344 VDPWR.n263 VDPWR.n261 0.6005
R11345 VDPWR.n5 VDPWR.n3 0.6005
R11346 VDPWR.n2207 VDPWR.n2205 0.52509
R11347 VDPWR.n467 VDPWR.n466 0.518882
R11348 VDPWR.n655 VDPWR.n654 0.511794
R11349 VDPWR.n3178 VDPWR.n116 0.511794
R11350 VDPWR.n2336 VDPWR.n2335 0.500125
R11351 VDPWR.n1594 VDPWR.n1593 0.500125
R11352 VDPWR.n1675 VDPWR.n1674 0.500125
R11353 VDPWR.n1596 VDPWR.n1090 0.500125
R11354 VDPWR.n2540 VDPWR.n2539 0.500125
R11355 VDPWR.n2504 VDPWR.n2501 0.500125
R11356 VDPWR.n142 VDPWR.n141 0.465384
R11357 VDPWR.n654 VDPWR 0.460219
R11358 VDPWR.n374 VDPWR 0.460219
R11359 VDPWR.n116 VDPWR 0.460219
R11360 VDPWR.n3091 VDPWR.n3090 0.457643
R11361 VDPWR.n376 VDPWR.n257 0.45408
R11362 VDPWR.n719 VDPWR.n704 0.405788
R11363 VDPWR.n649 VDPWR.n541 0.4005
R11364 VDPWR.n369 VDPWR.n261 0.4005
R11365 VDPWR.n111 VDPWR.n3 0.4005
R11366 VDPWR.n2253 VDPWR.n1046 0.3805
R11367 VDPWR.n1908 VDPWR.n1907 0.3805
R11368 VDPWR.n1590 VDPWR.n1589 0.3805
R11369 VDPWR.n1011 VDPWR.n943 0.3805
R11370 VDPWR.n3072 VDPWR.n3071 0.3805
R11371 VDPWR.n3069 VDPWR.n3068 0.3805
R11372 VDPWR.n2252 VDPWR.n1012 0.3805
R11373 VDPWR.n1192 VDPWR.n1162 0.3805
R11374 VDPWR.n1591 VDPWR.n1228 0.3805
R11375 VDPWR.n2333 VDPWR.n2332 0.3805
R11376 VDPWR.n2499 VDPWR.n871 0.3805
R11377 VDPWR.n2251 VDPWR.n2250 0.3805
R11378 VDPWR.n1673 VDPWR.n1246 0.3805
R11379 VDPWR.n1592 VDPWR.n1245 0.3805
R11380 VDPWR.n2334 VDPWR.n973 0.3805
R11381 VDPWR.n2506 VDPWR.n2505 0.3805
R11382 VDPWR.n780 VDPWR.n776 0.3805
R11383 VDPWR.n3109 VDPWR.n3108 0.3805
R11384 VDPWR.n2255 VDPWR.n2254 0.3805
R11385 VDPWR.n1906 VDPWR.n1905 0.3805
R11386 VDPWR.n1284 VDPWR.n1193 0.3805
R11387 VDPWR.n1010 VDPWR.n923 0.3805
R11388 VDPWR.n3070 VDPWR.n775 0.3805
R11389 VDPWR.n3111 VDPWR.n3110 0.3805
R11390 VDPWR.n2504 VDPWR.n2503 0.3805
R11391 VDPWR.n2539 VDPWR.n2538 0.3805
R11392 VDPWR.n2073 VDPWR.n1090 0.3805
R11393 VDPWR.n1674 VDPWR.n1116 0.3805
R11394 VDPWR.n1593 VDPWR.n1267 0.3805
R11395 VDPWR.n2335 VDPWR.n988 0.3805
R11396 VDPWR.n687 VDPWR.n672 0.379066
R11397 VDPWR.n444 VDPWR.n429 0.379066
R11398 VDPWR.n498 VDPWR.n483 0.379066
R11399 VDPWR.n721 VDPWR.n253 0.375001
R11400 VDPWR.n377 VDPWR 0.36983
R11401 VDPWR.n1435 VDPWR.n1323 0.369731
R11402 VDPWR.n1465 VDPWR.n1312 0.369731
R11403 VDPWR.n1466 VDPWR.n1311 0.369731
R11404 VDPWR.n1482 VDPWR.n1481 0.369731
R11405 VDPWR.n1397 VDPWR.n1396 0.369731
R11406 VDPWR.n1402 VDPWR.n1339 0.369731
R11407 VDPWR.n1405 VDPWR.n1404 0.369731
R11408 VDPWR.n1428 VDPWR.n1328 0.369731
R11409 VDPWR.n1575 VDPWR.n1521 0.369731
R11410 VDPWR.n1537 VDPWR.n1528 0.369731
R11411 VDPWR.n1727 VDPWR.n1726 0.369731
R11412 VDPWR.n1732 VDPWR.n1275 0.369731
R11413 VDPWR.n1735 VDPWR.n1734 0.369731
R11414 VDPWR.n1743 VDPWR.n1263 0.369731
R11415 VDPWR.n1769 VDPWR.n1768 0.369731
R11416 VDPWR.n1792 VDPWR.n1791 0.369731
R11417 VDPWR.n1798 VDPWR.n1797 0.369731
R11418 VDPWR.n1810 VDPWR.n1224 0.369731
R11419 VDPWR.n2016 VDPWR.n1156 0.369731
R11420 VDPWR.n1178 VDPWR.n1177 0.369731
R11421 VDPWR.n1153 VDPWR.n1151 0.369731
R11422 VDPWR.n2017 VDPWR.n1155 0.369731
R11423 VDPWR.n2040 VDPWR.n1134 0.369731
R11424 VDPWR.n2027 VDPWR.n2026 0.369731
R11425 VDPWR.n1640 VDPWR.n1639 0.369731
R11426 VDPWR.n2059 VDPWR.n2058 0.369731
R11427 VDPWR.n1649 VDPWR.n1628 0.369731
R11428 VDPWR.n1644 VDPWR.n1643 0.369731
R11429 VDPWR.n2136 VDPWR.n2135 0.369731
R11430 VDPWR.n2140 VDPWR.n2080 0.369731
R11431 VDPWR.n2142 VDPWR.n2141 0.369731
R11432 VDPWR.n2167 VDPWR.n2166 0.369731
R11433 VDPWR.n530 VDPWR.n515 0.360095
R11434 VDPWR.n703 VDPWR.n688 0.348599
R11435 VDPWR.n460 VDPWR.n445 0.348599
R11436 VDPWR.n514 VDPWR.n499 0.348599
R11437 VDPWR.n1028 VDPWR.n1026 0.317855
R11438 VDPWR.n1029 VDPWR.n1028 0.317855
R11439 VDPWR.n751 VDPWR.n739 0.310024
R11440 VDPWR.n605 VDPWR.n596 0.305262
R11441 VDPWR.n624 VDPWR.n623 0.305262
R11442 VDPWR.n574 VDPWR.n573 0.305262
R11443 VDPWR.n583 VDPWR.n582 0.305262
R11444 VDPWR.n559 VDPWR.n548 0.305262
R11445 VDPWR.n325 VDPWR.n316 0.305262
R11446 VDPWR.n344 VDPWR.n343 0.305262
R11447 VDPWR.n294 VDPWR.n293 0.305262
R11448 VDPWR.n303 VDPWR.n302 0.305262
R11449 VDPWR.n279 VDPWR.n268 0.305262
R11450 VDPWR.n750 VDPWR.n740 0.305262
R11451 VDPWR.n1936 VDPWR.n1928 0.305262
R11452 VDPWR.n2179 VDPWR.n1103 0.305262
R11453 VDPWR.n2884 VDPWR.n2883 0.305262
R11454 VDPWR.n2889 VDPWR.n2888 0.305262
R11455 VDPWR.n2763 VDPWR.n2762 0.305262
R11456 VDPWR.n2629 VDPWR.n2628 0.305262
R11457 VDPWR.n885 VDPWR.n884 0.305262
R11458 VDPWR.n3018 VDPWR.n917 0.305262
R11459 VDPWR.n2988 VDPWR.n2987 0.305262
R11460 VDPWR.n2412 VDPWR.n2411 0.305262
R11461 VDPWR.n2417 VDPWR.n2416 0.305262
R11462 VDPWR.n2420 VDPWR.n2349 0.305262
R11463 VDPWR.n2398 VDPWR.n2397 0.305262
R11464 VDPWR.n2404 VDPWR.n2357 0.305262
R11465 VDPWR.n2526 VDPWR.n2525 0.305262
R11466 VDPWR.n2524 VDPWR.n2434 0.305262
R11467 VDPWR.n2515 VDPWR.n2437 0.305262
R11468 VDPWR.n3095 VDPWR.n792 0.305262
R11469 VDPWR.n3080 VDPWR.n798 0.305262
R11470 VDPWR.n865 VDPWR.n864 0.305262
R11471 VDPWR.n831 VDPWR.n830 0.305262
R11472 VDPWR.n67 VDPWR.n58 0.305262
R11473 VDPWR.n86 VDPWR.n85 0.305262
R11474 VDPWR.n36 VDPWR.n35 0.305262
R11475 VDPWR.n45 VDPWR.n44 0.305262
R11476 VDPWR.n21 VDPWR.n10 0.305262
R11477 VDPWR.n2392 VDPWR.n2343 0.297373
R11478 VDPWR.n384 VDPWR.t772 0.27666
R11479 VDPWR.t772 VDPWR.n383 0.27666
R11480 VDPWR.n396 VDPWR.t119 0.27666
R11481 VDPWR.t119 VDPWR.n395 0.27666
R11482 VDPWR.n756 VDPWR.n721 0.262659
R11483 VDPWR.n738 VDPWR.n729 0.2565
R11484 VDPWR.n2773 VDPWR.n2771 0.25148
R11485 VDPWR.n2816 VDPWR.n982 0.246654
R11486 VDPWR.n256 VDPWR 0.245332
R11487 VDPWR.n2561 VDPWR 0.237784
R11488 VDPWR.n1886 VDPWR.n1884 0.231913
R11489 VDPWR.n1368 VDPWR.n1350 0.227049
R11490 VDPWR.n1391 VDPWR.n1341 0.227049
R11491 VDPWR.n1503 VDPWR.n1502 0.227049
R11492 VDPWR.n1516 VDPWR.n1292 0.227049
R11493 VDPWR.n1701 VDPWR.n1683 0.227049
R11494 VDPWR.n1721 VDPWR.n1277 0.227049
R11495 VDPWR.n2000 VDPWR.n1179 0.227049
R11496 VDPWR.n1995 VDPWR.n1994 0.227049
R11497 VDPWR.n2041 VDPWR.n1133 0.227049
R11498 VDPWR.n1603 VDPWR.n1602 0.227049
R11499 VDPWR.n1650 VDPWR.n1627 0.227049
R11500 VDPWR.n2108 VDPWR.n2090 0.227049
R11501 VDPWR.n2134 VDPWR.n2082 0.227049
R11502 VDPWR.n2212 VDPWR.n2211 0.227049
R11503 VDPWR.n1025 VDPWR.n1019 0.227049
R11504 VDPWR.n2270 VDPWR.n1066 0.227049
R11505 VDPWR.n2265 VDPWR.n2264 0.227049
R11506 VDPWR.n2953 VDPWR.n2952 0.227049
R11507 VDPWR.n2959 VDPWR.n929 0.227049
R11508 VDPWR.n2451 VDPWR.n2450 0.227049
R11509 VDPWR.n2485 VDPWR.n2484 0.227049
R11510 VDPWR.n1832 VDPWR 0.217591
R11511 VDPWR.n1839 VDPWR.n1221 0.21207
R11512 VDPWR.n2903 VDPWR.n953 0.21207
R11513 VDPWR.n2941 VDPWR.n937 0.21207
R11514 VDPWR.n2502 VDPWR 0.209323
R11515 VDPWR.n3166 VDPWR.n3165 0.209134
R11516 VDPWR.n3150 VDPWR.n3149 0.206276
R11517 VDPWR.n3107 VDPWR 0.206051
R11518 VDPWR.n2627 VDPWR.n878 0.203675
R11519 VDPWR.n2561 VDPWR 0.200023
R11520 VDPWR.n3116 VDPWR.n770 0.197315
R11521 VDPWR.n3103 VDPWR.n770 0.196829
R11522 VDPWR.n3107 VDPWR.n3106 0.196829
R11523 VDPWR.n2343 VDPWR.n779 0.195044
R11524 VDPWR.n2502 VDPWR.n778 0.195044
R11525 VDPWR.n2777 VDPWR.n1001 0.194439
R11526 VDPWR.n3176 VDPWR 0.189894
R11527 VDPWR.n1970 VDPWR.n1915 0.180304
R11528 VDPWR.n2624 VDPWR.n2622 0.180304
R11529 VDPWR.n1433 VDPWR 0.17983
R11530 VDPWR VDPWR.n2055 0.17983
R11531 VDPWR VDPWR.n1964 0.17983
R11532 VDPWR.n2746 VDPWR 0.17983
R11533 VDPWR VDPWR.n854 0.17983
R11534 VDPWR.n1362 VDPWR 0.179485
R11535 VDPWR.n1695 VDPWR 0.179485
R11536 VDPWR.n1884 VDPWR 0.179485
R11537 VDPWR VDPWR.n1609 0.179485
R11538 VDPWR.n1964 VDPWR 0.179485
R11539 VDPWR.n888 VDPWR 0.179485
R11540 VDPWR.n854 VDPWR 0.179485
R11541 VDPWR.n739 VDPWR.n728 0.176553
R11542 VDPWR VDPWR.n1361 0.172576
R11543 VDPWR VDPWR.n1694 0.172576
R11544 VDPWR.n1616 VDPWR 0.172576
R11545 VDPWR VDPWR.n2103 0.172576
R11546 VDPWR VDPWR.n2736 0.172576
R11547 VDPWR VDPWR.n2560 0.172576
R11548 VDPWR VDPWR.n2378 0.172576
R11549 VDPWR.n536 VDPWR 0.163379
R11550 VDPWR.n2932 VDPWR.n870 0.1603
R11551 VDPWR.n3067 VDPWR.n872 0.1603
R11552 VDPWR.n2844 VDPWR.n974 0.1603
R11553 VDPWR.n2755 VDPWR.n2719 0.1603
R11554 VDPWR.n2982 VDPWR.n2981 0.1603
R11555 VDPWR.n2805 VDPWR.n989 0.1603
R11556 VDPWR.n1765 VDPWR 0.158169
R11557 VDPWR.n1794 VDPWR 0.158169
R11558 VDPWR.n2460 VDPWR 0.158169
R11559 VDPWR.n203 VDPWR.n202 0.155911
R11560 VDPWR.n2177 VDPWR.n2176 0.152881
R11561 VDPWR.n3134 VDPWR.n3133 0.152187
R11562 VDPWR.n757 VDPWR.n756 0.150053
R11563 VDPWR.n3073 VDPWR.n3072 0.14385
R11564 VDPWR.n3068 VDPWR.n782 0.14385
R11565 VDPWR.n2507 VDPWR.n2499 0.14385
R11566 VDPWR.n2540 VDPWR.n2339 0.14385
R11567 VDPWR.n3113 VDPWR.n775 0.14385
R11568 VDPWR.n2538 VDPWR.n2537 0.14385
R11569 VDPWR.n2746 VDPWR.n2721 0.143027
R11570 VDPWR.n2290 VDPWR.n943 0.142675
R11571 VDPWR.n2332 VDPWR.n2331 0.142675
R11572 VDPWR.n2249 VDPWR.n973 0.142675
R11573 VDPWR.n2336 VDPWR.n1009 0.142675
R11574 VDPWR.n2256 VDPWR.n923 0.142675
R11575 VDPWR.n2159 VDPWR.n988 0.142675
R11576 VDPWR.n1362 VDPWR 0.14207
R11577 VDPWR.n1695 VDPWR 0.14207
R11578 VDPWR.n1609 VDPWR 0.14207
R11579 VDPWR VDPWR.n888 0.14207
R11580 VDPWR.n1433 VDPWR 0.141725
R11581 VDPWR.n1832 VDPWR 0.141725
R11582 VDPWR.n2055 VDPWR 0.141725
R11583 VDPWR.n1764 VDPWR 0.120408
R11584 VDPWR.n2104 VDPWR 0.120408
R11585 VDPWR VDPWR.n2476 0.120408
R11586 VDPWR.n1589 VDPWR.n1191 0.12035
R11587 VDPWR.n1820 VDPWR.n1228 0.12035
R11588 VDPWR.n1784 VDPWR.n1245 0.12035
R11589 VDPWR.n1714 VDPWR.n1594 0.12035
R11590 VDPWR.n1904 VDPWR.n1193 0.12035
R11591 VDPWR.n1754 VDPWR.n1267 0.12035
R11592 VDPWR.n587 VDPWR.n566 0.120292
R11593 VDPWR.n626 VDPWR.n567 0.120292
R11594 VDPWR.n619 VDPWR.n618 0.120292
R11595 VDPWR.n618 VDPWR.n592 0.120292
R11596 VDPWR.n614 VDPWR.n613 0.120292
R11597 VDPWR.n613 VDPWR.n612 0.120292
R11598 VDPWR.n609 VDPWR.n608 0.120292
R11599 VDPWR.n608 VDPWR.n607 0.120292
R11600 VDPWR.n604 VDPWR.n603 0.120292
R11601 VDPWR.n603 VDPWR.n597 0.120292
R11602 VDPWR.n599 VDPWR.n597 0.120292
R11603 VDPWR.n572 VDPWR.n568 0.120292
R11604 VDPWR.n585 VDPWR.n569 0.120292
R11605 VDPWR.n636 VDPWR.n563 0.120292
R11606 VDPWR.n637 VDPWR.n636 0.120292
R11607 VDPWR.n652 VDPWR.n538 0.120292
R11608 VDPWR.n648 VDPWR.n647 0.120292
R11609 VDPWR.n647 VDPWR.n542 0.120292
R11610 VDPWR.n558 VDPWR.n557 0.120292
R11611 VDPWR.n557 VDPWR.n549 0.120292
R11612 VDPWR.n552 VDPWR.n549 0.120292
R11613 VDPWR.n307 VDPWR.n286 0.120292
R11614 VDPWR.n346 VDPWR.n287 0.120292
R11615 VDPWR.n339 VDPWR.n338 0.120292
R11616 VDPWR.n338 VDPWR.n312 0.120292
R11617 VDPWR.n334 VDPWR.n333 0.120292
R11618 VDPWR.n333 VDPWR.n332 0.120292
R11619 VDPWR.n329 VDPWR.n328 0.120292
R11620 VDPWR.n328 VDPWR.n327 0.120292
R11621 VDPWR.n324 VDPWR.n323 0.120292
R11622 VDPWR.n323 VDPWR.n317 0.120292
R11623 VDPWR.n319 VDPWR.n317 0.120292
R11624 VDPWR.n292 VDPWR.n288 0.120292
R11625 VDPWR.n305 VDPWR.n289 0.120292
R11626 VDPWR.n356 VDPWR.n283 0.120292
R11627 VDPWR.n357 VDPWR.n356 0.120292
R11628 VDPWR.n372 VDPWR.n258 0.120292
R11629 VDPWR.n368 VDPWR.n367 0.120292
R11630 VDPWR.n367 VDPWR.n262 0.120292
R11631 VDPWR.n278 VDPWR.n277 0.120292
R11632 VDPWR.n277 VDPWR.n269 0.120292
R11633 VDPWR.n272 VDPWR.n269 0.120292
R11634 VDPWR.n1375 VDPWR.n1369 0.120292
R11635 VDPWR.n1388 VDPWR.n1342 0.120292
R11636 VDPWR.n1393 VDPWR.n1342 0.120292
R11637 VDPWR.n1394 VDPWR.n1393 0.120292
R11638 VDPWR.n1395 VDPWR.n1340 0.120292
R11639 VDPWR.n1400 VDPWR.n1340 0.120292
R11640 VDPWR.n1401 VDPWR.n1400 0.120292
R11641 VDPWR.n1407 VDPWR.n1338 0.120292
R11642 VDPWR.n1408 VDPWR.n1407 0.120292
R11643 VDPWR.n1409 VDPWR.n1408 0.120292
R11644 VDPWR.n1437 VDPWR.n1436 0.120292
R11645 VDPWR.n1437 VDPWR.n1322 0.120292
R11646 VDPWR.n1442 VDPWR.n1322 0.120292
R11647 VDPWR.n1443 VDPWR.n1442 0.120292
R11648 VDPWR.n1444 VDPWR.n1443 0.120292
R11649 VDPWR.n1464 VDPWR.n1313 0.120292
R11650 VDPWR VDPWR.n1464 0.120292
R11651 VDPWR.n1468 VDPWR.n1467 0.120292
R11652 VDPWR.n1468 VDPWR.n1310 0.120292
R11653 VDPWR.n1472 VDPWR.n1310 0.120292
R11654 VDPWR.n1473 VDPWR.n1472 0.120292
R11655 VDPWR.n1473 VDPWR.n1308 0.120292
R11656 VDPWR.n1477 VDPWR.n1308 0.120292
R11657 VDPWR.n1478 VDPWR.n1477 0.120292
R11658 VDPWR.n1479 VDPWR.n1478 0.120292
R11659 VDPWR.n1501 VDPWR.n1295 0.120292
R11660 VDPWR.n1508 VDPWR.n1295 0.120292
R11661 VDPWR.n1509 VDPWR.n1508 0.120292
R11662 VDPWR.n1510 VDPWR.n1509 0.120292
R11663 VDPWR.n1510 VDPWR.n1293 0.120292
R11664 VDPWR.n1514 VDPWR.n1293 0.120292
R11665 VDPWR.n1515 VDPWR.n1514 0.120292
R11666 VDPWR.n1574 VDPWR.n1573 0.120292
R11667 VDPWR.n1573 VDPWR.n1523 0.120292
R11668 VDPWR.n1569 VDPWR.n1523 0.120292
R11669 VDPWR.n1569 VDPWR.n1568 0.120292
R11670 VDPWR.n1568 VDPWR.n1525 0.120292
R11671 VDPWR.n1564 VDPWR.n1525 0.120292
R11672 VDPWR.n1564 VDPWR.n1563 0.120292
R11673 VDPWR.n1563 VDPWR.n1562 0.120292
R11674 VDPWR.n1562 VDPWR.n1527 0.120292
R11675 VDPWR.n1558 VDPWR.n1527 0.120292
R11676 VDPWR.n1703 VDPWR.n1702 0.120292
R11677 VDPWR.n1718 VDPWR.n1278 0.120292
R11678 VDPWR.n1723 VDPWR.n1278 0.120292
R11679 VDPWR.n1724 VDPWR.n1723 0.120292
R11680 VDPWR.n1725 VDPWR.n1276 0.120292
R11681 VDPWR.n1730 VDPWR.n1276 0.120292
R11682 VDPWR.n1731 VDPWR.n1730 0.120292
R11683 VDPWR.n1737 VDPWR.n1274 0.120292
R11684 VDPWR.n1738 VDPWR.n1737 0.120292
R11685 VDPWR.n1739 VDPWR.n1738 0.120292
R11686 VDPWR.n1772 VDPWR.n1256 0.120292
R11687 VDPWR.n1773 VDPWR.n1772 0.120292
R11688 VDPWR.n1774 VDPWR.n1773 0.120292
R11689 VDPWR.n1788 VDPWR.n1240 0.120292
R11690 VDPWR.n1793 VDPWR.n1240 0.120292
R11691 VDPWR.n1800 VDPWR.n1238 0.120292
R11692 VDPWR.n1801 VDPWR.n1800 0.120292
R11693 VDPWR.n1801 VDPWR.n1236 0.120292
R11694 VDPWR.n1806 VDPWR.n1236 0.120292
R11695 VDPWR.n1807 VDPWR.n1806 0.120292
R11696 VDPWR.n1808 VDPWR.n1807 0.120292
R11697 VDPWR.n1838 VDPWR.n1219 0.120292
R11698 VDPWR.n1843 VDPWR.n1219 0.120292
R11699 VDPWR.n1844 VDPWR.n1843 0.120292
R11700 VDPWR.n1845 VDPWR.n1844 0.120292
R11701 VDPWR.n1868 VDPWR.n1867 0.120292
R11702 VDPWR.n1869 VDPWR.n1868 0.120292
R11703 VDPWR.n1869 VDPWR.n1210 0.120292
R11704 VDPWR.n1878 VDPWR.n1210 0.120292
R11705 VDPWR.n1879 VDPWR.n1878 0.120292
R11706 VDPWR.n1880 VDPWR.n1879 0.120292
R11707 VDPWR.n1608 VDPWR.n1607 0.120292
R11708 VDPWR.n1656 VDPWR.n1626 0.120292
R11709 VDPWR.n1652 VDPWR.n1626 0.120292
R11710 VDPWR.n1652 VDPWR.n1651 0.120292
R11711 VDPWR.n1648 VDPWR.n1647 0.120292
R11712 VDPWR.n1647 VDPWR.n1629 0.120292
R11713 VDPWR.n1642 VDPWR.n1629 0.120292
R11714 VDPWR.n1641 VDPWR.n1631 0.120292
R11715 VDPWR.n1636 VDPWR.n1631 0.120292
R11716 VDPWR.n1636 VDPWR.n1635 0.120292
R11717 VDPWR.n2054 VDPWR.n1129 0.120292
R11718 VDPWR.n2044 VDPWR.n1129 0.120292
R11719 VDPWR.n2044 VDPWR.n2043 0.120292
R11720 VDPWR.n2043 VDPWR.n2042 0.120292
R11721 VDPWR.n2030 VDPWR.n1141 0.120292
R11722 VDPWR.n2025 VDPWR.n1141 0.120292
R11723 VDPWR.n2024 VDPWR.n2023 0.120292
R11724 VDPWR.n2023 VDPWR.n1152 0.120292
R11725 VDPWR.n2019 VDPWR.n1152 0.120292
R11726 VDPWR.n2019 VDPWR.n2018 0.120292
R11727 VDPWR.n2015 VDPWR.n2014 0.120292
R11728 VDPWR.n2014 VDPWR.n1157 0.120292
R11729 VDPWR.n2010 VDPWR.n1157 0.120292
R11730 VDPWR.n1999 VDPWR.n1998 0.120292
R11731 VDPWR.n1998 VDPWR.n1180 0.120292
R11732 VDPWR.n1993 VDPWR.n1180 0.120292
R11733 VDPWR.n1991 VDPWR.n1183 0.120292
R11734 VDPWR.n1985 VDPWR.n1984 0.120292
R11735 VDPWR.n1984 VDPWR.n1185 0.120292
R11736 VDPWR.n1962 VDPWR.n1923 0.120292
R11737 VDPWR.n1957 VDPWR.n1923 0.120292
R11738 VDPWR.n2114 VDPWR.n2109 0.120292
R11739 VDPWR.n2128 VDPWR.n2083 0.120292
R11740 VDPWR.n2132 VDPWR.n2083 0.120292
R11741 VDPWR.n2133 VDPWR.n2132 0.120292
R11742 VDPWR.n2138 VDPWR.n2081 0.120292
R11743 VDPWR.n2139 VDPWR.n2138 0.120292
R11744 VDPWR.n2144 VDPWR.n2143 0.120292
R11745 VDPWR.n2144 VDPWR.n2078 0.120292
R11746 VDPWR.n2148 VDPWR.n2078 0.120292
R11747 VDPWR.n2149 VDPWR.n2148 0.120292
R11748 VDPWR.n2182 VDPWR.n2181 0.120292
R11749 VDPWR.n2183 VDPWR.n1101 0.120292
R11750 VDPWR.n2189 VDPWR.n1101 0.120292
R11751 VDPWR.n2190 VDPWR.n2189 0.120292
R11752 VDPWR.n2234 VDPWR.n2198 0.120292
R11753 VDPWR.n2229 VDPWR.n2198 0.120292
R11754 VDPWR.n2229 VDPWR.n2228 0.120292
R11755 VDPWR.n2228 VDPWR.n2227 0.120292
R11756 VDPWR.n2224 VDPWR.n2223 0.120292
R11757 VDPWR.n2223 VDPWR.n2206 0.120292
R11758 VDPWR.n2218 VDPWR.n2206 0.120292
R11759 VDPWR.n2218 VDPWR.n2217 0.120292
R11760 VDPWR.n2312 VDPWR.n1027 0.120292
R11761 VDPWR.n2307 VDPWR.n1027 0.120292
R11762 VDPWR.n2307 VDPWR.n2306 0.120292
R11763 VDPWR.n2306 VDPWR.n1032 0.120292
R11764 VDPWR.n2301 VDPWR.n1032 0.120292
R11765 VDPWR.n2301 VDPWR.n2300 0.120292
R11766 VDPWR.n2300 VDPWR.n2299 0.120292
R11767 VDPWR.n2286 VDPWR.n1049 0.120292
R11768 VDPWR.n2280 VDPWR.n1049 0.120292
R11769 VDPWR.n2280 VDPWR.n2279 0.120292
R11770 VDPWR.n2279 VDPWR.n2278 0.120292
R11771 VDPWR.n2278 VDPWR.n1060 0.120292
R11772 VDPWR.n2273 VDPWR.n1060 0.120292
R11773 VDPWR.n2273 VDPWR.n2272 0.120292
R11774 VDPWR.n2269 VDPWR.n2268 0.120292
R11775 VDPWR.n2268 VDPWR.n1067 0.120292
R11776 VDPWR.n2764 VDPWR.n1004 0.120292
R11777 VDPWR.n2766 VDPWR.n2765 0.120292
R11778 VDPWR.n2766 VDPWR.n1002 0.120292
R11779 VDPWR.n2775 VDPWR.n1002 0.120292
R11780 VDPWR.n2778 VDPWR.n2775 0.120292
R11781 VDPWR.n2779 VDPWR.n2778 0.120292
R11782 VDPWR.n2786 VDPWR.n999 0.120292
R11783 VDPWR.n2787 VDPWR.n2786 0.120292
R11784 VDPWR.n2819 VDPWR.n2818 0.120292
R11785 VDPWR.n2826 VDPWR.n2825 0.120292
R11786 VDPWR.n2833 VDPWR.n2832 0.120292
R11787 VDPWR.n2856 VDPWR.n2855 0.120292
R11788 VDPWR.n2862 VDPWR.n966 0.120292
R11789 VDPWR.n2863 VDPWR.n2862 0.120292
R11790 VDPWR.n2864 VDPWR.n2863 0.120292
R11791 VDPWR.n2864 VDPWR.n963 0.120292
R11792 VDPWR.n2869 VDPWR.n963 0.120292
R11793 VDPWR.n2906 VDPWR.n2905 0.120292
R11794 VDPWR.n2906 VDPWR.n951 0.120292
R11795 VDPWR.n2911 VDPWR.n951 0.120292
R11796 VDPWR.n2912 VDPWR.n2911 0.120292
R11797 VDPWR.n2912 VDPWR.n949 0.120292
R11798 VDPWR.n2918 VDPWR.n949 0.120292
R11799 VDPWR.n2919 VDPWR.n2918 0.120292
R11800 VDPWR.n2920 VDPWR.n2919 0.120292
R11801 VDPWR.n2942 VDPWR.n938 0.120292
R11802 VDPWR.n2943 VDPWR.n2942 0.120292
R11803 VDPWR.n2949 VDPWR.n2948 0.120292
R11804 VDPWR.n2950 VDPWR.n2949 0.120292
R11805 VDPWR.n2955 VDPWR.n2954 0.120292
R11806 VDPWR.n2956 VDPWR.n2955 0.120292
R11807 VDPWR.n2956 VDPWR.n933 0.120292
R11808 VDPWR.n2961 VDPWR.n933 0.120292
R11809 VDPWR.n2715 VDPWR.n2544 0.120292
R11810 VDPWR.n2711 VDPWR.n2544 0.120292
R11811 VDPWR.n2711 VDPWR.n2710 0.120292
R11812 VDPWR.n2710 VDPWR.n2709 0.120292
R11813 VDPWR.n2709 VDPWR.n2580 0.120292
R11814 VDPWR.n2704 VDPWR.n2580 0.120292
R11815 VDPWR.n2704 VDPWR.n2703 0.120292
R11816 VDPWR.n2703 VDPWR.n2702 0.120292
R11817 VDPWR.n2702 VDPWR.n2584 0.120292
R11818 VDPWR.n2698 VDPWR.n2584 0.120292
R11819 VDPWR.n2698 VDPWR.n2697 0.120292
R11820 VDPWR.n2682 VDPWR.n2681 0.120292
R11821 VDPWR.n2681 VDPWR.n2680 0.120292
R11822 VDPWR.n2680 VDPWR.n2606 0.120292
R11823 VDPWR.n2674 VDPWR.n2606 0.120292
R11824 VDPWR.n2674 VDPWR.n2673 0.120292
R11825 VDPWR.n2673 VDPWR.n2672 0.120292
R11826 VDPWR.n2672 VDPWR.n2611 0.120292
R11827 VDPWR.n2667 VDPWR.n2611 0.120292
R11828 VDPWR.n2646 VDPWR.n2645 0.120292
R11829 VDPWR.n2645 VDPWR.n2644 0.120292
R11830 VDPWR.n2639 VDPWR.n2638 0.120292
R11831 VDPWR.n2638 VDPWR.n2622 0.120292
R11832 VDPWR.n3049 VDPWR.n3048 0.120292
R11833 VDPWR.n3048 VDPWR.n3047 0.120292
R11834 VDPWR.n3043 VDPWR.n895 0.120292
R11835 VDPWR.n3043 VDPWR.n3042 0.120292
R11836 VDPWR.n3042 VDPWR.n898 0.120292
R11837 VDPWR.n3028 VDPWR.n908 0.120292
R11838 VDPWR.n914 VDPWR.n908 0.120292
R11839 VDPWR.n3022 VDPWR.n914 0.120292
R11840 VDPWR.n3022 VDPWR.n3021 0.120292
R11841 VDPWR.n3021 VDPWR.n3020 0.120292
R11842 VDPWR.n3017 VDPWR.n3016 0.120292
R11843 VDPWR.n3016 VDPWR.n918 0.120292
R11844 VDPWR.n2384 VDPWR.n2367 0.120292
R11845 VDPWR.n2402 VDPWR.n2358 0.120292
R11846 VDPWR.n2407 VDPWR.n2354 0.120292
R11847 VDPWR.n2408 VDPWR.n2407 0.120292
R11848 VDPWR.n2414 VDPWR.n2413 0.120292
R11849 VDPWR.n2423 VDPWR.n2350 0.120292
R11850 VDPWR.n2522 VDPWR.n2435 0.120292
R11851 VDPWR.n2517 VDPWR.n2435 0.120292
R11852 VDPWR.n2517 VDPWR.n2516 0.120292
R11853 VDPWR.n2489 VDPWR.n2488 0.120292
R11854 VDPWR.n2488 VDPWR.n2487 0.120292
R11855 VDPWR.n2487 VDPWR.n2455 0.120292
R11856 VDPWR.n2482 VDPWR.n2481 0.120292
R11857 VDPWR.n2481 VDPWR.n2457 0.120292
R11858 VDPWR.n3088 VDPWR.n3087 0.120292
R11859 VDPWR.n3087 VDPWR.n3086 0.120292
R11860 VDPWR.n3086 VDPWR.n794 0.120292
R11861 VDPWR.n3082 VDPWR.n3081 0.120292
R11862 VDPWR.n861 VDPWR.n860 0.120292
R11863 VDPWR.n860 VDPWR.n816 0.120292
R11864 VDPWR.n49 VDPWR.n28 0.120292
R11865 VDPWR.n88 VDPWR.n29 0.120292
R11866 VDPWR.n81 VDPWR.n80 0.120292
R11867 VDPWR.n80 VDPWR.n54 0.120292
R11868 VDPWR.n76 VDPWR.n75 0.120292
R11869 VDPWR.n75 VDPWR.n74 0.120292
R11870 VDPWR.n71 VDPWR.n70 0.120292
R11871 VDPWR.n70 VDPWR.n69 0.120292
R11872 VDPWR.n66 VDPWR.n65 0.120292
R11873 VDPWR.n65 VDPWR.n59 0.120292
R11874 VDPWR.n61 VDPWR.n59 0.120292
R11875 VDPWR.n34 VDPWR.n30 0.120292
R11876 VDPWR.n47 VDPWR.n31 0.120292
R11877 VDPWR.n98 VDPWR.n25 0.120292
R11878 VDPWR.n99 VDPWR.n98 0.120292
R11879 VDPWR.n114 VDPWR.n0 0.120292
R11880 VDPWR.n110 VDPWR.n109 0.120292
R11881 VDPWR.n109 VDPWR.n4 0.120292
R11882 VDPWR.n20 VDPWR.n19 0.120292
R11883 VDPWR.n19 VDPWR.n11 0.120292
R11884 VDPWR.n14 VDPWR.n11 0.120292
R11885 VDPWR.n2335 VDPWR.n2334 0.120125
R11886 VDPWR.n2334 VDPWR.n2333 0.120125
R11887 VDPWR.n2333 VDPWR.n1011 0.120125
R11888 VDPWR.n1011 VDPWR.n1010 0.120125
R11889 VDPWR.n1593 VDPWR.n1592 0.120125
R11890 VDPWR.n1592 VDPWR.n1591 0.120125
R11891 VDPWR.n1591 VDPWR.n1590 0.120125
R11892 VDPWR.n1590 VDPWR.n1284 0.120125
R11893 VDPWR.n1674 VDPWR.n1673 0.120125
R11894 VDPWR.n1673 VDPWR.n1192 0.120125
R11895 VDPWR.n1907 VDPWR.n1192 0.120125
R11896 VDPWR.n1907 VDPWR.n1906 0.120125
R11897 VDPWR.n2251 VDPWR.n1090 0.120125
R11898 VDPWR.n2252 VDPWR.n2251 0.120125
R11899 VDPWR.n2253 VDPWR.n2252 0.120125
R11900 VDPWR.n2254 VDPWR.n2253 0.120125
R11901 VDPWR.n2539 VDPWR.n871 0.120125
R11902 VDPWR.n3069 VDPWR.n871 0.120125
R11903 VDPWR.n3071 VDPWR.n3069 0.120125
R11904 VDPWR.n3071 VDPWR.n3070 0.120125
R11905 VDPWR.n2505 VDPWR.n2504 0.120125
R11906 VDPWR.n2505 VDPWR.n776 0.120125
R11907 VDPWR.n3109 VDPWR.n776 0.120125
R11908 VDPWR.n3110 VDPWR.n3109 0.120125
R11909 VDPWR.n627 VDPWR.n566 0.11899
R11910 VDPWR.n347 VDPWR.n286 0.11899
R11911 VDPWR.n89 VDPWR.n28 0.11899
R11912 VDPWR.n3115 VDPWR.n771 0.116902
R11913 VDPWR.n2053 VDPWR.n2052 0.113774
R11914 VDPWR.n2052 VDPWR.n2047 0.113774
R11915 VDPWR.n757 VDPWR.n117 0.113371
R11916 VDPWR.n461 VDPWR.n403 0.1125
R11917 VDPWR.n1558 VDPWR.n1557 0.112479
R11918 VDPWR.n1076 VDPWR.n1067 0.112479
R11919 VDPWR.n2963 VDPWR.n2961 0.112479
R11920 VDPWR.n3010 VDPWR.n3009 0.112479
R11921 VDPWR.n849 VDPWR.n848 0.112479
R11922 VDPWR.n1974 VDPWR.n1046 0.1086
R11923 VDPWR.n2006 VDPWR.n1012 0.1086
R11924 VDPWR.n2250 VDPWR.n1091 0.1086
R11925 VDPWR.n1672 VDPWR.n1596 0.1086
R11926 VDPWR.n2255 VDPWR.n1089 0.1086
R11927 VDPWR.n2073 VDPWR.n2072 0.1086
R11928 VDPWR.n1444 VDPWR.n1319 0.107271
R11929 VDPWR.n1774 VDPWR.n1248 0.107271
R11930 VDPWR.n2039 VDPWR.n2038 0.107271
R11931 VDPWR.n2190 VDPWR.n1094 0.107271
R11932 VDPWR.n2833 VDPWR.n976 0.107271
R11933 VDPWR.n2667 VDPWR.n2666 0.107271
R11934 VDPWR.n3104 VDPWR.n779 0.10625
R11935 VDPWR.n3105 VDPWR.n778 0.10625
R11936 VDPWR.n2225 VDPWR.n2205 0.105418
R11937 VDPWR.n1062 VDPWR.n1059 0.105418
R11938 VDPWR.n1361 VDPWR 0.105238
R11939 VDPWR.n1694 VDPWR 0.105238
R11940 VDPWR.n1616 VDPWR 0.105238
R11941 VDPWR.n2103 VDPWR 0.105238
R11942 VDPWR.n2736 VDPWR 0.105238
R11943 VDPWR.n2560 VDPWR 0.105238
R11944 VDPWR.n2378 VDPWR 0.105238
R11945 VDPWR.n377 VDPWR.n254 0.103147
R11946 VDPWR.n1960 VDPWR.n1959 0.102087
R11947 VDPWR.n2891 VDPWR.n2890 0.102087
R11948 VDPWR.n3015 VDPWR.n3014 0.102087
R11949 VDPWR.n572 VDPWR 0.0981562
R11950 VDPWR.n292 VDPWR 0.0981562
R11951 VDPWR VDPWR.n1338 0.0981562
R11952 VDPWR.n1432 VDPWR 0.0981562
R11953 VDPWR.n1467 VDPWR 0.0981562
R11954 VDPWR.n1496 VDPWR 0.0981562
R11955 VDPWR VDPWR.n1274 0.0981562
R11956 VDPWR.n1759 VDPWR 0.0981562
R11957 VDPWR VDPWR.n1238 0.0981562
R11958 VDPWR.n1824 VDPWR 0.0981562
R11959 VDPWR.n1838 VDPWR 0.0981562
R11960 VDPWR VDPWR.n1641 0.0981562
R11961 VDPWR VDPWR.n2056 0.0981562
R11962 VDPWR VDPWR.n2054 0.0981562
R11963 VDPWR VDPWR.n2024 0.0981562
R11964 VDPWR.n2015 VDPWR 0.0981562
R11965 VDPWR VDPWR.n2002 0.0981562
R11966 VDPWR VDPWR.n1991 0.0981562
R11967 VDPWR VDPWR.n1962 0.0981562
R11968 VDPWR.n2143 VDPWR 0.0981562
R11969 VDPWR.n2169 VDPWR 0.0981562
R11970 VDPWR.n2175 VDPWR 0.0981562
R11971 VDPWR.n2181 VDPWR 0.0981562
R11972 VDPWR.n2224 VDPWR 0.0981562
R11973 VDPWR VDPWR.n2312 0.0981562
R11974 VDPWR VDPWR.n1004 0.0981562
R11975 VDPWR.n2825 VDPWR 0.0981562
R11976 VDPWR VDPWR.n966 0.0981562
R11977 VDPWR.n2646 VDPWR 0.0981562
R11978 VDPWR.n2382 VDPWR 0.0981562
R11979 VDPWR VDPWR.n2350 0.0981562
R11980 VDPWR VDPWR.n2522 0.0981562
R11981 VDPWR.n2440 VDPWR 0.0981562
R11982 VDPWR.n3088 VDPWR 0.0981562
R11983 VDPWR VDPWR.n3077 0.0981562
R11984 VDPWR VDPWR.n849 0.0981562
R11985 VDPWR.n34 VDPWR 0.0981562
R11986 VDPWR.n3103 VDPWR.n3102 0.0977722
R11987 VDPWR.n2508 VDPWR.n779 0.0977722
R11988 VDPWR.n2536 VDPWR.n2343 0.0977722
R11989 VDPWR.n3074 VDPWR.n770 0.0977722
R11990 VDPWR.n2832 VDPWR 0.0968542
R11991 VDPWR VDPWR.n3010 0.0968542
R11992 VDPWR.n628 VDPWR 0.0955521
R11993 VDPWR.n348 VDPWR 0.0955521
R11994 VDPWR.n90 VDPWR 0.0955521
R11995 VDPWR.n2695 VDPWR.n2589 0.0950946
R11996 VDPWR.n2690 VDPWR.n2592 0.0950946
R11997 VDPWR.n2665 VDPWR.n2615 0.0950946
R11998 VDPWR.n2660 VDPWR.n2618 0.0950946
R11999 VDPWR.n2509 VDPWR.n2444 0.0950946
R12000 VDPWR.n2494 VDPWR.n2446 0.0950946
R12001 VDPWR.n1490 VDPWR.n1489 0.0950946
R12002 VDPWR.n1494 VDPWR.n1299 0.0950946
R12003 VDPWR.n1454 VDPWR.n1453 0.0950946
R12004 VDPWR.n1458 VDPWR.n1316 0.0950946
R12005 VDPWR.n1421 VDPWR.n1420 0.0950946
R12006 VDPWR.n1425 VDPWR.n1330 0.0950946
R12007 VDPWR.n1373 VDPWR.n1371 0.0950946
R12008 VDPWR.n1386 VDPWR.n1345 0.0950946
R12009 VDPWR.n1556 VDPWR.n1530 0.0950946
R12010 VDPWR.n1546 VDPWR.n1544 0.0950946
R12011 VDPWR.n1586 VDPWR.n1585 0.0950946
R12012 VDPWR.n1579 VDPWR.n1290 0.0950946
R12013 VDPWR.n1818 VDPWR.n1817 0.0950946
R12014 VDPWR.n1822 VDPWR.n1226 0.0950946
R12015 VDPWR.n1782 VDPWR.n1781 0.0950946
R12016 VDPWR.n1786 VDPWR.n1243 0.0950946
R12017 VDPWR.n1752 VDPWR.n1751 0.0950946
R12018 VDPWR.n1756 VDPWR.n1265 0.0950946
R12019 VDPWR.n1712 VDPWR.n1711 0.0950946
R12020 VDPWR.n1716 VDPWR.n1281 0.0950946
R12021 VDPWR.n1889 VDPWR.n1887 0.0950946
R12022 VDPWR.n1900 VDPWR.n1195 0.0950946
R12023 VDPWR.n1856 VDPWR.n1855 0.0950946
R12024 VDPWR.n1862 VDPWR.n1861 0.0950946
R12025 VDPWR.n2008 VDPWR.n1160 0.0950946
R12026 VDPWR.n2004 VDPWR.n1164 0.0950946
R12027 VDPWR.n2037 VDPWR.n1136 0.0950946
R12028 VDPWR.n2032 VDPWR.n1139 0.0950946
R12029 VDPWR.n2070 VDPWR.n2069 0.0950946
R12030 VDPWR.n2063 VDPWR.n1123 0.0950946
R12031 VDPWR.n1670 VDPWR.n1669 0.0950946
R12032 VDPWR.n1662 VDPWR.n1661 0.0950946
R12033 VDPWR.n1955 VDPWR.n1930 0.0950946
R12034 VDPWR.n1945 VDPWR.n1943 0.0950946
R12035 VDPWR.n1978 VDPWR.n1188 0.0950946
R12036 VDPWR.n1972 VDPWR.n1910 0.0950946
R12037 VDPWR.n2329 VDPWR.n2328 0.0950946
R12038 VDPWR.n2321 VDPWR.n2320 0.0950946
R12039 VDPWR.n2247 VDPWR.n2246 0.0950946
R12040 VDPWR.n2239 VDPWR.n2238 0.0950946
R12041 VDPWR.n2157 VDPWR.n2156 0.0950946
R12042 VDPWR.n2162 VDPWR.n2161 0.0950946
R12043 VDPWR.n2112 VDPWR.n2110 0.0950946
R12044 VDPWR.n2126 VDPWR.n2086 0.0950946
R12045 VDPWR.n2261 VDPWR.n1078 0.0950946
R12046 VDPWR.n1088 VDPWR.n1082 0.0950946
R12047 VDPWR.n2294 VDPWR.n1043 0.0950946
R12048 VDPWR.n2288 VDPWR.n1048 0.0950946
R12049 VDPWR.n2880 VDPWR.n2878 0.0950946
R12050 VDPWR.n2898 VDPWR.n956 0.0950946
R12051 VDPWR.n2842 VDPWR.n2841 0.0950946
R12052 VDPWR.n2847 VDPWR.n2846 0.0950946
R12053 VDPWR.n2803 VDPWR.n2802 0.0950946
R12054 VDPWR.n2807 VDPWR.n986 0.0950946
R12055 VDPWR.n2753 VDPWR.n2752 0.0950946
R12056 VDPWR.n2757 VDPWR.n1007 0.0950946
R12057 VDPWR.n2966 VDPWR.n2964 0.0950946
R12058 VDPWR.n2977 VDPWR.n925 0.0950946
R12059 VDPWR.n2930 VDPWR.n2929 0.0950946
R12060 VDPWR.n2934 VDPWR.n941 0.0950946
R12061 VDPWR.n3036 VDPWR.n903 0.0950946
R12062 VDPWR.n3030 VDPWR.n906 0.0950946
R12063 VDPWR.n3065 VDPWR.n3064 0.0950946
R12064 VDPWR.n3057 VDPWR.n3056 0.0950946
R12065 VDPWR.n2465 VDPWR.n785 0.0950946
R12066 VDPWR.n3100 VDPWR.n784 0.0950946
R12067 VDPWR.n2571 VDPWR.n2549 0.0950946
R12068 VDPWR.n2717 VDPWR.n2542 0.0950946
R12069 VDPWR.n3008 VDPWR.n922 0.0950946
R12070 VDPWR.n3003 VDPWR.n2985 0.0950946
R12071 VDPWR.n2426 VDPWR.n2344 0.0950946
R12072 VDPWR.n2534 VDPWR.n2342 0.0950946
R12073 VDPWR.n2391 VDPWR.n2390 0.0950946
R12074 VDPWR.n2394 VDPWR.n2393 0.0950946
R12075 VDPWR.n847 VDPWR.n846 0.0950946
R12076 VDPWR.n839 VDPWR.n772 0.0950946
R12077 VDPWR.n3075 VDPWR.n802 0.0950946
R12078 VDPWR.n868 VDPWR.n804 0.0950946
R12079 VDPWR VDPWR.n2104 0.0930646
R12080 VDPWR.n586 VDPWR.n568 0.0916458
R12081 VDPWR.n306 VDPWR.n288 0.0916458
R12082 VDPWR.n48 VDPWR.n30 0.0916458
R12083 VDPWR.n3104 VDPWR.n3103 0.0913766
R12084 VDPWR.n3106 VDPWR.n3105 0.0913766
R12085 VDPWR.n3171 VDPWR.n759 0.08675
R12086 VDPWR.n1974 VDPWR.n1908 0.086275
R12087 VDPWR.n2006 VDPWR.n1162 0.086275
R12088 VDPWR.n1246 VDPWR.n1091 0.086275
R12089 VDPWR.n1675 VDPWR.n1672 0.086275
R12090 VDPWR.n1905 VDPWR.n1089 0.086275
R12091 VDPWR.n2072 VDPWR.n1116 0.086275
R12092 VDPWR.n3149 VDPWR.n3134 0.0848934
R12093 VDPWR.n3165 VDPWR.n3150 0.0844041
R12094 VDPWR.n1374 VDPWR.n1370 0.0838333
R12095 VDPWR.n1387 VDPWR.n1344 0.0838333
R12096 VDPWR.n1419 VDPWR.n1418 0.0838333
R12097 VDPWR.n1450 VDPWR.n1315 0.0838333
R12098 VDPWR.n1488 VDPWR.n1302 0.0838333
R12099 VDPWR.n1584 VDPWR.n1583 0.0838333
R12100 VDPWR.n1547 VDPWR.n1536 0.0838333
R12101 VDPWR.n1710 VDPWR.n1677 0.0838333
R12102 VDPWR.n1717 VDPWR.n1280 0.0838333
R12103 VDPWR.n1750 VDPWR.n1749 0.0838333
R12104 VDPWR.n1254 VDPWR.n1251 0.0838333
R12105 VDPWR.n1816 VDPWR.n1230 0.0838333
R12106 VDPWR.n1854 VDPWR.n1853 0.0838333
R12107 VDPWR.n1899 VDPWR.n1898 0.0838333
R12108 VDPWR.n1668 VDPWR.n1598 0.0838333
R12109 VDPWR.n1663 VDPWR.n1657 0.0838333
R12110 VDPWR.n2068 VDPWR.n2067 0.0838333
R12111 VDPWR.n1146 VDPWR.n1144 0.0838333
R12112 VDPWR.n2009 VDPWR.n1159 0.0838333
R12113 VDPWR.n1946 VDPWR.n1935 0.0838333
R12114 VDPWR.n2113 VDPWR.n2089 0.0838333
R12115 VDPWR.n2127 VDPWR.n2085 0.0838333
R12116 VDPWR.n2155 VDPWR.n2154 0.0838333
R12117 VDPWR.n2197 VDPWR.n1097 0.0838333
R12118 VDPWR.n2327 VDPWR.n1015 0.0838333
R12119 VDPWR.n2295 VDPWR.n1042 0.0838333
R12120 VDPWR.n1087 VDPWR.n1085 0.0838333
R12121 VDPWR.n2751 VDPWR.n2721 0.0838333
R12122 VDPWR.n2801 VDPWR.n2800 0.0838333
R12123 VDPWR.n2848 VDPWR.n970 0.0838333
R12124 VDPWR.n2881 VDPWR.n2877 0.0838333
R12125 VDPWR.n2928 VDPWR.n2927 0.0838333
R12126 VDPWR.n2976 VDPWR.n2975 0.0838333
R12127 VDPWR.n2570 VDPWR.n2569 0.0838333
R12128 VDPWR.n2716 VDPWR.n2543 0.0838333
R12129 VDPWR.n2654 VDPWR.n2653 0.0838333
R12130 VDPWR.n3063 VDPWR.n875 0.0838333
R12131 VDPWR.n3037 VDPWR.n902 0.0838333
R12132 VDPWR.n3002 VDPWR.n2986 0.0838333
R12133 VDPWR.n2389 VDPWR.n2365 0.0838333
R12134 VDPWR.n2395 VDPWR.n2361 0.0838333
R12135 VDPWR.n2496 VDPWR.n2495 0.0838333
R12136 VDPWR.n841 VDPWR.n840 0.0838333
R12137 VDPWR.n777 VDPWR 0.08275
R12138 VDPWR.n781 VDPWR 0.08275
R12139 VDPWR.n2500 VDPWR 0.08275
R12140 VDPWR.n3112 VDPWR 0.08275
R12141 VDPWR.n2340 VDPWR 0.08275
R12142 VDPWR VDPWR.n1915 0.082648
R12143 VDPWR VDPWR.n2624 0.082648
R12144 VDPWR VDPWR.n1764 0.082648
R12145 VDPWR.n1765 VDPWR 0.082648
R12146 VDPWR.n1794 VDPWR 0.082648
R12147 VDPWR.n2476 VDPWR 0.082648
R12148 VDPWR VDPWR.n2460 0.082648
R12149 VDPWR.n1427 VDPWR.n1426 0.0812292
R12150 VDPWR.n1460 VDPWR.n1459 0.0812292
R12151 VDPWR.n1483 VDPWR.n1298 0.0812292
R12152 VDPWR.n1578 VDPWR.n1289 0.0812292
R12153 VDPWR.n1551 VDPWR.n1550 0.0812292
R12154 VDPWR.n1758 VDPWR.n1757 0.0812292
R12155 VDPWR.n1787 VDPWR.n1242 0.0812292
R12156 VDPWR.n1811 VDPWR.n1225 0.0812292
R12157 VDPWR.n1863 VDPWR.n1214 0.0812292
R12158 VDPWR.n1891 VDPWR.n1198 0.0812292
R12159 VDPWR.n2057 VDPWR.n1124 0.0812292
R12160 VDPWR.n2031 VDPWR.n1140 0.0812292
R12161 VDPWR.n1174 VDPWR.n1165 0.0812292
R12162 VDPWR.n1913 VDPWR.n1912 0.0812292
R12163 VDPWR.n1950 VDPWR.n1949 0.0812292
R12164 VDPWR.n2168 VDPWR.n1111 0.0812292
R12165 VDPWR.n2241 VDPWR.n2240 0.0812292
R12166 VDPWR.n2322 VDPWR.n1020 0.0812292
R12167 VDPWR.n1054 VDPWR.n1053 0.0812292
R12168 VDPWR.n1084 VDPWR.n1083 0.0812292
R12169 VDPWR.n2809 VDPWR.n2808 0.0812292
R12170 VDPWR.n2849 VDPWR.n968 0.0812292
R12171 VDPWR.n960 VDPWR.n955 0.0812292
R12172 VDPWR.n2924 VDPWR.n940 0.0812292
R12173 VDPWR.n2968 VDPWR.n928 0.0812292
R12174 VDPWR.n2689 VDPWR.n2688 0.0812292
R12175 VDPWR.n3058 VDPWR.n880 0.0812292
R12176 VDPWR.n910 VDPWR.n909 0.0812292
R12177 VDPWR.n2996 VDPWR.n2995 0.0812292
R12178 VDPWR.n2529 VDPWR.n2346 0.0812292
R12179 VDPWR.n2493 VDPWR.n2449 0.0812292
R12180 VDPWR.n3099 VDPWR.n3098 0.0812292
R12181 VDPWR.n835 VDPWR.n829 0.0812292
R12182 VDPWR.n536 VDPWR 0.0800455
R12183 VDPWR.n1415 VDPWR.n1336 0.0760208
R12184 VDPWR.n1487 VDPWR.n1306 0.0760208
R12185 VDPWR.n1746 VDPWR.n1272 0.0760208
R12186 VDPWR.n1815 VDPWR.n1234 0.0760208
R12187 VDPWR.n1867 VDPWR.n1212 0.0760208
R12188 VDPWR.n2062 VDPWR.n1122 0.0760208
R12189 VDPWR.n1173 VDPWR.n1169 0.0760208
R12190 VDPWR.n1971 VDPWR.n1970 0.0760208
R12191 VDPWR.n2163 VDPWR.n1113 0.0760208
R12192 VDPWR.n2326 VDPWR.n1017 0.0760208
R12193 VDPWR.n2287 VDPWR.n2286 0.0760208
R12194 VDPWR.n2797 VDPWR.n994 0.0760208
R12195 VDPWR.n2893 VDPWR.n959 0.0760208
R12196 VDPWR.n2935 VDPWR.n938 0.0760208
R12197 VDPWR.n2602 VDPWR.n2601 0.0760208
R12198 VDPWR.n3062 VDPWR.n877 0.0760208
R12199 VDPWR.n3029 VDPWR.n3028 0.0760208
R12200 VDPWR.n862 VDPWR.n806 0.0760208
R12201 VDPWR.n1908 VDPWR.n1191 0.074525
R12202 VDPWR.n1820 VDPWR.n1162 0.074525
R12203 VDPWR.n1784 VDPWR.n1246 0.074525
R12204 VDPWR.n1714 VDPWR.n1675 0.074525
R12205 VDPWR.n1905 VDPWR.n1904 0.074525
R12206 VDPWR.n1754 VDPWR.n1116 0.074525
R12207 VDPWR.n753 VDPWR 0.0710357
R12208 VDPWR.n1381 VDPWR.n1348 0.0708125
R12209 VDPWR.n1452 VDPWR.n1447 0.0708125
R12210 VDPWR.n1709 VDPWR.n1681 0.0708125
R12211 VDPWR.n1780 VDPWR.n1250 0.0708125
R12212 VDPWR.n1845 VDPWR.n1217 0.0708125
R12213 VDPWR.n1667 VDPWR.n1600 0.0708125
R12214 VDPWR.n1143 VDPWR.n1135 0.0708125
R12215 VDPWR.n1187 VDPWR.n1185 0.0708125
R12216 VDPWR.n2121 VDPWR.n2119 0.0708125
R12217 VDPWR.n2245 VDPWR.n1096 0.0708125
R12218 VDPWR.n2299 VDPWR.n1037 0.0708125
R12219 VDPWR.n2750 VDPWR.n2725 0.0708125
R12220 VDPWR.n2840 VDPWR.n2838 0.0708125
R12221 VDPWR.n2920 VDPWR.n945 0.0708125
R12222 VDPWR.n2576 VDPWR.n2548 0.0708125
R12223 VDPWR.n2650 VDPWR.n2614 0.0708125
R12224 VDPWR.n901 VDPWR.n898 0.0708125
R12225 VDPWR.n3077 VDPWR.n3076 0.0708125
R12226 VDPWR.n2599 VDPWR.n2590 0.0680676
R12227 VDPWR.n2599 VDPWR.n2591 0.0680676
R12228 VDPWR.n2652 VDPWR.n2616 0.0680676
R12229 VDPWR.n2652 VDPWR.n2617 0.0680676
R12230 VDPWR.n2498 VDPWR.n2497 0.0680676
R12231 VDPWR.n2497 VDPWR.n2445 0.0680676
R12232 VDPWR.n1305 VDPWR.n1303 0.0680676
R12233 VDPWR.n1305 VDPWR.n1304 0.0680676
R12234 VDPWR.n1449 VDPWR.n1320 0.0680676
R12235 VDPWR.n1449 VDPWR.n1448 0.0680676
R12236 VDPWR.n1417 VDPWR.n1334 0.0680676
R12237 VDPWR.n1417 VDPWR.n1416 0.0680676
R12238 VDPWR.n1382 VDPWR.n1347 0.0680676
R12239 VDPWR.n1383 VDPWR.n1382 0.0680676
R12240 VDPWR.n1553 VDPWR.n1552 0.0680676
R12241 VDPWR.n1552 VDPWR.n1533 0.0680676
R12242 VDPWR.n1582 VDPWR.n1288 0.0680676
R12243 VDPWR.n1582 VDPWR.n1581 0.0680676
R12244 VDPWR.n1233 VDPWR.n1231 0.0680676
R12245 VDPWR.n1233 VDPWR.n1232 0.0680676
R12246 VDPWR.n1253 VDPWR.n1249 0.0680676
R12247 VDPWR.n1253 VDPWR.n1252 0.0680676
R12248 VDPWR.n1748 VDPWR.n1270 0.0680676
R12249 VDPWR.n1748 VDPWR.n1747 0.0680676
R12250 VDPWR.n1680 VDPWR.n1678 0.0680676
R12251 VDPWR.n1680 VDPWR.n1679 0.0680676
R12252 VDPWR.n1888 VDPWR.n1197 0.0680676
R12253 VDPWR.n1901 VDPWR.n1197 0.0680676
R12254 VDPWR.n1852 VDPWR.n1216 0.0680676
R12255 VDPWR.n1852 VDPWR.n1215 0.0680676
R12256 VDPWR.n1172 VDPWR.n1170 0.0680676
R12257 VDPWR.n1172 VDPWR.n1171 0.0680676
R12258 VDPWR.n1145 VDPWR.n1137 0.0680676
R12259 VDPWR.n1145 VDPWR.n1138 0.0680676
R12260 VDPWR.n2066 VDPWR.n1120 0.0680676
R12261 VDPWR.n2066 VDPWR.n2065 0.0680676
R12262 VDPWR.n1658 VDPWR.n1599 0.0680676
R12263 VDPWR.n1660 VDPWR.n1658 0.0680676
R12264 VDPWR.n1952 VDPWR.n1951 0.0680676
R12265 VDPWR.n1951 VDPWR.n1932 0.0680676
R12266 VDPWR.n1977 VDPWR.n1189 0.0680676
R12267 VDPWR.n1909 VDPWR.n1189 0.0680676
R12268 VDPWR.n1021 VDPWR.n1016 0.0680676
R12269 VDPWR.n1023 VDPWR.n1021 0.0680676
R12270 VDPWR.n2235 VDPWR.n1095 0.0680676
R12271 VDPWR.n2237 VDPWR.n2235 0.0680676
R12272 VDPWR.n2153 VDPWR.n2076 0.0680676
R12273 VDPWR.n2153 VDPWR.n1114 0.0680676
R12274 VDPWR.n2122 VDPWR.n2088 0.0680676
R12275 VDPWR.n2123 VDPWR.n2122 0.0680676
R12276 VDPWR.n2260 VDPWR.n1079 0.0680676
R12277 VDPWR.n1081 VDPWR.n1079 0.0680676
R12278 VDPWR.n2293 VDPWR.n1044 0.0680676
R12279 VDPWR.n1047 VDPWR.n1044 0.0680676
R12280 VDPWR.n2894 VDPWR.n958 0.0680676
R12281 VDPWR.n2895 VDPWR.n2894 0.0680676
R12282 VDPWR.n978 VDPWR.n977 0.0680676
R12283 VDPWR.n977 VDPWR.n971 0.0680676
R12284 VDPWR.n2799 VDPWR.n992 0.0680676
R12285 VDPWR.n2799 VDPWR.n2798 0.0680676
R12286 VDPWR.n2724 VDPWR.n2722 0.0680676
R12287 VDPWR.n2724 VDPWR.n2723 0.0680676
R12288 VDPWR.n2965 VDPWR.n927 0.0680676
R12289 VDPWR.n2978 VDPWR.n927 0.0680676
R12290 VDPWR.n2926 VDPWR.n946 0.0680676
R12291 VDPWR.n2926 VDPWR.n2925 0.0680676
R12292 VDPWR.n3035 VDPWR.n904 0.0680676
R12293 VDPWR.n905 VDPWR.n904 0.0680676
R12294 VDPWR.n881 VDPWR.n876 0.0680676
R12295 VDPWR.n883 VDPWR.n881 0.0680676
R12296 VDPWR.n786 VDPWR.n783 0.0680676
R12297 VDPWR.n3101 VDPWR.n786 0.0680676
R12298 VDPWR.n2575 VDPWR.n2573 0.0680676
R12299 VDPWR.n2575 VDPWR.n2574 0.0680676
R12300 VDPWR.n2994 VDPWR.n2983 0.0680676
R12301 VDPWR.n2994 VDPWR.n2984 0.0680676
R12302 VDPWR.n2345 VDPWR.n2341 0.0680676
R12303 VDPWR.n2535 VDPWR.n2345 0.0680676
R12304 VDPWR.n2364 VDPWR.n2363 0.0680676
R12305 VDPWR.n2363 VDPWR.n2362 0.0680676
R12306 VDPWR.n828 VDPWR.n773 0.0680676
R12307 VDPWR.n828 VDPWR.n774 0.0680676
R12308 VDPWR.n805 VDPWR.n803 0.0680676
R12309 VDPWR.n869 VDPWR.n805 0.0680676
R12310 VDPWR.n1409 VDPWR.n1333 0.0656042
R12311 VDPWR.n1739 VDPWR.n1269 0.0656042
R12312 VDPWR.n1635 VDPWR.n1119 0.0656042
R12313 VDPWR.n2149 VDPWR.n2075 0.0656042
R12314 VDPWR.n2787 VDPWR.n991 0.0656042
R12315 VDPWR.n2697 VDPWR.n2696 0.0656042
R12316 VDPWR.n2424 VDPWR.n2423 0.0656042
R12317 VDPWR.n718 VDPWR 0.06425
R12318 VDPWR.n702 VDPWR 0.06425
R12319 VDPWR.n686 VDPWR 0.06425
R12320 VDPWR.n670 VDPWR 0.06425
R12321 VDPWR.n529 VDPWR 0.06425
R12322 VDPWR.n513 VDPWR 0.06425
R12323 VDPWR.n497 VDPWR 0.06425
R12324 VDPWR.n481 VDPWR 0.06425
R12325 VDPWR.n465 VDPWR 0.06425
R12326 VDPWR.n389 VDPWR 0.06425
R12327 VDPWR.n401 VDPWR 0.06425
R12328 VDPWR.n459 VDPWR 0.06425
R12329 VDPWR.n443 VDPWR 0.06425
R12330 VDPWR.n427 VDPWR 0.06425
R12331 VDPWR.n3170 VDPWR 0.06425
R12332 VDPWR.n3164 VDPWR 0.06425
R12333 VDPWR.n3148 VDPWR 0.06425
R12334 VDPWR.n3132 VDPWR 0.06425
R12335 VDPWR.n256 VDPWR.n253 0.061697
R12336 VDPWR.n754 VDPWR 0.0615066
R12337 VDPWR.n620 VDPWR 0.0603958
R12338 VDPWR VDPWR.n619 0.0603958
R12339 VDPWR.n614 VDPWR 0.0603958
R12340 VDPWR.n609 VDPWR 0.0603958
R12341 VDPWR.n604 VDPWR 0.0603958
R12342 VDPWR.n580 VDPWR 0.0603958
R12343 VDPWR VDPWR.n579 0.0603958
R12344 VDPWR VDPWR.n563 0.0603958
R12345 VDPWR.n639 VDPWR 0.0603958
R12346 VDPWR VDPWR.n638 0.0603958
R12347 VDPWR.n648 VDPWR 0.0603958
R12348 VDPWR.n558 VDPWR 0.0603958
R12349 VDPWR.n340 VDPWR 0.0603958
R12350 VDPWR VDPWR.n339 0.0603958
R12351 VDPWR.n334 VDPWR 0.0603958
R12352 VDPWR.n329 VDPWR 0.0603958
R12353 VDPWR.n324 VDPWR 0.0603958
R12354 VDPWR.n300 VDPWR 0.0603958
R12355 VDPWR VDPWR.n299 0.0603958
R12356 VDPWR VDPWR.n283 0.0603958
R12357 VDPWR.n359 VDPWR 0.0603958
R12358 VDPWR VDPWR.n358 0.0603958
R12359 VDPWR.n368 VDPWR 0.0603958
R12360 VDPWR.n278 VDPWR 0.0603958
R12361 VDPWR.n1369 VDPWR 0.0603958
R12362 VDPWR.n1395 VDPWR 0.0603958
R12363 VDPWR.n1436 VDPWR 0.0603958
R12364 VDPWR.n1497 VDPWR 0.0603958
R12365 VDPWR.n1500 VDPWR 0.0603958
R12366 VDPWR.n1501 VDPWR 0.0603958
R12367 VDPWR.n1574 VDPWR 0.0603958
R12368 VDPWR.n1702 VDPWR 0.0603958
R12369 VDPWR.n1725 VDPWR 0.0603958
R12370 VDPWR.n1763 VDPWR 0.0603958
R12371 VDPWR VDPWR.n1256 0.0603958
R12372 VDPWR.n1831 VDPWR 0.0603958
R12373 VDPWR.n1837 VDPWR 0.0603958
R12374 VDPWR.n1883 VDPWR 0.0603958
R12375 VDPWR VDPWR.n1608 0.0603958
R12376 VDPWR.n1648 VDPWR 0.0603958
R12377 VDPWR.n2039 VDPWR 0.0603958
R12378 VDPWR.n1999 VDPWR 0.0603958
R12379 VDPWR VDPWR.n1992 0.0603958
R12380 VDPWR.n1985 VDPWR 0.0603958
R12381 VDPWR.n1965 VDPWR 0.0603958
R12382 VDPWR VDPWR.n1963 0.0603958
R12383 VDPWR.n1957 VDPWR 0.0603958
R12384 VDPWR.n2105 VDPWR 0.0603958
R12385 VDPWR.n2109 VDPWR 0.0603958
R12386 VDPWR VDPWR.n2081 0.0603958
R12387 VDPWR.n2170 VDPWR 0.0603958
R12388 VDPWR.n2174 VDPWR 0.0603958
R12389 VDPWR.n2183 VDPWR 0.0603958
R12390 VDPWR.n2217 VDPWR 0.0603958
R12391 VDPWR.n2214 VDPWR 0.0603958
R12392 VDPWR VDPWR.n2213 0.0603958
R12393 VDPWR VDPWR.n2318 0.0603958
R12394 VDPWR.n2314 VDPWR 0.0603958
R12395 VDPWR VDPWR.n2313 0.0603958
R12396 VDPWR.n2272 VDPWR 0.0603958
R12397 VDPWR.n2269 VDPWR 0.0603958
R12398 VDPWR.n2737 VDPWR 0.0603958
R12399 VDPWR.n2745 VDPWR 0.0603958
R12400 VDPWR.n2765 VDPWR 0.0603958
R12401 VDPWR VDPWR.n999 0.0603958
R12402 VDPWR.n2810 VDPWR 0.0603958
R12403 VDPWR.n2818 VDPWR 0.0603958
R12404 VDPWR.n2820 VDPWR 0.0603958
R12405 VDPWR VDPWR.n2826 0.0603958
R12406 VDPWR.n2827 VDPWR 0.0603958
R12407 VDPWR.n2831 VDPWR 0.0603958
R12408 VDPWR VDPWR.n2856 0.0603958
R12409 VDPWR.n2857 VDPWR 0.0603958
R12410 VDPWR VDPWR.n2869 0.0603958
R12411 VDPWR.n2870 VDPWR 0.0603958
R12412 VDPWR.n2870 VDPWR 0.0603958
R12413 VDPWR.n2876 VDPWR 0.0603958
R12414 VDPWR.n2882 VDPWR 0.0603958
R12415 VDPWR.n2900 VDPWR 0.0603958
R12416 VDPWR.n2901 VDPWR 0.0603958
R12417 VDPWR.n2905 VDPWR 0.0603958
R12418 VDPWR.n2948 VDPWR 0.0603958
R12419 VDPWR.n2954 VDPWR 0.0603958
R12420 VDPWR.n2568 VDPWR 0.0603958
R12421 VDPWR.n2604 VDPWR 0.0603958
R12422 VDPWR.n2682 VDPWR 0.0603958
R12423 VDPWR.n2640 VDPWR 0.0603958
R12424 VDPWR.n2640 VDPWR 0.0603958
R12425 VDPWR VDPWR.n2639 0.0603958
R12426 VDPWR.n2631 VDPWR 0.0603958
R12427 VDPWR VDPWR.n2630 0.0603958
R12428 VDPWR VDPWR.n3054 0.0603958
R12429 VDPWR.n3049 VDPWR 0.0603958
R12430 VDPWR.n3047 VDPWR 0.0603958
R12431 VDPWR.n895 VDPWR 0.0603958
R12432 VDPWR.n3017 VDPWR 0.0603958
R12433 VDPWR.n3011 VDPWR 0.0603958
R12434 VDPWR.n2379 VDPWR 0.0603958
R12435 VDPWR.n2383 VDPWR 0.0603958
R12436 VDPWR.n2384 VDPWR 0.0603958
R12437 VDPWR.n2388 VDPWR 0.0603958
R12438 VDPWR VDPWR.n2402 0.0603958
R12439 VDPWR.n2403 VDPWR 0.0603958
R12440 VDPWR VDPWR.n2354 0.0603958
R12441 VDPWR VDPWR.n2408 0.0603958
R12442 VDPWR.n2409 VDPWR 0.0603958
R12443 VDPWR.n2413 VDPWR 0.0603958
R12444 VDPWR VDPWR.n2414 0.0603958
R12445 VDPWR.n2415 VDPWR 0.0603958
R12446 VDPWR.n2529 VDPWR 0.0603958
R12447 VDPWR VDPWR.n2528 0.0603958
R12448 VDPWR VDPWR.n2527 0.0603958
R12449 VDPWR.n2523 VDPWR 0.0603958
R12450 VDPWR.n2439 VDPWR 0.0603958
R12451 VDPWR VDPWR.n2440 0.0603958
R12452 VDPWR.n2511 VDPWR 0.0603958
R12453 VDPWR.n2511 VDPWR 0.0603958
R12454 VDPWR.n2482 VDPWR 0.0603958
R12455 VDPWR VDPWR.n2457 0.0603958
R12456 VDPWR.n2477 VDPWR 0.0603958
R12457 VDPWR.n790 VDPWR 0.0603958
R12458 VDPWR.n3094 VDPWR 0.0603958
R12459 VDPWR VDPWR.n3093 0.0603958
R12460 VDPWR VDPWR.n794 0.0603958
R12461 VDPWR.n3082 VDPWR 0.0603958
R12462 VDPWR.n3078 VDPWR 0.0603958
R12463 VDPWR VDPWR.n861 0.0603958
R12464 VDPWR.n855 VDPWR 0.0603958
R12465 VDPWR VDPWR.n853 0.0603958
R12466 VDPWR.n850 VDPWR 0.0603958
R12467 VDPWR.n82 VDPWR 0.0603958
R12468 VDPWR VDPWR.n81 0.0603958
R12469 VDPWR.n76 VDPWR 0.0603958
R12470 VDPWR.n71 VDPWR 0.0603958
R12471 VDPWR.n66 VDPWR 0.0603958
R12472 VDPWR.n42 VDPWR 0.0603958
R12473 VDPWR VDPWR.n41 0.0603958
R12474 VDPWR VDPWR.n25 0.0603958
R12475 VDPWR.n101 VDPWR 0.0603958
R12476 VDPWR VDPWR.n100 0.0603958
R12477 VDPWR.n110 VDPWR 0.0603958
R12478 VDPWR.n20 VDPWR 0.0603958
R12479 VDPWR.n3115 VDPWR.n3114 0.0600933
R12480 VDPWR.n561 VDPWR 0.0590938
R12481 VDPWR.n281 VDPWR 0.0590938
R12482 VDPWR.n23 VDPWR 0.0590938
R12483 VDPWR.n3166 VDPWR.n759 0.0589638
R12484 VDPWR.n1911 VDPWR 0.0577917
R12485 VDPWR.n2758 VDPWR 0.0577917
R12486 VDPWR.n810 VDPWR 0.0577917
R12487 VDPWR.n2693 VDPWR.n2692 0.0574697
R12488 VDPWR.n2663 VDPWR.n2662 0.0574697
R12489 VDPWR.n1301 VDPWR.n1300 0.0574697
R12490 VDPWR.n1318 VDPWR.n1317 0.0574697
R12491 VDPWR.n1332 VDPWR.n1331 0.0574697
R12492 VDPWR.n1384 VDPWR.n1346 0.0574697
R12493 VDPWR.n1554 VDPWR.n1532 0.0574697
R12494 VDPWR.n1580 VDPWR.n1286 0.0574697
R12495 VDPWR.n1229 VDPWR.n1227 0.0574697
R12496 VDPWR.n1247 VDPWR.n1244 0.0574697
R12497 VDPWR.n1268 VDPWR.n1266 0.0574697
R12498 VDPWR.n1676 VDPWR.n1282 0.0574697
R12499 VDPWR.n1902 VDPWR.n1196 0.0574697
R12500 VDPWR.n1859 VDPWR.n1858 0.0574697
R12501 VDPWR.n1163 VDPWR.n1161 0.0574697
R12502 VDPWR.n2035 VDPWR.n2034 0.0574697
R12503 VDPWR.n2064 VDPWR.n1118 0.0574697
R12504 VDPWR.n1659 VDPWR.n1597 0.0574697
R12505 VDPWR.n1953 VDPWR.n1931 0.0574697
R12506 VDPWR.n1976 VDPWR.n1190 0.0574697
R12507 VDPWR.n1022 VDPWR.n1014 0.0574697
R12508 VDPWR.n2236 VDPWR.n1093 0.0574697
R12509 VDPWR.n2074 VDPWR.n1115 0.0574697
R12510 VDPWR.n2124 VDPWR.n2087 0.0574697
R12511 VDPWR.n2259 VDPWR.n2258 0.0574697
R12512 VDPWR.n2292 VDPWR.n1045 0.0574697
R12513 VDPWR.n2896 VDPWR.n957 0.0574697
R12514 VDPWR.n975 VDPWR.n972 0.0574697
R12515 VDPWR.n990 VDPWR.n987 0.0574697
R12516 VDPWR.n2720 VDPWR.n1008 0.0574697
R12517 VDPWR.n2979 VDPWR.n926 0.0574697
R12518 VDPWR.n944 VDPWR.n942 0.0574697
R12519 VDPWR.n3034 VDPWR.n3032 0.0574697
R12520 VDPWR.n882 VDPWR.n874 0.0574697
R12521 VDPWR.n2572 VDPWR.n2338 0.0574697
R12522 VDPWR.n2718 VDPWR.n2541 0.0574697
R12523 VDPWR.n3006 VDPWR.n3005 0.0574697
R12524 VDPWR.n1335 VDPWR.n1333 0.0551875
R12525 VDPWR.n1271 VDPWR.n1269 0.0551875
R12526 VDPWR.n1121 VDPWR.n1119 0.0551875
R12527 VDPWR.n2152 VDPWR.n2075 0.0551875
R12528 VDPWR.n993 VDPWR.n991 0.0551875
R12529 VDPWR.n2696 VDPWR.n2588 0.0551875
R12530 VDPWR.n2425 VDPWR.n2424 0.0551875
R12531 VDPWR.n752 VDPWR.n751 0.0540714
R12532 VDPWR.n466 VDPWR.n403 0.054
R12533 VDPWR.n1534 VDPWR 0.0538854
R12534 VDPWR.n2533 VDPWR 0.0538854
R12535 VDPWR VDPWR.n2467 0.0538854
R12536 VDPWR.n3176 VDPWR 0.0535303
R12537 VDPWR.n3116 VDPWR.n3115 0.0529556
R12538 VDPWR.n653 VDPWR 0.0525833
R12539 VDPWR.n373 VDPWR 0.0525833
R12540 VDPWR VDPWR.n1956 0.0525833
R12541 VDPWR.n2600 VDPWR 0.0525833
R12542 VDPWR.n2428 VDPWR 0.0525833
R12543 VDPWR.n2466 VDPWR 0.0525833
R12544 VDPWR.n115 VDPWR 0.0525833
R12545 VDPWR.n2290 VDPWR.n1046 0.0522
R12546 VDPWR.n2331 VDPWR.n1012 0.0522
R12547 VDPWR.n2250 VDPWR.n2249 0.0522
R12548 VDPWR.n1596 VDPWR.n1009 0.0522
R12549 VDPWR.n2256 VDPWR.n2255 0.0522
R12550 VDPWR.n2159 VDPWR.n2073 0.0522
R12551 VDPWR.n2507 VDPWR.n2506 0.051025
R12552 VDPWR VDPWR.n754 0.0500269
R12553 VDPWR.n1381 VDPWR.n1380 0.0499792
R12554 VDPWR.n1452 VDPWR.n1451 0.0499792
R12555 VDPWR.n1517 VDPWR.n1287 0.0499792
R12556 VDPWR.n1706 VDPWR.n1681 0.0499792
R12557 VDPWR.n1780 VDPWR.n1779 0.0499792
R12558 VDPWR.n1851 VDPWR.n1217 0.0499792
R12559 VDPWR.n1664 VDPWR.n1600 0.0499792
R12560 VDPWR.n1147 VDPWR.n1143 0.0499792
R12561 VDPWR VDPWR.n1187 0.0499792
R12562 VDPWR.n2121 VDPWR.n2120 0.0499792
R12563 VDPWR.n2245 VDPWR.n2244 0.0499792
R12564 VDPWR.n2296 VDPWR.n1037 0.0499792
R12565 VDPWR.n2748 VDPWR.n2725 0.0499792
R12566 VDPWR.n2840 VDPWR.n2839 0.0499792
R12567 VDPWR.n947 VDPWR.n945 0.0499792
R12568 VDPWR.n2577 VDPWR.n2576 0.0499792
R12569 VDPWR.n2651 VDPWR.n2650 0.0499792
R12570 VDPWR.n3038 VDPWR.n901 0.0499792
R12571 VDPWR.n2396 VDPWR.n2360 0.0499792
R12572 VDPWR.n2448 VDPWR.n2447 0.0499792
R12573 VDPWR.n3076 VDPWR.n801 0.0499792
R12574 VDPWR VDPWR.n2510 0.047375
R12575 VDPWR.n653 VDPWR.n652 0.0460729
R12576 VDPWR.n373 VDPWR.n372 0.0460729
R12577 VDPWR.n115 VDPWR.n114 0.0460729
R12578 VDPWR.n3108 VDPWR.n777 0.0460404
R12579 VDPWR.n781 VDPWR.n780 0.0460404
R12580 VDPWR.n3112 VDPWR.n3111 0.0460404
R12581 VDPWR.n2501 VDPWR.n2500 0.0454816
R12582 VDPWR.n1336 VDPWR.n1329 0.0447708
R12583 VDPWR.n1484 VDPWR.n1306 0.0447708
R12584 VDPWR.n1535 VDPWR.n1534 0.0447708
R12585 VDPWR.n1272 VDPWR.n1264 0.0447708
R12586 VDPWR.n1812 VDPWR.n1234 0.0447708
R12587 VDPWR.n1892 VDPWR.n1890 0.0447708
R12588 VDPWR.n2062 VDPWR.n2061 0.0447708
R12589 VDPWR.n1175 VDPWR.n1173 0.0447708
R12590 VDPWR.n1971 VDPWR.n1914 0.0447708
R12591 VDPWR.n1934 VDPWR.n1933 0.0447708
R12592 VDPWR.n2164 VDPWR.n2163 0.0447708
R12593 VDPWR.n2323 VDPWR.n1017 0.0447708
R12594 VDPWR.n2262 VDPWR.n1077 0.0447708
R12595 VDPWR.n994 VDPWR.n985 0.0447708
R12596 VDPWR.n2893 VDPWR.n2892 0.0447708
R12597 VDPWR.n2969 VDPWR.n2967 0.0447708
R12598 VDPWR.n2601 VDPWR.n2593 0.0447708
R12599 VDPWR.n3059 VDPWR.n877 0.0447708
R12600 VDPWR.n3029 VDPWR.n907 0.0447708
R12601 VDPWR.n2993 VDPWR.n2992 0.0447708
R12602 VDPWR.n2533 VDPWR.n2532 0.0447708
R12603 VDPWR.n2467 VDPWR.n787 0.0447708
R12604 VDPWR.n866 VDPWR.n806 0.0447708
R12605 VDPWR.n845 VDPWR.n844 0.0447708
R12606 VDPWR.n2503 VDPWR.n2340 0.0446687
R12607 VDPWR.n2590 VDPWR.n2589 0.0410405
R12608 VDPWR.n2592 VDPWR.n2591 0.0410405
R12609 VDPWR.n2616 VDPWR.n2615 0.0410405
R12610 VDPWR.n2618 VDPWR.n2617 0.0410405
R12611 VDPWR.n2498 VDPWR.n2444 0.0410405
R12612 VDPWR.n2494 VDPWR.n2445 0.0410405
R12613 VDPWR.n1489 VDPWR.n1303 0.0410405
R12614 VDPWR.n1304 VDPWR.n1299 0.0410405
R12615 VDPWR.n1453 VDPWR.n1320 0.0410405
R12616 VDPWR.n1448 VDPWR.n1316 0.0410405
R12617 VDPWR.n1420 VDPWR.n1334 0.0410405
R12618 VDPWR.n1416 VDPWR.n1330 0.0410405
R12619 VDPWR.n1371 VDPWR.n1347 0.0410405
R12620 VDPWR.n1383 VDPWR.n1345 0.0410405
R12621 VDPWR.n1553 VDPWR.n1530 0.0410405
R12622 VDPWR.n1544 VDPWR.n1533 0.0410405
R12623 VDPWR.n1585 VDPWR.n1288 0.0410405
R12624 VDPWR.n1581 VDPWR.n1579 0.0410405
R12625 VDPWR.n1817 VDPWR.n1231 0.0410405
R12626 VDPWR.n1232 VDPWR.n1226 0.0410405
R12627 VDPWR.n1781 VDPWR.n1249 0.0410405
R12628 VDPWR.n1252 VDPWR.n1243 0.0410405
R12629 VDPWR.n1751 VDPWR.n1270 0.0410405
R12630 VDPWR.n1747 VDPWR.n1265 0.0410405
R12631 VDPWR.n1711 VDPWR.n1678 0.0410405
R12632 VDPWR.n1679 VDPWR.n1281 0.0410405
R12633 VDPWR.n1889 VDPWR.n1888 0.0410405
R12634 VDPWR.n1901 VDPWR.n1900 0.0410405
R12635 VDPWR.n1855 VDPWR.n1216 0.0410405
R12636 VDPWR.n1862 VDPWR.n1215 0.0410405
R12637 VDPWR.n1170 VDPWR.n1160 0.0410405
R12638 VDPWR.n1171 VDPWR.n1164 0.0410405
R12639 VDPWR.n1137 VDPWR.n1136 0.0410405
R12640 VDPWR.n1139 VDPWR.n1138 0.0410405
R12641 VDPWR.n2069 VDPWR.n1120 0.0410405
R12642 VDPWR.n2065 VDPWR.n2063 0.0410405
R12643 VDPWR.n1669 VDPWR.n1599 0.0410405
R12644 VDPWR.n1662 VDPWR.n1660 0.0410405
R12645 VDPWR.n1952 VDPWR.n1930 0.0410405
R12646 VDPWR.n1943 VDPWR.n1932 0.0410405
R12647 VDPWR.n1978 VDPWR.n1977 0.0410405
R12648 VDPWR.n1910 VDPWR.n1909 0.0410405
R12649 VDPWR.n2328 VDPWR.n1016 0.0410405
R12650 VDPWR.n2321 VDPWR.n1023 0.0410405
R12651 VDPWR.n2246 VDPWR.n1095 0.0410405
R12652 VDPWR.n2238 VDPWR.n2237 0.0410405
R12653 VDPWR.n2156 VDPWR.n2076 0.0410405
R12654 VDPWR.n2162 VDPWR.n1114 0.0410405
R12655 VDPWR.n2110 VDPWR.n2088 0.0410405
R12656 VDPWR.n2123 VDPWR.n2086 0.0410405
R12657 VDPWR.n2261 VDPWR.n2260 0.0410405
R12658 VDPWR.n1082 VDPWR.n1081 0.0410405
R12659 VDPWR.n2294 VDPWR.n2293 0.0410405
R12660 VDPWR.n1048 VDPWR.n1047 0.0410405
R12661 VDPWR.n2878 VDPWR.n958 0.0410405
R12662 VDPWR.n2895 VDPWR.n956 0.0410405
R12663 VDPWR.n2841 VDPWR.n978 0.0410405
R12664 VDPWR.n2847 VDPWR.n971 0.0410405
R12665 VDPWR.n2802 VDPWR.n992 0.0410405
R12666 VDPWR.n2798 VDPWR.n986 0.0410405
R12667 VDPWR.n2752 VDPWR.n2722 0.0410405
R12668 VDPWR.n2723 VDPWR.n1007 0.0410405
R12669 VDPWR.n2966 VDPWR.n2965 0.0410405
R12670 VDPWR.n2978 VDPWR.n2977 0.0410405
R12671 VDPWR.n2929 VDPWR.n946 0.0410405
R12672 VDPWR.n2925 VDPWR.n941 0.0410405
R12673 VDPWR.n3036 VDPWR.n3035 0.0410405
R12674 VDPWR.n906 VDPWR.n905 0.0410405
R12675 VDPWR.n3064 VDPWR.n876 0.0410405
R12676 VDPWR.n3057 VDPWR.n883 0.0410405
R12677 VDPWR.n2465 VDPWR.n783 0.0410405
R12678 VDPWR.n3101 VDPWR.n3100 0.0410405
R12679 VDPWR.n2573 VDPWR.n2571 0.0410405
R12680 VDPWR.n2574 VDPWR.n2542 0.0410405
R12681 VDPWR.n2983 VDPWR.n922 0.0410405
R12682 VDPWR.n2985 VDPWR.n2984 0.0410405
R12683 VDPWR.n2426 VDPWR.n2341 0.0410405
R12684 VDPWR.n2535 VDPWR.n2534 0.0410405
R12685 VDPWR.n2390 VDPWR.n2364 0.0410405
R12686 VDPWR.n2394 VDPWR.n2362 0.0410405
R12687 VDPWR.n846 VDPWR.n773 0.0410405
R12688 VDPWR.n839 VDPWR.n774 0.0410405
R12689 VDPWR.n803 VDPWR.n802 0.0410405
R12690 VDPWR.n869 VDPWR.n868 0.0410405
R12691 VDPWR.n1589 VDPWR.n1588 0.04045
R12692 VDPWR.n1492 VDPWR.n1228 0.04045
R12693 VDPWR.n1456 VDPWR.n1245 0.04045
R12694 VDPWR.n1594 VDPWR.n1283 0.04045
R12695 VDPWR.n1531 VDPWR.n1193 0.04045
R12696 VDPWR.n1423 VDPWR.n1267 0.04045
R12697 VDPWR.n255 VDPWR.n254 0.0403788
R12698 VDPWR VDPWR.n376 0.0403708
R12699 VDPWR.n1426 VDPWR.n1329 0.0395625
R12700 VDPWR.n1459 VDPWR.n1313 0.0395625
R12701 VDPWR.n1484 VDPWR.n1483 0.0395625
R12702 VDPWR.n1578 VDPWR.n1577 0.0395625
R12703 VDPWR.n1551 VDPWR.n1535 0.0395625
R12704 VDPWR.n1757 VDPWR.n1264 0.0395625
R12705 VDPWR.n1788 VDPWR.n1787 0.0395625
R12706 VDPWR.n1812 VDPWR.n1811 0.0395625
R12707 VDPWR.n1864 VDPWR.n1863 0.0395625
R12708 VDPWR.n1892 VDPWR.n1891 0.0395625
R12709 VDPWR.n2061 VDPWR.n1124 0.0395625
R12710 VDPWR.n2031 VDPWR.n2030 0.0395625
R12711 VDPWR.n1175 VDPWR.n1174 0.0395625
R12712 VDPWR.n1914 VDPWR.n1913 0.0395625
R12713 VDPWR.n1950 VDPWR.n1934 0.0395625
R12714 VDPWR.n2164 VDPWR.n1111 0.0395625
R12715 VDPWR.n2240 VDPWR.n2234 0.0395625
R12716 VDPWR.n2323 VDPWR.n2322 0.0395625
R12717 VDPWR.n1055 VDPWR.n1054 0.0395625
R12718 VDPWR.n1083 VDPWR.n1077 0.0395625
R12719 VDPWR.n2808 VDPWR.n985 0.0395625
R12720 VDPWR.n2855 VDPWR.n968 0.0395625
R12721 VDPWR.n2892 VDPWR.n960 0.0395625
R12722 VDPWR.n2936 VDPWR.n940 0.0395625
R12723 VDPWR.n2969 VDPWR.n2968 0.0395625
R12724 VDPWR.n2689 VDPWR.n2593 0.0395625
R12725 VDPWR.n2659 VDPWR.n2658 0.0395625
R12726 VDPWR.n3059 VDPWR.n3058 0.0395625
R12727 VDPWR.n909 VDPWR.n907 0.0395625
R12728 VDPWR.n2995 VDPWR.n2993 0.0395625
R12729 VDPWR.n2532 VDPWR.n2346 0.0395625
R12730 VDPWR.n2489 VDPWR.n2449 0.0395625
R12731 VDPWR.n3099 VDPWR.n787 0.0395625
R12732 VDPWR.n867 VDPWR.n866 0.0395625
R12733 VDPWR.n844 VDPWR.n829 0.0395625
R12734 VDPWR.n580 VDPWR 0.0382604
R12735 VDPWR.n300 VDPWR 0.0382604
R12736 VDPWR.n42 VDPWR 0.0382604
R12737 VDPWR.n2492 VDPWR.n2491 0.0382581
R12738 VDPWR.n755 VDPWR 0.0376452
R12739 VDPWR VDPWR.n595 0.0369583
R12740 VDPWR VDPWR.n315 0.0369583
R12741 VDPWR VDPWR.n57 0.0369583
R12742 VDPWR.n2506 VDPWR 0.036925
R12743 VDPWR.n3108 VDPWR 0.0366988
R12744 VDPWR.n780 VDPWR 0.0366988
R12745 VDPWR.n3111 VDPWR 0.0366988
R12746 VDPWR VDPWR.n2501 0.0362546
R12747 VDPWR.n2503 VDPWR 0.0356084
R12748 VDPWR.n1380 VDPWR.n1344 0.0343542
R12749 VDPWR.n1451 VDPWR.n1450 0.0343542
R12750 VDPWR.n1548 VDPWR.n1547 0.0343542
R12751 VDPWR.n1706 VDPWR.n1280 0.0343542
R12752 VDPWR.n1779 VDPWR.n1254 0.0343542
R12753 VDPWR.n1854 VDPWR.n1851 0.0343542
R12754 VDPWR.n1898 VDPWR.n1897 0.0343542
R12755 VDPWR.n1664 VDPWR.n1663 0.0343542
R12756 VDPWR.n1147 VDPWR.n1146 0.0343542
R12757 VDPWR.n1947 VDPWR.n1946 0.0343542
R12758 VDPWR.n2120 VDPWR.n2085 0.0343542
R12759 VDPWR.n2244 VDPWR.n1097 0.0343542
R12760 VDPWR.n2296 VDPWR.n2295 0.0343542
R12761 VDPWR.n1087 VDPWR.n1086 0.0343542
R12762 VDPWR.n2839 VDPWR.n970 0.0343542
R12763 VDPWR.n2928 VDPWR.n947 0.0343542
R12764 VDPWR.n2975 VDPWR.n2974 0.0343542
R12765 VDPWR.n2577 VDPWR.n2543 0.0343542
R12766 VDPWR.n2653 VDPWR.n2651 0.0343542
R12767 VDPWR.n3038 VDPWR.n3037 0.0343542
R12768 VDPWR.n3002 VDPWR.n3001 0.0343542
R12769 VDPWR.n2396 VDPWR.n2395 0.0343542
R12770 VDPWR.n2496 VDPWR.n2448 0.0343542
R12771 VDPWR.n809 VDPWR.n801 0.0343542
R12772 VDPWR.n842 VDPWR.n841 0.0343542
R12773 VDPWR VDPWR.n1500 0.0330521
R12774 VDPWR VDPWR.n2745 0.0330521
R12775 VDPWR VDPWR.n2819 0.0330521
R12776 VDPWR.n2901 VDPWR 0.0330521
R12777 VDPWR VDPWR.n2382 0.0330521
R12778 VDPWR.n3094 VDPWR 0.0330521
R12779 VDPWR.n620 VDPWR 0.03175
R12780 VDPWR.n639 VDPWR 0.03175
R12781 VDPWR.n340 VDPWR 0.03175
R12782 VDPWR.n359 VDPWR 0.03175
R12783 VDPWR.n142 VDPWR.n138 0.03175
R12784 VDPWR.n173 VDPWR.n172 0.03175
R12785 VDPWR.n172 VDPWR.n151 0.03175
R12786 VDPWR.n168 VDPWR.n167 0.03175
R12787 VDPWR.n167 VDPWR.n166 0.03175
R12788 VDPWR.n163 VDPWR.n162 0.03175
R12789 VDPWR.n162 VDPWR.n161 0.03175
R12790 VDPWR.n158 VDPWR.n157 0.03175
R12791 VDPWR.n157 VDPWR.n156 0.03175
R12792 VDPWR.n201 VDPWR.n128 0.03175
R12793 VDPWR.n197 VDPWR.n196 0.03175
R12794 VDPWR.n196 VDPWR.n195 0.03175
R12795 VDPWR.n192 VDPWR.n191 0.03175
R12796 VDPWR.n191 VDPWR.n190 0.03175
R12797 VDPWR.n187 VDPWR.n186 0.03175
R12798 VDPWR.n186 VDPWR.n185 0.03175
R12799 VDPWR.n182 VDPWR.n181 0.03175
R12800 VDPWR.n181 VDPWR.n180 0.03175
R12801 VDPWR VDPWR.n1432 0.03175
R12802 VDPWR VDPWR.n1496 0.03175
R12803 VDPWR.n1497 VDPWR 0.03175
R12804 VDPWR.n1759 VDPWR 0.03175
R12805 VDPWR VDPWR.n1763 0.03175
R12806 VDPWR.n1824 VDPWR 0.03175
R12807 VDPWR VDPWR.n1883 0.03175
R12808 VDPWR.n2056 VDPWR 0.03175
R12809 VDPWR.n2002 VDPWR 0.03175
R12810 VDPWR.n1965 VDPWR 0.03175
R12811 VDPWR VDPWR.n2169 0.03175
R12812 VDPWR.n2170 VDPWR 0.03175
R12813 VDPWR.n2214 VDPWR 0.03175
R12814 VDPWR.n2318 VDPWR 0.03175
R12815 VDPWR.n2737 VDPWR 0.03175
R12816 VDPWR.n2810 VDPWR 0.03175
R12817 VDPWR VDPWR.n2876 0.03175
R12818 VDPWR VDPWR.n2900 0.03175
R12819 VDPWR VDPWR.n2598 0.03175
R12820 VDPWR VDPWR.n2604 0.03175
R12821 VDPWR.n2409 VDPWR 0.03175
R12822 VDPWR VDPWR.n2427 0.03175
R12823 VDPWR.n2528 VDPWR 0.03175
R12824 VDPWR.n2527 VDPWR 0.03175
R12825 VDPWR VDPWR.n2443 0.03175
R12826 VDPWR.n2477 VDPWR 0.03175
R12827 VDPWR VDPWR.n2464 0.03175
R12828 VDPWR VDPWR.n790 0.03175
R12829 VDPWR.n811 VDPWR 0.03175
R12830 VDPWR.n853 VDPWR 0.03175
R12831 VDPWR.n82 VDPWR 0.03175
R12832 VDPWR.n101 VDPWR 0.03175
R12833 VDPWR.n1555 VDPWR.n1554 0.0292489
R12834 VDPWR.n1545 VDPWR.n1532 0.0292489
R12835 VDPWR.n1196 VDPWR.n1194 0.0292489
R12836 VDPWR.n1903 VDPWR.n1902 0.0292489
R12837 VDPWR.n1954 VDPWR.n1953 0.0292489
R12838 VDPWR.n1944 VDPWR.n1931 0.0292489
R12839 VDPWR.n2259 VDPWR.n1080 0.0292489
R12840 VDPWR.n2258 VDPWR.n2257 0.0292489
R12841 VDPWR.n926 VDPWR.n924 0.0292489
R12842 VDPWR.n2980 VDPWR.n2979 0.0292489
R12843 VDPWR.n3034 VDPWR.n3033 0.0292489
R12844 VDPWR.n3032 VDPWR.n3031 0.0292489
R12845 VDPWR.n2931 VDPWR.n944 0.0292489
R12846 VDPWR.n2933 VDPWR.n942 0.0292489
R12847 VDPWR.n2292 VDPWR.n2291 0.0292489
R12848 VDPWR.n2289 VDPWR.n1045 0.0292489
R12849 VDPWR.n1976 VDPWR.n1975 0.0292489
R12850 VDPWR.n1973 VDPWR.n1190 0.0292489
R12851 VDPWR.n1858 VDPWR.n1857 0.0292489
R12852 VDPWR.n1860 VDPWR.n1859 0.0292489
R12853 VDPWR.n1587 VDPWR.n1286 0.0292489
R12854 VDPWR.n1580 VDPWR.n1285 0.0292489
R12855 VDPWR.n3066 VDPWR.n874 0.0292489
R12856 VDPWR.n882 VDPWR.n873 0.0292489
R12857 VDPWR.n2879 VDPWR.n957 0.0292489
R12858 VDPWR.n2897 VDPWR.n2896 0.0292489
R12859 VDPWR.n2330 VDPWR.n1014 0.0292489
R12860 VDPWR.n1022 VDPWR.n1013 0.0292489
R12861 VDPWR.n2007 VDPWR.n1161 0.0292489
R12862 VDPWR.n2005 VDPWR.n1163 0.0292489
R12863 VDPWR.n1819 VDPWR.n1229 0.0292489
R12864 VDPWR.n1821 VDPWR.n1227 0.0292489
R12865 VDPWR.n1491 VDPWR.n1301 0.0292489
R12866 VDPWR.n1493 VDPWR.n1300 0.0292489
R12867 VDPWR.n2664 VDPWR.n2663 0.0292489
R12868 VDPWR.n2662 VDPWR.n2661 0.0292489
R12869 VDPWR.n2843 VDPWR.n975 0.0292489
R12870 VDPWR.n2845 VDPWR.n972 0.0292489
R12871 VDPWR.n2248 VDPWR.n1093 0.0292489
R12872 VDPWR.n2236 VDPWR.n1092 0.0292489
R12873 VDPWR.n2036 VDPWR.n2035 0.0292489
R12874 VDPWR.n2034 VDPWR.n2033 0.0292489
R12875 VDPWR.n1783 VDPWR.n1247 0.0292489
R12876 VDPWR.n1785 VDPWR.n1244 0.0292489
R12877 VDPWR.n1455 VDPWR.n1318 0.0292489
R12878 VDPWR.n1457 VDPWR.n1317 0.0292489
R12879 VDPWR.n2754 VDPWR.n2720 0.0292489
R12880 VDPWR.n2756 VDPWR.n1008 0.0292489
R12881 VDPWR.n2111 VDPWR.n2087 0.0292489
R12882 VDPWR.n2125 VDPWR.n2124 0.0292489
R12883 VDPWR.n1671 VDPWR.n1597 0.0292489
R12884 VDPWR.n1659 VDPWR.n1595 0.0292489
R12885 VDPWR.n1713 VDPWR.n1676 0.0292489
R12886 VDPWR.n1715 VDPWR.n1282 0.0292489
R12887 VDPWR.n1372 VDPWR.n1346 0.0292489
R12888 VDPWR.n1385 VDPWR.n1384 0.0292489
R12889 VDPWR.n2541 VDPWR.n2337 0.0292489
R12890 VDPWR.n2572 VDPWR.n2337 0.0292489
R12891 VDPWR.n3007 VDPWR.n3006 0.0292489
R12892 VDPWR.n3005 VDPWR.n3004 0.0292489
R12893 VDPWR.n2694 VDPWR.n2693 0.0292489
R12894 VDPWR.n2692 VDPWR.n2691 0.0292489
R12895 VDPWR.n2804 VDPWR.n990 0.0292489
R12896 VDPWR.n2806 VDPWR.n987 0.0292489
R12897 VDPWR.n2158 VDPWR.n2074 0.0292489
R12898 VDPWR.n2160 VDPWR.n1115 0.0292489
R12899 VDPWR.n2071 VDPWR.n1118 0.0292489
R12900 VDPWR.n2064 VDPWR.n1117 0.0292489
R12901 VDPWR.n1753 VDPWR.n1268 0.0292489
R12902 VDPWR.n1755 VDPWR.n1266 0.0292489
R12903 VDPWR.n1422 VDPWR.n1332 0.0292489
R12904 VDPWR.n1424 VDPWR.n1331 0.0292489
R12905 VDPWR.n586 VDPWR.n585 0.0291458
R12906 VDPWR.n306 VDPWR.n305 0.0291458
R12907 VDPWR.n1419 VDPWR.n1335 0.0291458
R12908 VDPWR.n1479 VDPWR.n1302 0.0291458
R12909 VDPWR.n1750 VDPWR.n1271 0.0291458
R12910 VDPWR.n1808 VDPWR.n1230 0.0291458
R12911 VDPWR.n2068 VDPWR.n1121 0.0291458
R12912 VDPWR.n2010 VDPWR.n2009 0.0291458
R12913 VDPWR.n2155 VDPWR.n2152 0.0291458
R12914 VDPWR.n2213 VDPWR.n1015 0.0291458
R12915 VDPWR.n2801 VDPWR.n993 0.0291458
R12916 VDPWR.n2882 VDPWR.n2881 0.0291458
R12917 VDPWR.n2630 VDPWR.n875 0.0291458
R12918 VDPWR.n48 VDPWR.n47 0.0291458
R12919 VDPWR.n753 VDPWR.n752 0.0281786
R12920 VDPWR.n1979 VDPWR 0.0265417
R12921 VDPWR.n2747 VDPWR 0.0265417
R12922 VDPWR VDPWR.n809 0.0265417
R12923 VDPWR.n202 VDPWR.n127 0.0249565
R12924 VDPWR.n727 VDPWR.n725 0.0247347
R12925 VDPWR.n1375 VDPWR.n1374 0.0239375
R12926 VDPWR.n1703 VDPWR.n1677 0.0239375
R12927 VDPWR.n1607 VDPWR.n1598 0.0239375
R12928 VDPWR.n2114 VDPWR.n2113 0.0239375
R12929 VDPWR VDPWR.n2831 0.0239375
R12930 VDPWR.n2569 VDPWR.n2568 0.0239375
R12931 VDPWR.n3011 VDPWR 0.0239375
R12932 VDPWR.n2367 VDPWR.n2365 0.0239375
R12933 VDPWR.n655 VDPWR 0.0236148
R12934 VDPWR VDPWR.n3178 0.0236148
R12935 VDPWR.n728 VDPWR.n723 0.0234592
R12936 VDPWR.n1010 VDPWR 0.022975
R12937 VDPWR.n1284 VDPWR 0.022975
R12938 VDPWR.n1906 VDPWR 0.022975
R12939 VDPWR.n2254 VDPWR 0.022975
R12940 VDPWR.n3070 VDPWR 0.022975
R12941 VDPWR.n3110 VDPWR 0.022975
R12942 VDPWR VDPWR.n567 0.0226354
R12943 VDPWR VDPWR.n592 0.0226354
R12944 VDPWR.n612 VDPWR 0.0226354
R12945 VDPWR.n607 VDPWR 0.0226354
R12946 VDPWR.n599 VDPWR 0.0226354
R12947 VDPWR VDPWR.n569 0.0226354
R12948 VDPWR.n579 VDPWR 0.0226354
R12949 VDPWR.n629 VDPWR 0.0226354
R12950 VDPWR VDPWR.n637 0.0226354
R12951 VDPWR.n638 VDPWR 0.0226354
R12952 VDPWR VDPWR.n538 0.0226354
R12953 VDPWR VDPWR.n542 0.0226354
R12954 VDPWR VDPWR.n547 0.0226354
R12955 VDPWR.n552 VDPWR 0.0226354
R12956 VDPWR VDPWR.n287 0.0226354
R12957 VDPWR VDPWR.n312 0.0226354
R12958 VDPWR.n332 VDPWR 0.0226354
R12959 VDPWR.n327 VDPWR 0.0226354
R12960 VDPWR.n319 VDPWR 0.0226354
R12961 VDPWR VDPWR.n289 0.0226354
R12962 VDPWR.n299 VDPWR 0.0226354
R12963 VDPWR.n349 VDPWR 0.0226354
R12964 VDPWR VDPWR.n357 0.0226354
R12965 VDPWR.n358 VDPWR 0.0226354
R12966 VDPWR VDPWR.n258 0.0226354
R12967 VDPWR VDPWR.n262 0.0226354
R12968 VDPWR VDPWR.n267 0.0226354
R12969 VDPWR.n272 VDPWR 0.0226354
R12970 VDPWR VDPWR.n1394 0.0226354
R12971 VDPWR.n1401 VDPWR 0.0226354
R12972 VDPWR.n1427 VDPWR 0.0226354
R12973 VDPWR.n1515 VDPWR 0.0226354
R12974 VDPWR.n1517 VDPWR 0.0226354
R12975 VDPWR.n1577 VDPWR 0.0226354
R12976 VDPWR.n1522 VDPWR 0.0226354
R12977 VDPWR VDPWR.n1529 0.0226354
R12978 VDPWR.n1548 VDPWR 0.0226354
R12979 VDPWR VDPWR.n1724 0.0226354
R12980 VDPWR.n1731 VDPWR 0.0226354
R12981 VDPWR VDPWR.n1758 0.0226354
R12982 VDPWR VDPWR.n1793 0.0226354
R12983 VDPWR VDPWR.n1831 0.0226354
R12984 VDPWR VDPWR.n1837 0.0226354
R12985 VDPWR.n1864 VDPWR 0.0226354
R12986 VDPWR VDPWR.n1212 0.0226354
R12987 VDPWR.n1880 VDPWR 0.0226354
R12988 VDPWR.n1885 VDPWR 0.0226354
R12989 VDPWR.n1897 VDPWR 0.0226354
R12990 VDPWR.n1651 VDPWR 0.0226354
R12991 VDPWR.n1642 VDPWR 0.0226354
R12992 VDPWR.n2057 VDPWR 0.0226354
R12993 VDPWR.n2042 VDPWR 0.0226354
R12994 VDPWR.n2025 VDPWR 0.0226354
R12995 VDPWR.n2018 VDPWR 0.0226354
R12996 VDPWR.n1993 VDPWR 0.0226354
R12997 VDPWR.n1992 VDPWR 0.0226354
R12998 VDPWR.n1963 VDPWR 0.0226354
R12999 VDPWR VDPWR.n1929 0.0226354
R13000 VDPWR.n1947 VDPWR 0.0226354
R13001 VDPWR.n2105 VDPWR 0.0226354
R13002 VDPWR.n2133 VDPWR 0.0226354
R13003 VDPWR.n2139 VDPWR 0.0226354
R13004 VDPWR VDPWR.n2168 0.0226354
R13005 VDPWR VDPWR.n2174 0.0226354
R13006 VDPWR.n2175 VDPWR 0.0226354
R13007 VDPWR VDPWR.n2182 0.0226354
R13008 VDPWR.n2227 VDPWR 0.0226354
R13009 VDPWR.n2314 VDPWR 0.0226354
R13010 VDPWR.n2313 VDPWR 0.0226354
R13011 VDPWR.n1055 VDPWR 0.0226354
R13012 VDPWR.n2287 VDPWR 0.0226354
R13013 VDPWR.n2263 VDPWR 0.0226354
R13014 VDPWR.n1086 VDPWR 0.0226354
R13015 VDPWR.n2748 VDPWR 0.0226354
R13016 VDPWR.n2759 VDPWR 0.0226354
R13017 VDPWR VDPWR.n2764 0.0226354
R13018 VDPWR.n2779 VDPWR 0.0226354
R13019 VDPWR VDPWR.n2809 0.0226354
R13020 VDPWR.n2820 VDPWR 0.0226354
R13021 VDPWR.n2827 VDPWR 0.0226354
R13022 VDPWR.n2857 VDPWR 0.0226354
R13023 VDPWR.n2936 VDPWR 0.0226354
R13024 VDPWR VDPWR.n2935 0.0226354
R13025 VDPWR.n2943 VDPWR 0.0226354
R13026 VDPWR.n2962 VDPWR 0.0226354
R13027 VDPWR.n2974 VDPWR 0.0226354
R13028 VDPWR VDPWR.n2588 0.0226354
R13029 VDPWR.n2688 VDPWR 0.0226354
R13030 VDPWR.n2655 VDPWR 0.0226354
R13031 VDPWR.n2658 VDPWR 0.0226354
R13032 VDPWR.n2644 VDPWR 0.0226354
R13033 VDPWR.n3054 VDPWR 0.0226354
R13034 VDPWR.n3020 VDPWR 0.0226354
R13035 VDPWR VDPWR.n918 0.0226354
R13036 VDPWR VDPWR.n921 0.0226354
R13037 VDPWR.n3001 VDPWR 0.0226354
R13038 VDPWR.n2379 VDPWR 0.0226354
R13039 VDPWR VDPWR.n2383 0.0226354
R13040 VDPWR.n2403 VDPWR 0.0226354
R13041 VDPWR.n2415 VDPWR 0.0226354
R13042 VDPWR VDPWR.n2425 0.0226354
R13043 VDPWR.n2429 VDPWR 0.0226354
R13044 VDPWR.n2523 VDPWR 0.0226354
R13045 VDPWR.n2516 VDPWR 0.0226354
R13046 VDPWR VDPWR.n2439 0.0226354
R13047 VDPWR VDPWR.n2455 0.0226354
R13048 VDPWR.n2468 VDPWR 0.0226354
R13049 VDPWR.n3093 VDPWR 0.0226354
R13050 VDPWR.n3081 VDPWR 0.0226354
R13051 VDPWR.n3078 VDPWR 0.0226354
R13052 VDPWR.n862 VDPWR 0.0226354
R13053 VDPWR VDPWR.n816 0.0226354
R13054 VDPWR.n855 VDPWR 0.0226354
R13055 VDPWR.n850 VDPWR 0.0226354
R13056 VDPWR VDPWR.n827 0.0226354
R13057 VDPWR.n842 VDPWR 0.0226354
R13058 VDPWR VDPWR.n29 0.0226354
R13059 VDPWR VDPWR.n54 0.0226354
R13060 VDPWR.n74 VDPWR 0.0226354
R13061 VDPWR.n69 VDPWR 0.0226354
R13062 VDPWR.n61 VDPWR 0.0226354
R13063 VDPWR VDPWR.n31 0.0226354
R13064 VDPWR.n41 VDPWR 0.0226354
R13065 VDPWR.n91 VDPWR 0.0226354
R13066 VDPWR VDPWR.n99 0.0226354
R13067 VDPWR.n100 VDPWR 0.0226354
R13068 VDPWR VDPWR.n0 0.0226354
R13069 VDPWR VDPWR.n4 0.0226354
R13070 VDPWR VDPWR.n9 0.0226354
R13071 VDPWR.n14 VDPWR 0.0226354
R13072 VDPWR.n248 VDPWR.n121 0.0226154
R13073 VDPWR.n243 VDPWR.n242 0.0226154
R13074 VDPWR.n238 VDPWR.n237 0.0226154
R13075 VDPWR.n233 VDPWR.n232 0.0226154
R13076 VDPWR.n228 VDPWR.n227 0.0226154
R13077 VDPWR.n223 VDPWR.n222 0.0226154
R13078 VDPWR.n218 VDPWR.n217 0.0226154
R13079 VDPWR.n213 VDPWR.n212 0.0226154
R13080 VDPWR.n208 VDPWR.n207 0.0226154
R13081 VDPWR.n3105 VDPWR.n3104 0.0218125
R13082 VDPWR VDPWR.n1183 0.0213333
R13083 VDPWR.n2950 VDPWR 0.0213333
R13084 VDPWR.n2659 VDPWR 0.0213333
R13085 VDPWR.n2631 VDPWR 0.0213333
R13086 VDPWR.n867 VDPWR 0.0213333
R13087 VDPWR VDPWR.n1495 0.0200312
R13088 VDPWR VDPWR.n1823 0.0200312
R13089 VDPWR.n2003 VDPWR 0.0200312
R13090 VDPWR.n2319 VDPWR 0.0200312
R13091 VDPWR VDPWR.n2899 0.0200312
R13092 VDPWR.n3055 VDPWR 0.0200312
R13093 VDPWR VDPWR.n788 0.0200312
R13094 VDPWR VDPWR.n248 0.0185288
R13095 VDPWR.n243 VDPWR 0.0185288
R13096 VDPWR.n238 VDPWR 0.0185288
R13097 VDPWR.n233 VDPWR 0.0185288
R13098 VDPWR.n223 VDPWR 0.0185288
R13099 VDPWR.n218 VDPWR 0.0185288
R13100 VDPWR.n213 VDPWR 0.0185288
R13101 VDPWR.n208 VDPWR 0.0185288
R13102 VDPWR.n2932 VDPWR.n943 0.018125
R13103 VDPWR.n2332 VDPWR.n872 0.018125
R13104 VDPWR.n2844 VDPWR.n973 0.018125
R13105 VDPWR.n2755 VDPWR.n2336 0.018125
R13106 VDPWR.n2981 VDPWR.n923 0.018125
R13107 VDPWR.n2805 VDPWR.n988 0.018125
R13108 VDPWR.n3072 VDPWR.n870 0.01695
R13109 VDPWR.n3068 VDPWR.n3067 0.01695
R13110 VDPWR.n2499 VDPWR.n974 0.01695
R13111 VDPWR.n2719 VDPWR.n2540 0.01695
R13112 VDPWR.n2982 VDPWR.n775 0.01695
R13113 VDPWR.n2538 VDPWR.n989 0.01695
R13114 VDPWR VDPWR.n137 0.016125
R13115 VDPWR.n149 VDPWR 0.016125
R13116 VDPWR.n150 VDPWR 0.016125
R13117 VDPWR.n174 VDPWR 0.016125
R13118 VDPWR VDPWR.n173 0.016125
R13119 VDPWR.n168 VDPWR 0.016125
R13120 VDPWR.n163 VDPWR 0.016125
R13121 VDPWR.n158 VDPWR 0.016125
R13122 VDPWR VDPWR.n127 0.016125
R13123 VDPWR.n197 VDPWR 0.016125
R13124 VDPWR.n192 VDPWR 0.016125
R13125 VDPWR.n187 VDPWR 0.016125
R13126 VDPWR.n182 VDPWR 0.016125
R13127 VDPWR.n177 VDPWR 0.016125
R13128 VDPWR VDPWR.n1522 0.016125
R13129 VDPWR.n1890 VDPWR 0.016125
R13130 VDPWR.n1933 VDPWR 0.016125
R13131 VDPWR VDPWR.n2262 0.016125
R13132 VDPWR.n2967 VDPWR 0.016125
R13133 VDPWR.n2992 VDPWR 0.016125
R13134 VDPWR.n845 VDPWR 0.016125
R13135 VDPWR.n203 VDPWR 0.0137212
R13136 VDPWR.n1370 VDPWR.n1348 0.0135208
R13137 VDPWR.n1447 VDPWR.n1319 0.0135208
R13138 VDPWR.n1710 VDPWR.n1709 0.0135208
R13139 VDPWR.n1250 VDPWR.n1248 0.0135208
R13140 VDPWR.n1668 VDPWR.n1667 0.0135208
R13141 VDPWR.n2038 VDPWR.n1135 0.0135208
R13142 VDPWR.n2119 VDPWR.n2089 0.0135208
R13143 VDPWR.n1096 VDPWR.n1094 0.0135208
R13144 VDPWR.n2751 VDPWR.n2750 0.0135208
R13145 VDPWR.n2838 VDPWR.n976 0.0135208
R13146 VDPWR.n2570 VDPWR.n2548 0.0135208
R13147 VDPWR.n2666 VDPWR.n2614 0.0135208
R13148 VDPWR.n2389 VDPWR.n2388 0.0135208
R13149 VDPWR.n2510 VDPWR.n2443 0.0135208
R13150 VDPWR.n3117 VDPWR 0.0122968
R13151 VDPWR.n1584 VDPWR 0.0122188
R13152 VDPWR VDPWR.n1979 0.0122188
R13153 VDPWR VDPWR.n2747 0.0122188
R13154 VDPWR VDPWR.n249 0.0115577
R13155 VDPWR VDPWR.n121 0.0115577
R13156 VDPWR.n122 VDPWR 0.0115577
R13157 VDPWR.n242 VDPWR 0.0115577
R13158 VDPWR VDPWR.n241 0.0115577
R13159 VDPWR.n237 VDPWR 0.0115577
R13160 VDPWR VDPWR.n236 0.0115577
R13161 VDPWR.n232 VDPWR 0.0115577
R13162 VDPWR VDPWR.n231 0.0115577
R13163 VDPWR.n227 VDPWR 0.0115577
R13164 VDPWR VDPWR.n226 0.0115577
R13165 VDPWR.n222 VDPWR 0.0115577
R13166 VDPWR VDPWR.n221 0.0115577
R13167 VDPWR.n217 VDPWR 0.0115577
R13168 VDPWR VDPWR.n216 0.0115577
R13169 VDPWR.n212 VDPWR 0.0115577
R13170 VDPWR VDPWR.n211 0.0115577
R13171 VDPWR.n207 VDPWR 0.0115577
R13172 VDPWR.n252 VDPWR 0.0115577
R13173 VDPWR VDPWR.n1287 0.0109167
R13174 VDPWR VDPWR.n2360 0.0109167
R13175 VDPWR.n2447 VDPWR 0.0109167
R13176 VDPWR VDPWR.n3107 0.00972152
R13177 VDPWR.n3106 VDPWR 0.00972152
R13178 VDPWR VDPWR.n778 0.00972152
R13179 VDPWR VDPWR.n2502 0.00972152
R13180 VDPWR.n375 VDPWR.n254 0.00887356
R13181 VDPWR.n137 VDPWR 0.00865217
R13182 VDPWR VDPWR.n149 0.00865217
R13183 VDPWR VDPWR.n150 0.00865217
R13184 VDPWR.n174 VDPWR 0.00865217
R13185 VDPWR.n177 VDPWR 0.00865217
R13186 VDPWR.n1418 VDPWR.n1415 0.0083125
R13187 VDPWR.n1488 VDPWR.n1487 0.0083125
R13188 VDPWR.n1557 VDPWR.n1529 0.0083125
R13189 VDPWR.n1749 VDPWR.n1746 0.0083125
R13190 VDPWR.n1816 VDPWR.n1815 0.0083125
R13191 VDPWR.n1886 VDPWR.n1885 0.0083125
R13192 VDPWR.n2067 VDPWR.n1122 0.0083125
R13193 VDPWR.n1169 VDPWR.n1159 0.0083125
R13194 VDPWR.n1956 VDPWR.n1929 0.0083125
R13195 VDPWR.n2154 VDPWR.n1113 0.0083125
R13196 VDPWR.n2327 VDPWR.n2326 0.0083125
R13197 VDPWR.n2263 VDPWR.n1076 0.0083125
R13198 VDPWR.n2800 VDPWR.n2797 0.0083125
R13199 VDPWR.n2877 VDPWR.n959 0.0083125
R13200 VDPWR.n2963 VDPWR.n2962 0.0083125
R13201 VDPWR.n2602 VDPWR.n2600 0.0083125
R13202 VDPWR.n3063 VDPWR.n3062 0.0083125
R13203 VDPWR.n3009 VDPWR.n921 0.0083125
R13204 VDPWR.n2429 VDPWR.n2428 0.0083125
R13205 VDPWR.n2468 VDPWR.n2466 0.0083125
R13206 VDPWR.n848 VDPWR.n827 0.0083125
R13207 VDPWR.n202 VDPWR.n201 0.00729348
R13208 VDPWR.n2598 VDPWR 0.00701042
R13209 VDPWR.n2427 VDPWR 0.00701042
R13210 VDPWR.n2464 VDPWR 0.00701042
R13211 VDPWR VDPWR.n151 0.00627446
R13212 VDPWR.n166 VDPWR 0.00627446
R13213 VDPWR.n161 VDPWR 0.00627446
R13214 VDPWR.n156 VDPWR 0.00627446
R13215 VDPWR VDPWR.n128 0.00627446
R13216 VDPWR.n195 VDPWR 0.00627446
R13217 VDPWR.n190 VDPWR 0.00627446
R13218 VDPWR.n185 VDPWR 0.00627446
R13219 VDPWR.n180 VDPWR 0.00627446
R13220 VDPWR VDPWR.n252 0.00626923
R13221 VDPWR.n138 VDPWR 0.00593478
R13222 VDPWR.n228 VDPWR.n203 0.00530769
R13223 VDPWR.n3073 VDPWR.n777 0.0052
R13224 VDPWR.n782 VDPWR.n781 0.0052
R13225 VDPWR.n2500 VDPWR.n2339 0.0052
R13226 VDPWR.n3113 VDPWR.n3112 0.0052
R13227 VDPWR.n2537 VDPWR.n2340 0.0052
R13228 VDPWR.n249 VDPWR 0.00458654
R13229 VDPWR VDPWR.n122 0.00458654
R13230 VDPWR.n241 VDPWR 0.00458654
R13231 VDPWR.n236 VDPWR 0.00458654
R13232 VDPWR.n231 VDPWR 0.00458654
R13233 VDPWR.n226 VDPWR 0.00458654
R13234 VDPWR.n221 VDPWR 0.00458654
R13235 VDPWR.n216 VDPWR 0.00458654
R13236 VDPWR.n211 VDPWR 0.00458654
R13237 VDPWR.n629 VDPWR.n628 0.00310417
R13238 VDPWR.n349 VDPWR.n348 0.00310417
R13239 VDPWR.n1388 VDPWR.n1387 0.00310417
R13240 VDPWR.n1460 VDPWR.n1315 0.00310417
R13241 VDPWR.n1495 VDPWR.n1298 0.00310417
R13242 VDPWR.n1583 VDPWR.n1289 0.00310417
R13243 VDPWR.n1550 VDPWR.n1536 0.00310417
R13244 VDPWR.n1718 VDPWR.n1717 0.00310417
R13245 VDPWR.n1251 VDPWR.n1242 0.00310417
R13246 VDPWR.n1823 VDPWR.n1225 0.00310417
R13247 VDPWR.n1853 VDPWR.n1214 0.00310417
R13248 VDPWR.n1899 VDPWR.n1198 0.00310417
R13249 VDPWR.n1657 VDPWR.n1656 0.00310417
R13250 VDPWR.n1144 VDPWR.n1140 0.00310417
R13251 VDPWR.n2003 VDPWR.n1165 0.00310417
R13252 VDPWR.n1912 VDPWR.n1911 0.00310417
R13253 VDPWR.n1949 VDPWR.n1935 0.00310417
R13254 VDPWR.n2128 VDPWR.n2127 0.00310417
R13255 VDPWR.n2241 VDPWR.n2197 0.00310417
R13256 VDPWR.n2319 VDPWR.n1020 0.00310417
R13257 VDPWR.n1053 VDPWR.n1042 0.00310417
R13258 VDPWR.n1085 VDPWR.n1084 0.00310417
R13259 VDPWR.n2759 VDPWR.n2758 0.00310417
R13260 VDPWR.n2849 VDPWR.n2848 0.00310417
R13261 VDPWR.n2899 VDPWR.n955 0.00310417
R13262 VDPWR.n2927 VDPWR.n2924 0.00310417
R13263 VDPWR.n2976 VDPWR.n928 0.00310417
R13264 VDPWR.n2716 VDPWR.n2715 0.00310417
R13265 VDPWR.n2655 VDPWR.n2654 0.00310417
R13266 VDPWR.n3055 VDPWR.n880 0.00310417
R13267 VDPWR.n910 VDPWR.n902 0.00310417
R13268 VDPWR.n2996 VDPWR.n2986 0.00310417
R13269 VDPWR.n2361 VDPWR.n2358 0.00310417
R13270 VDPWR.n2495 VDPWR.n2493 0.00310417
R13271 VDPWR.n3098 VDPWR.n788 0.00310417
R13272 VDPWR.n811 VDPWR.n810 0.00310417
R13273 VDPWR.n840 VDPWR.n835 0.00310417
R13274 VDPWR.n91 VDPWR.n90 0.00310417
R13275 VDPWR.n627 VDPWR.n626 0.00180208
R13276 VDPWR.n595 VDPWR 0.00180208
R13277 VDPWR.n561 VDPWR.n547 0.00180208
R13278 VDPWR.n347 VDPWR.n346 0.00180208
R13279 VDPWR.n315 VDPWR 0.00180208
R13280 VDPWR.n281 VDPWR.n267 0.00180208
R13281 VDPWR.n89 VDPWR.n88 0.00180208
R13282 VDPWR.n57 VDPWR 0.00180208
R13283 VDPWR.n23 VDPWR.n9 0.00180208
R13284 VDPWR.n728 VDPWR.n727 0.00177551
R13285 VDPWR.n257 VDPWR.n255 0.00105731
R13286 muxtest_0.x2.x2.GP1.n2 muxtest_0.x2.x2.GP1.t4 450.938
R13287 muxtest_0.x2.x2.GP1.n2 muxtest_0.x2.x2.GP1.t5 445.666
R13288 muxtest_0.x2.x2.GP1.n4 muxtest_0.x2.x2.GP1.n3 195.832
R13289 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n0 96.8352
R13290 muxtest_0.x2.x2.GP1.n3 muxtest_0.x2.x2.GP1.t3 26.5955
R13291 muxtest_0.x2.x2.GP1.n3 muxtest_0.x2.x2.GP1.t2 26.5955
R13292 muxtest_0.x2.x2.GP1.n0 muxtest_0.x2.x2.GP1.t1 24.9236
R13293 muxtest_0.x2.x2.GP1.n0 muxtest_0.x2.x2.GP1.t0 24.9236
R13294 muxtest_0.x2.x2.GP1.n5 muxtest_0.x2.x2.GP1.n4 13.1346
R13295 muxtest_0.x2.x2.GP1.n4 muxtest_0.x2.x2.GP1 12.2007
R13296 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n1 11.2645
R13297 muxtest_0.x2.x2.GP1.n1 muxtest_0.x2.x2.GP1 6.1445
R13298 muxtest_0.x2.x2.GP1.n1 muxtest_0.x2.x2.GP1 4.65505
R13299 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n2 3.07707
R13300 muxtest_0.x2.x2.GP1.n5 muxtest_0.x2.x2.GP1 2.0485
R13301 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n5 1.55202
R13302 ua[3].n10 ua[3].t4 26.3998
R13303 ua[3].n6 ua[3].t6 23.6581
R13304 ua[3].n1 ua[3].t3 23.6581
R13305 ua[3].n10 ua[3].t5 23.5483
R13306 ua[3].n8 ua[3].t8 23.3739
R13307 ua[3].n3 ua[3].t2 23.3739
R13308 ua[3].n11 ua[3].t10 12.9758
R13309 ua[3].n11 ua[3].t11 10.8618
R13310 ua[3].n6 ua[3].t1 10.7528
R13311 ua[3].n1 ua[3].t9 10.7528
R13312 ua[3].n5 ua[3].t0 10.6417
R13313 ua[3].n0 ua[3].t7 10.6417
R13314 ua[3].n15 ua[3] 4.48702
R13315 ua[3].n12 ua[3].n10 3.06895
R13316 ua[3].n12 ua[3].n11 2.14822
R13317 ua[3].n14 ua[3] 1.938
R13318 ua[3].n7 ua[3].n6 1.30064
R13319 ua[3].n2 ua[3].n1 1.30064
R13320 ua[3].n13 ua[3].n12 1.12636
R13321 ua[3] ua[3].n9 0.983856
R13322 ua[3] ua[3].n4 0.966624
R13323 ua[3].n8 ua[3].n7 0.726502
R13324 ua[3].n3 ua[3].n2 0.726502
R13325 ua[3].n17 ua[3].n16 0.683625
R13326 ua[3].n7 ua[3].n5 0.512491
R13327 ua[3].n2 ua[3].n0 0.512491
R13328 ua[3].n15 ua[3] 0.398
R13329 ua[3] ua[3].n15 0.398
R13330 ua[3].n16 ua[3] 0.37425
R13331 ua[3].n9 ua[3].n5 0.359663
R13332 ua[3].n4 ua[3].n0 0.359663
R13333 ua[3].n16 ua[3] 0.2705
R13334 ua[3].n9 ua[3].n8 0.216071
R13335 ua[3].n4 ua[3].n3 0.216071
R13336 ua[3].n14 ua[3].n13 0.148615
R13337 ua[3] ua[3].n14 0.146333
R13338 ua[3].n17 ua[3] 0.124875
R13339 ua[3].n13 ua[3] 0.0655
R13340 ua[3] ua[3].n17 0.063
R13341 ua[2].n6 ua[2].t2 23.6581
R13342 ua[2].n15 ua[2].t6 23.6581
R13343 ua[2].n22 ua[2].t4 23.6581
R13344 ua[2].n1 ua[2].t9 23.6581
R13345 ua[2].n5 ua[2].t3 23.3739
R13346 ua[2].n14 ua[2].t7 23.3739
R13347 ua[2].n21 ua[2].t5 23.3739
R13348 ua[2].n0 ua[2].t8 23.3739
R13349 ua[2].n28 ua[2] 21.5313
R13350 ua[2].n6 ua[2].t15 10.7528
R13351 ua[2].n15 ua[2].t1 10.7528
R13352 ua[2].n22 ua[2].t10 10.7528
R13353 ua[2].n1 ua[2].t12 10.7528
R13354 ua[2].n8 ua[2].t14 10.6417
R13355 ua[2].n17 ua[2].t0 10.6417
R13356 ua[2].n24 ua[2].t11 10.6417
R13357 ua[2].n3 ua[2].t13 10.6417
R13358 ua[2].n7 ua[2].n6 1.30064
R13359 ua[2].n16 ua[2].n15 1.30064
R13360 ua[2].n23 ua[2].n22 1.30064
R13361 ua[2].n2 ua[2].n1 1.30064
R13362 ua[2] ua[2].n4 0.983856
R13363 ua[2].n10 ua[2].n9 0.956356
R13364 ua[2].n26 ua[2].n25 0.946356
R13365 ua[2].n19 ua[2].n18 0.927606
R13366 ua[2].n7 ua[2].n5 0.726502
R13367 ua[2].n16 ua[2].n14 0.726502
R13368 ua[2].n23 ua[2].n21 0.726502
R13369 ua[2].n2 ua[2].n0 0.726502
R13370 ua[2].n11 ua[2] 0.681056
R13371 ua[2].n20 ua[2].n13 0.54925
R13372 ua[2].n27 ua[2].n20 0.54425
R13373 ua[2].n28 ua[2].n27 0.53675
R13374 ua[2].n8 ua[2].n7 0.512491
R13375 ua[2].n17 ua[2].n16 0.512491
R13376 ua[2].n24 ua[2].n23 0.512491
R13377 ua[2].n3 ua[2].n2 0.512491
R13378 ua[2].n9 ua[2].n8 0.359663
R13379 ua[2].n18 ua[2].n17 0.359663
R13380 ua[2].n25 ua[2].n24 0.359663
R13381 ua[2].n4 ua[2].n3 0.359663
R13382 ua[2].n9 ua[2].n5 0.216071
R13383 ua[2].n18 ua[2].n14 0.216071
R13384 ua[2].n25 ua[2].n21 0.216071
R13385 ua[2].n4 ua[2].n0 0.216071
R13386 ua[2].n20 ua[2] 0.18675
R13387 ua[2].n13 ua[2] 0.18425
R13388 ua[2].n27 ua[2] 0.16425
R13389 ua[2] ua[2].n28 0.163
R13390 ua[2].n12 ua[2] 0.135115
R13391 ua[2].n19 ua[2] 0.05675
R13392 ua[2] ua[2].n19 0.0561931
R13393 ua[2].n12 ua[2].n11 0.0530774
R13394 ua[2].n26 ua[2] 0.038
R13395 ua[2] ua[2].n26 0.0376287
R13396 ua[2].n10 ua[2] 0.028
R13397 ua[2] ua[2].n10 0.0266905
R13398 ua[2].n11 ua[2] 0.01175
R13399 ua[2].n13 ua[2].n12 0.006125
R13400 ringtest_0.x4.clknet_0_clk.n33 ringtest_0.x4.clknet_0_clk.n31 333.392
R13401 ringtest_0.x4.clknet_0_clk.n38 ringtest_0.x4.clknet_0_clk.n26 301.392
R13402 ringtest_0.x4.clknet_0_clk.n37 ringtest_0.x4.clknet_0_clk.n27 301.392
R13403 ringtest_0.x4.clknet_0_clk.n36 ringtest_0.x4.clknet_0_clk.n28 301.392
R13404 ringtest_0.x4.clknet_0_clk.n35 ringtest_0.x4.clknet_0_clk.n29 301.392
R13405 ringtest_0.x4.clknet_0_clk.n34 ringtest_0.x4.clknet_0_clk.n30 301.392
R13406 ringtest_0.x4.clknet_0_clk.n33 ringtest_0.x4.clknet_0_clk.n32 301.392
R13407 ringtest_0.x4.clknet_0_clk.n39 ringtest_0.x4.clknet_0_clk.n25 297.863
R13408 ringtest_0.x4.clknet_0_clk.n2 ringtest_0.x4.clknet_0_clk.n0 248.638
R13409 ringtest_0.x4.clknet_0_clk.n2 ringtest_0.x4.clknet_0_clk.n1 203.463
R13410 ringtest_0.x4.clknet_0_clk.n4 ringtest_0.x4.clknet_0_clk.n3 203.463
R13411 ringtest_0.x4.clknet_0_clk.n8 ringtest_0.x4.clknet_0_clk.n7 203.463
R13412 ringtest_0.x4.clknet_0_clk.n24 ringtest_0.x4.clknet_0_clk.n23 203.463
R13413 ringtest_0.x4.clknet_0_clk.n6 ringtest_0.x4.clknet_0_clk.n5 202.456
R13414 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n41 199.607
R13415 ringtest_0.x4.clknet_0_clk.n21 ringtest_0.x4.clknet_0_clk.n9 188.201
R13416 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.t46 184.768
R13417 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.t43 184.768
R13418 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.t42 184.768
R13419 ringtest_0.x4.clknet_0_clk.n15 ringtest_0.x4.clknet_0_clk.t45 184.768
R13420 ringtest_0.x4.clknet_0_clk.n10 ringtest_0.x4.clknet_0_clk.t41 184.768
R13421 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.t37 184.768
R13422 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.t40 184.768
R13423 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.t39 184.768
R13424 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n18 173.609
R13425 ringtest_0.x4.clknet_0_clk.n14 ringtest_0.x4.clknet_0_clk.n13 171.375
R13426 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.t38 146.208
R13427 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.t35 146.208
R13428 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.t34 146.208
R13429 ringtest_0.x4.clknet_0_clk.n15 ringtest_0.x4.clknet_0_clk.t36 146.208
R13430 ringtest_0.x4.clknet_0_clk.n10 ringtest_0.x4.clknet_0_clk.t33 146.208
R13431 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.t44 146.208
R13432 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.t32 146.208
R13433 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.t47 146.208
R13434 ringtest_0.x4.clknet_0_clk.n4 ringtest_0.x4.clknet_0_clk.n2 45.177
R13435 ringtest_0.x4.clknet_0_clk.n22 ringtest_0.x4.clknet_0_clk.n8 45.177
R13436 ringtest_0.x4.clknet_0_clk.n24 ringtest_0.x4.clknet_0_clk.n22 45.177
R13437 ringtest_0.x4.clknet_0_clk.n6 ringtest_0.x4.clknet_0_clk.n4 44.0476
R13438 ringtest_0.x4.clknet_0_clk.n8 ringtest_0.x4.clknet_0_clk.n6 44.0476
R13439 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.n17 40.6397
R13440 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.n16 40.6397
R13441 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.n15 40.6397
R13442 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.n10 40.6397
R13443 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.n11 40.6397
R13444 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.n12 40.6397
R13445 ringtest_0.x4.clknet_0_clk.n0 ringtest_0.x4.clknet_0_clk.t2 40.0005
R13446 ringtest_0.x4.clknet_0_clk.n0 ringtest_0.x4.clknet_0_clk.t15 40.0005
R13447 ringtest_0.x4.clknet_0_clk.n1 ringtest_0.x4.clknet_0_clk.t4 40.0005
R13448 ringtest_0.x4.clknet_0_clk.n1 ringtest_0.x4.clknet_0_clk.t6 40.0005
R13449 ringtest_0.x4.clknet_0_clk.n3 ringtest_0.x4.clknet_0_clk.t8 40.0005
R13450 ringtest_0.x4.clknet_0_clk.n3 ringtest_0.x4.clknet_0_clk.t10 40.0005
R13451 ringtest_0.x4.clknet_0_clk.n5 ringtest_0.x4.clknet_0_clk.t5 40.0005
R13452 ringtest_0.x4.clknet_0_clk.n5 ringtest_0.x4.clknet_0_clk.t7 40.0005
R13453 ringtest_0.x4.clknet_0_clk.n7 ringtest_0.x4.clknet_0_clk.t9 40.0005
R13454 ringtest_0.x4.clknet_0_clk.n7 ringtest_0.x4.clknet_0_clk.t11 40.0005
R13455 ringtest_0.x4.clknet_0_clk.n9 ringtest_0.x4.clknet_0_clk.t0 40.0005
R13456 ringtest_0.x4.clknet_0_clk.n9 ringtest_0.x4.clknet_0_clk.t13 40.0005
R13457 ringtest_0.x4.clknet_0_clk.n23 ringtest_0.x4.clknet_0_clk.t14 40.0005
R13458 ringtest_0.x4.clknet_0_clk.n23 ringtest_0.x4.clknet_0_clk.t12 40.0005
R13459 ringtest_0.x4.clknet_0_clk.n41 ringtest_0.x4.clknet_0_clk.t1 40.0005
R13460 ringtest_0.x4.clknet_0_clk.n41 ringtest_0.x4.clknet_0_clk.t3 40.0005
R13461 ringtest_0.x4.clknet_0_clk.n38 ringtest_0.x4.clknet_0_clk.n37 32.0005
R13462 ringtest_0.x4.clknet_0_clk.n37 ringtest_0.x4.clknet_0_clk.n36 32.0005
R13463 ringtest_0.x4.clknet_0_clk.n35 ringtest_0.x4.clknet_0_clk.n34 32.0005
R13464 ringtest_0.x4.clknet_0_clk.n34 ringtest_0.x4.clknet_0_clk.n33 32.0005
R13465 ringtest_0.x4.clknet_0_clk.n36 ringtest_0.x4.clknet_0_clk.n35 31.2005
R13466 ringtest_0.x4.clknet_0_clk.n31 ringtest_0.x4.clknet_0_clk.t27 27.5805
R13467 ringtest_0.x4.clknet_0_clk.n31 ringtest_0.x4.clknet_0_clk.t24 27.5805
R13468 ringtest_0.x4.clknet_0_clk.n26 ringtest_0.x4.clknet_0_clk.t23 27.5805
R13469 ringtest_0.x4.clknet_0_clk.n26 ringtest_0.x4.clknet_0_clk.t21 27.5805
R13470 ringtest_0.x4.clknet_0_clk.n25 ringtest_0.x4.clknet_0_clk.t26 27.5805
R13471 ringtest_0.x4.clknet_0_clk.n25 ringtest_0.x4.clknet_0_clk.t28 27.5805
R13472 ringtest_0.x4.clknet_0_clk.n27 ringtest_0.x4.clknet_0_clk.t25 27.5805
R13473 ringtest_0.x4.clknet_0_clk.n27 ringtest_0.x4.clknet_0_clk.t22 27.5805
R13474 ringtest_0.x4.clknet_0_clk.n28 ringtest_0.x4.clknet_0_clk.t18 27.5805
R13475 ringtest_0.x4.clknet_0_clk.n28 ringtest_0.x4.clknet_0_clk.t20 27.5805
R13476 ringtest_0.x4.clknet_0_clk.n29 ringtest_0.x4.clknet_0_clk.t30 27.5805
R13477 ringtest_0.x4.clknet_0_clk.n29 ringtest_0.x4.clknet_0_clk.t16 27.5805
R13478 ringtest_0.x4.clknet_0_clk.n30 ringtest_0.x4.clknet_0_clk.t17 27.5805
R13479 ringtest_0.x4.clknet_0_clk.n30 ringtest_0.x4.clknet_0_clk.t19 27.5805
R13480 ringtest_0.x4.clknet_0_clk.n32 ringtest_0.x4.clknet_0_clk.t29 27.5805
R13481 ringtest_0.x4.clknet_0_clk.n32 ringtest_0.x4.clknet_0_clk.t31 27.5805
R13482 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n14 25.9814
R13483 ringtest_0.x4.clknet_0_clk.n22 ringtest_0.x4.clknet_0_clk.n21 15.262
R13484 ringtest_0.x4.clknet_0_clk.n20 ringtest_0.x4.clknet_0_clk.n19 14.7771
R13485 ringtest_0.x4.clknet_0_clk.n40 ringtest_0.x4.clknet_0_clk.n24 13.177
R13486 ringtest_0.x4.clknet_0_clk.n39 ringtest_0.x4.clknet_0_clk.n38 10.4484
R13487 ringtest_0.x4.clknet_0_clk.n19 ringtest_0.x4.clknet_0_clk 10.3624
R13488 ringtest_0.x4.clknet_0_clk.n21 ringtest_0.x4.clknet_0_clk.n20 9.3005
R13489 ringtest_0.x4.clknet_0_clk.n19 ringtest_0.x4.clknet_0_clk 3.45447
R13490 ringtest_0.x4.clknet_0_clk.n40 ringtest_0.x4.clknet_0_clk 3.13183
R13491 ringtest_0.x4.clknet_0_clk.n14 ringtest_0.x4.clknet_0_clk 2.23542
R13492 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n39 1.75844
R13493 ringtest_0.x4.clknet_0_clk.n20 ringtest_0.x4.clknet_0_clk 1.5927
R13494 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n40 0.604792
R13495 ringtest_0.x4.net6.n3 ringtest_0.x4.net6.t13 323.342
R13496 ringtest_0.x4.net6.n0 ringtest_0.x4.net6.t4 323.342
R13497 ringtest_0.x4.net6.n1 ringtest_0.x4.net6.t2 260.322
R13498 ringtest_0.x4.net6.n8 ringtest_0.x4.net6.t5 241.536
R13499 ringtest_0.x4.net6.n17 ringtest_0.x4.net6.t1 222.679
R13500 ringtest_0.x4.net6.n12 ringtest_0.x4.net6.t14 212.081
R13501 ringtest_0.x4.net6.n13 ringtest_0.x4.net6.t7 212.081
R13502 ringtest_0.x4.net6.n3 ringtest_0.x4.net6.t6 194.809
R13503 ringtest_0.x4.net6.n0 ringtest_0.x4.net6.t8 194.809
R13504 ringtest_0.x4.net6.n5 ringtest_0.x4.net6.t10 183.505
R13505 ringtest_0.x4.net6.n1 ringtest_0.x4.net6.t12 175.169
R13506 ringtest_0.x4.net6.n8 ringtest_0.x4.net6.t11 169.237
R13507 ringtest_0.x4.net6 ringtest_0.x4.net6.n3 158.133
R13508 ringtest_0.x4.net6 ringtest_0.x4.net6.n0 158.133
R13509 ringtest_0.x4.net6 ringtest_0.x4.net6.n8 157.555
R13510 ringtest_0.x4.net6.n15 ringtest_0.x4.net6.n14 155.52
R13511 ringtest_0.x4.net6.n6 ringtest_0.x4.net6.n5 153.863
R13512 ringtest_0.x4.net6.n2 ringtest_0.x4.net6.n1 152
R13513 ringtest_0.x4.net6.n12 ringtest_0.x4.net6.t9 139.78
R13514 ringtest_0.x4.net6.n13 ringtest_0.x4.net6.t15 139.78
R13515 ringtest_0.x4.net6.n18 ringtest_0.x4.net6.t0 129.078
R13516 ringtest_0.x4.net6.n5 ringtest_0.x4.net6.t3 114.532
R13517 ringtest_0.x4.net6.n18 ringtest_0.x4.net6.n17 96.7191
R13518 ringtest_0.x4.net6.n11 ringtest_0.x4.net6 55.2785
R13519 ringtest_0.x4.net6.n14 ringtest_0.x4.net6.n13 37.246
R13520 ringtest_0.x4.net6.n14 ringtest_0.x4.net6.n12 24.1005
R13521 ringtest_0.x4.net6.n10 ringtest_0.x4.net6.n9 21.4124
R13522 ringtest_0.x4.net6.n16 ringtest_0.x4.net6.n15 21.1949
R13523 ringtest_0.x4.net6.n4 ringtest_0.x4.net6.n2 20.043
R13524 ringtest_0.x4.net6.n7 ringtest_0.x4.net6.n6 15.2615
R13525 ringtest_0.x4.net6.n17 ringtest_0.x4.net6.n16 12.4213
R13526 ringtest_0.x4.net6.n9 ringtest_0.x4.net6 12.3175
R13527 ringtest_0.x4.net6.n16 ringtest_0.x4.net6.n11 8.09819
R13528 ringtest_0.x4.net6.n11 ringtest_0.x4.net6.n10 7.53948
R13529 ringtest_0.x4.net6.n4 ringtest_0.x4.net6 7.39885
R13530 ringtest_0.x4.net6 ringtest_0.x4.net6.n18 5.84085
R13531 ringtest_0.x4.net6.n15 ringtest_0.x4.net6 5.4405
R13532 ringtest_0.x4.net6.n9 ringtest_0.x4.net6 4.10616
R13533 ringtest_0.x4.net6.n7 ringtest_0.x4.net6.n4 2.60421
R13534 ringtest_0.x4.net6.n10 ringtest_0.x4.net6.n7 2.43577
R13535 ringtest_0.x4.net6.n6 ringtest_0.x4.net6 1.97868
R13536 ringtest_0.x4.net6.n2 ringtest_0.x4.net6 1.55726
R13537 ringtest_0.x4.clknet_1_1__leaf_clk.n29 ringtest_0.x4.clknet_1_1__leaf_clk.n27 333.392
R13538 ringtest_0.x4.clknet_1_1__leaf_clk.n29 ringtest_0.x4.clknet_1_1__leaf_clk.n28 301.392
R13539 ringtest_0.x4.clknet_1_1__leaf_clk.n31 ringtest_0.x4.clknet_1_1__leaf_clk.n30 301.392
R13540 ringtest_0.x4.clknet_1_1__leaf_clk.n33 ringtest_0.x4.clknet_1_1__leaf_clk.n32 301.392
R13541 ringtest_0.x4.clknet_1_1__leaf_clk.n35 ringtest_0.x4.clknet_1_1__leaf_clk.n34 301.392
R13542 ringtest_0.x4.clknet_1_1__leaf_clk.n37 ringtest_0.x4.clknet_1_1__leaf_clk.n36 301.392
R13543 ringtest_0.x4.clknet_1_1__leaf_clk.n39 ringtest_0.x4.clknet_1_1__leaf_clk.n38 301.392
R13544 ringtest_0.x4.clknet_1_1__leaf_clk.n40 ringtest_0.x4.clknet_1_1__leaf_clk.n26 297.863
R13545 ringtest_0.x4.clknet_1_1__leaf_clk.n18 ringtest_0.x4.clknet_1_1__leaf_clk.t36 294.557
R13546 ringtest_0.x4.clknet_1_1__leaf_clk.n15 ringtest_0.x4.clknet_1_1__leaf_clk.t33 294.557
R13547 ringtest_0.x4.clknet_1_1__leaf_clk.n13 ringtest_0.x4.clknet_1_1__leaf_clk.t34 294.557
R13548 ringtest_0.x4.clknet_1_1__leaf_clk.n11 ringtest_0.x4.clknet_1_1__leaf_clk.t41 294.557
R13549 ringtest_0.x4.clknet_1_1__leaf_clk.n10 ringtest_0.x4.clknet_1_1__leaf_clk.t32 294.557
R13550 ringtest_0.x4.clknet_1_1__leaf_clk.n2 ringtest_0.x4.clknet_1_1__leaf_clk.n0 248.638
R13551 ringtest_0.x4.clknet_1_1__leaf_clk.n18 ringtest_0.x4.clknet_1_1__leaf_clk.t39 211.01
R13552 ringtest_0.x4.clknet_1_1__leaf_clk.n15 ringtest_0.x4.clknet_1_1__leaf_clk.t40 211.01
R13553 ringtest_0.x4.clknet_1_1__leaf_clk.n13 ringtest_0.x4.clknet_1_1__leaf_clk.t38 211.01
R13554 ringtest_0.x4.clknet_1_1__leaf_clk.n11 ringtest_0.x4.clknet_1_1__leaf_clk.t35 211.01
R13555 ringtest_0.x4.clknet_1_1__leaf_clk.n10 ringtest_0.x4.clknet_1_1__leaf_clk.t37 211.01
R13556 ringtest_0.x4.clknet_1_1__leaf_clk.n2 ringtest_0.x4.clknet_1_1__leaf_clk.n1 203.463
R13557 ringtest_0.x4.clknet_1_1__leaf_clk.n4 ringtest_0.x4.clknet_1_1__leaf_clk.n3 203.463
R13558 ringtest_0.x4.clknet_1_1__leaf_clk.n8 ringtest_0.x4.clknet_1_1__leaf_clk.n7 203.463
R13559 ringtest_0.x4.clknet_1_1__leaf_clk.n25 ringtest_0.x4.clknet_1_1__leaf_clk.n24 203.463
R13560 ringtest_0.x4.clknet_1_1__leaf_clk.n6 ringtest_0.x4.clknet_1_1__leaf_clk.n5 202.456
R13561 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n42 199.607
R13562 ringtest_0.x4.clknet_1_1__leaf_clk.n22 ringtest_0.x4.clknet_1_1__leaf_clk.n9 188.201
R13563 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n13 156.207
R13564 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n10 156.207
R13565 ringtest_0.x4.clknet_1_1__leaf_clk.n19 ringtest_0.x4.clknet_1_1__leaf_clk.n18 153.097
R13566 ringtest_0.x4.clknet_1_1__leaf_clk.n16 ringtest_0.x4.clknet_1_1__leaf_clk.n15 152.296
R13567 ringtest_0.x4.clknet_1_1__leaf_clk.n12 ringtest_0.x4.clknet_1_1__leaf_clk.n11 152.296
R13568 ringtest_0.x4.clknet_1_1__leaf_clk.n4 ringtest_0.x4.clknet_1_1__leaf_clk.n2 45.177
R13569 ringtest_0.x4.clknet_1_1__leaf_clk.n23 ringtest_0.x4.clknet_1_1__leaf_clk.n8 45.177
R13570 ringtest_0.x4.clknet_1_1__leaf_clk.n25 ringtest_0.x4.clknet_1_1__leaf_clk.n23 45.177
R13571 ringtest_0.x4.clknet_1_1__leaf_clk.n6 ringtest_0.x4.clknet_1_1__leaf_clk.n4 44.0476
R13572 ringtest_0.x4.clknet_1_1__leaf_clk.n8 ringtest_0.x4.clknet_1_1__leaf_clk.n6 44.0476
R13573 ringtest_0.x4.clknet_1_1__leaf_clk.n0 ringtest_0.x4.clknet_1_1__leaf_clk.t13 40.0005
R13574 ringtest_0.x4.clknet_1_1__leaf_clk.n0 ringtest_0.x4.clknet_1_1__leaf_clk.t14 40.0005
R13575 ringtest_0.x4.clknet_1_1__leaf_clk.n1 ringtest_0.x4.clknet_1_1__leaf_clk.t15 40.0005
R13576 ringtest_0.x4.clknet_1_1__leaf_clk.n1 ringtest_0.x4.clknet_1_1__leaf_clk.t12 40.0005
R13577 ringtest_0.x4.clknet_1_1__leaf_clk.n3 ringtest_0.x4.clknet_1_1__leaf_clk.t11 40.0005
R13578 ringtest_0.x4.clknet_1_1__leaf_clk.n3 ringtest_0.x4.clknet_1_1__leaf_clk.t10 40.0005
R13579 ringtest_0.x4.clknet_1_1__leaf_clk.n5 ringtest_0.x4.clknet_1_1__leaf_clk.t6 40.0005
R13580 ringtest_0.x4.clknet_1_1__leaf_clk.n5 ringtest_0.x4.clknet_1_1__leaf_clk.t8 40.0005
R13581 ringtest_0.x4.clknet_1_1__leaf_clk.n7 ringtest_0.x4.clknet_1_1__leaf_clk.t2 40.0005
R13582 ringtest_0.x4.clknet_1_1__leaf_clk.n7 ringtest_0.x4.clknet_1_1__leaf_clk.t4 40.0005
R13583 ringtest_0.x4.clknet_1_1__leaf_clk.n9 ringtest_0.x4.clknet_1_1__leaf_clk.t5 40.0005
R13584 ringtest_0.x4.clknet_1_1__leaf_clk.n9 ringtest_0.x4.clknet_1_1__leaf_clk.t7 40.0005
R13585 ringtest_0.x4.clknet_1_1__leaf_clk.n24 ringtest_0.x4.clknet_1_1__leaf_clk.t1 40.0005
R13586 ringtest_0.x4.clknet_1_1__leaf_clk.n24 ringtest_0.x4.clknet_1_1__leaf_clk.t9 40.0005
R13587 ringtest_0.x4.clknet_1_1__leaf_clk.n42 ringtest_0.x4.clknet_1_1__leaf_clk.t3 40.0005
R13588 ringtest_0.x4.clknet_1_1__leaf_clk.n42 ringtest_0.x4.clknet_1_1__leaf_clk.t0 40.0005
R13589 ringtest_0.x4.clknet_1_1__leaf_clk.n21 ringtest_0.x4.clknet_1_1__leaf_clk 34.5053
R13590 ringtest_0.x4.clknet_1_1__leaf_clk.n14 ringtest_0.x4.clknet_1_1__leaf_clk 33.8485
R13591 ringtest_0.x4.clknet_1_1__leaf_clk.n31 ringtest_0.x4.clknet_1_1__leaf_clk.n29 32.0005
R13592 ringtest_0.x4.clknet_1_1__leaf_clk.n33 ringtest_0.x4.clknet_1_1__leaf_clk.n31 32.0005
R13593 ringtest_0.x4.clknet_1_1__leaf_clk.n37 ringtest_0.x4.clknet_1_1__leaf_clk.n35 32.0005
R13594 ringtest_0.x4.clknet_1_1__leaf_clk.n39 ringtest_0.x4.clknet_1_1__leaf_clk.n37 32.0005
R13595 ringtest_0.x4.clknet_1_1__leaf_clk.n35 ringtest_0.x4.clknet_1_1__leaf_clk.n33 31.2005
R13596 ringtest_0.x4.clknet_1_1__leaf_clk.n27 ringtest_0.x4.clknet_1_1__leaf_clk.t19 27.5805
R13597 ringtest_0.x4.clknet_1_1__leaf_clk.n27 ringtest_0.x4.clknet_1_1__leaf_clk.t20 27.5805
R13598 ringtest_0.x4.clknet_1_1__leaf_clk.n28 ringtest_0.x4.clknet_1_1__leaf_clk.t21 27.5805
R13599 ringtest_0.x4.clknet_1_1__leaf_clk.n28 ringtest_0.x4.clknet_1_1__leaf_clk.t18 27.5805
R13600 ringtest_0.x4.clknet_1_1__leaf_clk.n30 ringtest_0.x4.clknet_1_1__leaf_clk.t17 27.5805
R13601 ringtest_0.x4.clknet_1_1__leaf_clk.n30 ringtest_0.x4.clknet_1_1__leaf_clk.t16 27.5805
R13602 ringtest_0.x4.clknet_1_1__leaf_clk.n32 ringtest_0.x4.clknet_1_1__leaf_clk.t28 27.5805
R13603 ringtest_0.x4.clknet_1_1__leaf_clk.n32 ringtest_0.x4.clknet_1_1__leaf_clk.t30 27.5805
R13604 ringtest_0.x4.clknet_1_1__leaf_clk.n34 ringtest_0.x4.clknet_1_1__leaf_clk.t24 27.5805
R13605 ringtest_0.x4.clknet_1_1__leaf_clk.n34 ringtest_0.x4.clknet_1_1__leaf_clk.t26 27.5805
R13606 ringtest_0.x4.clknet_1_1__leaf_clk.n36 ringtest_0.x4.clknet_1_1__leaf_clk.t27 27.5805
R13607 ringtest_0.x4.clknet_1_1__leaf_clk.n36 ringtest_0.x4.clknet_1_1__leaf_clk.t29 27.5805
R13608 ringtest_0.x4.clknet_1_1__leaf_clk.n26 ringtest_0.x4.clknet_1_1__leaf_clk.t25 27.5805
R13609 ringtest_0.x4.clknet_1_1__leaf_clk.n26 ringtest_0.x4.clknet_1_1__leaf_clk.t22 27.5805
R13610 ringtest_0.x4.clknet_1_1__leaf_clk.n38 ringtest_0.x4.clknet_1_1__leaf_clk.t23 27.5805
R13611 ringtest_0.x4.clknet_1_1__leaf_clk.n38 ringtest_0.x4.clknet_1_1__leaf_clk.t31 27.5805
R13612 ringtest_0.x4.clknet_1_1__leaf_clk.n23 ringtest_0.x4.clknet_1_1__leaf_clk.n22 15.262
R13613 ringtest_0.x4.clknet_1_1__leaf_clk.n20 ringtest_0.x4.clknet_1_1__leaf_clk.n19 13.8005
R13614 ringtest_0.x4.clknet_1_1__leaf_clk.n41 ringtest_0.x4.clknet_1_1__leaf_clk.n25 13.177
R13615 ringtest_0.x4.clknet_1_1__leaf_clk.n14 ringtest_0.x4.clknet_1_1__leaf_clk.n12 11.6482
R13616 ringtest_0.x4.clknet_1_1__leaf_clk.n22 ringtest_0.x4.clknet_1_1__leaf_clk.n21 10.8268
R13617 ringtest_0.x4.clknet_1_1__leaf_clk.n40 ringtest_0.x4.clknet_1_1__leaf_clk.n39 10.4484
R13618 ringtest_0.x4.clknet_1_1__leaf_clk.n17 ringtest_0.x4.clknet_1_1__leaf_clk.n16 9.3005
R13619 ringtest_0.x4.clknet_1_1__leaf_clk.n20 ringtest_0.x4.clknet_1_1__leaf_clk.n17 8.37704
R13620 ringtest_0.x4.clknet_1_1__leaf_clk.n21 ringtest_0.x4.clknet_1_1__leaf_clk 5.19349
R13621 ringtest_0.x4.clknet_1_1__leaf_clk.n17 ringtest_0.x4.clknet_1_1__leaf_clk.n14 3.99105
R13622 ringtest_0.x4.clknet_1_1__leaf_clk.n41 ringtest_0.x4.clknet_1_1__leaf_clk 3.13183
R13623 ringtest_0.x4.clknet_1_1__leaf_clk.n19 ringtest_0.x4.clknet_1_1__leaf_clk 3.10907
R13624 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n40 1.75844
R13625 ringtest_0.x4.clknet_1_1__leaf_clk.n16 ringtest_0.x4.clknet_1_1__leaf_clk 1.67435
R13626 ringtest_0.x4.clknet_1_1__leaf_clk.n12 ringtest_0.x4.clknet_1_1__leaf_clk 1.67435
R13627 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n20 0.693495
R13628 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n41 0.604792
R13629 ui_in[1].n10 ui_in[1].t8 327.99
R13630 ui_in[1].n3 ui_in[1].t1 293.969
R13631 ui_in[1].n6 ui_in[1].t7 256.07
R13632 ui_in[1].n0 ui_in[1].t0 212.081
R13633 ui_in[1].n1 ui_in[1].t2 212.081
R13634 ui_in[1].n10 ui_in[1].t9 199.457
R13635 ui_in[1].n2 ui_in[1].n1 182.929
R13636 ui_in[1] ui_in[1].n3 154.065
R13637 ui_in[1].n11 ui_in[1].n10 152
R13638 ui_in[1].n7 ui_in[1].n6 152
R13639 ui_in[1].n6 ui_in[1].t3 150.03
R13640 ui_in[1].n0 ui_in[1].t5 139.78
R13641 ui_in[1].n1 ui_in[1].t6 139.78
R13642 ui_in[1].n3 ui_in[1].t4 138.338
R13643 ui_in[1].n1 ui_in[1].n0 61.346
R13644 ui_in[1].n16 ui_in[1] 30.7401
R13645 ui_in[1].n5 ui_in[1] 17.455
R13646 ui_in[1].n14 ui_in[1].n13 14.6836
R13647 ui_in[1].n13 ui_in[1].n12 14.6704
R13648 ui_in[1].n4 ui_in[1] 13.8328
R13649 ui_in[1].n14 ui_in[1].n2 10.6811
R13650 ui_in[1].n7 ui_in[1].n5 10.4374
R13651 ui_in[1].n9 ui_in[1].n8 8.15776
R13652 ui_in[1].n12 ui_in[1] 6.61383
R13653 ui_in[1].n2 ui_in[1] 6.1445
R13654 ui_in[1].n4 ui_in[1] 5.16179
R13655 ui_in[1].n11 ui_in[1] 4.90717
R13656 ui_in[1].n9 ui_in[1].n4 4.65206
R13657 ui_in[1].n15 ui_in[1] 4.54217
R13658 ui_in[1].n8 ui_in[1] 3.93896
R13659 ui_in[1].n12 ui_in[1].n11 2.98717
R13660 ui_in[1].n5 ui_in[1] 2.16665
R13661 ui_in[1].n8 ui_in[1].n7 1.57588
R13662 ui_in[1].n13 ui_in[1].n9 0.79438
R13663 ui_in[1].n15 ui_in[1] 0.606561
R13664 ui_in[1] ui_in[1].n14 0.248606
R13665 ui_in[1] ui_in[1].n15 0.222091
R13666 ui_in[1] ui_in[1].n16 0.122375
R13667 ui_in[1].n16 ui_in[1] 0.121168
R13668 muxtest_0.x1.x3.GP1.n3 muxtest_0.x1.x3.GP1.t4 450.938
R13669 muxtest_0.x1.x3.GP1.n2 muxtest_0.x1.x3.GP1.t6 450.938
R13670 muxtest_0.x1.x3.GP1.n3 muxtest_0.x1.x3.GP1.t5 445.666
R13671 muxtest_0.x1.x3.GP1.n2 muxtest_0.x1.x3.GP1.t7 445.666
R13672 muxtest_0.x1.x3.GP1.n6 muxtest_0.x1.x3.GP1.n5 195.832
R13673 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n0 96.8352
R13674 muxtest_0.x1.x3.GP1.n5 muxtest_0.x1.x3.GP1.t2 26.5955
R13675 muxtest_0.x1.x3.GP1.n5 muxtest_0.x1.x3.GP1.t3 26.5955
R13676 muxtest_0.x1.x3.GP1.n0 muxtest_0.x1.x3.GP1.t1 24.9236
R13677 muxtest_0.x1.x3.GP1.n0 muxtest_0.x1.x3.GP1.t0 24.9236
R13678 muxtest_0.x1.x3.GP1.n4 muxtest_0.x1.x3.GP1 13.257
R13679 muxtest_0.x1.x3.GP1.n7 muxtest_0.x1.x3.GP1.n6 13.1346
R13680 muxtest_0.x1.x3.GP1.n6 muxtest_0.x1.x3.GP1 11.8965
R13681 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n1 11.2645
R13682 muxtest_0.x1.x3.GP1.n1 muxtest_0.x1.x3.GP1 6.1445
R13683 muxtest_0.x1.x3.GP1.n4 muxtest_0.x1.x3.GP1 5.31412
R13684 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n4 5.26828
R13685 muxtest_0.x1.x3.GP1.n1 muxtest_0.x1.x3.GP1 4.65505
R13686 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n2 3.07895
R13687 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n3 2.90754
R13688 muxtest_0.x1.x3.GP1.n7 muxtest_0.x1.x3.GP1 2.0485
R13689 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n7 1.55202
R13690 muxtest_0.x1.x3.GP4.n3 muxtest_0.x1.x3.GP4.t5 450.938
R13691 muxtest_0.x1.x3.GP4.n2 muxtest_0.x1.x3.GP4.t7 450.938
R13692 muxtest_0.x1.x3.GP4.n3 muxtest_0.x1.x3.GP4.t4 445.666
R13693 muxtest_0.x1.x3.GP4.n2 muxtest_0.x1.x3.GP4.t6 445.666
R13694 muxtest_0.x1.x3.GP4.n7 muxtest_0.x1.x3.GP4.n6 208.965
R13695 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n0 96.8352
R13696 muxtest_0.x1.x3.GP4.n6 muxtest_0.x1.x3.GP4.t2 26.5955
R13697 muxtest_0.x1.x3.GP4.n6 muxtest_0.x1.x3.GP4.t3 26.5955
R13698 muxtest_0.x1.x3.GP4.n0 muxtest_0.x1.x3.GP4.t1 24.9236
R13699 muxtest_0.x1.x3.GP4.n0 muxtest_0.x1.x3.GP4.t0 24.9236
R13700 muxtest_0.x1.x3.GP4.n4 muxtest_0.x1.x3.x4.GP 10.9863
R13701 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n5 10.2405
R13702 muxtest_0.x1.x1.gpo3 muxtest_0.x1.x3.GP4.n4 9.34192
R13703 muxtest_0.x1.x3.GP4.n5 muxtest_0.x1.x1.gpo3 7.73829
R13704 muxtest_0.x1.x3.GP4.n1 muxtest_0.x1.x1.x14.Y 6.1445
R13705 muxtest_0.x1.x3.GP4.n4 muxtest_0.x1.x2.x4.GP 5.84951
R13706 muxtest_0.x1.x3.GP4.n1 muxtest_0.x1.x1.x14.Y 4.65505
R13707 muxtest_0.x1.x2.x4.GP muxtest_0.x1.x3.GP4.n3 2.95993
R13708 muxtest_0.x1.x3.x4.GP muxtest_0.x1.x3.GP4.n2 2.95993
R13709 muxtest_0.x1.x3.GP4.n7 muxtest_0.x1.x1.x14.Y 2.0485
R13710 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n7 1.55202
R13711 muxtest_0.x1.x3.GP4.n5 muxtest_0.x1.x3.GP4.n1 1.0245
R13712 ringtest_0.x4._11_ ringtest_0.x4._11_.n0 623.909
R13713 ringtest_0.x4._11_.n24 ringtest_0.x4._11_.t6 334.723
R13714 ringtest_0.x4._11_.n5 ringtest_0.x4._11_.t5 334.723
R13715 ringtest_0.x4._11_.n18 ringtest_0.x4._11_.t19 261.887
R13716 ringtest_0.x4._11_.n14 ringtest_0.x4._11_.t14 256.07
R13717 ringtest_0.x4._11_.n8 ringtest_0.x4._11_.t10 241.536
R13718 ringtest_0.x4._11_.n3 ringtest_0.x4._11_.t13 241.536
R13719 ringtest_0.x4._11_.n1 ringtest_0.x4._11_.t12 231.835
R13720 ringtest_0.x4._11_.n21 ringtest_0.x4._11_.t8 230.363
R13721 ringtest_0.x4._11_ ringtest_0.x4._11_.n30 216.464
R13722 ringtest_0.x4._11_.n24 ringtest_0.x4._11_.t20 206.19
R13723 ringtest_0.x4._11_.n5 ringtest_0.x4._11_.t17 206.19
R13724 ringtest_0.x4._11_.n11 ringtest_0.x4._11_.t11 183.505
R13725 ringtest_0.x4._11_.n8 ringtest_0.x4._11_.t21 169.237
R13726 ringtest_0.x4._11_.n3 ringtest_0.x4._11_.t7 169.237
R13727 ringtest_0.x4._11_.n21 ringtest_0.x4._11_.t16 158.064
R13728 ringtest_0.x4._11_ ringtest_0.x4._11_.n3 157.555
R13729 ringtest_0.x4._11_ ringtest_0.x4._11_.n8 157.166
R13730 ringtest_0.x4._11_.n1 ringtest_0.x4._11_.t9 157.07
R13731 ringtest_0.x4._11_.n18 ringtest_0.x4._11_.t15 155.847
R13732 ringtest_0.x4._11_.n22 ringtest_0.x4._11_.n21 154.048
R13733 ringtest_0.x4._11_.n12 ringtest_0.x4._11_.n11 153.863
R13734 ringtest_0.x4._11_.n19 ringtest_0.x4._11_.n18 153.13
R13735 ringtest_0.x4._11_.n25 ringtest_0.x4._11_.n24 152
R13736 ringtest_0.x4._11_.n15 ringtest_0.x4._11_.n14 152
R13737 ringtest_0.x4._11_.n6 ringtest_0.x4._11_.n5 152
R13738 ringtest_0.x4._11_.n2 ringtest_0.x4._11_.n1 152
R13739 ringtest_0.x4._11_.n14 ringtest_0.x4._11_.t4 150.03
R13740 ringtest_0.x4._11_.n11 ringtest_0.x4._11_.t18 114.532
R13741 ringtest_0.x4._11_.n27 ringtest_0.x4._11_.n26 41.0809
R13742 ringtest_0.x4._11_.n30 ringtest_0.x4._11_.t0 38.5719
R13743 ringtest_0.x4._11_.n30 ringtest_0.x4._11_.t1 38.5719
R13744 ringtest_0.x4._11_.n0 ringtest_0.x4._11_.t3 26.5955
R13745 ringtest_0.x4._11_.n0 ringtest_0.x4._11_.t2 26.5955
R13746 ringtest_0.x4._11_.n17 ringtest_0.x4._11_.n16 25.2401
R13747 ringtest_0.x4._11_.n20 ringtest_0.x4._11_.n19 22.3199
R13748 ringtest_0.x4._11_.n10 ringtest_0.x4._11_.n9 21.8442
R13749 ringtest_0.x4._11_.n10 ringtest_0.x4._11_.n7 20.8523
R13750 ringtest_0.x4._11_.n28 ringtest_0.x4._11_.n27 13.7699
R13751 ringtest_0.x4._11_.n28 ringtest_0.x4._11_.n2 12.7179
R13752 ringtest_0.x4._11_.n4 ringtest_0.x4._11_ 12.3175
R13753 ringtest_0.x4._11_.n9 ringtest_0.x4._11_ 11.4531
R13754 ringtest_0.x4._11_.n7 ringtest_0.x4._11_.n4 11.4418
R13755 ringtest_0.x4._11_.n23 ringtest_0.x4._11_.n20 10.8618
R13756 ringtest_0.x4._11_.n7 ringtest_0.x4._11_.n6 10.3976
R13757 ringtest_0.x4._11_.n25 ringtest_0.x4._11_ 9.6005
R13758 ringtest_0.x4._11_.n29 ringtest_0.x4._11_ 9.6005
R13759 ringtest_0.x4._11_ ringtest_0.x4._11_.n22 9.39918
R13760 ringtest_0.x4._11_.n13 ringtest_0.x4._11_.n12 9.3005
R13761 ringtest_0.x4._11_.n29 ringtest_0.x4._11_.n28 9.3005
R13762 ringtest_0.x4._11_.n23 ringtest_0.x4._11_ 8.80957
R13763 ringtest_0.x4._11_.n6 ringtest_0.x4._11_ 8.22907
R13764 ringtest_0.x4._11_.n15 ringtest_0.x4._11_ 7.6805
R13765 ringtest_0.x4._11_.n16 ringtest_0.x4._11_.n15 4.6085
R13766 ringtest_0.x4._11_.n16 ringtest_0.x4._11_ 4.58918
R13767 ringtest_0.x4._11_.n22 ringtest_0.x4._11_ 4.3525
R13768 ringtest_0.x4._11_.n4 ringtest_0.x4._11_ 4.10616
R13769 ringtest_0.x4._11_.n9 ringtest_0.x4._11_ 3.81804
R13770 ringtest_0.x4._11_.n26 ringtest_0.x4._11_ 3.62717
R13771 ringtest_0.x4._11_.n19 ringtest_0.x4._11_ 3.2005
R13772 ringtest_0.x4._11_ ringtest_0.x4._11_.n29 3.2005
R13773 ringtest_0.x4._11_.n17 ringtest_0.x4._11_.n13 2.49494
R13774 ringtest_0.x4._11_.n2 ringtest_0.x4._11_ 2.3045
R13775 ringtest_0.x4._11_.n12 ringtest_0.x4._11_ 1.97868
R13776 ringtest_0.x4._11_.n13 ringtest_0.x4._11_.n10 1.71582
R13777 ringtest_0.x4._11_.n27 ringtest_0.x4._11_.n23 1.38649
R13778 ringtest_0.x4._11_.n26 ringtest_0.x4._11_.n25 1.2805
R13779 ringtest_0.x4._11_.n20 ringtest_0.x4._11_.n17 1.24753
R13780 ui_in[0].n5 ui_in[0].t7 327.99
R13781 ui_in[0].n9 ui_in[0].t4 293.969
R13782 ui_in[0].n3 ui_in[0].t5 261.887
R13783 ui_in[0].n0 ui_in[0].t8 212.081
R13784 ui_in[0].n1 ui_in[0].t6 212.081
R13785 ui_in[0].n5 ui_in[0].t1 199.457
R13786 ui_in[0].n2 ui_in[0].n1 183.185
R13787 ui_in[0].n3 ui_in[0].t9 155.847
R13788 ui_in[0] ui_in[0].n9 154.065
R13789 ui_in[0].n4 ui_in[0].n3 153.506
R13790 ui_in[0].n6 ui_in[0].n5 152
R13791 ui_in[0].n0 ui_in[0].t3 139.78
R13792 ui_in[0].n1 ui_in[0].t0 139.78
R13793 ui_in[0].n9 ui_in[0].t2 138.338
R13794 ui_in[0].n1 ui_in[0].n0 61.346
R13795 ui_in[0].n13 ui_in[0] 38.2119
R13796 ui_in[0].n10 ui_in[0] 13.4199
R13797 ui_in[0].n11 ui_in[0].n8 11.7395
R13798 ui_in[0].n12 ui_in[0].n11 11.5949
R13799 ui_in[0].n8 ui_in[0].n4 10.4004
R13800 ui_in[0].n12 ui_in[0].n2 9.68118
R13801 ui_in[0].n6 ui_in[0] 9.6005
R13802 ui_in[0].n2 ui_in[0] 5.8885
R13803 ui_in[0].n10 ui_in[0] 5.57469
R13804 ui_in[0].n13 ui_in[0] 4.74482
R13805 ui_in[0].n8 ui_in[0].n7 4.6505
R13806 ui_in[0].n11 ui_in[0].n10 4.6505
R13807 ui_in[0].n7 ui_in[0].n6 2.98717
R13808 ui_in[0].n4 ui_in[0] 2.82403
R13809 ui_in[0].n7 ui_in[0] 1.9205
R13810 ui_in[0] ui_in[0].n12 0.559212
R13811 ui_in[0] ui_in[0].n13 0.02675
R13812 muxtest_0.R3R4.n5 muxtest_0.R3R4.t3 26.3998
R13813 muxtest_0.R3R4.n0 muxtest_0.R3R4.t6 26.3998
R13814 muxtest_0.R3R4.n5 muxtest_0.R3R4.t2 23.5483
R13815 muxtest_0.R3R4.n0 muxtest_0.R3R4.t5 23.5483
R13816 muxtest_0.R3R4.n6 muxtest_0.R3R4.t9 12.9758
R13817 muxtest_0.R3R4.n1 muxtest_0.R3R4.t0 12.9758
R13818 muxtest_0.R3R4.n6 muxtest_0.R3R4.t8 10.8618
R13819 muxtest_0.R3R4.n1 muxtest_0.R3R4.t1 10.8618
R13820 muxtest_0.R3R4.n4 muxtest_0.R3R4.t7 10.5285
R13821 muxtest_0.R3R4.n11 muxtest_0.R3R4.n10 7.08509
R13822 muxtest_0.R3R4.n7 muxtest_0.R3R4.n5 3.06895
R13823 muxtest_0.R3R4.n2 muxtest_0.R3R4.n0 3.06895
R13824 muxtest_0.R3R4.n7 muxtest_0.R3R4.n6 2.14822
R13825 muxtest_0.R3R4.n2 muxtest_0.R3R4.n1 2.14822
R13826 muxtest_0.R3R4.n8 muxtest_0.R3R4.n7 1.12636
R13827 muxtest_0.R3R4.n3 muxtest_0.R3R4.n2 1.12636
R13828 muxtest_0.R3R4.n4 muxtest_0.R3R4.t4 1.06523
R13829 muxtest_0.R3R4.n12 muxtest_0.R3R4 0.893
R13830 muxtest_0.R3R4.n9 muxtest_0.R3R4 0.670143
R13831 muxtest_0.R3R4.n12 muxtest_0.R3R4.n11 0.40675
R13832 muxtest_0.R3R4.n10 muxtest_0.R3R4.n9 0.223714
R13833 muxtest_0.R3R4.n11 muxtest_0.R3R4.n4 0.183423
R13834 muxtest_0.R3R4 muxtest_0.R3R4.n3 0.148615
R13835 muxtest_0.R3R4.n9 muxtest_0.R3R4.n8 0.132418
R13836 muxtest_0.R3R4.n12 muxtest_0.R3R4 0.08425
R13837 muxtest_0.R3R4.n8 muxtest_0.R3R4 0.0655
R13838 muxtest_0.R3R4.n3 muxtest_0.R3R4 0.0655
R13839 muxtest_0.R3R4 muxtest_0.R3R4.n12 0.04425
R13840 muxtest_0.R3R4.n10 muxtest_0.R3R4 0.00907843
R13841 ui_in[4].n26 ui_in[4].t3 327.99
R13842 ui_in[4].n10 ui_in[4].t0 327.99
R13843 ui_in[4].n19 ui_in[4].t1 293.969
R13844 ui_in[4].n3 ui_in[4].t19 293.969
R13845 ui_in[4].n22 ui_in[4].t14 256.07
R13846 ui_in[4].n6 ui_in[4].t12 256.07
R13847 ui_in[4].n16 ui_in[4].t9 212.081
R13848 ui_in[4].n17 ui_in[4].t15 212.081
R13849 ui_in[4].n0 ui_in[4].t6 212.081
R13850 ui_in[4].n1 ui_in[4].t4 212.081
R13851 ui_in[4].n26 ui_in[4].t8 199.457
R13852 ui_in[4].n10 ui_in[4].t5 199.457
R13853 ui_in[4].n18 ui_in[4].n17 182.929
R13854 ui_in[4].n2 ui_in[4].n1 182.929
R13855 ui_in[4] ui_in[4].n19 154.065
R13856 ui_in[4] ui_in[4].n3 154.065
R13857 ui_in[4].n27 ui_in[4].n26 152
R13858 ui_in[4].n23 ui_in[4].n22 152
R13859 ui_in[4].n11 ui_in[4].n10 152
R13860 ui_in[4].n7 ui_in[4].n6 152
R13861 ui_in[4].n22 ui_in[4].t11 150.03
R13862 ui_in[4].n6 ui_in[4].t7 150.03
R13863 ui_in[4].n16 ui_in[4].t18 139.78
R13864 ui_in[4].n17 ui_in[4].t2 139.78
R13865 ui_in[4].n0 ui_in[4].t16 139.78
R13866 ui_in[4].n1 ui_in[4].t10 139.78
R13867 ui_in[4].n19 ui_in[4].t17 138.338
R13868 ui_in[4].n3 ui_in[4].t13 138.338
R13869 ui_in[4].n17 ui_in[4].n16 61.346
R13870 ui_in[4].n1 ui_in[4].n0 61.346
R13871 ui_in[4].n31 ui_in[4] 29.9743
R13872 ui_in[4].n21 ui_in[4] 17.455
R13873 ui_in[4].n5 ui_in[4] 17.455
R13874 ui_in[4].n30 ui_in[4].n29 14.6836
R13875 ui_in[4].n14 ui_in[4].n13 14.6836
R13876 ui_in[4].n29 ui_in[4].n28 14.6704
R13877 ui_in[4].n13 ui_in[4].n12 14.6704
R13878 ui_in[4].n20 ui_in[4] 13.8328
R13879 ui_in[4].n4 ui_in[4] 13.8328
R13880 ui_in[4].n31 ui_in[4] 12.499
R13881 ui_in[4].n30 ui_in[4].n18 10.6811
R13882 ui_in[4].n14 ui_in[4].n2 10.6811
R13883 ui_in[4].n23 ui_in[4].n21 10.4374
R13884 ui_in[4].n7 ui_in[4].n5 10.4374
R13885 ui_in[4].n25 ui_in[4].n24 8.15776
R13886 ui_in[4].n9 ui_in[4].n8 8.15776
R13887 ui_in[4].n28 ui_in[4] 6.61383
R13888 ui_in[4].n12 ui_in[4] 6.61383
R13889 ui_in[4].n18 ui_in[4] 6.1445
R13890 ui_in[4].n2 ui_in[4] 6.1445
R13891 ui_in[4].n20 ui_in[4] 5.16179
R13892 ui_in[4].n4 ui_in[4] 5.16179
R13893 ui_in[4].n27 ui_in[4] 4.90717
R13894 ui_in[4].n11 ui_in[4] 4.90717
R13895 ui_in[4].n25 ui_in[4].n20 4.65206
R13896 ui_in[4].n9 ui_in[4].n4 4.65206
R13897 ui_in[4].n24 ui_in[4] 3.93896
R13898 ui_in[4].n8 ui_in[4] 3.93896
R13899 ui_in[4].n28 ui_in[4].n27 2.98717
R13900 ui_in[4].n12 ui_in[4].n11 2.98717
R13901 ui_in[4].n21 ui_in[4] 2.16665
R13902 ui_in[4].n5 ui_in[4] 2.16665
R13903 ui_in[4].n24 ui_in[4].n23 1.57588
R13904 ui_in[4].n8 ui_in[4].n7 1.57588
R13905 ui_in[4].n29 ui_in[4].n25 0.79438
R13906 ui_in[4].n13 ui_in[4].n9 0.79438
R13907 ui_in[4] ui_in[4].n15 0.287559
R13908 ui_in[4] ui_in[4].n31 0.28675
R13909 ui_in[4] ui_in[4].n30 0.248606
R13910 ui_in[4] ui_in[4].n14 0.248606
R13911 ui_in[4].n15 ui_in[4] 0.11603
R13912 ui_in[4].n15 ui_in[4] 0.0460882
R13913 muxtest_0.R1R2.n0 muxtest_0.R1R2.t1 26.3998
R13914 muxtest_0.R1R2.n0 muxtest_0.R1R2.t0 23.5483
R13915 muxtest_0.R1R2.n1 muxtest_0.R1R2.t5 12.9758
R13916 muxtest_0.R1R2.n4 muxtest_0.R1R2.t3 10.8648
R13917 muxtest_0.R1R2.n1 muxtest_0.R1R2.t4 10.8618
R13918 muxtest_0.R1R2.n4 muxtest_0.R1R2.t2 10.5295
R13919 muxtest_0.R1R2.n2 muxtest_0.R1R2.n0 3.06895
R13920 muxtest_0.R1R2.n2 muxtest_0.R1R2.n1 2.14822
R13921 muxtest_0.R1R2.n3 muxtest_0.R1R2.n2 1.12636
R13922 muxtest_0.R1R2.n5 muxtest_0.R1R2 0.96675
R13923 muxtest_0.R1R2.n5 muxtest_0.R1R2.n4 0.494965
R13924 muxtest_0.R1R2 muxtest_0.R1R2.n3 0.132418
R13925 muxtest_0.R1R2.n5 muxtest_0.R1R2 0.06925
R13926 muxtest_0.R1R2.n3 muxtest_0.R1R2 0.0655
R13927 muxtest_0.R1R2 muxtest_0.R1R2.n5 0.04425
R13928 a_19289_13081.n0 a_19289_13081.t12 1681.78
R13929 a_19289_13081.n2 a_19289_13081.t7 1681.21
R13930 a_19289_13081.n1 a_19289_13081.t13 1681.21
R13931 a_19289_13081.n0 a_19289_13081.t2 1681.21
R13932 a_19289_13081.n13 a_19289_13081.t14 1681.21
R13933 a_19289_13081.n11 a_19289_13081.t10 1681.21
R13934 a_19289_13081.n9 a_19289_13081.t17 1681.21
R13935 a_19289_13081.n7 a_19289_13081.t9 1681.21
R13936 a_19289_13081.n3 a_19289_13081.t4 703.317
R13937 a_19289_13081.n7 a_19289_13081.t6 702.768
R13938 a_19289_13081.n5 a_19289_13081.t11 702.747
R13939 a_19289_13081.n4 a_19289_13081.t5 702.747
R13940 a_19289_13081.n3 a_19289_13081.t15 702.747
R13941 a_19289_13081.n12 a_19289_13081.t3 702.747
R13942 a_19289_13081.n10 a_19289_13081.t8 702.747
R13943 a_19289_13081.n8 a_19289_13081.t16 702.747
R13944 a_19289_13081.n6 a_19289_13081.t0 30.088
R13945 a_19289_13081.t1 a_19289_13081.n15 26.0464
R13946 a_19289_13081.n15 a_19289_13081.n2 20.0759
R13947 a_19289_13081.n6 a_19289_13081.n5 0.875353
R13948 a_19289_13081.n1 a_19289_13081.n0 0.576859
R13949 a_19289_13081.n2 a_19289_13081.n1 0.576859
R13950 a_19289_13081.n4 a_19289_13081.n3 0.570292
R13951 a_19289_13081.n5 a_19289_13081.n4 0.570292
R13952 a_19289_13081.n15 a_19289_13081.n14 0.267403
R13953 a_19289_13081.n14 a_19289_13081.n6 0.10833
R13954 a_19289_13081.n14 a_19289_13081.n13 0.0744583
R13955 a_19289_13081.n8 a_19289_13081.n7 0.0205
R13956 a_19289_13081.n9 a_19289_13081.n8 0.0205
R13957 a_19289_13081.n10 a_19289_13081.n9 0.0205
R13958 a_19289_13081.n11 a_19289_13081.n10 0.0205
R13959 a_19289_13081.n12 a_19289_13081.n11 0.0205
R13960 a_19289_13081.n13 a_19289_13081.n12 0.0205
R13961 ringtest_0.drv_out.n7 ringtest_0.drv_out.t21 184.768
R13962 ringtest_0.drv_out.n6 ringtest_0.drv_out.t20 184.768
R13963 ringtest_0.drv_out.n5 ringtest_0.drv_out.t23 184.768
R13964 ringtest_0.drv_out.n4 ringtest_0.drv_out.t22 184.768
R13965 ringtest_0.drv_out.n8 ringtest_0.drv_out.n7 171.375
R13966 ringtest_0.drv_out.n7 ringtest_0.drv_out.t25 146.208
R13967 ringtest_0.drv_out.n6 ringtest_0.drv_out.t24 146.208
R13968 ringtest_0.drv_out.n5 ringtest_0.drv_out.t27 146.208
R13969 ringtest_0.drv_out.n4 ringtest_0.drv_out.t26 146.208
R13970 ringtest_0.drv_out.n7 ringtest_0.drv_out.n6 40.6397
R13971 ringtest_0.drv_out.n6 ringtest_0.drv_out.n5 40.6397
R13972 ringtest_0.drv_out.n5 ringtest_0.drv_out.n4 40.6397
R13973 ringtest_0.drv_out.n0 ringtest_0.drv_out.t19 26.3998
R13974 ringtest_0.drv_out.n21 ringtest_0.drv_out.n20 26.0838
R13975 ringtest_0.drv_out.n21 ringtest_0.drv_out.n17 26.0838
R13976 ringtest_0.drv_out.n21 ringtest_0.drv_out.n19 26.0838
R13977 ringtest_0.drv_out.n21 ringtest_0.drv_out.n18 26.0838
R13978 ringtest_0.drv_out.n16 ringtest_0.drv_out.n12 24.902
R13979 ringtest_0.drv_out.n16 ringtest_0.drv_out.n14 24.902
R13980 ringtest_0.drv_out.n16 ringtest_0.drv_out.n13 24.902
R13981 ringtest_0.drv_out.n16 ringtest_0.drv_out.n15 24.902
R13982 ringtest_0.drv_out.n0 ringtest_0.drv_out.t0 23.5483
R13983 ringtest_0.drv_out.n1 ringtest_0.drv_out.t1 12.9758
R13984 ringtest_0.drv_out ringtest_0.drv_out.n8 12.3171
R13985 ringtest_0.drv_out.n1 ringtest_0.drv_out.t2 10.8618
R13986 ringtest_0.drv_out.n20 ringtest_0.drv_out.t10 6.6005
R13987 ringtest_0.drv_out.n20 ringtest_0.drv_out.t5 6.6005
R13988 ringtest_0.drv_out.n17 ringtest_0.drv_out.t6 6.6005
R13989 ringtest_0.drv_out.n17 ringtest_0.drv_out.t8 6.6005
R13990 ringtest_0.drv_out.n19 ringtest_0.drv_out.t3 6.6005
R13991 ringtest_0.drv_out.n19 ringtest_0.drv_out.t4 6.6005
R13992 ringtest_0.drv_out.n18 ringtest_0.drv_out.t7 6.6005
R13993 ringtest_0.drv_out.n18 ringtest_0.drv_out.t9 6.6005
R13994 ringtest_0.drv_out.n11 ringtest_0.drv_out 5.69273
R13995 ringtest_0.drv_out.n12 ringtest_0.drv_out.t17 3.61217
R13996 ringtest_0.drv_out.n12 ringtest_0.drv_out.t12 3.61217
R13997 ringtest_0.drv_out.n14 ringtest_0.drv_out.t13 3.61217
R13998 ringtest_0.drv_out.n14 ringtest_0.drv_out.t15 3.61217
R13999 ringtest_0.drv_out.n13 ringtest_0.drv_out.t14 3.61217
R14000 ringtest_0.drv_out.n13 ringtest_0.drv_out.t16 3.61217
R14001 ringtest_0.drv_out.n15 ringtest_0.drv_out.t18 3.61217
R14002 ringtest_0.drv_out.n15 ringtest_0.drv_out.t11 3.61217
R14003 ringtest_0.drv_out.n2 ringtest_0.drv_out.n0 3.06895
R14004 ringtest_0.drv_out.n11 ringtest_0.drv_out 2.87193
R14005 ringtest_0.drv_out.n8 ringtest_0.drv_out 2.23542
R14006 ringtest_0.drv_out.n2 ringtest_0.drv_out.n1 2.14822
R14007 ringtest_0.drv_out.n10 ringtest_0.drv_out 1.7806
R14008 ringtest_0.drv_out ringtest_0.drv_out.n10 1.54574
R14009 ringtest_0.drv_out.n9 ringtest_0.drv_out 1.25273
R14010 ringtest_0.drv_out.n3 ringtest_0.drv_out.n2 1.12636
R14011 ringtest_0.drv_out ringtest_0.drv_out.n22 0.461707
R14012 ringtest_0.drv_out.n9 ringtest_0.drv_out 0.316378
R14013 ringtest_0.drv_out ringtest_0.drv_out.n11 0.188041
R14014 ringtest_0.drv_out ringtest_0.drv_out.n3 0.138152
R14015 ringtest_0.drv_out.n22 ringtest_0.drv_out.n16 0.0921193
R14016 ringtest_0.drv_out.n22 ringtest_0.drv_out.n21 0.069392
R14017 ringtest_0.drv_out.n3 ringtest_0.drv_out 0.0655
R14018 ringtest_0.drv_out.n10 ringtest_0.drv_out.n9 0.0596216
R14019 ringtest_0.x4.net3.t3 ringtest_0.x4.net3.t4 395.01
R14020 ringtest_0.x4.net3 ringtest_0.x4.net3.t3 320.745
R14021 ringtest_0.x4.net3.n3 ringtest_0.x4.net3.t6 260.322
R14022 ringtest_0.x4.net3.n0 ringtest_0.x4.net3.t7 229.369
R14023 ringtest_0.x4.net3.n7 ringtest_0.x4.net3.t1 222.68
R14024 ringtest_0.x4.net3.n3 ringtest_0.x4.net3.t5 175.169
R14025 ringtest_0.x4.net3.n0 ringtest_0.x4.net3.t2 157.07
R14026 ringtest_0.x4.net3.n4 ringtest_0.x4.net3.n3 152
R14027 ringtest_0.x4.net3.n1 ringtest_0.x4.net3.n0 152
R14028 ringtest_0.x4.net3.n8 ringtest_0.x4.net3.t0 132.322
R14029 ringtest_0.x4.net3.n8 ringtest_0.x4.net3.n7 95.0273
R14030 ringtest_0.x4.net3.n5 ringtest_0.x4.net3 25.2581
R14031 ringtest_0.x4.net3.n5 ringtest_0.x4.net3 20.1696
R14032 ringtest_0.x4.net3.n7 ringtest_0.x4.net3.n6 12.7813
R14033 ringtest_0.x4.net3.n1 ringtest_0.x4.net3 12.0005
R14034 ringtest_0.x4.net3 ringtest_0.x4.net3.n4 11.2497
R14035 ringtest_0.x4.net3.n6 ringtest_0.x4.net3.n2 9.79203
R14036 ringtest_0.x4.net3.n6 ringtest_0.x4.net3.n5 5.9277
R14037 ringtest_0.x4.net3.n2 ringtest_0.x4.net3 4.53383
R14038 ringtest_0.x4.net3 ringtest_0.x4.net3.n8 2.70465
R14039 ringtest_0.x4.net3.n2 ringtest_0.x4.net3.n1 1.6005
R14040 ringtest_0.x4.net3.n4 ringtest_0.x4.net3 1.55726
R14041 ui_in[2].n2 ui_in[2].t0 450.938
R14042 ui_in[2].n2 ui_in[2].t6 445.666
R14043 ui_in[2].n0 ui_in[2].t7 377.486
R14044 ui_in[2].n0 ui_in[2].t1 374.202
R14045 ui_in[2].n5 ui_in[2].t2 212.081
R14046 ui_in[2].n6 ui_in[2].t3 212.081
R14047 ui_in[2].n7 ui_in[2].n6 183.441
R14048 ui_in[2].n5 ui_in[2].t4 139.78
R14049 ui_in[2].n6 ui_in[2].t5 139.78
R14050 ui_in[2].n6 ui_in[2].n5 61.346
R14051 ui_in[2].n4 ui_in[2].n1 12.4088
R14052 ui_in[2] ui_in[2].n7 11.4331
R14053 ui_in[2].n4 ui_in[2].n3 9.10647
R14054 ui_in[2].n8 ui_in[2].n4 8.98648
R14055 ui_in[2].n7 ui_in[2] 5.6325
R14056 ui_in[2].n8 ui_in[2] 5.02323
R14057 ui_in[2].n3 ui_in[2].n2 3.1748
R14058 ui_in[2] ui_in[2].n0 2.04102
R14059 ui_in[2] ui_in[2].n8 0.888758
R14060 ui_in[2].n1 ui_in[2] 0.412375
R14061 ui_in[2].n3 ui_in[2] 0.063625
R14062 ui_in[2].n1 ui_in[2] 0.061125
R14063 ringtest_0.x3.x2.GP4.n2 ringtest_0.x3.x2.GP4.t5 450.938
R14064 ringtest_0.x3.x2.GP4.n2 ringtest_0.x3.x2.GP4.t4 445.666
R14065 ringtest_0.x3.x2.GP4.n5 ringtest_0.x3.x2.GP4.n4 208.965
R14066 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n0 96.8352
R14067 ringtest_0.x3.x2.GP4.n4 ringtest_0.x3.x2.GP4.t3 26.5955
R14068 ringtest_0.x3.x2.GP4.n4 ringtest_0.x3.x2.GP4.t2 26.5955
R14069 ringtest_0.x3.x2.GP4.n0 ringtest_0.x3.x2.GP4.t1 24.9236
R14070 ringtest_0.x3.x2.GP4.n0 ringtest_0.x3.x2.GP4.t0 24.9236
R14071 ringtest_0.x3.x1.gpo3 ringtest_0.x3.x2.x4.GP 16.5032
R14072 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n3 10.2405
R14073 ringtest_0.x3.x2.GP4.n3 ringtest_0.x3.x1.gpo3 7.76481
R14074 ringtest_0.x3.x2.GP4.n1 ringtest_0.x3.x1.x14.Y 6.1445
R14075 ringtest_0.x3.x2.GP4.n1 ringtest_0.x3.x1.x14.Y 4.65505
R14076 ringtest_0.x3.x2.x4.GP ringtest_0.x3.x2.GP4.n2 2.95993
R14077 ringtest_0.x3.x2.GP4.n5 ringtest_0.x3.x1.x14.Y 2.0485
R14078 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n5 1.55202
R14079 ringtest_0.x3.x2.GP4.n3 ringtest_0.x3.x2.GP4.n1 1.0245
R14080 ringtest_0.counter7.n0 ringtest_0.counter7.t5 368.521
R14081 ringtest_0.counter7.n1 ringtest_0.counter7.t4 216.155
R14082 ringtest_0.counter7.n1 ringtest_0.counter7 78.8791
R14083 ringtest_0.counter7.n4 ringtest_0.counter7.t0 26.3998
R14084 ringtest_0.counter7.n4 ringtest_0.counter7.t1 23.5483
R14085 ringtest_0.counter7.n3 ringtest_0.counter7.n2 18.2765
R14086 ringtest_0.counter7.n5 ringtest_0.counter7.t3 12.9758
R14087 ringtest_0.counter7.n5 ringtest_0.counter7.t2 10.8618
R14088 ringtest_0.counter7 ringtest_0.counter7.n0 10.5563
R14089 ringtest_0.counter7.n0 ringtest_0.counter7 5.48477
R14090 ringtest_0.counter7.n2 ringtest_0.counter7 4.18512
R14091 ringtest_0.counter7.n6 ringtest_0.counter7.n4 3.06895
R14092 ringtest_0.counter7.n6 ringtest_0.counter7.n5 2.14822
R14093 ringtest_0.counter7 ringtest_0.counter7.n6 1.27287
R14094 ringtest_0.counter7.n3 ringtest_0.counter7 1.27059
R14095 ringtest_0.counter7.n2 ringtest_0.counter7.n1 0.985115
R14096 ringtest_0.counter7 ringtest_0.counter7.n3 0.647091
R14097 ua[1].n6 ua[1].t12 23.6581
R14098 ua[1].n12 ua[1].t7 23.6581
R14099 ua[1].n19 ua[1].t2 23.6581
R14100 ua[1].n1 ua[1].t1 23.6581
R14101 ua[1].n5 ua[1].t4 23.3739
R14102 ua[1].n11 ua[1].t13 23.3739
R14103 ua[1].n18 ua[1].t3 23.3739
R14104 ua[1].n0 ua[1].t0 23.3739
R14105 ua[1].n25 ua[1] 15.3856
R14106 ua[1].n6 ua[1].t8 10.7528
R14107 ua[1].n12 ua[1].t11 10.7528
R14108 ua[1].n19 ua[1].t15 10.7528
R14109 ua[1].n1 ua[1].t5 10.7528
R14110 ua[1].n8 ua[1].t9 10.6417
R14111 ua[1].n14 ua[1].t10 10.6417
R14112 ua[1].n21 ua[1].t14 10.6417
R14113 ua[1].n3 ua[1].t6 10.6417
R14114 ua[1].n7 ua[1].n6 1.30064
R14115 ua[1].n13 ua[1].n12 1.30064
R14116 ua[1].n20 ua[1].n19 1.30064
R14117 ua[1].n2 ua[1].n1 1.30064
R14118 ua[1] ua[1].n4 0.983856
R14119 ua[1].n23 ua[1].n22 0.946356
R14120 ua[1].n16 ua[1].n15 0.927606
R14121 ua[1].n10 ua[1].n9 0.925106
R14122 ua[1].n17 ua[1] 0.748625
R14123 ua[1].n7 ua[1].n5 0.726502
R14124 ua[1].n13 ua[1].n11 0.726502
R14125 ua[1].n20 ua[1].n18 0.726502
R14126 ua[1].n2 ua[1].n0 0.726502
R14127 ua[1].n24 ua[1].n17 0.54425
R14128 ua[1].n25 ua[1] 0.532375
R14129 ua[1].n8 ua[1].n7 0.512491
R14130 ua[1].n14 ua[1].n13 0.512491
R14131 ua[1].n21 ua[1].n20 0.512491
R14132 ua[1].n3 ua[1].n2 0.512491
R14133 ua[1].n9 ua[1].n8 0.359663
R14134 ua[1].n15 ua[1].n14 0.359663
R14135 ua[1].n22 ua[1].n21 0.359663
R14136 ua[1].n4 ua[1].n3 0.359663
R14137 ua[1].n9 ua[1].n5 0.216071
R14138 ua[1].n15 ua[1].n11 0.216071
R14139 ua[1].n22 ua[1].n18 0.216071
R14140 ua[1].n4 ua[1].n0 0.216071
R14141 ua[1].n17 ua[1] 0.20175
R14142 ua[1].n24 ua[1] 0.17925
R14143 ua[1] ua[1].n25 0.178
R14144 ua[1].n24 ua[1] 0.063
R14145 ua[1].n10 ua[1] 0.05925
R14146 ua[1].n16 ua[1] 0.05675
R14147 ua[1] ua[1].n16 0.0561931
R14148 ua[1] ua[1].n10 0.0561872
R14149 ua[1].n23 ua[1] 0.038
R14150 ua[1] ua[1].n23 0.0376287
R14151 ua[1] ua[1].n24 0.004875
R14152 ringtest_0.x4.clknet_1_0__leaf_clk.n25 ringtest_0.x4.clknet_1_0__leaf_clk.n23 333.392
R14153 ringtest_0.x4.clknet_1_0__leaf_clk.n25 ringtest_0.x4.clknet_1_0__leaf_clk.n24 301.392
R14154 ringtest_0.x4.clknet_1_0__leaf_clk.n27 ringtest_0.x4.clknet_1_0__leaf_clk.n26 301.392
R14155 ringtest_0.x4.clknet_1_0__leaf_clk.n29 ringtest_0.x4.clknet_1_0__leaf_clk.n28 301.392
R14156 ringtest_0.x4.clknet_1_0__leaf_clk.n22 ringtest_0.x4.clknet_1_0__leaf_clk.n4 301.392
R14157 ringtest_0.x4.clknet_1_0__leaf_clk.n31 ringtest_0.x4.clknet_1_0__leaf_clk.n30 301.392
R14158 ringtest_0.x4.clknet_1_0__leaf_clk.n21 ringtest_0.x4.clknet_1_0__leaf_clk.n5 297.863
R14159 ringtest_0.x4.clknet_1_0__leaf_clk.n2 ringtest_0.x4.clknet_1_0__leaf_clk.t32 294.557
R14160 ringtest_0.x4.clknet_1_0__leaf_clk.n0 ringtest_0.x4.clknet_1_0__leaf_clk.t38 294.557
R14161 ringtest_0.x4.clknet_1_0__leaf_clk.n41 ringtest_0.x4.clknet_1_0__leaf_clk.t35 294.557
R14162 ringtest_0.x4.clknet_1_0__leaf_clk.n38 ringtest_0.x4.clknet_1_0__leaf_clk.t33 294.557
R14163 ringtest_0.x4.clknet_1_0__leaf_clk.n36 ringtest_0.x4.clknet_1_0__leaf_clk.t36 294.557
R14164 ringtest_0.x4.clknet_1_0__leaf_clk.n34 ringtest_0.x4.clknet_1_0__leaf_clk.n33 287.303
R14165 ringtest_0.x4.clknet_1_0__leaf_clk.n8 ringtest_0.x4.clknet_1_0__leaf_clk.n6 248.638
R14166 ringtest_0.x4.clknet_1_0__leaf_clk.n2 ringtest_0.x4.clknet_1_0__leaf_clk.t37 211.01
R14167 ringtest_0.x4.clknet_1_0__leaf_clk.n0 ringtest_0.x4.clknet_1_0__leaf_clk.t41 211.01
R14168 ringtest_0.x4.clknet_1_0__leaf_clk.n41 ringtest_0.x4.clknet_1_0__leaf_clk.t34 211.01
R14169 ringtest_0.x4.clknet_1_0__leaf_clk.n38 ringtest_0.x4.clknet_1_0__leaf_clk.t40 211.01
R14170 ringtest_0.x4.clknet_1_0__leaf_clk.n36 ringtest_0.x4.clknet_1_0__leaf_clk.t39 211.01
R14171 ringtest_0.x4.clknet_1_0__leaf_clk.n8 ringtest_0.x4.clknet_1_0__leaf_clk.n7 203.463
R14172 ringtest_0.x4.clknet_1_0__leaf_clk.n10 ringtest_0.x4.clknet_1_0__leaf_clk.n9 203.463
R14173 ringtest_0.x4.clknet_1_0__leaf_clk.n14 ringtest_0.x4.clknet_1_0__leaf_clk.n13 203.463
R14174 ringtest_0.x4.clknet_1_0__leaf_clk.n16 ringtest_0.x4.clknet_1_0__leaf_clk.n15 203.463
R14175 ringtest_0.x4.clknet_1_0__leaf_clk.n18 ringtest_0.x4.clknet_1_0__leaf_clk.n17 203.463
R14176 ringtest_0.x4.clknet_1_0__leaf_clk.n12 ringtest_0.x4.clknet_1_0__leaf_clk.n11 202.456
R14177 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n19 199.607
R14178 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n2 156.207
R14179 ringtest_0.x4.clknet_1_0__leaf_clk.n37 ringtest_0.x4.clknet_1_0__leaf_clk.n36 153.097
R14180 ringtest_0.x4.clknet_1_0__leaf_clk.n39 ringtest_0.x4.clknet_1_0__leaf_clk.n38 152.296
R14181 ringtest_0.x4.clknet_1_0__leaf_clk.n1 ringtest_0.x4.clknet_1_0__leaf_clk.n0 152
R14182 ringtest_0.x4.clknet_1_0__leaf_clk.n42 ringtest_0.x4.clknet_1_0__leaf_clk.n41 152
R14183 ringtest_0.x4.clknet_1_0__leaf_clk.n10 ringtest_0.x4.clknet_1_0__leaf_clk.n8 45.177
R14184 ringtest_0.x4.clknet_1_0__leaf_clk.n16 ringtest_0.x4.clknet_1_0__leaf_clk.n14 45.177
R14185 ringtest_0.x4.clknet_1_0__leaf_clk.n18 ringtest_0.x4.clknet_1_0__leaf_clk.n16 45.177
R14186 ringtest_0.x4.clknet_1_0__leaf_clk.n12 ringtest_0.x4.clknet_1_0__leaf_clk.n10 44.0476
R14187 ringtest_0.x4.clknet_1_0__leaf_clk.n14 ringtest_0.x4.clknet_1_0__leaf_clk.n12 44.0476
R14188 ringtest_0.x4.clknet_1_0__leaf_clk.n6 ringtest_0.x4.clknet_1_0__leaf_clk.t8 40.0005
R14189 ringtest_0.x4.clknet_1_0__leaf_clk.n6 ringtest_0.x4.clknet_1_0__leaf_clk.t11 40.0005
R14190 ringtest_0.x4.clknet_1_0__leaf_clk.n7 ringtest_0.x4.clknet_1_0__leaf_clk.t13 40.0005
R14191 ringtest_0.x4.clknet_1_0__leaf_clk.n7 ringtest_0.x4.clknet_1_0__leaf_clk.t15 40.0005
R14192 ringtest_0.x4.clknet_1_0__leaf_clk.n9 ringtest_0.x4.clknet_1_0__leaf_clk.t10 40.0005
R14193 ringtest_0.x4.clknet_1_0__leaf_clk.n9 ringtest_0.x4.clknet_1_0__leaf_clk.t12 40.0005
R14194 ringtest_0.x4.clknet_1_0__leaf_clk.n11 ringtest_0.x4.clknet_1_0__leaf_clk.t14 40.0005
R14195 ringtest_0.x4.clknet_1_0__leaf_clk.n11 ringtest_0.x4.clknet_1_0__leaf_clk.t9 40.0005
R14196 ringtest_0.x4.clknet_1_0__leaf_clk.n13 ringtest_0.x4.clknet_1_0__leaf_clk.t1 40.0005
R14197 ringtest_0.x4.clknet_1_0__leaf_clk.n13 ringtest_0.x4.clknet_1_0__leaf_clk.t4 40.0005
R14198 ringtest_0.x4.clknet_1_0__leaf_clk.n15 ringtest_0.x4.clknet_1_0__leaf_clk.t6 40.0005
R14199 ringtest_0.x4.clknet_1_0__leaf_clk.n15 ringtest_0.x4.clknet_1_0__leaf_clk.t7 40.0005
R14200 ringtest_0.x4.clknet_1_0__leaf_clk.n17 ringtest_0.x4.clknet_1_0__leaf_clk.t3 40.0005
R14201 ringtest_0.x4.clknet_1_0__leaf_clk.n17 ringtest_0.x4.clknet_1_0__leaf_clk.t5 40.0005
R14202 ringtest_0.x4.clknet_1_0__leaf_clk.n19 ringtest_0.x4.clknet_1_0__leaf_clk.t0 40.0005
R14203 ringtest_0.x4.clknet_1_0__leaf_clk.n19 ringtest_0.x4.clknet_1_0__leaf_clk.t2 40.0005
R14204 ringtest_0.x4.clknet_1_0__leaf_clk.n27 ringtest_0.x4.clknet_1_0__leaf_clk.n25 32.0005
R14205 ringtest_0.x4.clknet_1_0__leaf_clk.n29 ringtest_0.x4.clknet_1_0__leaf_clk.n27 32.0005
R14206 ringtest_0.x4.clknet_1_0__leaf_clk.n32 ringtest_0.x4.clknet_1_0__leaf_clk.n22 32.0005
R14207 ringtest_0.x4.clknet_1_0__leaf_clk.n32 ringtest_0.x4.clknet_1_0__leaf_clk.n31 32.0005
R14208 ringtest_0.x4.clknet_1_0__leaf_clk.n31 ringtest_0.x4.clknet_1_0__leaf_clk.n29 31.2005
R14209 ringtest_0.x4.clknet_1_0__leaf_clk.n35 ringtest_0.x4.clknet_1_0__leaf_clk.n34 28.6283
R14210 ringtest_0.x4.clknet_1_0__leaf_clk.n3 ringtest_0.x4.clknet_1_0__leaf_clk 28.0697
R14211 ringtest_0.x4.clknet_1_0__leaf_clk.n23 ringtest_0.x4.clknet_1_0__leaf_clk.t19 27.5805
R14212 ringtest_0.x4.clknet_1_0__leaf_clk.n23 ringtest_0.x4.clknet_1_0__leaf_clk.t22 27.5805
R14213 ringtest_0.x4.clknet_1_0__leaf_clk.n24 ringtest_0.x4.clknet_1_0__leaf_clk.t24 27.5805
R14214 ringtest_0.x4.clknet_1_0__leaf_clk.n24 ringtest_0.x4.clknet_1_0__leaf_clk.t26 27.5805
R14215 ringtest_0.x4.clknet_1_0__leaf_clk.n26 ringtest_0.x4.clknet_1_0__leaf_clk.t21 27.5805
R14216 ringtest_0.x4.clknet_1_0__leaf_clk.n26 ringtest_0.x4.clknet_1_0__leaf_clk.t23 27.5805
R14217 ringtest_0.x4.clknet_1_0__leaf_clk.n28 ringtest_0.x4.clknet_1_0__leaf_clk.t25 27.5805
R14218 ringtest_0.x4.clknet_1_0__leaf_clk.n28 ringtest_0.x4.clknet_1_0__leaf_clk.t20 27.5805
R14219 ringtest_0.x4.clknet_1_0__leaf_clk.n4 ringtest_0.x4.clknet_1_0__leaf_clk.t30 27.5805
R14220 ringtest_0.x4.clknet_1_0__leaf_clk.n4 ringtest_0.x4.clknet_1_0__leaf_clk.t16 27.5805
R14221 ringtest_0.x4.clknet_1_0__leaf_clk.n5 ringtest_0.x4.clknet_1_0__leaf_clk.t27 27.5805
R14222 ringtest_0.x4.clknet_1_0__leaf_clk.n5 ringtest_0.x4.clknet_1_0__leaf_clk.t29 27.5805
R14223 ringtest_0.x4.clknet_1_0__leaf_clk.n33 ringtest_0.x4.clknet_1_0__leaf_clk.t17 27.5805
R14224 ringtest_0.x4.clknet_1_0__leaf_clk.n33 ringtest_0.x4.clknet_1_0__leaf_clk.t18 27.5805
R14225 ringtest_0.x4.clknet_1_0__leaf_clk.n30 ringtest_0.x4.clknet_1_0__leaf_clk.t28 27.5805
R14226 ringtest_0.x4.clknet_1_0__leaf_clk.n30 ringtest_0.x4.clknet_1_0__leaf_clk.t31 27.5805
R14227 ringtest_0.x4.clknet_1_0__leaf_clk.n43 ringtest_0.x4.clknet_1_0__leaf_clk.n42 27.3319
R14228 ringtest_0.x4.clknet_1_0__leaf_clk.n40 ringtest_0.x4.clknet_1_0__leaf_clk.n39 21.4985
R14229 ringtest_0.x4.clknet_1_0__leaf_clk.n3 ringtest_0.x4.clknet_1_0__leaf_clk.n1 21.401
R14230 ringtest_0.x4.clknet_1_0__leaf_clk.n34 ringtest_0.x4.clknet_1_0__leaf_clk.n32 14.0898
R14231 ringtest_0.x4.clknet_1_0__leaf_clk.n20 ringtest_0.x4.clknet_1_0__leaf_clk.n18 13.177
R14232 ringtest_0.x4.clknet_1_0__leaf_clk.n40 ringtest_0.x4.clknet_1_0__leaf_clk.n37 11.0654
R14233 ringtest_0.x4.clknet_1_0__leaf_clk.n22 ringtest_0.x4.clknet_1_0__leaf_clk.n21 10.4484
R14234 ringtest_0.x4.clknet_1_0__leaf_clk.n43 ringtest_0.x4.clknet_1_0__leaf_clk.n40 7.18319
R14235 ringtest_0.x4.clknet_1_0__leaf_clk.n35 ringtest_0.x4.clknet_1_0__leaf_clk.n3 5.63649
R14236 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n20 3.13183
R14237 ringtest_0.x4.clknet_1_0__leaf_clk.n37 ringtest_0.x4.clknet_1_0__leaf_clk 3.10907
R14238 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n43 2.66671
R14239 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n35 2.66671
R14240 ringtest_0.x4.clknet_1_0__leaf_clk.n42 ringtest_0.x4.clknet_1_0__leaf_clk 2.01193
R14241 ringtest_0.x4.clknet_1_0__leaf_clk.n21 ringtest_0.x4.clknet_1_0__leaf_clk 1.75844
R14242 ringtest_0.x4.clknet_1_0__leaf_clk.n39 ringtest_0.x4.clknet_1_0__leaf_clk 1.67435
R14243 ringtest_0.x4.clknet_1_0__leaf_clk.n1 ringtest_0.x4.clknet_1_0__leaf_clk 1.37896
R14244 ringtest_0.x4.clknet_1_0__leaf_clk.n20 ringtest_0.x4.clknet_1_0__leaf_clk 0.604792
R14245 ringtest_0.counter3.n0 ringtest_0.counter3.t3 368.521
R14246 ringtest_0.counter3.n1 ringtest_0.counter3.t2 216.155
R14247 ringtest_0.counter3.n1 ringtest_0.counter3 78.8791
R14248 ringtest_0.counter3.n4 ringtest_0.counter3.t1 26.3998
R14249 ringtest_0.counter3.n4 ringtest_0.counter3.t0 23.5483
R14250 ringtest_0.counter3.n3 ringtest_0.counter3.n2 17.5689
R14251 ringtest_0.counter3.n5 ringtest_0.counter3.t5 12.9693
R14252 ringtest_0.counter3.n5 ringtest_0.counter3.t4 10.8444
R14253 ringtest_0.counter3 ringtest_0.counter3.n0 10.5563
R14254 ringtest_0.counter3.n0 ringtest_0.counter3 5.48477
R14255 ringtest_0.counter3.n2 ringtest_0.counter3 4.18512
R14256 ringtest_0.counter3.n6 ringtest_0.counter3.n4 3.06895
R14257 ringtest_0.counter3.n6 ringtest_0.counter3.n5 2.14822
R14258 ringtest_0.counter3.n3 ringtest_0.counter3 1.28175
R14259 ringtest_0.counter3 ringtest_0.counter3.n6 1.25828
R14260 ringtest_0.counter3.n2 ringtest_0.counter3.n1 0.985115
R14261 ringtest_0.counter3 ringtest_0.counter3.n3 0.688
R14262 muxtest_0.x1.x3.GP2.n3 muxtest_0.x1.x3.GP2.t4 450.938
R14263 muxtest_0.x1.x3.GP2.n2 muxtest_0.x1.x3.GP2.t7 450.938
R14264 muxtest_0.x1.x3.GP2.n3 muxtest_0.x1.x3.GP2.t5 445.666
R14265 muxtest_0.x1.x3.GP2.n2 muxtest_0.x1.x3.GP2.t6 445.666
R14266 muxtest_0.x1.x3.GP2.n6 muxtest_0.x1.x3.GP2.n5 195.958
R14267 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n0 96.8352
R14268 muxtest_0.x1.x3.GP2.n5 muxtest_0.x1.x3.GP2.t2 26.5955
R14269 muxtest_0.x1.x3.GP2.n5 muxtest_0.x1.x3.GP2.t3 26.5955
R14270 muxtest_0.x1.x3.GP2.n0 muxtest_0.x1.x3.GP2.t0 24.9236
R14271 muxtest_0.x1.x3.GP2.n0 muxtest_0.x1.x3.GP2.t1 24.9236
R14272 muxtest_0.x1.x3.GP2.n4 muxtest_0.x1.x3.GP2 14.8953
R14273 muxtest_0.x1.x3.GP2.n7 muxtest_0.x1.x3.GP2.n6 13.0077
R14274 muxtest_0.x1.x3.GP2.n6 muxtest_0.x1.x3.GP2 11.8741
R14275 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n1 11.2645
R14276 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n4 8.64182
R14277 muxtest_0.x1.x3.GP2.n1 muxtest_0.x1.x3.GP2 6.1445
R14278 muxtest_0.x1.x3.GP2.n4 muxtest_0.x1.x3.GP2 5.75481
R14279 muxtest_0.x1.x3.GP2.n1 muxtest_0.x1.x3.GP2 4.65505
R14280 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n2 3.12276
R14281 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n3 2.94361
R14282 muxtest_0.x1.x3.GP2.n7 muxtest_0.x1.x3.GP2 2.0485
R14283 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n7 1.55202
R14284 muxtest_0.R5R6.n0 muxtest_0.R5R6.t0 26.3998
R14285 muxtest_0.R5R6.n0 muxtest_0.R5R6.t1 23.5483
R14286 muxtest_0.R5R6.n1 muxtest_0.R5R6.t4 12.9758
R14287 muxtest_0.R5R6.n1 muxtest_0.R5R6.t5 10.8618
R14288 muxtest_0.R5R6.n4 muxtest_0.R5R6.t3 10.55
R14289 muxtest_0.R5R6.n2 muxtest_0.R5R6.n0 3.06895
R14290 muxtest_0.R5R6.n2 muxtest_0.R5R6.n1 2.14822
R14291 muxtest_0.R5R6.n3 muxtest_0.R5R6.n2 1.12636
R14292 muxtest_0.R5R6.n4 muxtest_0.R5R6.t2 1.11543
R14293 muxtest_0.R5R6 muxtest_0.R5R6.n4 0.694875
R14294 muxtest_0.R5R6 muxtest_0.R5R6.n3 0.132418
R14295 muxtest_0.R5R6.n3 muxtest_0.R5R6 0.0655
R14296 ringtest_0.x4._16_.n12 ringtest_0.x4._16_.t1 339.418
R14297 ringtest_0.x4._16_ ringtest_0.x4._16_.t0 269.426
R14298 ringtest_0.x4._16_.n1 ringtest_0.x4._16_.t7 264.029
R14299 ringtest_0.x4._16_ ringtest_0.x4._16_.n5 241.976
R14300 ringtest_0.x4._16_.n3 ringtest_0.x4._16_.t3 241.536
R14301 ringtest_0.x4._16_.n5 ringtest_0.x4._16_.t8 241.536
R14302 ringtest_0.x4._16_.n1 ringtest_0.x4._16_.t2 206.19
R14303 ringtest_0.x4._16_.n4 ringtest_0.x4._16_.n3 171.332
R14304 ringtest_0.x4._16_.n3 ringtest_0.x4._16_.t9 169.237
R14305 ringtest_0.x4._16_.n5 ringtest_0.x4._16_.t4 169.237
R14306 ringtest_0.x4._16_.n2 ringtest_0.x4._16_.n1 160.96
R14307 ringtest_0.x4._16_.n9 ringtest_0.x4._16_.n8 153.165
R14308 ringtest_0.x4._16_.n8 ringtest_0.x4._16_.t6 144.548
R14309 ringtest_0.x4._16_.n8 ringtest_0.x4._16_.t5 128.482
R14310 ringtest_0.x4._16_.n7 ringtest_0.x4._16_.n2 21.45
R14311 ringtest_0.x4._16_.n7 ringtest_0.x4._16_.n6 16.7975
R14312 ringtest_0.x4._16_.n10 ringtest_0.x4._16_ 15.8161
R14313 ringtest_0.x4._16_.n11 ringtest_0.x4._16_.n10 14.0946
R14314 ringtest_0.x4._16_ ringtest_0.x4._16_.n0 11.2645
R14315 ringtest_0.x4._16_ ringtest_0.x4._16_.n9 9.55788
R14316 ringtest_0.x4._16_.n6 ringtest_0.x4._16_ 6.4005
R14317 ringtest_0.x4._16_.n0 ringtest_0.x4._16_ 6.1445
R14318 ringtest_0.x4._16_.n2 ringtest_0.x4._16_ 5.4405
R14319 ringtest_0.x4._16_.n0 ringtest_0.x4._16_ 4.63498
R14320 ringtest_0.x4._16_.n4 ringtest_0.x4._16_ 4.44132
R14321 ringtest_0.x4._16_.n11 ringtest_0.x4._16_ 4.3525
R14322 ringtest_0.x4._16_.n13 ringtest_0.x4._16_.n12 4.0914
R14323 ringtest_0.x4._16_ ringtest_0.x4._16_.n13 3.61789
R14324 ringtest_0.x4._16_.n9 ringtest_0.x4._16_ 3.29747
R14325 ringtest_0.x4._16_.n13 ringtest_0.x4._16_.n11 2.3045
R14326 ringtest_0.x4._16_.n12 ringtest_0.x4._16_ 1.74382
R14327 ringtest_0.x4._16_.n6 ringtest_0.x4._16_.n4 1.50638
R14328 ringtest_0.x4._16_.n10 ringtest_0.x4._16_.n7 1.38649
R14329 muxtest_0.x2.x2.GP2.n2 muxtest_0.x2.x2.GP2.t4 450.938
R14330 muxtest_0.x2.x2.GP2.n2 muxtest_0.x2.x2.GP2.t5 445.666
R14331 muxtest_0.x2.x2.GP2.n4 muxtest_0.x2.x2.GP2.n3 195.958
R14332 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n0 96.8352
R14333 muxtest_0.x2.x2.GP2.n3 muxtest_0.x2.x2.GP2.t3 26.5955
R14334 muxtest_0.x2.x2.GP2.n3 muxtest_0.x2.x2.GP2.t2 26.5955
R14335 muxtest_0.x2.x2.GP2.n0 muxtest_0.x2.x2.GP2.t0 24.9236
R14336 muxtest_0.x2.x2.GP2.n0 muxtest_0.x2.x2.GP2.t1 24.9236
R14337 muxtest_0.x2.x2.GP2.n5 muxtest_0.x2.x2.GP2.n4 13.0077
R14338 muxtest_0.x2.x2.GP2.n4 muxtest_0.x2.x2.GP2 11.995
R14339 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n1 11.2645
R14340 muxtest_0.x2.x2.GP2.n1 muxtest_0.x2.x2.GP2 6.1445
R14341 muxtest_0.x2.x2.GP2.n1 muxtest_0.x2.x2.GP2 4.65505
R14342 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n2 3.12839
R14343 muxtest_0.x2.x2.GP2.n5 muxtest_0.x2.x2.GP2 2.0485
R14344 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n5 1.55202
R14345 muxtest_0.R6R7.n0 muxtest_0.R6R7.t1 26.3998
R14346 muxtest_0.R6R7.n0 muxtest_0.R6R7.t0 23.5483
R14347 muxtest_0.R6R7.n4 muxtest_0.R6R7.t4 17.4454
R14348 muxtest_0.R6R7.n1 muxtest_0.R6R7.t3 12.9758
R14349 muxtest_0.R6R7.n1 muxtest_0.R6R7.t2 10.8618
R14350 muxtest_0.R6R7.n4 muxtest_0.R6R7.t5 10.5739
R14351 muxtest_0.R6R7.n2 muxtest_0.R6R7.n0 3.06895
R14352 muxtest_0.R6R7.n2 muxtest_0.R6R7.n1 2.14822
R14353 muxtest_0.R6R7.n3 muxtest_0.R6R7.n2 1.12636
R14354 muxtest_0.R6R7.n5 muxtest_0.R6R7 1.11925
R14355 muxtest_0.R6R7.n5 muxtest_0.R6R7.n4 0.370193
R14356 muxtest_0.R6R7 muxtest_0.R6R7.n3 0.138152
R14357 muxtest_0.R6R7.n5 muxtest_0.R6R7 0.073
R14358 muxtest_0.R6R7.n3 muxtest_0.R6R7 0.0655
R14359 muxtest_0.R6R7 muxtest_0.R6R7.n5 0.04925
R14360 ua[0].n6 ua[0].t3 26.3998
R14361 ua[0].n0 ua[0].t5 26.3998
R14362 ua[0].n6 ua[0].t2 23.5483
R14363 ua[0].n0 ua[0].t6 23.5483
R14364 ua[0].n7 ua[0].t0 12.9758
R14365 ua[0].n1 ua[0].t7 12.9758
R14366 ua[0].n5 ua[0] 12.8371
R14367 ua[0].n7 ua[0].t1 10.8618
R14368 ua[0].n1 ua[0].t8 10.8618
R14369 ua[0].n4 ua[0].t4 10.5739
R14370 ua[0].n8 ua[0].n6 3.06895
R14371 ua[0].n2 ua[0].n0 3.06895
R14372 ua[0].n8 ua[0].n7 2.14822
R14373 ua[0].n2 ua[0].n1 2.14822
R14374 ua[0].n4 ua[0] 1.39577
R14375 ua[0].n9 ua[0].n8 1.12636
R14376 ua[0].n3 ua[0].n2 1.12636
R14377 ua[0].n5 ua[0].n4 0.545106
R14378 ua[0] ua[0].n9 0.138152
R14379 ua[0] ua[0].n3 0.134513
R14380 ua[0].n9 ua[0] 0.0655
R14381 ua[0].n3 ua[0] 0.0655
R14382 ua[0] ua[0].n5 0.0579534
R14383 ua[0].n5 ua[0] 0.0532872
R14384 muxtest_0.R7R8.n5 muxtest_0.R7R8.t5 26.3998
R14385 muxtest_0.R7R8.n0 muxtest_0.R7R8.t4 26.3998
R14386 muxtest_0.R7R8.n5 muxtest_0.R7R8.t6 23.5483
R14387 muxtest_0.R7R8.n0 muxtest_0.R7R8.t3 23.5483
R14388 muxtest_0.R7R8.n6 muxtest_0.R7R8.t8 12.9758
R14389 muxtest_0.R7R8.n1 muxtest_0.R7R8.t1 12.9758
R14390 muxtest_0.R7R8.n6 muxtest_0.R7R8.t7 10.8618
R14391 muxtest_0.R7R8.n1 muxtest_0.R7R8.t0 10.8618
R14392 muxtest_0.R7R8.n4 muxtest_0.R7R8.t9 10.5709
R14393 muxtest_0.R7R8.n9 muxtest_0.R7R8 8.65896
R14394 muxtest_0.R7R8.n7 muxtest_0.R7R8.n5 3.06895
R14395 muxtest_0.R7R8.n2 muxtest_0.R7R8.n0 3.06895
R14396 muxtest_0.R7R8.n7 muxtest_0.R7R8.n6 2.14822
R14397 muxtest_0.R7R8.n2 muxtest_0.R7R8.n1 2.14822
R14398 muxtest_0.R7R8.n8 muxtest_0.R7R8.n7 1.12636
R14399 muxtest_0.R7R8.n3 muxtest_0.R7R8.n2 1.12636
R14400 muxtest_0.R7R8.n4 muxtest_0.R7R8.t2 1.01856
R14401 muxtest_0.R7R8 muxtest_0.R7R8.n9 0.32175
R14402 muxtest_0.R7R8.n9 muxtest_0.R7R8.n4 0.230945
R14403 muxtest_0.R7R8 muxtest_0.R7R8.n3 0.148615
R14404 muxtest_0.R7R8 muxtest_0.R7R8.n8 0.134513
R14405 muxtest_0.R7R8.n8 muxtest_0.R7R8 0.0655
R14406 muxtest_0.R7R8.n3 muxtest_0.R7R8 0.0655
R14407 ui_in[3].n18 ui_in[3].t0 327.99
R14408 ui_in[3].n5 ui_in[3].t19 327.99
R14409 ui_in[3].n22 ui_in[3].t4 293.969
R14410 ui_in[3].n9 ui_in[3].t17 293.969
R14411 ui_in[3].n16 ui_in[3].t11 261.887
R14412 ui_in[3].n3 ui_in[3].t10 261.887
R14413 ui_in[3].n13 ui_in[3].t5 212.081
R14414 ui_in[3].n14 ui_in[3].t8 212.081
R14415 ui_in[3].n0 ui_in[3].t18 212.081
R14416 ui_in[3].n1 ui_in[3].t3 212.081
R14417 ui_in[3].n18 ui_in[3].t14 199.457
R14418 ui_in[3].n5 ui_in[3].t9 199.457
R14419 ui_in[3].n15 ui_in[3].n14 183.185
R14420 ui_in[3].n2 ui_in[3].n1 183.185
R14421 ui_in[3].n16 ui_in[3].t7 155.847
R14422 ui_in[3].n3 ui_in[3].t6 155.847
R14423 ui_in[3] ui_in[3].n22 154.065
R14424 ui_in[3] ui_in[3].n9 154.065
R14425 ui_in[3].n17 ui_in[3].n16 153.506
R14426 ui_in[3].n4 ui_in[3].n3 153.506
R14427 ui_in[3].n19 ui_in[3].n18 152
R14428 ui_in[3].n6 ui_in[3].n5 152
R14429 ui_in[3].n13 ui_in[3].t13 139.78
R14430 ui_in[3].n14 ui_in[3].t16 139.78
R14431 ui_in[3].n0 ui_in[3].t2 139.78
R14432 ui_in[3].n1 ui_in[3].t12 139.78
R14433 ui_in[3].n22 ui_in[3].t1 138.338
R14434 ui_in[3].n9 ui_in[3].t15 138.338
R14435 ui_in[3].n14 ui_in[3].n13 61.346
R14436 ui_in[3].n1 ui_in[3].n0 61.346
R14437 ui_in[3].n26 ui_in[3] 35.166
R14438 ui_in[3].n23 ui_in[3] 13.4199
R14439 ui_in[3].n10 ui_in[3] 13.4199
R14440 ui_in[3].n26 ui_in[3] 12.2088
R14441 ui_in[3].n24 ui_in[3].n21 11.7395
R14442 ui_in[3].n11 ui_in[3].n8 11.7395
R14443 ui_in[3].n25 ui_in[3].n24 11.5949
R14444 ui_in[3].n12 ui_in[3].n11 11.5949
R14445 ui_in[3].n21 ui_in[3].n17 10.4004
R14446 ui_in[3].n8 ui_in[3].n4 10.4004
R14447 ui_in[3].n25 ui_in[3].n15 9.68118
R14448 ui_in[3].n12 ui_in[3].n2 9.68118
R14449 ui_in[3].n19 ui_in[3] 9.6005
R14450 ui_in[3].n6 ui_in[3] 9.6005
R14451 ui_in[3].n15 ui_in[3] 5.8885
R14452 ui_in[3].n2 ui_in[3] 5.8885
R14453 ui_in[3].n23 ui_in[3] 5.57469
R14454 ui_in[3].n10 ui_in[3] 5.57469
R14455 ui_in[3].n21 ui_in[3].n20 4.6505
R14456 ui_in[3].n24 ui_in[3].n23 4.6505
R14457 ui_in[3].n8 ui_in[3].n7 4.6505
R14458 ui_in[3].n11 ui_in[3].n10 4.6505
R14459 ui_in[3].n20 ui_in[3].n19 2.98717
R14460 ui_in[3].n7 ui_in[3].n6 2.98717
R14461 ui_in[3].n17 ui_in[3] 2.82403
R14462 ui_in[3].n4 ui_in[3] 2.82403
R14463 ui_in[3].n20 ui_in[3] 1.9205
R14464 ui_in[3].n7 ui_in[3] 1.9205
R14465 ui_in[3] ui_in[3].n25 0.559212
R14466 ui_in[3] ui_in[3].n12 0.559212
R14467 ui_in[3] ui_in[3].n26 0.47425
R14468 ringtest_0.x3.x2.GP1.n2 ringtest_0.x3.x2.GP1.t5 450.938
R14469 ringtest_0.x3.x2.GP1.n2 ringtest_0.x3.x2.GP1.t4 445.666
R14470 ringtest_0.x3.x2.GP1.n4 ringtest_0.x3.x2.GP1.n3 195.832
R14471 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n0 96.8352
R14472 ringtest_0.x3.x2.GP1.n3 ringtest_0.x3.x2.GP1.t3 26.5955
R14473 ringtest_0.x3.x2.GP1.n3 ringtest_0.x3.x2.GP1.t2 26.5955
R14474 ringtest_0.x3.x2.GP1.n0 ringtest_0.x3.x2.GP1.t1 24.9236
R14475 ringtest_0.x3.x2.GP1.n0 ringtest_0.x3.x2.GP1.t0 24.9236
R14476 ringtest_0.x3.x2.GP1.n5 ringtest_0.x3.x2.GP1.n4 13.1346
R14477 ringtest_0.x3.x2.GP1.n4 ringtest_0.x3.x2.GP1 12.2007
R14478 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n1 11.2645
R14479 ringtest_0.x3.x2.GP1.n1 ringtest_0.x3.x2.GP1 6.1445
R14480 ringtest_0.x3.x2.GP1.n1 ringtest_0.x3.x2.GP1 4.65505
R14481 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n2 3.07707
R14482 ringtest_0.x3.x2.GP1.n5 ringtest_0.x3.x2.GP1 2.0485
R14483 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n5 1.55202
R14484 ringtest_0.ring_out.n0 ringtest_0.ring_out.t13 844.321
R14485 ringtest_0.ring_out.n0 ringtest_0.ring_out.t12 354.322
R14486 ringtest_0.ring_out.n3 ringtest_0.ring_out.n1 243.68
R14487 ringtest_0.ring_out.n8 ringtest_0.ring_out.t10 212.081
R14488 ringtest_0.ring_out.n7 ringtest_0.ring_out.t11 212.081
R14489 ringtest_0.ring_out.n5 ringtest_0.ring_out.n4 206.249
R14490 ringtest_0.ring_out.n3 ringtest_0.ring_out.n2 205.28
R14491 ringtest_0.ring_out.n9 ringtest_0.ring_out.n8 184.806
R14492 ringtest_0.ring_out.n8 ringtest_0.ring_out.t14 139.78
R14493 ringtest_0.ring_out.n7 ringtest_0.ring_out.t15 139.78
R14494 ringtest_0.ring_out.n8 ringtest_0.ring_out.n7 61.346
R14495 ringtest_0.ring_out.n1 ringtest_0.ring_out.t2 26.5955
R14496 ringtest_0.ring_out.n1 ringtest_0.ring_out.t1 26.5955
R14497 ringtest_0.ring_out.n2 ringtest_0.ring_out.t7 26.5955
R14498 ringtest_0.ring_out.n2 ringtest_0.ring_out.t8 26.5955
R14499 ringtest_0.ring_out.n11 ringtest_0.ring_out.t5 26.3998
R14500 ringtest_0.ring_out ringtest_0.ring_out.n3 24.9955
R14501 ringtest_0.ring_out.n4 ringtest_0.ring_out.t9 24.9236
R14502 ringtest_0.ring_out.n4 ringtest_0.ring_out.t0 24.9236
R14503 ringtest_0.ring_out.n11 ringtest_0.ring_out.t6 23.5483
R14504 ringtest_0.ring_out.n10 ringtest_0.ring_out.n9 21.363
R14505 ringtest_0.ring_out ringtest_0.ring_out.n5 14.8576
R14506 ringtest_0.ring_out.n12 ringtest_0.ring_out.t4 12.9758
R14507 ringtest_0.ring_out.n6 ringtest_0.ring_out 10.9719
R14508 ringtest_0.ring_out.n12 ringtest_0.ring_out.t3 10.8618
R14509 ringtest_0.ring_out.n10 ringtest_0.ring_out.n6 9.53262
R14510 ringtest_0.ring_out.n6 ringtest_0.ring_out 4.57193
R14511 ringtest_0.ring_out.n13 ringtest_0.ring_out.n11 3.06895
R14512 ringtest_0.ring_out.n9 ringtest_0.ring_out 2.32777
R14513 ringtest_0.ring_out.n13 ringtest_0.ring_out.n12 2.14822
R14514 ringtest_0.ring_out ringtest_0.ring_out.n13 1.12636
R14515 ringtest_0.ring_out.n5 ringtest_0.ring_out 0.686214
R14516 ringtest_0.ring_out ringtest_0.ring_out.n10 0.631142
R14517 ringtest_0.ring_out ringtest_0.ring_out.n0 0.354518
R14518 ringtest_0.x3.x2.GP2.n2 ringtest_0.x3.x2.GP2.t4 450.938
R14519 ringtest_0.x3.x2.GP2.n2 ringtest_0.x3.x2.GP2.t5 445.666
R14520 ringtest_0.x3.x2.GP2.n4 ringtest_0.x3.x2.GP2.n3 195.958
R14521 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n0 96.8352
R14522 ringtest_0.x3.x2.GP2.n3 ringtest_0.x3.x2.GP2.t3 26.5955
R14523 ringtest_0.x3.x2.GP2.n3 ringtest_0.x3.x2.GP2.t2 26.5955
R14524 ringtest_0.x3.x2.GP2.n0 ringtest_0.x3.x2.GP2.t1 24.9236
R14525 ringtest_0.x3.x2.GP2.n0 ringtest_0.x3.x2.GP2.t0 24.9236
R14526 ringtest_0.x3.x2.GP2.n5 ringtest_0.x3.x2.GP2.n4 13.0077
R14527 ringtest_0.x3.x2.GP2.n4 ringtest_0.x3.x2.GP2 11.995
R14528 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n1 11.2645
R14529 ringtest_0.x3.x2.GP2.n1 ringtest_0.x3.x2.GP2 6.1445
R14530 ringtest_0.x3.x2.GP2.n1 ringtest_0.x3.x2.GP2 4.65505
R14531 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n2 3.12839
R14532 ringtest_0.x3.x2.GP2.n5 ringtest_0.x3.x2.GP2 2.0485
R14533 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n5 1.55202
R14534 muxtest_0.x2.x2.GP4.n2 muxtest_0.x2.x2.GP4.t4 450.938
R14535 muxtest_0.x2.x2.GP4.n2 muxtest_0.x2.x2.GP4.t5 445.666
R14536 muxtest_0.x2.x2.GP4.n5 muxtest_0.x2.x2.GP4.n4 208.965
R14537 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n0 96.8352
R14538 muxtest_0.x2.x2.GP4.n4 muxtest_0.x2.x2.GP4.t3 26.5955
R14539 muxtest_0.x2.x2.GP4.n4 muxtest_0.x2.x2.GP4.t2 26.5955
R14540 muxtest_0.x2.x2.GP4.n0 muxtest_0.x2.x2.GP4.t1 24.9236
R14541 muxtest_0.x2.x2.GP4.n0 muxtest_0.x2.x2.GP4.t0 24.9236
R14542 muxtest_0.x2.x1.gpo3 muxtest_0.x2.x2.x4.GP 16.5032
R14543 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n3 10.2405
R14544 muxtest_0.x2.x2.GP4.n3 muxtest_0.x2.x1.gpo3 7.76481
R14545 muxtest_0.x2.x2.GP4.n1 muxtest_0.x2.x1.x14.Y 6.1445
R14546 muxtest_0.x2.x2.GP4.n1 muxtest_0.x2.x1.x14.Y 4.65505
R14547 muxtest_0.x2.x2.x4.GP muxtest_0.x2.x2.GP4.n2 2.95993
R14548 muxtest_0.x2.x2.GP4.n5 muxtest_0.x2.x1.x14.Y 2.0485
R14549 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n5 1.55202
R14550 muxtest_0.x2.x2.GP4.n3 muxtest_0.x2.x2.GP4.n1 1.0245
R14551 muxtest_0.R4R5.n0 muxtest_0.R4R5.t1 26.3998
R14552 muxtest_0.R4R5.n0 muxtest_0.R4R5.t2 23.5483
R14553 muxtest_0.R4R5.n1 muxtest_0.R4R5.t5 12.9758
R14554 muxtest_0.R4R5.n1 muxtest_0.R4R5.t4 10.8618
R14555 muxtest_0.R4R5.n4 muxtest_0.R4R5.t0 10.8231
R14556 muxtest_0.R4R5.n4 muxtest_0.R4R5.t3 10.5739
R14557 muxtest_0.R4R5.n2 muxtest_0.R4R5.n0 3.06895
R14558 muxtest_0.R4R5.n2 muxtest_0.R4R5.n1 2.14822
R14559 muxtest_0.R4R5.n3 muxtest_0.R4R5.n2 1.12636
R14560 muxtest_0.R4R5 muxtest_0.R4R5.n4 0.790021
R14561 muxtest_0.R4R5 muxtest_0.R4R5.n3 0.134513
R14562 muxtest_0.R4R5.n3 muxtest_0.R4R5 0.0655
R14563 muxtest_0.R2R3.n0 muxtest_0.R2R3.t0 26.3998
R14564 muxtest_0.R2R3.n0 muxtest_0.R2R3.t1 23.5483
R14565 muxtest_0.R2R3.n1 muxtest_0.R2R3.t3 12.9758
R14566 muxtest_0.R2R3.n1 muxtest_0.R2R3.t2 10.8618
R14567 muxtest_0.R2R3.n4 muxtest_0.R2R3.t4 10.8167
R14568 muxtest_0.R2R3.n4 muxtest_0.R2R3.t5 10.5739
R14569 muxtest_0.R2R3.n2 muxtest_0.R2R3.n0 3.06895
R14570 muxtest_0.R2R3.n2 muxtest_0.R2R3.n1 2.14822
R14571 muxtest_0.R2R3.n3 muxtest_0.R2R3.n2 1.12636
R14572 muxtest_0.R2R3 muxtest_0.R2R3.n4 0.71627
R14573 muxtest_0.R2R3 muxtest_0.R2R3.n3 0.138152
R14574 muxtest_0.R2R3.n3 muxtest_0.R2R3 0.0655
R14575 ui_in[6].n0 ui_in[6].t0 212.081
R14576 ui_in[6].n1 ui_in[6].t1 212.081
R14577 ui_in[6] ui_in[6].n2 152.512
R14578 ui_in[6].n0 ui_in[6].t2 139.78
R14579 ui_in[6].n1 ui_in[6].t3 139.78
R14580 ui_in[6].n2 ui_in[6].n0 30.6732
R14581 ui_in[6].n2 ui_in[6].n1 30.6732
R14582 ui_in[6].n3 ui_in[6] 16.4378
R14583 ui_in[6] ui_in[6].n3 0.7505
R14584 ui_in[6].n3 ui_in[6] 0.0808571
R14585 ui_in[5].n0 ui_in[5].t0 260.322
R14586 ui_in[5].n0 ui_in[5].t1 175.169
R14587 ui_in[5].n1 ui_in[5].n0 153.13
R14588 ui_in[5].n3 ui_in[5] 19.5879
R14589 ui_in[5] ui_in[5].n1 9.86591
R14590 ui_in[5].n3 ui_in[5].n2 4.07076
R14591 ui_in[5].n1 ui_in[5] 3.2005
R14592 ui_in[5].n2 ui_in[5] 0.960321
R14593 ui_in[5].n2 ui_in[5] 0.392836
R14594 ui_in[5] ui_in[5].n3 0.0499792
C0 muxtest_0.R7R8 muxtest_0.x2.x2.GN3 0.01204f
C1 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GP3 2.78e-20
C2 a_22392_5990# ringtest_0.x4._16_ 1.01e-19
C3 ringtest_0.ring_out ui_in[6] 0.550306f
C4 ringtest_0.x4._11_ ringtest_0.counter3 1.13e-19
C5 muxtest_0.x1.x4.A a_12849_23648# 1.34e-19
C6 uio_in[1] uio_in[0] 0.033505f
C7 ringtest_0.x4.clknet_1_1__leaf_clk a_24800_5334# 0.033626f
C8 ringtest_0.x4.clknet_0_clk a_23619_6788# 9.48e-20
C9 ringtest_0.x4._13_ a_21951_5878# 7.99e-20
C10 muxtest_0.x2.x1.nSEL1 VDPWR 0.649185f
C11 a_21981_8976# ringtest_0.x4._01_ 0.00226f
C12 ringtest_0.x4.net3 a_22399_8976# 4.27e-20
C13 ringtest_0.x4.clknet_1_0__leaf_clk a_21591_6128# 0.001585f
C14 ringtest_0.x4._00_ ringtest_0.x4._11_ 0.003231f
C15 a_26627_4246# a_26817_4566# 0.011458f
C16 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A 0.429373f
C17 a_27065_5156# a_27303_4246# 3.93e-20
C18 a_13025_23980# ui_in[3] 0.279858f
C19 ringtest_0.x4.net1 a_21780_8964# 1.42e-19
C20 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A 5.04e-19
C21 ringtest_0.x4.net7 a_26007_6788# 0.003849f
C22 a_24527_5340# a_25225_5334# 0.192206f
C23 a_21840_5308# a_21587_5334# 3.39e-19
C24 a_21399_5340# a_21798_5712# 8.12e-19
C25 a_24968_5308# a_25393_5308# 1.28e-19
C26 a_24361_5340# a_26201_5340# 0.002059f
C27 a_21948_5156# ringtest_0.x4.counter[2] 1.99e-20
C28 a_19114_31955# muxtest_0.x1.x3.GN2 0.106131f
C29 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._23_ 0.071442f
C30 ringtest_0.x4._11_ ringtest_0.x4.net10 0.36244f
C31 ringtest_0.x4.clknet_1_1__leaf_clk a_26367_4790# 0.031849f
C32 a_24336_6544# ringtest_0.x4._19_ 0.457296f
C33 VDPWR ua[0] 3.15952f
C34 a_12849_23648# muxtest_0.x2.x2.GP2 3.07e-19
C35 ringtest_0.x4.clknet_0_clk a_25225_5334# 0.013741f
C36 muxtest_0.x1.x3.GP3 ui_in[0] 2.74e-19
C37 ringtest_0.x4._15_ ringtest_0.x4.net5 0.016962f
C38 ringtest_0.x4._03_ a_22765_4478# 1.19e-19
C39 ringtest_0.x4.net4 a_22983_5654# 5.3e-19
C40 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2 2.14737f
C41 ringtest_0.drv_out VDPWR 16.4224f
C42 muxtest_0.x2.nselect2 ui_in[4] 0.001201f
C43 a_17231_12017# ui_in[4] 0.125445f
C44 ringtest_0.x4._11_ a_22775_5878# 8.02e-19
C45 ringtest_0.x4._24_ a_27065_5334# 0.013075f
C46 a_15575_12017# a_15749_12123# 0.006584f
C47 ringtest_0.x3.x1.nSEL1 a_16155_12151# 9.57e-19
C48 ringtest_0.x4._11_ a_24627_6200# 4.38e-19
C49 a_22541_5058# ringtest_0.x4.net5 0.13266f
C50 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN1 0.034862f
C51 ringtest_0.x4._08_ ringtest_0.x4._07_ 9.41e-21
C52 muxtest_0.R3R4 ua[3] 0.039417f
C53 ringtest_0.x4._11_ ringtest_0.x4.counter[4] 6.77e-20
C54 ringtest_0.x4._18_ a_23993_5654# 6.01e-19
C55 a_13675_24012# VDPWR 8.97e-19
C56 ringtest_0.x4.net8 a_26895_3867# 7.5e-19
C57 a_22392_5990# a_22649_6244# 0.036838f
C58 muxtest_0.x2.x2.GN3 VDPWR 0.650589f
C59 a_21951_5878# ringtest_0.x4.net8 0.001542f
C60 a_23879_6940# a_24715_5334# 2.19e-20
C61 ringtest_0.x4.net9 a_25977_4220# 9.8e-19
C62 a_22052_8875# ringtest_0.x4._10_ 2.11e-19
C63 a_23949_6654# a_23770_5308# 8.51e-20
C64 ringtest_0.x4._01_ a_22228_8598# 5.75e-19
C65 muxtest_0.x1.x3.GN4 muxtest_0.R2R3 0.127088f
C66 ringtest_0.x4.net9 a_25719_4790# 0.001933f
C67 muxtest_0.x1.x3.GN4 ui_in[1] 0.059771f
C68 a_24329_6640# ringtest_0.x4._16_ 1.49e-19
C69 ringtest_0.x4.net4 a_22486_4246# 0.003167f
C70 ringtest_0.x4._07_ a_25336_4902# 0.004454f
C71 a_24336_6544# ringtest_0.x4.net9 1.52e-20
C72 ringtest_0.x4._22_ a_25168_5156# 0.002895f
C73 ringtest_0.x3.x2.GP2 ui_in[3] 5.28e-19
C74 ringtest_0.x4._24_ a_26627_4246# 0.085832f
C75 muxtest_0.R3R4 m3_13316_18955# 1.46e-19
C76 ringtest_0.x4.net7 a_25977_4220# 0.023542f
C77 ringtest_0.x4._00_ a_22399_9142# 0.139872f
C78 ringtest_0.x4._18_ ringtest_0.x4._04_ 0.003255f
C79 ringtest_0.x4._24_ a_27149_5156# 8.56e-19
C80 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN4 9.02e-19
C81 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN3 0.012418f
C82 ringtest_0.x4._23_ a_26367_4790# 0.031117f
C83 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN2 0.154394f
C84 ringtest_0.x4._07_ VDPWR 0.322336f
C85 a_24336_6544# ringtest_0.x4.net7 0.027472f
C86 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.001676f
C87 ringtest_0.x4._06_ a_24361_5340# 0.091082f
C88 ringtest_0.x4.clknet_1_1__leaf_clk a_25593_5156# 0.044904f
C89 ringtest_0.x4.net8 a_26808_5308# 8.61e-20
C90 ringtest_0.x4._16_ a_24545_5878# 0.036674f
C91 ringtest_0.x4._11_ a_25393_5308# 1.18e-19
C92 ringtest_0.x4._17_ a_24336_6544# 0.050404f
C93 a_25055_3867# VDPWR 0.315151f
C94 a_16155_12151# ringtest_0.x3.x2.GN3 5.17e-20
C95 ringtest_0.x3.x2.GN2 a_16707_12151# 3.11e-20
C96 ringtest_0.x4.net2 ringtest_0.x4._03_ 5.34e-20
C97 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN3 0.002857f
C98 ringtest_0.x4._08_ a_26201_5340# 0.097891f
C99 muxtest_0.x2.x1.nSEL1 a_12849_23648# 7.84e-19
C100 a_25364_5878# ringtest_0.x4._16_ 0.001016f
C101 a_24264_6788# VDPWR 7.65e-20
C102 muxtest_0.x2.x1.nSEL0 ua[3] 7.05e-20
C103 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ui_in[6] 0.108977f
C104 ringtest_0.x4.net6 a_26367_5340# 1.27e-19
C105 ringtest_0.x4._03_ a_23381_4818# 2.2e-20
C106 ringtest_0.x4._15_ a_24527_5340# 0.027322f
C107 a_21509_4790# a_23809_4790# 1.62e-21
C108 a_21845_8816# a_21395_6940# 6.92e-20
C109 a_25225_5334# a_25168_5156# 7.26e-19
C110 a_27273_4220# a_27489_3702# 1.29e-21
C111 a_26817_4566# a_26721_4246# 1.26e-19
C112 muxtest_0.x1.x4.A muxtest_0.x1.x5.A 2.05508f
C113 ringtest_0.x4.clknet_0_clk ringtest_0.x4._15_ 4.05e-19
C114 a_16203_12091# VDPWR 0.192568f
C115 muxtest_0.x1.x3.GP1 muxtest_0.R7R8 4.13739f
C116 a_21561_8830# ringtest_0.x4._12_ 0.036321f
C117 ringtest_0.x4.net8 a_23381_4584# 9.57e-20
C118 ringtest_0.x4._11_ a_27191_4790# 9.67e-22
C119 ringtest_0.x4.net9 a_25677_5156# 8.89e-19
C120 ringtest_0.x4.net11 a_26895_3867# 3.2e-20
C121 ringtest_0.x4._11_ a_26808_4902# 8.51e-19
C122 ringtest_0.x4.counter[1] ua[1] 3.21e-19
C123 ringtest_0.x4._16_ a_24317_4942# 1.3e-19
C124 a_16707_12151# ui_in[3] 0.001558f
C125 a_24045_6654# ringtest_0.x4.net8 1.55e-19
C126 ringtest_0.x3.x2.GN2 ui_in[3] 0.114345f
C127 a_27233_5308# a_27065_5334# 0.310858f
C128 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._04_ 1.67e-21
C129 a_22265_5308# a_23899_5334# 2.67e-21
C130 a_22765_5308# a_22795_5334# 0.025037f
C131 a_24968_5308# a_24715_5334# 3.39e-19
C132 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A 0.159172f
C133 a_26201_5340# VDPWR 0.714632f
C134 ringtest_0.x4._05_ a_24883_6800# 0.114695f
C135 a_24465_6800# a_24287_6422# 9.73e-19
C136 ringtest_0.x4.net6 a_22765_4478# 5.34e-20
C137 ringtest_0.x4._16_ a_23151_5334# 0.010038f
C138 ringtest_0.x4._18_ ringtest_0.x4.net4 3.06e-19
C139 ringtest_0.counter7 ringtest_0.x4.net4 6.88e-20
C140 ringtest_0.drv_out a_23879_6940# 0.318051f
C141 ringtest_0.x4.net7 a_25677_5156# 0.002598f
C142 ringtest_0.x4._23_ a_25593_5156# 0.001187f
C143 a_25593_5156# a_26367_4790# 2.56e-19
C144 a_24729_4790# a_26555_4790# 4.76e-21
C145 a_23949_6654# ringtest_0.x4.net6 1.76e-19
C146 ringtest_0.x4.counter[5] VDPWR 0.450193f
C147 a_12849_23648# muxtest_0.x2.x2.GN3 0.104151f
C148 a_13025_23980# muxtest_0.x2.x2.GN1 3.78e-20
C149 ringtest_0.x4._21_ ringtest_0.x4._07_ 4.77e-20
C150 a_22224_6244# ringtest_0.x4._14_ 5.19e-22
C151 ringtest_0.x4.net7 a_23899_5334# 0.006434f
C152 ringtest_0.x4.net9 ringtest_0.x4.counter[9] 5.19e-19
C153 a_26749_6422# a_26808_5308# 2.48e-20
C154 ringtest_0.x4._25_ a_26201_5340# 1.01e-19
C155 m2_15612_11606# ui_in[3] 0.130999f
C156 ringtest_0.x3.nselect2 a_16579_11759# 1.29e-19
C157 a_22164_4362# VDPWR 0.108977f
C158 ringtest_0.counter3 ringtest_0.x4.counter[4] 0.07836f
C159 ringtest_0.x4.net8 ringtest_0.x4.counter[6] 0.079257f
C160 ringtest_0.x4.net8 a_24699_6200# 0.003186f
C161 ringtest_0.x4._17_ a_23899_5334# 9.12e-21
C162 a_27233_5058# VDPWR 0.462064f
C163 a_22224_6244# a_22319_6244# 0.007724f
C164 a_22392_5990# a_22733_6244# 9.73e-19
C165 ringtest_0.counter3 a_23399_3867# 0.110188f
C166 a_23529_6422# VDPWR 0.185924f
C167 ringtest_0.x4.net4 a_22295_3867# 0.202764f
C168 ringtest_0.x4._12_ a_21049_8598# 0.090947f
C169 muxtest_0.x1.x3.GP1 muxtest_0.R5R6 0.122287f
C170 ringtest_0.x4._19_ ringtest_0.x4._16_ 0.001191f
C171 a_23770_5308# ringtest_0.x4._20_ 3.36e-20
C172 ringtest_0.x4._18_ a_23837_5878# 0.002103f
C173 ringtest_0.x4.net6 a_24004_6128# 0.074355f
C174 ringtest_0.counter7 ringtest_0.x4._22_ 1.31e-20
C175 a_21672_5334# a_21509_4790# 4.57e-19
C176 a_21233_5340# a_21948_5156# 0.001041f
C177 a_21840_5308# ringtest_0.x4._03_ 0.009555f
C178 a_25977_4220# a_26627_4246# 0.010893f
C179 a_22765_4478# a_22939_4584# 0.006584f
C180 a_22021_4220# a_22486_4246# 0.005941f
C181 ringtest_0.x4.net8 a_24479_4790# 0.002158f
C182 ringtest_0.x4._11_ a_25083_4790# 0.016192f
C183 muxtest_0.x1.x3.GP1 VDPWR 3.2848f
C184 a_21465_9294# ringtest_0.x4.net3 9.98e-20
C185 a_24699_6200# a_24729_4790# 5.07e-21
C186 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN3 0.08518f
C187 ringtest_0.x4.net9 a_27149_5334# 1.06e-19
C188 a_21465_9294# a_21845_9116# 0.048748f
C189 a_21561_9116# a_21852_9416# 0.194892f
C190 ringtest_0.counter7 a_24135_3867# 2.81e-20
C191 ringtest_0.x4.net8 a_23809_4790# 7.44e-19
C192 a_20318_32213# VDPWR 0.217349f
C193 ringtest_0.x4._11_ a_21948_5156# 0.00274f
C194 a_22265_5308# a_22097_5334# 0.310858f
C195 ringtest_0.ring_out ui_in[4] 0.016625f
C196 muxtest_0.x1.x1.nSEL0 a_19666_31955# 1.91e-20
C197 ringtest_0.x4._16_ a_22265_5308# 7.03e-19
C198 ringtest_0.x4._06_ VDPWR 0.276236f
C199 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.025028f
C200 a_24336_6544# a_24536_6699# 0.074815f
C201 a_24329_6640# a_24465_6800# 0.136009f
C202 a_24045_6654# ringtest_0.x4._05_ 9.72e-20
C203 a_24070_5852# VDPWR 0.084816f
C204 a_25168_5156# a_25263_5156# 0.007724f
C205 a_21395_6940# a_21399_5340# 1.82e-21
C206 ringtest_0.x4.net6 a_23381_4818# 4.93e-21
C207 ringtest_0.x4.net9 ringtest_0.x4._16_ 0.243936f
C208 a_24763_6143# ringtest_0.x4._22_ 0.155189f
C209 a_21845_8816# VDPWR 0.446206f
C210 ringtest_0.x4._04_ ringtest_0.x4._02_ 1.6e-19
C211 a_23809_4790# a_24729_4790# 2.37e-21
C212 ringtest_0.x4._15_ a_22983_5654# 1.54e-19
C213 ringtest_0.x4.net2 a_21055_5334# 0.002977f
C214 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._02_ 0.254839f
C215 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ui_in[6] 6.29e-19
C216 a_21675_4790# a_21948_5156# 0.081834f
C217 a_23399_3867# ringtest_0.x4.counter[4] 0.001146f
C218 a_26640_5334# a_26201_4790# 1.73e-19
C219 a_23891_4790# VDPWR 2.86e-19
C220 ringtest_0.x4.net7 ringtest_0.x4._16_ 5.07e-19
C221 a_22164_4362# ringtest_0.x4.counter[2] 6.46e-19
C222 a_24465_6800# a_24545_5878# 1.71e-20
C223 a_22373_5156# VDPWR 0.183311f
C224 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._22_ 0.031888f
C225 ringtest_0.x3.x1.nSEL0 VDPWR 0.5228f
C226 ringtest_0.x4.net3 a_21981_8976# 2.06e-19
C227 a_26640_5334# a_26555_5334# 0.037333f
C228 a_26808_5308# a_26766_5712# 4.62e-19
C229 ringtest_0.x4._17_ ringtest_0.x4._16_ 0.048058f
C230 a_21845_9116# a_21981_8976# 5.28e-20
C231 a_21852_9416# ringtest_0.x4._01_ 8.68e-20
C232 a_22052_9116# a_22052_8875# 0.013851f
C233 ringtest_0.drv_out a_25925_6788# 1.34e-19
C234 ringtest_0.x4._05_ a_24699_6200# 3.16e-19
C235 muxtest_0.x2.x1.nSEL1 m2_11882_23495# 0.00815f
C236 ringtest_0.x3.x2.GN4 ringtest_0.counter3 0.237196f
C237 a_21767_5334# VDPWR 0.003619f
C238 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP2 0.068989f
C239 ringtest_0.x4.net1 a_21845_8816# 0.002755f
C240 ringtest_0.ring_out ringtest_0.x3.x2.GP1 4.09516f
C241 ringtest_0.x4.net2 a_21981_9142# 3.46e-19
C242 a_12977_24040# muxtest_0.x2.x2.GP3 4.39e-19
C243 a_22224_6244# a_21509_4790# 5.5e-20
C244 ringtest_0.x4._09_ a_26555_4790# 0.129132f
C245 a_26201_4790# a_26735_5156# 0.002698f
C246 a_21785_5878# a_21948_5156# 8.98e-19
C247 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP3 0.004298f
C248 ringtest_0.x4._07_ a_24968_5308# 0.011124f
C249 ringtest_0.x4._22_ a_24800_5334# 0.006172f
C250 ringtest_0.x4.net5 a_22765_4478# 0.081136f
C251 ringtest_0.x4.clknet_1_0__leaf_clk a_22116_4902# 0.001507f
C252 ringtest_0.x4.net6 ringtest_0.x4._20_ 0.00624f
C253 muxtest_0.x2.nselect2 muxtest_0.x2.x2.GN4 1.53e-20
C254 a_23349_6422# a_23529_6422# 0.185422f
C255 a_22201_8964# VDPWR 0.002269f
C256 ringtest_0.x4._20_ a_24895_4790# 0.003428f
C257 a_26269_4612# VDPWR 0.001259f
C258 ringtest_0.x4.net10 a_26808_4902# 1.26e-19
C259 a_13025_23980# ua[3] 9.59e-19
C260 ringtest_0.x4._21_ ringtest_0.x4._06_ 0.224771f
C261 ringtest_0.counter7 ua[3] 1.17e-19
C262 ringtest_0.x4.net4 ringtest_0.x4._02_ 1.19e-19
C263 a_22817_6146# ringtest_0.x4._16_ 0.001048f
C264 ringtest_0.x3.x1.nSEL1 ui_in[4] 0.272823f
C265 a_24070_5852# ringtest_0.x4._21_ 0.114705f
C266 a_22139_5878# a_22319_6244# 0.001229f
C267 a_27489_3702# ringtest_0.x4.counter[8] 0.006251f
C268 a_24004_6128# a_23932_6128# 0.005941f
C269 muxtest_0.x1.x4.A a_13501_23906# 0.001685f
C270 a_21395_6940# a_21951_5878# 1.63e-19
C271 ringtest_0.x4.clknet_1_1__leaf_clk a_25225_5334# 0.024694f
C272 ringtest_0.x4.net6 a_21840_5308# 6.4e-20
C273 ringtest_0.drv_out ringtest_0.x4._11_ 1.2e-19
C274 ringtest_0.x4.clknet_0_clk a_24685_6788# 4.62e-19
C275 ringtest_0.x4._23_ ringtest_0.x4._22_ 0.511385f
C276 ringtest_0.x4._13_ a_22224_6244# 5.02e-20
C277 a_22499_4790# VDPWR 4.65e-19
C278 ringtest_0.x4._22_ a_26367_4790# 3.15e-20
C279 a_27065_5334# a_27149_5334# 0.008508f
C280 ringtest_0.x4._24_ ringtest_0.x4.net8 1.23e-20
C281 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._04_ 0.005301f
C282 a_22021_4220# a_22295_3867# 4.71e-19
C283 a_25364_5878# a_26201_4790# 6.92e-20
C284 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A 0.429199f
C285 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 5.02073f
C286 muxtest_0.x2.x2.GN1 ui_in[3] 0.021261f
C287 a_23879_6940# ringtest_0.x4._06_ 1.96e-20
C288 ringtest_0.x4.net7 a_26201_6788# 5.71e-19
C289 ringtest_0.x4._17_ a_22649_6244# 1.03e-20
C290 a_23879_6940# a_24070_5852# 3.15e-19
C291 a_21672_5334# a_21798_5712# 0.005525f
C292 a_24527_5340# a_26367_5340# 0.001861f
C293 a_19666_31955# muxtest_0.x1.x3.GN2 1.61e-19
C294 ringtest_0.x4.net6 a_26569_6422# 2.84e-19
C295 ringtest_0.x4._17_ a_26201_6788# 3.01e-19
C296 a_21399_5340# VDPWR 0.341027f
C297 a_25364_5878# a_26555_5334# 9.53e-19
C298 muxtest_0.x1.x1.nSEL1 a_18662_32213# 0.193944f
C299 ringtest_0.x4.net4 a_22116_4902# 0.007782f
C300 ringtest_0.x4.clknet_1_1__leaf_clk a_26640_5156# 3.02e-19
C301 ringtest_0.x4._05_ a_25421_6641# 0.121098f
C302 muxtest_0.x2.x2.GP2 ua[2] 0.349855f
C303 a_24465_6800# ringtest_0.x4._19_ 0.040707f
C304 ringtest_0.x4._18_ ringtest_0.x4._15_ 0.045245f
C305 ringtest_0.counter7 ringtest_0.x4._15_ 0.003538f
C306 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.001676f
C307 a_24968_5308# ringtest_0.x4.counter[5] 2.7e-21
C308 ringtest_0.x4.net2 ringtest_0.x4.net5 7.09e-21
C309 muxtest_0.x1.x3.GN4 ui_in[0] 0.218694f
C310 muxtest_0.x1.x1.nSEL1 m2_18699_31802# 0.00815f
C311 ringtest_0.x4.net5 a_23963_4790# 1.04e-20
C312 a_17405_12123# ui_in[4] 8.84e-19
C313 ringtest_0.x4._15_ a_27191_5712# 6.51e-20
C314 ringtest_0.x3.x2.GN3 ui_in[4] 0.273713f
C315 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GP1 1.21e-19
C316 ringtest_0.x4._11_ ringtest_0.x4._07_ 0.161717f
C317 a_16027_11759# ringtest_0.x3.x2.GN2 0.106178f
C318 a_21863_4790# a_22043_5156# 0.001229f
C319 a_23381_4818# ringtest_0.x4.net5 4.5e-19
C320 muxtest_0.x1.x3.GN3 muxtest_0.R1R2 4.03753f
C321 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ui_in[6] 3.49e-19
C322 muxtest_0.R7R8 muxtest_0.R4R5 0.286971f
C323 a_22817_6146# a_22649_6244# 0.310858f
C324 a_22224_6244# ringtest_0.x4.net8 4.11e-20
C325 uio_in[6] uio_in[5] 0.031023f
C326 ringtest_0.x4.net9 a_27273_4220# 0.001158f
C327 ringtest_0.x4._01_ ringtest_0.x4._10_ 0.002197f
C328 a_24045_6654# a_24361_5340# 1.16e-21
C329 ringtest_0.x4.net4 ringtest_0.x4._04_ 0.689049f
C330 ringtest_0.x4.net9 a_26766_4790# 0.002793f
C331 ringtest_0.x4._15_ a_24763_6143# 1.57e-19
C332 muxtest_0.x1.x3.GN1 muxtest_0.R3R4 3.99705f
C333 a_24536_6699# ringtest_0.x4._16_ 1.35e-21
C334 ringtest_0.x4._07_ a_25761_5058# 3.3e-20
C335 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR 0.639695f
C336 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP3 0.09552f
C337 a_24465_6800# ringtest_0.x4.net9 0.004659f
C338 ringtest_0.x4._22_ a_25593_5156# 6.29e-19
C339 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net4 0.158995f
C340 ringtest_0.x4.clknet_0_clk a_23949_6654# 0.002548f
C341 ringtest_0.x4.net6 a_22392_5990# 3.85e-19
C342 ringtest_0.x4.net2 a_21007_3867# 0.223155f
C343 ringtest_0.x4._24_ a_26749_6422# 0.197975f
C344 ringtest_0.x4._24_ ringtest_0.x4.net11 0.002712f
C345 a_16027_11759# ui_in[3] 0.246189f
C346 ringtest_0.x4.net6 a_24287_6422# 1.73e-19
C347 ringtest_0.x4._23_ a_26640_5156# 0.011058f
C348 a_26808_4902# a_27191_4790# 4.67e-20
C349 ringtest_0.x4._05_ ringtest_0.x4._24_ 2.08e-20
C350 a_26367_4790# a_26640_5156# 0.078545f
C351 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._15_ 0.471647f
C352 ringtest_0.x4._14_ a_22097_5334# 2.97e-21
C353 a_24465_6800# ringtest_0.x4.net7 0.035198f
C354 ringtest_0.x4.clknet_1_1__leaf_clk a_25263_5156# 0.001835f
C355 ringtest_0.x4._06_ a_24968_5308# 0.001008f
C356 ringtest_0.x4._16_ ringtest_0.x4._14_ 0.202586f
C357 ringtest_0.x4.net8 a_27233_5308# 4.93e-20
C358 ringtest_0.x4._11_ a_26201_5340# 3.54e-20
C359 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP1 0.001426f
C360 a_24699_6200# a_24361_5340# 0.001396f
C361 ringtest_0.x4._17_ a_24465_6800# 0.016441f
C362 a_26895_3867# VDPWR 0.303091f
C363 a_21951_5878# VDPWR 0.304738f
C364 ringtest_0.x4._08_ a_26808_5308# 0.047112f
C365 ringtest_0.x4.net5 ringtest_0.x4._20_ 8.42e-21
C366 a_24883_6800# VDPWR 0.085296f
C367 muxtest_0.x1.x3.GP2 muxtest_0.R1R2 0.153531f
C368 ringtest_0.x4.clknet_0_clk a_24004_6128# 2.03e-19
C369 a_21509_4790# a_21863_4790# 0.062224f
C370 ringtest_0.x4._15_ a_24800_5334# 0.026278f
C371 muxtest_0.R5R6 muxtest_0.R4R5 2.29244f
C372 ringtest_0.x4._22_ a_25441_4612# 0.002353f
C373 a_21785_8054# ringtest_0.x4._10_ 0.107891f
C374 ringtest_0.x4._13_ a_22139_5878# 5.97e-20
C375 a_22052_8875# a_21395_6940# 2.84e-19
C376 VDPWR ua[1] 17.382101f
C377 ringtest_0.drv_out ringtest_0.counter3 1.91048f
C378 a_25225_5334# a_25593_5156# 3.78e-19
C379 a_26555_5334# a_26735_5334# 0.001229f
C380 a_16755_12091# VDPWR 0.26222f
C381 a_22224_6244# a_22390_4566# 4.44e-21
C382 ringtest_0.x4.net8 a_25977_4220# 0.004343f
C383 a_21852_8720# ringtest_0.x4._12_ 0.206007f
C384 ringtest_0.x4._11_ a_22164_4362# 1e-19
C385 muxtest_0.x1.x3.GP1 muxtest_0.x1.x5.A 0.353808f
C386 muxtest_0.R4R5 VDPWR 1.56678f
C387 ringtest_0.x4.net9 a_26201_4790# 0.11266f
C388 ringtest_0.x4.net11 a_27815_3867# 0.003661f
C389 ringtest_0.x4.net8 a_25719_4790# 5.67e-20
C390 ringtest_0.x4._11_ a_27233_5058# 5.38e-21
C391 ua[0] ua[2] 4.5205f
C392 a_24336_6544# ringtest_0.x4.net8 4.93e-19
C393 ringtest_0.x4.net2 ringtest_0.x4._12_ 0.10227f
C394 a_24800_5334# a_24926_5712# 0.005525f
C395 ringtest_0.x4._11_ a_23529_6422# 0.001495f
C396 a_19114_31955# muxtest_0.x1.x3.GP1 9.8e-19
C397 a_26808_5308# VDPWR 0.182123f
C398 ua[3] ui_in[3] 0.553118f
C399 ringtest_0.x4._15_ ringtest_0.x4._23_ 0.683594f
C400 a_24329_6640# a_24712_6422# 0.001632f
C401 ringtest_0.x4.net6 a_25149_4220# 0.211407f
C402 ringtest_0.x4._24_ ringtest_0.x4._09_ 0.151845f
C403 a_18662_32213# muxtest_0.x1.x3.GN1 0.128677f
C404 ringtest_0.x4._15_ a_26367_4790# 0.036316f
C405 muxtest_0.R7R8 ui_in[2] 0.054741f
C406 a_24895_4790# a_25149_4220# 0.002313f
C407 ringtest_0.x4.net7 a_26201_4790# 0.007864f
C408 a_24329_6640# ringtest_0.x4.net6 0.001597f
C409 a_13501_23906# a_13675_24012# 0.006584f
C410 muxtest_0.x1.x3.GN1 m2_18699_31802# 0.06935f
C411 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.025028f
C412 a_13501_23906# muxtest_0.x2.x2.GN3 1.07e-20
C413 muxtest_0.x2.x2.GN1 a_12425_24040# 1.22e-20
C414 a_12019_24012# muxtest_0.x2.x2.GN2 8.86e-19
C415 a_22116_4902# a_22021_4220# 1.66e-20
C416 muxtest_0.x2.x2.GN3 ua[2] 0.429994f
C417 a_21675_4790# a_22164_4362# 0.010312f
C418 a_24329_6640# a_24895_4790# 4.79e-20
C419 ringtest_0.x4._24_ a_26766_5712# 9.29e-19
C420 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP2 1.19e-20
C421 a_27065_5334# a_27273_4220# 9.49e-21
C422 ringtest_0.x4.net8 a_24986_5878# 1.76e-19
C423 ringtest_0.x3.nselect2 a_17231_12017# 9.77e-20
C424 a_23381_4584# VDPWR 0.2419f
C425 a_27233_5308# ringtest_0.x4.net11 1.16e-19
C426 ringtest_0.x4._11_ ringtest_0.x4._06_ 0.020042f
C427 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GN4 3.13e-20
C428 a_21675_9686# VDPWR 0.262851f
C429 a_22224_6244# a_22350_5878# 0.005525f
C430 a_21785_8054# a_21867_8054# 0.005167f
C431 a_21951_5878# ringtest_0.x4._21_ 2.75e-21
C432 a_26555_4790# VDPWR 0.079695f
C433 ringtest_0.x4.net9 a_27303_4246# 0.005829f
C434 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ui_in[6] 1.67e-19
C435 ringtest_0.x4._11_ a_24070_5852# 0.002559f
C436 ringtest_0.x4._19_ a_23770_5308# 8.51e-20
C437 muxtest_0.x1.x3.GP3 muxtest_0.R3R4 0.384927f
C438 a_24045_6654# VDPWR 0.175351f
C439 ringtest_0.x4.net6 a_24545_5878# 0.00514f
C440 a_21845_8816# ringtest_0.x4._11_ 9.54e-19
C441 ringtest_0.x4._12_ a_22399_8976# 0.023132f
C442 a_21852_8720# a_22245_8054# 0.011211f
C443 muxtest_0.x2.x2.GP2 m3_13302_19985# 0.005314f
C444 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR 0.637448f
C445 ringtest_0.x4.net6 a_25364_5878# 0.047825f
C446 ringtest_0.x4.net2 a_22245_8054# 3.45e-20
C447 ringtest_0.x4.counter[2] ua[1] 3.21e-19
C448 a_22097_5334# a_21509_4790# 0.002525f
C449 a_23381_4584# a_23467_4584# 0.006584f
C450 a_26627_4246# a_27273_4220# 0.016298f
C451 ringtest_0.x4._11_ a_23891_4790# 0.002312f
C452 a_25364_5878# a_24895_4790# 1.98e-20
C453 ringtest_0.x4.net11 a_25977_4220# 1.29e-21
C454 ringtest_0.x4._16_ a_21509_4790# 1.96e-20
C455 a_21852_9416# a_21845_9116# 0.966391f
C456 a_21465_9294# a_21981_9142# 1.28e-19
C457 a_21233_5340# a_21767_5334# 0.002698f
C458 ringtest_0.counter7 a_25975_3867# 8.66e-19
C459 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GP1 6.21e-20
C460 a_22392_5990# ringtest_0.x4.net5 1.47e-21
C461 ringtest_0.x4._11_ a_22373_5156# 0.045224f
C462 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP3 0.001226f
C463 muxtest_0.x1.x5.GN a_19242_32347# 1.08e-19
C464 muxtest_0.x1.x1.nSEL1 a_18836_32319# 0.00175f
C465 muxtest_0.R5R6 ui_in[2] 2.39e-19
C466 ringtest_0.x4.net1 a_21675_9686# 0.073427f
C467 a_22265_5308# a_23770_5308# 1e-20
C468 a_23879_6940# a_24883_6800# 8.9e-19
C469 ringtest_0.x4._15_ a_25593_5156# 1.98e-20
C470 ringtest_0.x4.net8 a_23899_5334# 2.79e-20
C471 ringtest_0.x4.net6 a_24551_4790# 7.29e-19
C472 ringtest_0.x4._11_ a_21767_5334# 3.45e-19
C473 ringtest_0.x4._16_ a_22765_5308# 0.243866f
C474 a_24336_6544# ringtest_0.x4._05_ 0.181338f
C475 ringtest_0.x4.counter[6] VDPWR 0.462317f
C476 a_24536_6699# a_24465_6800# 0.239923f
C477 a_24699_6200# VDPWR 0.2552f
C478 VDPWR ui_in[2] 4.46272f
C479 muxtest_0.R3R4 muxtest_0.R1R2 0.184502f
C480 a_21395_6940# a_21672_5334# 7.35e-19
C481 ringtest_0.x4.net6 a_24317_4942# 0.173962f
C482 muxtest_0.x2.x2.GN2 ui_in[4] 0.108808f
C483 ringtest_0.drv_out a_25393_5308# 1.4e-22
C484 a_22052_8875# VDPWR 0.271061f
C485 a_24317_4942# a_24895_4790# 0.00145f
C486 ringtest_0.x4.net9 ringtest_0.x4.counter[8] 2.39e-19
C487 ringtest_0.x4.net6 a_23151_5334# 7.79e-20
C488 ringtest_0.x4._15_ a_23993_5654# 0.004604f
C489 ringtest_0.x4.net8 ringtest_0.x4.counter[9] 1.68e-20
C490 ringtest_0.x4.net3 ringtest_0.x4._14_ 0.471315f
C491 a_27065_5334# a_26201_4790# 1.29e-19
C492 a_22116_4902# a_22541_5058# 1.28e-19
C493 a_27233_5308# ringtest_0.x4._09_ 5.87e-19
C494 a_21675_4790# a_22373_5156# 0.195152f
C495 ringtest_0.x4.net7 a_23770_5308# 0.142058f
C496 a_22399_8976# a_22245_8054# 6.31e-19
C497 a_21785_5878# a_24070_5852# 1.55e-21
C498 a_24479_4790# VDPWR 4.84e-19
C499 ringtest_0.x4._11_ a_26269_4612# 0.006396f
C500 ringtest_0.x4.clknet_0_clk a_26569_6422# 2.96e-20
C501 ringtest_0.x4._17_ a_23770_5308# 1.33e-19
C502 a_21465_8830# a_21780_8964# 7.84e-20
C503 a_23809_4790# VDPWR 0.211123f
C504 muxtest_0.x1.x3.GN3 muxtest_0.R6R7 0.260987f
C505 a_26201_5340# ringtest_0.x4.net10 4.73e-19
C506 ringtest_0.x4.clknet_1_0__leaf_clk a_21561_8830# 0.044938f
C507 a_21981_9142# a_21981_8976# 0.013661f
C508 ringtest_0.x4.net4 a_22021_4220# 0.021386f
C509 a_24045_6654# ringtest_0.x4._21_ 9.57e-19
C510 ringtest_0.x4._15_ ringtest_0.x4._04_ 3.75e-19
C511 a_22795_5334# VDPWR 0.261491f
C512 ringtest_0.x4._15_ a_25441_4612# 3.42e-21
C513 ringtest_0.x4.net1 a_22052_8875# 1.33e-19
C514 ringtest_0.x4._11_ a_22499_4790# 5.7e-19
C515 ringtest_0.drv_out ringtest_0.x3.x2.GN4 0.071598f
C516 a_26201_4790# a_26627_4246# 9.12e-19
C517 ringtest_0.x4._09_ a_25977_4220# 1.89e-19
C518 muxtest_0.x1.x4.A ua[0] 4.51511f
C519 a_21425_9686# a_21675_9686# 0.025037f
C520 a_21785_5878# a_22373_5156# 0.001131f
C521 ringtest_0.x4.net8 a_27149_5334# 2.29e-20
C522 ringtest_0.x4._04_ a_22541_5058# 7.11e-19
C523 ringtest_0.x4._07_ a_25393_5308# 0.008579f
C524 ringtest_0.x4._19_ ringtest_0.x4.net6 0.04173f
C525 a_21233_5340# a_21399_5340# 0.968904f
C526 ringtest_0.x4._22_ a_25225_5334# 1.1e-21
C527 ringtest_0.x4.net5 a_25149_4220# 1.18e-20
C528 ringtest_0.x4.clknet_1_0__leaf_clk a_22541_5058# 1.1e-19
C529 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.001676f
C530 ringtest_0.x4._18_ a_23949_6654# 0.006776f
C531 a_23879_6940# a_24045_6654# 0.017149f
C532 a_16579_11759# ringtest_0.x3.x2.GP2 3.07e-19
C533 a_21803_8598# VDPWR 0.004522f
C534 ringtest_0.x4._20_ a_25168_5156# 9.2e-20
C535 a_22649_6244# a_22765_5308# 0.001534f
C536 m3_13302_19985# ua[0] 0.003764f
C537 ringtest_0.x4._11_ a_21399_5340# 0.008371f
C538 ringtest_0.x4.net10 a_27233_5058# 0.008159f
C539 muxtest_0.x2.x2.GN1 ua[3] 4.69116f
C540 muxtest_0.x1.x4.A a_13675_24012# 2.9e-19
C541 ringtest_0.counter3 m3_17036_9140# 2.1e-20
C542 ringtest_0.x4.net8 ringtest_0.x4._16_ 0.193029f
C543 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN3 8.22e-19
C544 a_24699_6200# ringtest_0.x4._21_ 0.001146f
C545 ringtest_0.x4.counter[4] ringtest_0.x4.counter[5] 0.068962f
C546 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[6] 5.64e-20
C547 a_25421_6641# VDPWR 0.209324f
C548 ringtest_0.x4.clknet_1_1__leaf_clk a_26367_5340# 0.026802f
C549 ringtest_0.x4.clknet_0_clk a_24287_6422# 2.01e-19
C550 ringtest_0.x4.net6 a_22265_5308# 6.37e-19
C551 muxtest_0.x1.x3.GP2 muxtest_0.R6R7 4.11376f
C552 muxtest_0.x2.x2.GP2 ua[0] 4.069f
C553 ringtest_0.x4.net3 ringtest_0.x4._10_ 0.003052f
C554 ringtest_0.x4.net11 ringtest_0.x4.counter[9] 0.066386f
C555 ringtest_0.x4._22_ a_26640_5156# 0.004398f
C556 a_21587_5334# a_21509_4790# 2.5e-19
C557 ringtest_0.x4.net6 ringtest_0.x4.net9 0.566537f
C558 ringtest_0.x4.clknet_1_0__leaf_clk a_21049_8598# 3.26e-19
C559 ringtest_0.x4._23_ a_25975_3867# 2.99e-20
C560 muxtest_0.x2.x2.GN3 m3_13302_19985# 0.087318f
C561 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR 0.637284f
C562 ringtest_0.x4._16_ a_24729_4790# 1.25e-20
C563 a_21399_5340# a_21675_4790# 6.25e-19
C564 ringtest_0.counter7 m3_17032_8096# 6.07e-21
C565 ringtest_0.x4.net11 a_27491_4566# 0.001149f
C566 ringtest_0.x4._24_ ringtest_0.x4._08_ 0.423487f
C567 ringtest_0.x4.net9 a_24895_4790# 0.017191f
C568 ringtest_0.x4._15_ ringtest_0.x4.net4 0.003757f
C569 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP1 4.57902f
C570 ringtest_0.x4._00_ a_21845_8816# 8.76e-20
C571 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GN4 0.190572f
C572 ringtest_0.x4._18_ a_24004_6128# 5.77e-19
C573 a_23879_6940# a_24699_6200# 6.61e-19
C574 a_19794_32347# VDPWR 0.001496f
C575 ringtest_0.x4._21_ a_23809_4790# 0.087922f
C576 a_25393_5308# a_26201_5340# 4.62e-19
C577 a_20318_32213# muxtest_0.x1.x3.GN2 7.58e-21
C578 muxtest_0.x1.x3.GN1 a_18836_32319# 0.001144f
C579 a_25421_6641# ringtest_0.x4._25_ 6.03e-21
C580 ringtest_0.x4._17_ a_24712_6422# 0.002153f
C581 a_21672_5334# VDPWR 0.259474f
C582 ringtest_0.x4.net6 ringtest_0.x4.net7 0.905861f
C583 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP2 2.65608f
C584 muxtest_0.x1.x1.nSEL1 a_19290_32287# 0.041068f
C585 ringtest_0.x4.net4 a_22541_5058# 0.020834f
C586 ringtest_0.x4.clknet_1_1__leaf_clk a_27065_5156# 2.2e-19
C587 ringtest_0.ring_out ringtest_0.x3.nselect2 0.006614f
C588 ringtest_0.x4.net7 a_24895_4790# 0.030766f
C589 a_23949_6654# ringtest_0.x4.clknet_1_1__leaf_clk 1.77e-20
C590 ringtest_0.x4._17_ ringtest_0.x4.net6 0.277113f
C591 ringtest_0.x4.net3 a_21509_4790# 0.005671f
C592 ringtest_0.x4.net2 ringtest_0.counter7 6.88e-20
C593 muxtest_0.R7R8 muxtest_0.x2.x2.GP3 0.17349f
C594 ringtest_0.x4._17_ a_24895_4790# 6.74e-21
C595 a_16579_11759# a_16707_12151# 0.004764f
C596 a_16579_11759# ringtest_0.x3.x2.GN2 1.63e-19
C597 a_21785_5878# a_21399_5340# 1.36e-19
C598 a_21951_5878# a_21233_5340# 9.16e-19
C599 ringtest_0.x4._18_ a_23381_4818# 1.7e-19
C600 ringtest_0.x4._23_ a_26367_5340# 0.031087f
C601 a_22097_5334# a_22390_4566# 3.78e-21
C602 ringtest_0.x4._24_ VDPWR 0.6956f
C603 a_26367_5340# a_26367_4790# 0.027195f
C604 a_26201_5340# a_26808_4902# 1.99e-20
C605 ringtest_0.x4._11_ a_21951_5878# 0.082924f
C606 ringtest_0.x4._16_ a_22390_4566# 3.76e-19
C607 a_22649_6244# ringtest_0.x4.net8 3.5e-19
C608 muxtest_0.x1.x5.A muxtest_0.R4R5 4.5151f
C609 ringtest_0.x4.net3 a_21867_8054# 1.25e-19
C610 a_24336_6544# a_24361_5340# 1.6e-20
C611 a_24329_6640# a_24527_5340# 3.93e-19
C612 ringtest_0.x4._15_ a_23837_5878# 9.44e-19
C613 ringtest_0.x4._15_ ringtest_0.x4._22_ 0.422897f
C614 ringtest_0.x4._11_ a_24883_6800# 7.39e-21
C615 ringtest_0.x4._05_ ringtest_0.x4._16_ 0.001611f
C616 ringtest_0.x4.net3 ringtest_0.x4._13_ 0.031667f
C617 ringtest_0.x4._07_ a_25083_4790# 0.128255f
C618 ringtest_0.x3.x2.GP2 m3_17032_8096# 0.005314f
C619 ringtest_0.x4.clknet_0_clk a_24329_6640# 0.043419f
C620 ringtest_0.x4.net6 a_22817_6146# 0.129987f
C621 ringtest_0.x4.clknet_1_1__leaf_clk a_24004_6128# 0.007927f
C622 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP2 0.059353f
C623 a_21465_9294# ringtest_0.x4._12_ 6.08e-20
C624 a_23891_4790# ringtest_0.x4.counter[4] 4.37e-20
C625 ringtest_0.x4._14_ ringtest_0.x4._03_ 0.071143f
C626 ringtest_0.x4._24_ ringtest_0.x4._25_ 0.095329f
C627 ringtest_0.x4._09_ a_27491_4566# 0.002954f
C628 a_25083_4790# a_25055_3867# 7.39e-20
C629 a_25593_5156# a_25975_3867# 3.85e-20
C630 a_16579_11759# ui_in[3] 0.086353f
C631 ringtest_0.x4.net7 a_27169_6641# 2.85e-19
C632 ringtest_0.x4._23_ a_27065_5156# 0.006274f
C633 a_27233_5058# a_27191_4790# 7.84e-20
C634 a_26808_4902# a_27233_5058# 1.28e-19
C635 a_26367_4790# a_27065_5156# 0.194892f
C636 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ui_in[4] 2.42e-19
C637 ringtest_0.x4._06_ a_25393_5308# 1.75e-19
C638 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.025028f
C639 a_23879_6940# a_25421_6641# 1.59e-19
C640 a_24699_6200# a_24968_5308# 1e-18
C641 a_27815_3867# VDPWR 0.276039f
C642 ringtest_0.x3.x2.GP3 ringtest_0.counter7 0.165274f
C643 a_11845_23906# muxtest_0.x2.x2.GN2 0.039612f
C644 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN3 0.012418f
C645 a_22224_6244# VDPWR 0.255338f
C646 ringtest_0.x4._08_ a_27233_5308# 0.004928f
C647 ringtest_0.x4.clknet_1_1__leaf_clk a_23381_4818# 2.67e-20
C648 a_22350_5878# ringtest_0.x4._16_ 2.63e-21
C649 a_27149_5334# ringtest_0.x4._09_ 1.2e-19
C650 a_26007_6788# VDPWR 0.001434f
C651 ringtest_0.x4.clknet_0_clk a_25364_5878# 0.316676f
C652 muxtest_0.x2.x2.GP3 VDPWR 1.78328f
C653 ringtest_0.x3.x1.nSEL0 a_15575_12017# 0.081627f
C654 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.nselect2 0.047548f
C655 ringtest_0.x4._15_ a_25225_5334# 0.0351f
C656 muxtest_0.R7R8 muxtest_0.R2R3 0.215077f
C657 ringtest_0.x4._22_ a_26173_4612# 0.001961f
C658 ringtest_0.x4._01_ a_21395_6940# 3.77e-19
C659 muxtest_0.R7R8 ui_in[1] 4.98e-22
C660 a_21785_5878# a_21951_5878# 0.966818f
C661 a_16155_12151# VDPWR 2.96e-19
C662 ringtest_0.x3.x2.GN1 VDPWR 1.47002f
C663 a_21981_8976# ringtest_0.x4._12_ 0.039032f
C664 ringtest_0.x4._11_ a_23381_4584# 0.002917f
C665 a_22265_5308# ringtest_0.x4.net5 6.71e-21
C666 muxtest_0.x1.x3.GP1 muxtest_0.x1.x4.A 0.354981f
C667 muxtest_0.x2.x2.GN3 ua[0] 0.214839f
C668 ringtest_0.x4._11_ a_26555_4790# 2.79e-20
C669 ringtest_0.x3.x2.GN4 m3_17036_9140# 7.17e-19
C670 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR 0.637855f
C671 ringtest_0.x3.x2.GN2 m3_17032_8096# 0.016745f
C672 ringtest_0.x4._17_ a_23932_6128# 0.002503f
C673 a_24465_6800# ringtest_0.x4.net8 0.00192f
C674 muxtest_0.x1.x5.GN muxtest_0.R7R8 0.558172f
C675 ringtest_0.x4._11_ a_24045_6654# 1.82e-19
C676 a_24361_5340# a_23899_5334# 1.44e-19
C677 a_19666_31955# muxtest_0.x1.x3.GP1 1.19e-20
C678 ringtest_0.x4.clknet_1_1__leaf_clk a_26375_4612# 5.67e-20
C679 a_27233_5308# VDPWR 0.48745f
C680 a_24536_6699# a_24712_6422# 0.007724f
C681 ringtest_0.x4._15_ a_22021_4220# 3.5e-20
C682 ringtest_0.x4.net6 a_26627_4246# 5.59e-20
C683 a_19290_32287# muxtest_0.x1.x3.GN1 1.45e-19
C684 ringtest_0.x4._15_ a_26640_5156# 0.001788f
C685 a_25168_5156# a_25149_4220# 1.83e-19
C686 VDPWR ui_in[6] 1.10022f
C687 muxtest_0.x1.x5.A ui_in[2] 5.67943f
C688 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x3.nselect2 2.88e-20
C689 a_12977_24040# muxtest_0.x2.x2.GN4 3.22e-19
C690 muxtest_0.x2.x2.GN3 a_13675_24012# 1.07e-20
C691 a_24536_6699# ringtest_0.x4.net6 6.81e-19
C692 a_25336_4902# a_25719_4790# 4.67e-20
C693 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP3 0.031766f
C694 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GN4 8.84e-19
C695 a_21948_5156# a_22164_4362# 0.003601f
C696 ua[3] ua[6] 0.008019f
C697 muxtest_0.x2.x2.GP1 ui_in[4] 0.001143f
C698 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._20_ 0.0051f
C699 a_24329_6640# a_25168_5156# 7.91e-22
C700 a_19114_31955# ui_in[2] 8.66e-20
C701 a_12297_23648# ui_in[4] 0.03417f
C702 ringtest_0.x3.nselect2 ringtest_0.x3.x2.GN3 7.39e-21
C703 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN4 2.26e-20
C704 a_21780_9142# VDPWR 4.59e-19
C705 a_25977_4220# VDPWR 0.419035f
C706 a_21785_8054# a_21395_6940# 5.68e-19
C707 ringtest_0.x4._11_ ringtest_0.x4.counter[6] 0.002692f
C708 ringtest_0.x4._10_ a_21939_8054# 5.49e-20
C709 a_21561_9116# VDPWR 0.19379f
C710 a_25719_4790# VDPWR 2.75e-19
C711 ringtest_0.x4._11_ a_24699_6200# 0.042839f
C712 uio_in[0] ui_in[7] 0.031023f
C713 ringtest_0.x4._19_ a_24527_5340# 4.93e-21
C714 a_21509_4790# ringtest_0.x4._03_ 0.095111f
C715 a_24336_6544# VDPWR 0.321592f
C716 ringtest_0.x4.net2 ringtest_0.x4._02_ 0.035742f
C717 ringtest_0.x4.net3 ringtest_0.x4.counter[1] 0.103986f
C718 muxtest_0.x1.x3.GN4 muxtest_0.R3R4 0.237766f
C719 muxtest_0.R2R3 VDPWR 1.6072f
C720 ringtest_0.x4.clknet_0_clk ringtest_0.x4._19_ 0.038005f
C721 a_21465_8830# a_21845_8816# 0.048748f
C722 VDPWR ui_in[1] 2.66846f
C723 ringtest_0.x4._04_ a_22765_4478# 1.25e-20
C724 ringtest_0.x4.net3 a_22390_4566# 9.94e-20
C725 ringtest_0.counter3 ua[1] 4.52195f
C726 muxtest_0.x1.x5.GN muxtest_0.R5R6 7.03e-21
C727 a_25761_5058# ringtest_0.x4.counter[6] 4.54e-21
C728 ringtest_0.x4.net8 a_26201_4790# 3.27e-19
C729 ringtest_0.x4._23_ a_26375_4612# 1.08e-20
C730 ringtest_0.x4._11_ a_24479_4790# 0.001677f
C731 a_21981_9142# a_22201_9142# 4.62e-19
C732 ringtest_0.x4.net11 a_27273_4220# 0.088145f
C733 a_21845_9116# a_22052_9116# 0.273138f
C734 a_21561_9116# a_21803_9508# 0.008508f
C735 a_21852_9416# a_21981_9142# 0.110715f
C736 ringtest_0.counter7 a_27489_3702# 3.7e-19
C737 a_21233_5340# a_22795_5334# 2.77e-19
C738 ringtest_0.x4._18_ a_22392_5990# 1.41e-19
C739 ringtest_0.x4.net1 a_21780_9142# 2.14e-19
C740 ringtest_0.x4._11_ a_23809_4790# 0.222369f
C741 ringtest_0.x4._14_ a_21055_5334# 6.31e-19
C742 ringtest_0.x4.clknet_1_1__leaf_clk a_26569_6422# 7.87e-19
C743 muxtest_0.x1.x5.GN VDPWR 3.74211f
C744 ringtest_0.x4.net1 a_21561_9116# 0.017118f
C745 a_22111_10993# a_21852_9416# 4.65e-23
C746 ringtest_0.x4._06_ a_24715_5334# 0.114717f
C747 a_24986_5878# VDPWR 1.76e-19
C748 ringtest_0.x4.net10 a_26895_3867# 2.65e-20
C749 ringtest_0.x4.net8 a_26555_5334# 1.28e-19
C750 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[4] 8.27e-22
C751 ringtest_0.x4._11_ a_22795_5334# 2.49e-20
C752 ringtest_0.x4._16_ a_24361_5340# 1.57e-19
C753 a_12849_23648# muxtest_0.x2.x2.GP3 0.00144f
C754 ringtest_0.x4.net9 a_24527_5340# 0.002182f
C755 a_24465_6800# ringtest_0.x4._05_ 0.001005f
C756 a_16707_12151# ringtest_0.x3.x2.GP3 4.39e-19
C757 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.001676f
C758 a_22139_5878# VDPWR 0.093135f
C759 a_25336_4902# a_25677_5156# 9.73e-19
C760 ua[2] ua[1] 1.12657f
C761 a_24729_4790# a_26201_4790# 0.003146f
C762 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP3 0.004296f
C763 ringtest_0.x4._15_ a_22541_5058# 2.99e-20
C764 muxtest_0.x2.nselect2 a_13025_23980# 6.01e-20
C765 muxtest_0.x1.x1.nSEL0 ui_in[2] 0.131256f
C766 ringtest_0.x4._01_ VDPWR 0.468919f
C767 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net9 0.132797f
C768 ringtest_0.x4._15_ a_24926_5712# 0.002542f
C769 ringtest_0.x4._07_ a_25055_3867# 7.51e-19
C770 ringtest_0.x4._22_ a_25975_3867# 2.78e-19
C771 ringtest_0.x4._14_ a_22939_4584# 5.76e-19
C772 ringtest_0.x4.net7 a_24527_5340# 0.456298f
C773 ringtest_0.x4._04_ a_24004_6128# 3.15e-21
C774 a_21007_3867# ringtest_0.x4.counter[0] 0.109791f
C775 a_25677_5156# VDPWR 0.004788f
C776 ringtest_0.x4._17_ a_24527_5340# 1.22e-20
C777 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net7 0.043959f
C778 a_21863_4790# VDPWR 0.083158f
C779 muxtest_0.x1.x3.GN2 muxtest_0.R4R5 0.116214f
C780 a_26808_5308# ringtest_0.x4.net10 2.56e-19
C781 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR 0.637064f
C782 ringtest_0.x4.clknet_1_0__leaf_clk a_21852_8720# 0.083453f
C783 a_24336_6544# ringtest_0.x4._21_ 0.001538f
C784 ringtest_0.x4.net4 a_22765_4478# 0.130038f
C785 ringtest_0.x4.counter[4] ua[1] 3.21e-19
C786 ringtest_0.x4._11_ a_25421_6641# 0.004334f
C787 ringtest_0.x3.x2.GP3 ui_in[3] 2.82e-19
C788 ringtest_0.x4.net2 ringtest_0.x4._04_ 4.09e-22
C789 ringtest_0.x4.clknet_0_clk ringtest_0.x4._17_ 0.029087f
C790 a_23899_5334# VDPWR 0.206364f
C791 ringtest_0.x4.net6 a_26721_4246# 7.2e-20
C792 ringtest_0.x4._15_ a_26173_4612# 0.006963f
C793 ringtest_0.x4.net1 ringtest_0.x4._01_ 1.96e-19
C794 a_25925_6788# ringtest_0.x4._24_ 4.18e-19
C795 ringtest_0.x4._23_ a_26569_6422# 0.213625f
C796 ringtest_0.x4.net2 ringtest_0.x4.clknet_1_0__leaf_clk 0.026712f
C797 ringtest_0.x4._09_ a_27273_4220# 0.17213f
C798 ringtest_0.x4._00_ a_21675_9686# 0.07841f
C799 a_21425_9686# a_21561_9116# 7.31e-19
C800 a_26749_6422# a_26201_4790# 3.35e-21
C801 ringtest_0.x4._09_ a_26766_4790# 3.07e-19
C802 a_26201_4790# ringtest_0.x4.net11 3.07e-19
C803 ringtest_0.x4._02_ a_21840_5308# 4.65e-19
C804 ringtest_0.x4._22_ a_26367_5340# 4.96e-21
C805 a_21233_5340# a_21672_5334# 0.273138f
C806 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x3.nselect2 5.69e-21
C807 ringtest_0.x4._08_ a_27149_5334# 2.34e-19
C808 ringtest_0.x4.counter[9] VDPWR 0.449609f
C809 ringtest_0.x4._18_ a_24329_6640# 6.58e-19
C810 a_21785_8054# VDPWR 0.266078f
C811 a_23879_6940# a_24336_6544# 0.016444f
C812 ringtest_0.x4.net8 a_23770_5308# 2.76e-19
C813 ringtest_0.x4._20_ a_25593_5156# 1.2e-20
C814 ringtest_0.x4.clknet_1_0__leaf_clk a_22181_5334# 3.7e-19
C815 ringtest_0.x4._11_ a_21672_5334# 0.003174f
C816 ringtest_0.x4._07_ ringtest_0.x4.counter[5] 1.62e-19
C817 a_27491_4566# VDPWR 0.003335f
C818 ringtest_0.counter3 m3_17046_7066# 8.01e-20
C819 ringtest_0.x4.clknet_0_clk a_22817_6146# 3.43e-19
C820 ringtest_0.drv_out m3_17036_9140# 0.132758f
C821 muxtest_0.R7R8 ui_in[4] 0.104361f
C822 a_25055_3867# ringtest_0.x4.counter[5] 0.1107f
C823 ringtest_0.x4.clknet_1_1__leaf_clk a_26640_5334# 0.001015f
C824 ringtest_0.x4.net6 a_22765_5308# 0.080758f
C825 ringtest_0.x4.clknet_0_clk a_26095_6788# 9.17e-20
C826 a_12019_24012# VDPWR 9.09e-19
C827 ringtest_0.x4._11_ ringtest_0.x4._24_ 4.57e-19
C828 ringtest_0.x4.clknet_1_0__leaf_clk a_22399_8976# 0.018091f
C829 a_23949_6654# a_23837_5878# 2.76e-20
C830 ringtest_0.x4._23_ a_27489_3702# 9.55e-20
C831 a_27273_4220# a_27659_4246# 0.006406f
C832 ringtest_0.x4._14_ ringtest_0.x4.net5 0.258421f
C833 a_24329_6640# a_24763_6143# 0.00484f
C834 ringtest_0.x4._16_ a_25336_4902# 8.82e-22
C835 a_27149_5334# VDPWR 0.00533f
C836 a_21399_5340# a_21948_5156# 0.002f
C837 a_21672_5334# a_21675_4790# 0.004962f
C838 ringtest_0.x4.net9 a_25168_5156# 0.003585f
C839 ringtest_0.x4.net11 a_27303_4246# 0.01512f
C840 a_26808_4902# a_26895_3867# 2.21e-20
C841 ringtest_0.x4.net1 a_21785_8054# 0.232539f
C842 ringtest_0.x4.net6 ringtest_0.x4._13_ 2.81e-21
C843 a_25925_6788# a_26007_6788# 0.005781f
C844 ringtest_0.x4.net2 ringtest_0.x4.net4 8.49e-21
C845 a_22097_5334# a_22223_5712# 0.006169f
C846 a_25225_5334# a_26367_5340# 8.68e-20
C847 ringtest_0.x4.clknet_1_1__leaf_clk a_25149_4220# 1.84e-19
C848 a_22097_5334# VDPWR 0.228175f
C849 ringtest_0.x4.net4 a_23381_4818# 4.87e-19
C850 muxtest_0.x1.x1.nSEL1 a_19842_32287# 1.59e-19
C851 ringtest_0.x4._16_ VDPWR 2.17996f
C852 a_26201_4790# ringtest_0.x4._09_ 0.098799f
C853 ringtest_0.x4.net7 a_25168_5156# 0.005696f
C854 ringtest_0.x4._03_ a_22390_4566# 9.33e-19
C855 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk 0.228247f
C856 a_22695_8304# VDPWR 0.006514f
C857 ringtest_0.x3.x2.GN4 ua[1] 0.446629f
C858 muxtest_0.x1.x3.GN2 ui_in[2] 0.001516f
C859 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.025028f
C860 a_24763_6143# a_24545_5878# 0.004465f
C861 ringtest_0.x4._06_ ringtest_0.x4._07_ 5.11e-20
C862 a_11845_23906# a_12297_23648# 0.002207f
C863 a_16755_12091# ringtest_0.x3.x2.GN4 0.003699f
C864 a_24004_6128# a_23837_5878# 0.046138f
C865 a_17231_12017# ringtest_0.x3.x2.GN2 7.58e-21
C866 a_21785_5878# a_21672_5334# 0.002054f
C867 ringtest_0.x3.x2.GN1 a_15749_12123# 0.001144f
C868 ringtest_0.x4._04_ a_21840_5308# 8.38e-20
C869 ringtest_0.x4._14_ a_21007_3867# 0.001394f
C870 ringtest_0.x4._23_ a_26640_5334# 0.012578f
C871 ringtest_0.x4.clknet_1_0__leaf_clk a_21840_5308# 0.01796f
C872 a_26367_5340# a_26640_5156# 1.54e-19
C873 a_26808_5308# a_26808_4902# 0.012451f
C874 a_26640_5334# a_26367_4790# 1.54e-19
C875 ringtest_0.x4._18_ a_23151_5334# 2.06e-20
C876 ringtest_0.x4._16_ a_23467_4584# 8.82e-20
C877 ringtest_0.x4._11_ a_22224_6244# 0.054008f
C878 a_21852_9416# ui_in[5] 4.56e-21
C879 muxtest_0.x1.x4.A muxtest_0.R4R5 0.003925f
C880 a_24465_6800# a_24361_5340# 5.48e-20
C881 ringtest_0.x4.net3 a_21395_6940# 0.011213f
C882 a_24536_6699# a_24527_5340# 8.21e-21
C883 a_24329_6640# a_24800_5334# 8.34e-21
C884 ringtest_0.x4._11_ a_26007_6788# 2.28e-19
C885 ringtest_0.x4.clknet_1_1__leaf_clk a_24545_5878# 3.57e-20
C886 ringtest_0.x4.net11 ringtest_0.x4.counter[8] 0.024563f
C887 VDPWR ui_in[4] 9.60897f
C888 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR 0.636224f
C889 ringtest_0.x4.clknet_0_clk a_24536_6699# 0.004436f
C890 ringtest_0.x4.clknet_1_1__leaf_clk a_25364_5878# 1.80017f
C891 a_21425_9686# a_21785_8054# 2.44e-21
C892 ringtest_0.x4.net6 ringtest_0.x4.net8 0.806426f
C893 a_21852_9416# ringtest_0.x4._12_ 0.003541f
C894 ringtest_0.x4._09_ a_27303_4246# 0.07143f
C895 muxtest_0.x2.nselect2 ui_in[3] 1.88e-19
C896 ringtest_0.x4.net8 a_24895_4790# 0.003497f
C897 ringtest_0.x4._23_ a_25149_4220# 2.79e-19
C898 a_17231_12017# ui_in[3] 0.220366f
C899 a_23809_4790# ringtest_0.x4.counter[4] 2.6e-19
C900 ringtest_0.x4._23_ a_26735_5156# 8.32e-19
C901 a_26808_4902# a_26555_4790# 3.39e-19
C902 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP1 8.08e-19
C903 muxtest_0.R7R8 ui_in[0] 2.25e-21
C904 ringtest_0.x4.net10 a_26817_4566# 8.38e-19
C905 ringtest_0.x4._06_ a_26201_5340# 4.19e-21
C906 ringtest_0.x4.net6 a_24729_4790# 0.083542f
C907 ringtest_0.x4._18_ ringtest_0.x4._19_ 0.036736f
C908 a_12473_23980# muxtest_0.x2.x2.GN2 0.017071f
C909 a_22649_6244# VDPWR 0.169689f
C910 a_24729_4790# a_24895_4790# 0.966391f
C911 ringtest_0.x4.clknet_1_1__leaf_clk a_24317_4942# 0.050301f
C912 ringtest_0.x4._21_ ringtest_0.x4._16_ 0.249175f
C913 a_26201_6788# VDPWR 0.002272f
C914 ringtest_0.x4._16_ ringtest_0.x4.counter[2] 3.86e-19
C915 ringtest_0.x4.net4 a_21840_5308# 5.24e-19
C916 ringtest_0.x4.clknet_1_1__leaf_clk a_23151_5334# 8.24e-20
C917 ringtest_0.x3.x1.nSEL0 a_16203_12091# 0.001174f
C918 ringtest_0.x4._15_ a_26367_5340# 0.058771f
C919 a_21509_4790# ringtest_0.x4.net5 8.46e-19
C920 ringtest_0.x4._03_ a_22074_4790# 0.001074f
C921 ringtest_0.x4._22_ a_26375_4612# 2.76e-20
C922 ringtest_0.x3.x2.GP1 VDPWR 1.86466f
C923 ringtest_0.x4._04_ a_22392_5990# 0.04931f
C924 a_21785_5878# a_22224_6244# 0.269567f
C925 a_23467_4818# VDPWR 0.00273f
C926 ringtest_0.x4._18_ a_22265_5308# 3.26e-20
C927 ringtest_0.x4._11_ a_25977_4220# 0.19543f
C928 a_22765_5308# ringtest_0.x4.net5 0.001034f
C929 ringtest_0.x4._23_ a_25364_5878# 0.042503f
C930 ringtest_0.x4.clknet_1_0__leaf_clk a_22392_5990# 5.16e-19
C931 a_21852_9416# a_22245_8054# 6.42e-21
C932 muxtest_0.x1.x3.GN1 ua[3] 4.34e-20
C933 ringtest_0.x3.x2.GN4 m3_17046_7066# 0.084813f
C934 ringtest_0.x4._11_ a_25719_4790# 2.44e-19
C935 a_23837_5878# ringtest_0.x4._20_ 6.22e-20
C936 a_25364_5878# a_26367_4790# 2.14e-19
C937 a_19114_31955# ui_in[1] 0.03417f
C938 a_23879_6940# ringtest_0.x4._16_ 4.51e-19
C939 ringtest_0.x4._22_ ringtest_0.x4._20_ 2.69e-20
C940 ringtest_0.counter7 ringtest_0.x4.net9 0.006102f
C941 a_24361_5340# a_26555_5334# 2.33e-21
C942 ringtest_0.x4._11_ a_24336_6544# 3.7e-19
C943 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A 4.01025f
C944 a_21587_5334# VDPWR 0.075425f
C945 a_19242_32347# muxtest_0.x1.x3.GN3 5.17e-20
C946 muxtest_0.x1.x3.GN2 a_19794_32347# 3.11e-20
C947 ringtest_0.x4._15_ a_22765_4478# 1.84e-19
C948 ringtest_0.ring_out ringtest_0.x3.x2.GP2 0.080385f
C949 ringtest_0.x4.net6 a_26749_6422# 7.38e-20
C950 a_19842_32287# muxtest_0.x1.x3.GN1 1.69e-20
C951 a_25761_5058# a_25977_4220# 0.001105f
C952 muxtest_0.x1.x5.GN a_19114_31955# 3.56e-19
C953 muxtest_0.x1.x4.A ui_in[2] 4.96786f
C954 ringtest_0.x4._05_ ringtest_0.x4.net6 0.03493f
C955 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._19_ 0.060342f
C956 a_23949_6654# ringtest_0.x4._15_ 1.78e-19
C957 a_25761_5058# a_25719_4790# 7.84e-20
C958 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ui_in[4] 4.96e-21
C959 ringtest_0.x4._18_ ringtest_0.x4.net7 0.004371f
C960 ringtest_0.counter7 ringtest_0.x4.net7 6.88e-20
C961 a_22541_5058# a_22765_4478# 0.001036f
C962 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.001676f
C963 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 3.14e-21
C964 ringtest_0.x4._24_ ringtest_0.x4.net10 0.13484f
C965 a_19666_31955# ui_in[2] 0.009143f
C966 VDPWR ui_in[0] 1.24711f
C967 a_22139_5878# a_21233_5340# 3.23e-19
C968 ringtest_0.x4._17_ ringtest_0.x4._18_ 0.181987f
C969 muxtest_0.R3R4 muxtest_0.x2.x2.GN2 0.015374f
C970 ringtest_0.x4.net9 a_24763_6143# 0.122363f
C971 a_12849_23648# ui_in[4] 0.261734f
C972 ringtest_0.x4.net3 VDPWR 2.1402f
C973 a_27273_4220# VDPWR 0.230416f
C974 a_24070_5852# ringtest_0.x4._06_ 0.004838f
C975 a_21845_9116# VDPWR 0.721856f
C976 a_26766_4790# VDPWR -4.73e-35
C977 a_22649_6244# ringtest_0.x4._21_ 8.88e-21
C978 ringtest_0.x4.net8 a_23932_6128# 0.001644f
C979 ringtest_0.x4._11_ a_22139_5878# 0.020189f
C980 a_27659_4246# ringtest_0.x4.counter[8] 1.28e-20
C981 ringtest_0.x4._19_ a_24800_5334# 6.46e-21
C982 a_24465_6800# VDPWR 0.191062f
C983 ringtest_0.x4._01_ ringtest_0.x4._11_ 0.20957f
C984 ringtest_0.x4._12_ ringtest_0.x4._10_ 0.002721f
C985 ringtest_0.x4.net4 a_22392_5990# 0.034264f
C986 ringtest_0.x4.net7 a_24763_6143# 1.85e-20
C987 ringtest_0.x4._15_ a_24004_6128# 5.11e-20
C988 a_21561_8830# a_21852_8720# 0.192341f
C989 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net9 0.461828f
C990 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR 0.636188f
C991 ringtest_0.x4._23_ a_26913_4566# 2.44e-19
C992 a_25149_4220# a_25441_4612# 0.001675f
C993 ringtest_0.x4._17_ a_24763_6143# 2.72e-19
C994 muxtest_0.x1.x1.nSEL0 ui_in[1] 0.137587f
C995 a_25364_5878# a_25593_5156# 0.001605f
C996 a_26749_6422# a_27169_6641# 0.017591f
C997 ringtest_0.drv_out ua[1] 4.52048f
C998 ringtest_0.x4.net2 a_21561_8830# 0.00144f
C999 a_21465_9294# ringtest_0.x4.clknet_1_0__leaf_clk 0.007095f
C1000 ringtest_0.counter7 ringtest_0.x4.counter[0] 0.003899f
C1001 ringtest_0.x4._08_ a_26201_4790# 1.13e-19
C1002 a_22052_9116# a_21981_9142# 0.239923f
C1003 ringtest_0.x4._18_ a_22817_6146# 0.001543f
C1004 ringtest_0.x4.net1 ringtest_0.x4.net3 0.313425f
C1005 ringtest_0.x4.net8 ringtest_0.x4.net5 0.002187f
C1006 ringtest_0.x4._11_ a_21863_4790# 4.78e-19
C1007 ringtest_0.ring_out a_16707_12151# 2.99e-20
C1008 a_22111_10993# a_22052_9116# 2.02e-20
C1009 a_23770_5308# a_24361_5340# 0.044245f
C1010 ringtest_0.x4.net1 a_21845_9116# 0.003904f
C1011 ringtest_0.x4._19_ ringtest_0.x4._23_ 2.58e-20
C1012 ringtest_0.ring_out ringtest_0.x3.x2.GN2 0.23158f
C1013 ringtest_0.x4.net10 a_27815_3867# 0.219068f
C1014 ringtest_0.x4.net8 a_24895_5334# 4.84e-19
C1015 ringtest_0.x4.net6 ringtest_0.x4._09_ 1.5e-20
C1016 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net7 0.397702f
C1017 ringtest_0.x4._15_ a_23963_4790# 2.18e-19
C1018 ringtest_0.x4._11_ a_23899_5334# 0.07562f
C1019 muxtest_0.x2.x2.GP3 ua[2] 0.357853f
C1020 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x5.GN 0.043714f
C1021 ringtest_0.x4._16_ a_24968_5308# 0.001117f
C1022 ringtest_0.x4.net9 a_24800_5334# 6.38e-21
C1023 a_22733_6244# VDPWR 0.004177f
C1024 ringtest_0.x4._08_ a_26555_5334# 0.134213f
C1025 a_25168_5156# a_25294_4790# 0.005525f
C1026 ringtest_0.x4.clknet_0_clk a_22765_5308# 4.87e-21
C1027 ringtest_0.x4._15_ a_23381_4818# 0.22097f
C1028 ringtest_0.x4._17_ ringtest_0.x4.clknet_1_1__leaf_clk 0.044595f
C1029 ringtest_0.x4._23_ a_26735_5334# 8.32e-19
C1030 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN2 0.154394f
C1031 ringtest_0.x3.x2.GN3 ringtest_0.counter7 0.005062f
C1032 muxtest_0.R7R8 muxtest_0.x2.x2.GN4 3.97956f
C1033 a_22541_5058# a_23381_4818# 7.43e-20
C1034 a_21675_4790# a_21863_4790# 0.097994f
C1035 ringtest_0.x4._14_ a_22486_4246# 0.003598f
C1036 ringtest_0.x4.net7 a_24800_5334# 0.034093f
C1037 a_26201_4790# VDPWR 0.667506f
C1038 a_21785_5878# a_22139_5878# 0.062224f
C1039 ringtest_0.x4._10_ a_22245_8054# 0.423817f
C1040 a_21785_8054# ringtest_0.x4._11_ 0.005192f
C1041 uio_in[5] uio_in[4] 0.031023f
C1042 ringtest_0.ring_out ui_in[3] 3.69e-19
C1043 muxtest_0.x1.x3.GP3 ua[3] 0.023203f
C1044 ringtest_0.x4.net3 ringtest_0.x4.counter[2] 7.38e-19
C1045 a_11845_23906# VDPWR 0.211573f
C1046 ringtest_0.x4._23_ ringtest_0.x4.net9 0.065132f
C1047 ringtest_0.x4._17_ a_24800_5334# 9.6e-21
C1048 a_22457_5156# VDPWR 0.004797f
C1049 ringtest_0.x4.net9 a_26367_4790# 0.047741f
C1050 ua[3] ua[5] 0.008019f
C1051 a_23899_5654# a_23899_5334# 6.96e-20
C1052 a_27065_5334# a_27191_5712# 0.006169f
C1053 a_27233_5308# ringtest_0.x4.net10 0.084593f
C1054 ringtest_0.x4.clknet_1_0__leaf_clk a_21981_8976# 0.024273f
C1055 a_24465_6800# ringtest_0.x4._21_ 1.21e-19
C1056 a_26555_5334# VDPWR 0.078044f
C1057 ringtest_0.x4._15_ a_26375_4612# 0.002119f
C1058 ringtest_0.x4.net2 a_21049_8598# 0.07281f
C1059 a_19842_32287# muxtest_0.x1.x3.GP3 4.69e-19
C1060 muxtest_0.x2.x1.nSEL1 ui_in[2] 8.19e-21
C1061 a_19666_31955# a_19794_32347# 0.004764f
C1062 ringtest_0.x4.net7 ringtest_0.x4._23_ 0.074369f
C1063 a_21425_9686# a_21845_9116# 0.001828f
C1064 ringtest_0.x4._24_ a_26808_4902# 0.014122f
C1065 ringtest_0.x4._00_ a_21561_9116# 0.001635f
C1066 ringtest_0.x4.net7 a_26367_4790# 0.001362f
C1067 a_21233_5340# a_22097_5334# 0.032244f
C1068 ringtest_0.x4.net5 a_22390_4566# 0.075434f
C1069 ringtest_0.x4._02_ a_22265_5308# 1.8e-19
C1070 ringtest_0.counter7 a_26627_4246# 1.91e-19
C1071 ringtest_0.x4._17_ ringtest_0.x4._23_ 0.082072f
C1072 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ui_in[4] 4.96e-21
C1073 ringtest_0.x4._04_ a_23151_5334# 2.55e-19
C1074 ringtest_0.x4._15_ ringtest_0.x4._20_ 0.093509f
C1075 ringtest_0.x4._16_ a_21233_5340# 0.001516f
C1076 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP2 2.65608f
C1077 ringtest_0.x4._18_ a_24536_6699# 5.4e-20
C1078 ringtest_0.x4.net10 a_25977_4220# 0.158335f
C1079 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 7.08e-21
C1080 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.025028f
C1081 muxtest_0.R1R2 ua[3] 0.017912f
C1082 ringtest_0.x4.net8 a_24527_5340# 0.031957f
C1083 a_23879_6940# a_24465_6800# 0.013455f
C1084 ringtest_0.x4._11_ a_22097_5334# 0.017838f
C1085 a_27303_4246# VDPWR 0.283149f
C1086 ringtest_0.x3.x1.nSEL1 a_16707_12151# 4.08e-19
C1087 ringtest_0.x4._11_ ringtest_0.x4._16_ 0.223435f
C1088 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN2 0.209956f
C1089 a_22373_5156# a_22499_4790# 0.006169f
C1090 a_15575_12017# ringtest_0.x3.x2.GN1 0.12869f
C1091 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net8 8.45e-19
C1092 ringtest_0.x4._11_ a_22695_8304# 0.002858f
C1093 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A a_15575_12017# 6.58e-22
C1094 ringtest_0.x4.clknet_1_1__leaf_clk a_27065_5334# 1.84e-19
C1095 muxtest_0.x2.x2.GN4 VDPWR 1.23441f
C1096 ringtest_0.x4.net6 a_24361_5340# 0.0618f
C1097 a_21007_3867# ringtest_0.x4.counter[1] 0.057818f
C1098 ringtest_0.x4._22_ a_25149_4220# 0.106132f
C1099 a_24361_5340# a_24895_4790# 0.003047f
C1100 a_24527_5340# a_24729_4790# 0.003672f
C1101 muxtest_0.x1.x3.GN2 muxtest_0.R2R3 3.99837f
C1102 ringtest_0.x4.net3 a_21375_3867# 0.233128f
C1103 ringtest_0.x4.clknet_1_0__leaf_clk a_22228_8598# 0.002447f
C1104 a_24329_6640# ringtest_0.x4._22_ 1.01e-19
C1105 muxtest_0.x1.x3.GN2 ui_in[1] 0.108644f
C1106 ringtest_0.x4._03_ VDPWR 0.393273f
C1107 a_24536_6699# a_24763_6143# 3.7e-19
C1108 a_22265_5308# a_22116_4902# 0.001344f
C1109 ringtest_0.x4.net9 a_25593_5156# 0.031858f
C1110 a_22097_5334# a_21675_4790# 0.003824f
C1111 a_21672_5334# a_21948_5156# 4.47e-19
C1112 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR 0.638508f
C1113 ringtest_0.x4.counter[5] ua[1] 3.21e-19
C1114 ringtest_0.x4.clknet_0_clk a_24729_4790# 1.17e-21
C1115 ringtest_0.x4._00_ ringtest_0.x4._01_ 0.014628f
C1116 a_25925_6788# a_26201_6788# 0.00119f
C1117 m2_11882_23495# ui_in[4] 0.183786f
C1118 ringtest_0.x4._16_ a_21675_4790# 2.51e-21
C1119 ringtest_0.x3.x1.nSEL1 m2_15612_11606# 0.00815f
C1120 a_22765_5308# a_22983_5654# 0.007234f
C1121 a_26201_5340# a_26808_5308# 0.141453f
C1122 ringtest_0.x3.x1.nSEL1 ui_in[3] 0.168464f
C1123 ringtest_0.x4._15_ a_26569_6422# 0.001697f
C1124 a_23770_5308# VDPWR 0.17068f
C1125 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN2 7.45e-19
C1126 a_24045_6654# a_24264_6788# 0.006169f
C1127 ringtest_0.x4._16_ a_23899_5654# 0.001343f
C1128 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN1 0.034842f
C1129 ringtest_0.x4.net7 a_25593_5156# 0.040127f
C1130 ringtest_0.x4._03_ a_23467_4584# 5.07e-20
C1131 ringtest_0.x4.counter[8] VDPWR 0.228646f
C1132 a_12473_23980# muxtest_0.x2.x2.GP1 2.33e-21
C1133 a_24536_6699# ringtest_0.x4.clknet_1_1__leaf_clk 4.65e-20
C1134 a_21939_8054# VDPWR 3.14e-19
C1135 ringtest_0.x4.net4 a_23151_5334# 6.79e-19
C1136 ringtest_0.x4._22_ a_24545_5878# 9.75e-19
C1137 ringtest_0.x3.x2.GN3 a_16707_12151# 0.001073f
C1138 ringtest_0.x3.x2.GN2 a_17405_12123# 8.14e-21
C1139 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN4 0.001072f
C1140 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GN3 0.067463f
C1141 a_12297_23648# a_12473_23980# 0.185422f
C1142 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP3 0.005595f
C1143 a_21785_5878# a_22097_5334# 0.001393f
C1144 a_24699_6200# ringtest_0.x4._07_ 0.096566f
C1145 ringtest_0.x4._04_ a_22265_5308# 0.008333f
C1146 a_22074_4790# ringtest_0.x4.net5 3e-19
C1147 a_25364_5878# ringtest_0.x4._22_ 8.12e-19
C1148 ringtest_0.x4._14_ a_22295_3867# 4.42e-19
C1149 a_25225_5334# a_25149_4220# 3.32e-21
C1150 muxtest_0.x2.nselect2 ua[3] 0.005153f
C1151 a_21785_5878# ringtest_0.x4._16_ 6.86e-20
C1152 ringtest_0.x4.clknet_1_0__leaf_clk a_22265_5308# 0.002373f
C1153 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A a_16203_12091# 2.34e-20
C1154 a_26640_5334# a_26640_5156# 0.013839f
C1155 a_26367_5340# a_27065_5156# 1.3e-19
C1156 a_27065_5334# a_26367_4790# 1.3e-19
C1157 a_25055_3867# ringtest_0.x4.counter[6] 4.98e-19
C1158 ringtest_0.x4._11_ a_22649_6244# 0.043928f
C1159 ringtest_0.x4.net9 a_25441_4612# 6.97e-19
C1160 a_21951_5878# a_24070_5852# 8.39e-21
C1161 ringtest_0.x4._17_ a_23993_5654# 3.09e-20
C1162 a_22052_9116# ui_in[5] 1.46e-21
C1163 ringtest_0.x4._05_ a_24527_5340# 2.65e-21
C1164 ui_in[6] uio_in[0] 0.001316f
C1165 muxtest_0.x1.x3.GP1 muxtest_0.R4R5 0.123828f
C1166 ringtest_0.x4._11_ a_26201_6788# 0.005861f
C1167 ringtest_0.x4.clknet_0_clk a_26749_6422# 1.5e-20
C1168 muxtest_0.x2.x2.GP3 m3_13302_19985# 0.002824f
C1169 ringtest_0.x4._13_ a_21591_6128# 0.01129f
C1170 ringtest_0.ring_out a_17377_14114# 0.105448f
C1171 muxtest_0.x1.x3.GN3 muxtest_0.R7R8 0.129382f
C1172 ringtest_0.x4.net1 a_21939_8054# 0.002601f
C1173 ringtest_0.x4.clknet_0_clk ringtest_0.x4._05_ 0.067252f
C1174 a_22052_9116# ringtest_0.x4._12_ 5.69e-20
C1175 ringtest_0.x4._07_ a_23809_4790# 1.81e-20
C1176 a_17405_12123# ui_in[3] 1.4e-19
C1177 ringtest_0.x3.x2.GN3 ui_in[3] 0.254198f
C1178 ringtest_0.x4.net8 a_25168_5156# 0.001808f
C1179 ringtest_0.x4._23_ a_26627_4246# 0.04546f
C1180 ringtest_0.x4.net7 a_25441_4612# 0.006602f
C1181 ringtest_0.x4.net6 ringtest_0.x4._08_ 5.42e-20
C1182 ringtest_0.drv_out a_25421_6641# 0.012863f
C1183 ringtest_0.x4._11_ a_23467_4818# 0.003027f
C1184 ringtest_0.x4._17_ ringtest_0.x4._04_ 6.62e-21
C1185 a_26367_4790# a_26627_4246# 0.008374f
C1186 ringtest_0.x4.net10 ringtest_0.x4.counter[9] 0.092658f
C1187 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP3 0.031766f
C1188 a_21233_5340# a_21587_5334# 0.062224f
C1189 a_22392_5990# a_22541_5058# 8.5e-21
C1190 a_21951_5878# a_22373_5156# 0.001133f
C1191 a_26640_5156# a_26735_5156# 0.007724f
C1192 a_22224_6244# a_21948_5156# 9.19e-21
C1193 a_26367_4790# a_27149_5156# 6.32e-19
C1194 a_23899_5334# ringtest_0.x4.counter[4] 4.47e-20
C1195 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._17_ 3.38e-20
C1196 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ui_in[4] 4.1e-20
C1197 ringtest_0.x4.net10 a_27491_4566# 0.002502f
C1198 ringtest_0.x4.clknet_1_1__leaf_clk a_25294_4790# 4.82e-19
C1199 ringtest_0.x4.net6 a_25336_4902# 6.78e-21
C1200 ringtest_0.x4._11_ a_21587_5334# 2.52e-19
C1201 ringtest_0.x4._21_ a_23770_5308# 0.005326f
C1202 a_12849_23648# muxtest_0.x2.x2.GN4 6.84e-19
C1203 a_25364_5878# a_25225_5334# 5.73e-19
C1204 muxtest_0.R3R4 muxtest_0.x2.x2.GP1 0.011522f
C1205 a_13025_23980# muxtest_0.x2.x2.GN2 5.62e-20
C1206 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.001676f
C1207 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 1.11e-20
C1208 a_24895_4790# a_25336_4902# 0.110715f
C1209 a_24729_4790# a_25168_5156# 0.273138f
C1210 a_19114_31955# ui_in[0] 0.246193f
C1211 a_24712_6422# VDPWR 0.004407f
C1212 ringtest_0.counter3 ringtest_0.x4._16_ 1.05e-19
C1213 ringtest_0.x4.net4 a_22265_5308# 0.110738f
C1214 ringtest_0.x4.counter[5] ringtest_0.x4.counter[6] 0.070133f
C1215 ringtest_0.x4._15_ a_26640_5334# 0.001174f
C1216 ringtest_0.x3.x1.nSEL0 a_16755_12091# 1.21e-20
C1217 ringtest_0.x4.net3 a_21233_5340# 0.023332f
C1218 ringtest_0.x4._22_ a_26913_4566# 3.67e-19
C1219 ringtest_0.x4.net6 VDPWR 3.11824f
C1220 muxtest_0.x1.x4.A muxtest_0.R2R3 4.52053f
C1221 ringtest_0.x4._04_ a_22817_6146# 0.003723f
C1222 ringtest_0.x4.net10 a_27149_5334# 3.67e-19
C1223 a_21785_5878# a_22649_6244# 0.030894f
C1224 a_24895_4790# VDPWR 0.323392f
C1225 ringtest_0.x4.net3 ringtest_0.x4._11_ 0.005186f
C1226 ringtest_0.x4._18_ a_22765_5308# 0.002375f
C1227 muxtest_0.x1.x3.GP2 muxtest_0.R7R8 0.131352f
C1228 ringtest_0.x4._11_ a_27273_4220# 2.01e-20
C1229 a_23879_6940# a_23770_5308# 4.81e-21
C1230 ringtest_0.x4._19_ ringtest_0.x4._22_ 7e-20
C1231 ringtest_0.x4.clknet_1_0__leaf_clk a_22817_6146# 1.77e-20
C1232 muxtest_0.x1.x3.GN3 muxtest_0.R5R6 4.12612f
C1233 a_21845_9116# ringtest_0.x4._11_ 8.58e-21
C1234 ringtest_0.x4._11_ a_26766_4790# 4.03e-21
C1235 a_25364_5878# a_26640_5156# 6.58e-20
C1236 a_27169_6641# ringtest_0.x4._08_ 0.109717f
C1237 a_19666_31955# ui_in[1] 0.261734f
C1238 a_24361_5340# a_24895_5334# 0.001632f
C1239 ringtest_0.x4._11_ a_24465_6800# 5.19e-20
C1240 a_24045_6654# a_24070_5852# 0.006438f
C1241 a_21465_9294# a_21561_8830# 6.79e-19
C1242 a_21561_9116# a_21465_8830# 6.79e-19
C1243 a_23949_6654# a_24004_6128# 3.4e-19
C1244 muxtest_0.x1.x5.GN muxtest_0.x1.x4.A 4.14763f
C1245 a_21055_5334# VDPWR 0.006911f
C1246 muxtest_0.x1.x3.GN3 VDPWR 0.766397f
C1247 ringtest_0.x4._15_ a_25149_4220# 1.2e-20
C1248 ringtest_0.x4._19_ a_23619_6788# 8.17e-20
C1249 ringtest_0.x4.net6 ringtest_0.x4._25_ 2.22e-20
C1250 ringtest_0.x4._17_ ringtest_0.x4.net4 9.08e-20
C1251 ringtest_0.x4.net2 a_21507_9686# 0.00492f
C1252 muxtest_0.x1.x5.GN a_19666_31955# 3.51e-19
C1253 a_21509_4790# a_22295_3867# 8.97e-21
C1254 a_24329_6640# ringtest_0.x4._15_ 3.85e-20
C1255 ringtest_0.x4._14_ ringtest_0.x4._02_ 0.166596f
C1256 muxtest_0.x1.x3.GP1 ui_in[2] 5.64e-19
C1257 ringtest_0.x4.net3 a_21675_4790# 0.00115f
C1258 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GP1 6.21e-20
C1259 ringtest_0.x4._16_ a_22775_5878# 4.87e-20
C1260 a_16579_11759# ringtest_0.x3.x2.GP3 0.00144f
C1261 ringtest_0.x4.net9 ringtest_0.x4._22_ 0.369389f
C1262 a_13501_23906# ui_in[4] 0.125445f
C1263 ui_in[4] ua[2] 0.936267f
C1264 muxtest_0.x2.x1.nSEL0 a_12297_23648# 0.03096f
C1265 a_21951_5878# a_21399_5340# 5.5e-20
C1266 muxtest_0.x1.x1.nSEL0 ui_in[0] 0.325407f
C1267 a_22939_4584# VDPWR 3.83e-21
C1268 a_24699_6200# ringtest_0.x4._06_ 0.003245f
C1269 ringtest_0.x4._16_ a_23399_3867# 3.59e-21
C1270 a_27169_6641# VDPWR 0.28996f
C1271 a_21981_9142# VDPWR 0.211499f
C1272 ringtest_0.x4._11_ a_22733_6244# 0.002344f
C1273 a_22111_10993# VDPWR 0.305606f
C1274 ringtest_0.x4.clknet_1_1__leaf_clk a_22765_5308# 1.5e-19
C1275 ringtest_0.x4.net4 a_22817_6146# 7.5e-19
C1276 muxtest_0.x1.x3.GP2 muxtest_0.R5R6 0.312699f
C1277 muxtest_0.x2.x2.GP3 ua[0] 0.050476f
C1278 ringtest_0.x4.net7 ringtest_0.x4._22_ 0.179589f
C1279 ringtest_0.x4.net3 a_21785_5878# 1.48e-19
C1280 ringtest_0.x3.nselect2 VDPWR 1.23654f
C1281 ringtest_0.x4.net6 ringtest_0.x4._21_ 0.083542f
C1282 ringtest_0.x4._15_ a_25364_5878# 0.047247f
C1283 a_21561_8830# a_21981_8976# 0.036838f
C1284 a_21845_8816# a_22052_8875# 0.260055f
C1285 a_21465_8830# ringtest_0.x4._01_ 1.56e-19
C1286 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B a_17377_14114# 0.110771f
C1287 ringtest_0.x4._17_ a_23837_5878# 0.060488f
C1288 ringtest_0.x4._23_ a_26721_4246# 0.038842f
C1289 ringtest_0.x4._17_ ringtest_0.x4._22_ 1.76e-19
C1290 a_22390_4566# a_22486_4246# 0.002032f
C1291 ringtest_0.x4._11_ a_26201_4790# 0.012822f
C1292 a_11845_23906# m2_11882_23495# 0.01297f
C1293 ringtest_0.x4._14_ a_22116_4902# 1.1e-19
C1294 ringtest_0.x4.clknet_1_0__leaf_clk a_22201_9142# 0.002297f
C1295 ringtest_0.x3.x2.GP1 ringtest_0.counter3 5.62e-21
C1296 muxtest_0.x1.x3.GP2 VDPWR 3.26769f
C1297 a_27169_6641# ringtest_0.x4._25_ 0.227897f
C1298 a_26367_4790# a_26721_4246# 1.65e-19
C1299 a_21845_9116# a_22399_9142# 0.062224f
C1300 ringtest_0.x4.net2 a_21852_8720# 8.79e-19
C1301 ringtest_0.x4._18_ ringtest_0.x4.net8 0.01511f
C1302 a_22052_9116# a_22228_9508# 0.007724f
C1303 a_21852_9416# ringtest_0.x4.clknet_1_0__leaf_clk 0.470509f
C1304 a_21981_9142# a_21803_9508# 9.73e-19
C1305 ringtest_0.counter7 ringtest_0.x4.net8 6.32e-19
C1306 ringtest_0.x4.net7 a_23619_6788# 5.91e-19
C1307 ringtest_0.x4._11_ a_22457_5156# 0.002515f
C1308 a_24070_5852# a_23809_4790# 7.94e-19
C1309 ringtest_0.x4.net1 a_21981_9142# 0.002441f
C1310 a_24361_5340# a_24527_5340# 0.961627f
C1311 ringtest_0.drv_out ringtest_0.x3.x2.GN1 3.11e-19
C1312 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 2.86851f
C1313 ringtest_0.x4._17_ a_23619_6788# 7.93e-19
C1314 a_22111_10993# ringtest_0.x4.net1 0.10983f
C1315 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ui_in[4] 0.008686f
C1316 ringtest_0.x4.net9 a_25225_5334# 0.002503f
C1317 a_23932_6128# VDPWR 0.011634f
C1318 a_25761_5058# a_26201_4790# 0.001745f
C1319 ringtest_0.x4.clknet_0_clk a_24361_5340# 0.009291f
C1320 ringtest_0.x4._15_ a_24317_4942# 2.8e-19
C1321 a_23879_6940# ringtest_0.x4.net6 8.49e-19
C1322 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 1.99e-20
C1323 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.025028f
C1324 ua[0] ui_in[6] 0.619336f
C1325 a_23949_6654# ringtest_0.x4._20_ 1.63e-20
C1326 a_23809_4790# a_23891_4790# 0.005167f
C1327 a_22817_6146# a_23837_5878# 3.28e-20
C1328 ringtest_0.x4._04_ ringtest_0.x4._14_ 4.63e-22
C1329 a_22649_6244# a_22775_5878# 0.006169f
C1330 a_21395_6940# ringtest_0.x4.clknet_0_clk 0.317755f
C1331 a_15575_12017# ui_in[4] 0.02803f
C1332 ringtest_0.x4._24_ a_26201_5340# 0.031818f
C1333 ringtest_0.x4.net8 a_24763_6143# 0.003744f
C1334 a_21948_5156# a_21863_4790# 0.037333f
C1335 a_21675_4790# a_22457_5156# 3.14e-19
C1336 ringtest_0.x3.x1.nSEL1 a_16027_11759# 0.073392f
C1337 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A a_16755_12091# 9.97e-21
C1338 ringtest_0.x4.net7 a_25225_5334# 0.054488f
C1339 a_22265_5308# a_22021_4220# 2.52e-20
C1340 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._14_ 0.088295f
C1341 muxtest_0.R7R8 muxtest_0.R3R4 5.65992f
C1342 ringtest_0.x4._12_ a_21395_6940# 4.42e-19
C1343 a_12473_23980# VDPWR 0.193262f
C1344 ringtest_0.x4.net3 ringtest_0.counter3 6.21e-20
C1345 ringtest_0.x4._17_ a_25225_5334# 8.73e-21
C1346 ringtest_0.x4.clknet_1_0__leaf_clk a_22319_6244# 4.17e-19
C1347 muxtest_0.x1.x3.GN4 ua[3] 0.014367f
C1348 a_21132_8918# ringtest_0.x4._12_ 0.001776f
C1349 a_21852_8720# a_22399_8976# 0.099725f
C1350 a_21465_8830# a_21785_8054# 3.66e-19
C1351 a_22052_8875# a_22201_8964# 0.005525f
C1352 ringtest_0.x4.net5 VDPWR 0.923749f
C1353 ringtest_0.x4.net9 a_26640_5156# 0.023502f
C1354 ringtest_0.x3.x2.GP3 m3_17032_8096# 0.002824f
C1355 a_12977_24040# ui_in[3] 0.001558f
C1356 a_24895_5334# VDPWR 0.004219f
C1357 muxtest_0.x1.x3.GN4 a_20492_32319# 0.001562f
C1358 muxtest_0.x2.x2.GN2 ui_in[3] 0.11443f
C1359 ringtest_0.x4._02_ a_21509_4790# 3.71e-19
C1360 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net8 0.073766f
C1361 ringtest_0.x4.net2 a_22399_8976# 1.01e-21
C1362 a_21233_5340# ringtest_0.x4._03_ 0.001727f
C1363 ringtest_0.x4._15_ a_26913_4566# 0.001637f
C1364 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP3 0.075682f
C1365 muxtest_0.R2R3 ua[0] 2.39e-19
C1366 ringtest_0.counter7 ringtest_0.x4.counter[1] 0.003115f
C1367 a_24004_6128# ringtest_0.x4._20_ 4.3e-20
C1368 a_19842_32287# muxtest_0.x1.x3.GN4 0.003645f
C1369 ringtest_0.x4._24_ a_27233_5058# 0.009415f
C1370 ringtest_0.x4._00_ a_21845_9116# 0.118744f
C1371 ringtest_0.x4._11_ ringtest_0.x4._03_ 0.00174f
C1372 ringtest_0.x4._19_ ringtest_0.x4._15_ 6.2e-22
C1373 ringtest_0.x4.net7 a_26640_5156# 4.39e-19
C1374 ringtest_0.x4._02_ a_22765_5308# 7.66e-20
C1375 ringtest_0.x4.net5 a_23467_4584# 0.001706f
C1376 ringtest_0.x4.clknet_1_0__leaf_clk a_22043_5156# 5.04e-19
C1377 ringtest_0.counter7 ringtest_0.x4.net11 1.31e-19
C1378 ringtest_0.x4.clknet_1_1__leaf_clk a_24729_4790# 0.319108f
C1379 ringtest_0.x4.net10 a_27273_4220# 0.104575f
C1380 ringtest_0.x4._18_ ringtest_0.x4._05_ 1.11e-19
C1381 ringtest_0.x4.net8 a_24800_5334# 0.003635f
C1382 ringtest_0.x4._20_ a_23963_4790# 0.001506f
C1383 muxtest_0.x1.x3.GN2 ui_in[0] 0.114399f
C1384 ringtest_0.x4._11_ a_23770_5308# 0.058411f
C1385 a_21007_3867# VDPWR 0.25802f
C1386 ringtest_0.x3.x2.GN4 ui_in[4] 0.059808f
C1387 a_16027_11759# ringtest_0.x3.x2.GN3 6.68e-19
C1388 ringtest_0.x4._08_ a_24527_5340# 8.29e-20
C1389 a_16203_12091# ringtest_0.x3.x2.GN1 1.46e-19
C1390 ringtest_0.x4._13_ ringtest_0.x4._02_ 0.053355f
C1391 a_23381_4818# ringtest_0.x4._20_ 3.41e-19
C1392 ringtest_0.x4.net4 ringtest_0.x4._14_ 0.209869f
C1393 ringtest_0.x4._11_ a_21939_8054# 2.12e-19
C1394 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.173286f
C1395 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x1.nSEL0 1.14e-19
C1396 ringtest_0.x4.net6 a_24968_5308# 0.012704f
C1397 ringtest_0.x4._03_ a_21675_4790# 0.260627f
C1398 a_21509_4790# a_22116_4902# 0.141453f
C1399 muxtest_0.x1.x4.A ui_in[4] 0.034362f
C1400 ringtest_0.x4._15_ a_22265_5308# 1.37e-19
C1401 ringtest_0.x4._22_ a_26627_4246# 0.140356f
C1402 a_24968_5308# a_24895_4790# 0.001607f
C1403 a_24361_5340# a_25168_5156# 4.58e-19
C1404 a_24800_5334# a_24729_4790# 2.14e-19
C1405 a_24527_5340# a_25336_4902# 6.74e-19
C1406 ringtest_0.x4._15_ ringtest_0.x4.net9 0.08758f
C1407 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._10_ 0.006812f
C1408 muxtest_0.R3R4 VDPWR 3.2635f
C1409 ringtest_0.x4._16_ a_25083_4790# 1.98e-21
C1410 ringtest_0.x4._23_ ringtest_0.x4.net8 0.011201f
C1411 ringtest_0.x4._05_ a_24763_6143# 2.43e-19
C1412 a_22097_5334# a_21948_5156# 0.001152f
C1413 a_22265_5308# a_22541_5058# 0.007214f
C1414 ringtest_0.x4.net8 a_26367_4790# 1.04e-19
C1415 ringtest_0.x4.clknet_0_clk a_25336_4902# 8.09e-19
C1416 ringtest_0.x4._16_ a_21948_5156# 2.79e-19
C1417 ringtest_0.x4._21_ ringtest_0.x4.net5 2.83e-22
C1418 a_21672_5334# a_21767_5334# 0.007724f
C1419 a_23770_5308# a_23899_5654# 0.010132f
C1420 a_21840_5308# a_22181_5334# 9.73e-19
C1421 a_26201_5340# a_27233_5308# 0.048748f
C1422 a_26367_5340# a_26640_5334# 0.078545f
C1423 a_24527_5340# VDPWR 0.300379f
C1424 ringtest_0.x4.net7 ringtest_0.x4._15_ 0.590844f
C1425 ringtest_0.x4.clknet_1_1__leaf_clk a_26749_6422# 3.65e-19
C1426 ringtest_0.x4.net6 a_25925_6788# 0.157729f
C1427 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net11 1.82e-20
C1428 VDPWR ui_in[5] 0.255037f
C1429 ringtest_0.x4._04_ a_21509_4790# 2.08e-19
C1430 a_21785_5878# ringtest_0.x4._03_ 4.31e-20
C1431 ringtest_0.x4.net7 a_25263_5156# 5.23e-19
C1432 ringtest_0.x4._23_ a_24729_4790# 3.56e-21
C1433 a_13025_23980# muxtest_0.x2.x2.GP1 2.87e-20
C1434 ringtest_0.x4._17_ ringtest_0.x4._15_ 0.083602f
C1435 ringtest_0.x4._05_ ringtest_0.x4.clknet_1_1__leaf_clk 0.143201f
C1436 ringtest_0.x4.clknet_0_clk VDPWR 2.53166f
C1437 muxtest_0.x2.x2.GP2 ui_in[4] 4.34e-19
C1438 a_24729_4790# a_26367_4790# 8.05e-21
C1439 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP1 8.08e-19
C1440 ringtest_0.x4.clknet_1_0__leaf_clk a_21509_4790# 0.293401f
C1441 ua[3] ua[4] 0.008019f
C1442 ringtest_0.counter7 ringtest_0.x4._09_ 5.27e-21
C1443 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 5.48e-19
C1444 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y 0.001676f
C1445 muxtest_0.x2.x1.nSEL1 a_12019_24012# 0.00175f
C1446 a_12473_23980# a_12849_23648# 3.02e-19
C1447 ringtest_0.x4._12_ VDPWR 0.307826f
C1448 ringtest_0.x4._04_ a_22765_5308# 0.171873f
C1449 ringtest_0.x4.counter[9] ua[0] 0.004138f
C1450 ringtest_0.x4.net10 a_26201_4790# 0.001924f
C1451 a_27191_5712# ringtest_0.x4._09_ 1.66e-19
C1452 ringtest_0.x4.net7 a_24926_5712# 2.79e-19
C1453 ringtest_0.x4.clknet_1_0__leaf_clk a_22765_5308# 1.95e-19
C1454 a_27233_5308# a_27233_5058# 0.026048f
C1455 ringtest_0.x4._05_ a_24800_5334# 6.05e-21
C1456 ringtest_0.x4.net6 a_21233_5340# 1.88e-19
C1457 ringtest_0.x4._13_ ringtest_0.x4._04_ 1.41e-19
C1458 ringtest_0.x4.clknet_1_0__leaf_clk a_21867_8054# 2.61e-19
C1459 ringtest_0.x4.net1 ui_in[5] 0.067291f
C1460 a_26555_5334# ringtest_0.x4.net10 6.3e-20
C1461 muxtest_0.x2.x1.nSEL0 VDPWR 0.523833f
C1462 ringtest_0.x4._22_ a_25294_4790# 6.82e-19
C1463 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A 0.429924f
C1464 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._13_ 0.02176f
C1465 ringtest_0.x4.counter[6] ua[1] 3.21e-19
C1466 ringtest_0.x4._11_ ringtest_0.x4.net6 2.01574f
C1467 ringtest_0.x3.x2.GN1 m3_17036_9140# 6.03e-20
C1468 ringtest_0.x4.net1 ringtest_0.x4._12_ 0.312817f
C1469 ringtest_0.x4.net7 a_26173_4612# 6.49e-19
C1470 ringtest_0.x4.net8 a_25593_5156# 0.007067f
C1471 ringtest_0.x4._11_ a_24895_4790# 0.042209f
C1472 ringtest_0.x4._23_ a_26749_6422# 0.007723f
C1473 ringtest_0.x4._23_ ringtest_0.x4.net11 0.257634f
C1474 a_26640_5156# a_26627_4246# 2.47e-19
C1475 a_19114_31955# muxtest_0.x1.x3.GN3 6.68e-19
C1476 a_21233_5340# a_21055_5334# 5.87e-19
C1477 a_26749_6422# a_26367_4790# 3.03e-21
C1478 muxtest_0.R4R5 ui_in[2] 6.76e-20
C1479 a_26808_4902# a_26766_4790# 4.62e-19
C1480 a_22224_6244# a_22373_5156# 1.06e-19
C1481 a_26367_4790# ringtest_0.x4.net11 2.58e-19
C1482 a_18662_32213# VDPWR 0.213938f
C1483 ringtest_0.x4._05_ ringtest_0.x4._23_ 9.36e-20
C1484 a_21399_5340# a_21672_5334# 0.078737f
C1485 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._09_ 0.003413f
C1486 ringtest_0.x4.net4 a_21509_4790# 0.008383f
C1487 ringtest_0.x4.net10 a_27303_4246# 0.001384f
C1488 ringtest_0.x4.net6 a_25761_5058# 3.96e-21
C1489 m2_18699_31802# VDPWR 0.140918f
C1490 a_13501_23906# muxtest_0.x2.x2.GN4 0.134079f
C1491 muxtest_0.x2.x2.GN2 a_12425_24040# 0.002418f
C1492 muxtest_0.x2.x2.GN4 ua[2] 0.446579f
C1493 a_25364_5878# a_26367_5340# 0.008007f
C1494 ringtest_0.x4._21_ a_24527_5340# 0.002388f
C1495 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN2 0.065156f
C1496 a_23949_6654# a_24329_6640# 0.048635f
C1497 a_22245_8054# VDPWR 0.292813f
C1498 a_24895_4790# a_25761_5058# 0.034054f
C1499 a_24729_4790# a_25593_5156# 0.032244f
C1500 a_25336_4902# a_25168_5156# 0.239923f
C1501 a_19666_31955# ui_in[0] 0.086357f
C1502 ringtest_0.x4.net4 a_22765_5308# 0.005124f
C1503 muxtest_0.x2.x1.nSEL1 ui_in[4] 0.275874f
C1504 muxtest_0.x1.x3.GP3 muxtest_0.R1R2 4.25867f
C1505 ringtest_0.x3.x1.nSEL0 a_16155_12151# 2.51e-19
C1506 ringtest_0.x4.clknet_0_clk ringtest_0.x4._21_ 4.86e-19
C1507 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN1 0.004375f
C1508 ringtest_0.x4._15_ a_27065_5334# 2.78e-19
C1509 ringtest_0.x4._22_ a_26721_4246# 0.063386f
C1510 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 5.04e-19
C1511 ringtest_0.x4._14_ a_22021_4220# 0.134293f
C1512 ringtest_0.x4._04_ ringtest_0.x4.net8 7.52e-21
C1513 muxtest_0.x1.x3.GP1 muxtest_0.R2R3 0.127193f
C1514 a_25168_5156# VDPWR 0.256044f
C1515 a_21007_3867# a_21375_3867# 2.48e-19
C1516 ringtest_0.x4._18_ a_24361_5340# 5.99e-21
C1517 ringtest_0.x4.net8 a_25441_4612# 0.001229f
C1518 ringtest_0.x4._11_ a_22939_4584# 8.14e-19
C1519 a_23879_6940# a_24527_5340# 4.98e-20
C1520 ringtest_0.x4.net4 ringtest_0.x4._13_ 0.050083f
C1521 muxtest_0.x1.x3.GP1 ui_in[1] 8.43e-19
C1522 muxtest_0.x1.x3.GP2 muxtest_0.x1.x5.A 0.350698f
C1523 ringtest_0.x4.net3 a_21465_8830# 0.115857f
C1524 a_24336_6544# ringtest_0.x4._06_ 1.63e-21
C1525 a_20318_32213# ui_in[1] 0.125445f
C1526 ringtest_0.x4.net1 a_22245_8054# 4.64e-19
C1527 ringtest_0.x4.clknet_0_clk a_23349_6422# 2.32e-20
C1528 a_25225_5334# a_25351_5712# 0.006169f
C1529 a_24527_5340# a_25309_5334# 3.14e-19
C1530 a_21425_9686# ringtest_0.x4._12_ 1.27e-21
C1531 a_21852_9416# a_21561_8830# 1.53e-19
C1532 a_21561_9116# a_21845_8816# 9.64e-20
C1533 ringtest_0.x4.clknet_0_clk a_23879_6940# 1.74729f
C1534 a_24329_6640# a_24004_6128# 0.001895f
C1535 ringtest_0.x4.net6 a_21785_5878# 0.006287f
C1536 a_22983_5654# VDPWR 0.001324f
C1537 ringtest_0.x4._15_ a_26627_4246# 0.087822f
C1538 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP1 0.041018f
C1539 ringtest_0.x4._19_ a_24685_6788# 2.79e-19
C1540 ringtest_0.x4.net10 ringtest_0.x4.counter[8] 0.009948f
C1541 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN3 4.01e-20
C1542 ringtest_0.x4.net2 a_21465_9294# 0.092265f
C1543 ringtest_0.drv_out ui_in[4] 1.17e-19
C1544 ringtest_0.x4._23_ ringtest_0.x4._09_ 0.130147f
C1545 muxtest_0.x1.x5.GN a_20318_32213# 1.19e-19
C1546 ringtest_0.ring_out a_16579_11759# 5.47e-20
C1547 ringtest_0.x4._09_ a_26367_4790# 0.413296f
C1548 a_24536_6699# ringtest_0.x4._15_ 1.61e-21
C1549 a_26201_4790# a_26808_4902# 0.141453f
C1550 ui_in[6] ui_in[7] 0.03107f
C1551 ringtest_0.x4.net3 a_21948_5156# 3.32e-20
C1552 a_24763_6143# a_24361_5340# 0.004179f
C1553 a_13675_24012# ui_in[4] 8.84e-19
C1554 ringtest_0.x4._16_ ringtest_0.x4._07_ 0.003808f
C1555 ringtest_0.x4._06_ a_24986_5878# 6.53e-20
C1556 muxtest_0.x2.x2.GN3 ui_in[4] 0.273874f
C1557 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y 0.174714f
C1558 a_21591_6128# VDPWR 0.006535f
C1559 ringtest_0.x4._23_ a_26766_5712# 9.59e-19
C1560 muxtest_0.x2.x1.nSEL0 a_12849_23648# 1.91e-20
C1561 a_24004_6128# a_24545_5878# 4.72e-19
C1562 a_21951_5878# a_21672_5334# 0.001124f
C1563 ringtest_0.x4.clknet_1_0__leaf_clk a_21798_5712# 0.001807f
C1564 a_22486_4246# VDPWR 0.012117f
C1565 a_22228_9508# VDPWR 0.005789f
C1566 ringtest_0.x4.net9 a_25975_3867# 7.77e-19
C1567 ringtest_0.x4._11_ a_23932_6128# 0.002546f
C1568 ringtest_0.x4._15_ ringtest_0.x4._14_ 1.65e-19
C1569 ringtest_0.x4.clknet_1_1__leaf_clk a_24361_5340# 0.670964f
C1570 ringtest_0.x4.net4 ringtest_0.x4.net8 0.001699f
C1571 a_21852_8720# a_21981_8976# 0.124967f
C1572 a_21845_8816# ringtest_0.x4._01_ 0.092611f
C1573 ringtest_0.x4._24_ a_26895_3867# 0.00116f
C1574 muxtest_0.x2.x2.GP1 ui_in[3] 9.65e-19
C1575 ringtest_0.counter3 ringtest_0.x4.net6 1.1e-21
C1576 muxtest_0.x1.x3.GN1 muxtest_0.R6R7 0.254376f
C1577 ringtest_0.x4.net7 a_25975_3867# 4.41e-19
C1578 a_25977_4220# a_26269_4612# 0.001675f
C1579 ringtest_0.x4._23_ a_27659_4246# 0.009249f
C1580 ringtest_0.x4._14_ a_22541_5058# 1.14e-20
C1581 a_26640_5156# a_26721_4246# 7.6e-20
C1582 a_22052_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.040993f
C1583 a_12297_23648# ui_in[3] 0.246189f
C1584 ringtest_0.x4.net2 a_21981_8976# 8.2e-21
C1585 a_21981_9142# a_22399_9142# 3.39e-19
C1586 ringtest_0.x4.net7 a_24685_6788# 0.002551f
C1587 ringtest_0.drv_out ringtest_0.x3.x2.GP1 0.125793f
C1588 ringtest_0.x4._11_ ringtest_0.x4.net5 0.388184f
C1589 a_24004_6128# a_24317_4942# 2.49e-20
C1590 ringtest_0.x4.net1 a_22228_9508# 4.16e-19
C1591 a_24361_5340# a_24800_5334# 0.260055f
C1592 a_24527_5340# a_24968_5308# 0.110715f
C1593 ringtest_0.x4._06_ a_23899_5334# 2.02e-19
C1594 a_24070_5852# a_23899_5334# 1.06e-19
C1595 ringtest_0.x4.net9 a_26367_5340# 0.001054f
C1596 a_23949_6654# ringtest_0.x4._19_ 0.065395f
C1597 ringtest_0.counter3 a_21055_5334# 1.26e-20
C1598 ringtest_0.x4._08_ a_27191_5712# 7.43e-19
C1599 a_25593_5156# ringtest_0.x4._09_ 1.4e-19
C1600 ringtest_0.x4.clknet_0_clk a_24968_5308# 3.18e-19
C1601 a_21509_4790# a_22021_4220# 2.64e-19
C1602 ringtest_0.x4.net4 a_21798_5712# 1.81e-19
C1603 a_12977_24040# ua[3] 1.48e-19
C1604 ringtest_0.x4.net6 ringtest_0.x4.net10 1.08e-19
C1605 muxtest_0.x2.x2.GN2 ua[3] 0.234749f
C1606 ringtest_0.x4._15_ a_25351_5712# 0.00162f
C1607 ringtest_0.x4.net8 a_23837_5878# 0.057781f
C1608 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN4 0.011047f
C1609 a_16203_12091# ui_in[4] 0.254026f
C1610 ringtest_0.x4._24_ a_26808_5308# 0.015657f
C1611 ringtest_0.x4.net8 ringtest_0.x4._22_ 0.137056f
C1612 ringtest_0.x3.x1.nSEL1 a_16579_11759# 7.84e-19
C1613 a_21675_4790# ringtest_0.x4.net5 8.3e-19
C1614 a_22116_4902# a_22074_4790# 4.62e-19
C1615 ringtest_0.x4.net7 a_26367_5340# 2.99e-20
C1616 ringtest_0.x4._23_ a_24361_5340# 1.94e-21
C1617 a_21675_10006# VDPWR 5.43e-19
C1618 ringtest_0.x4._04_ a_22350_5878# 2.91e-19
C1619 muxtest_0.x1.x5.A muxtest_0.R3R4 4.07e-21
C1620 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.173286f
C1621 muxtest_0.x1.x3.GN3 a_13501_23906# 1.84e-20
C1622 a_21951_5878# a_22224_6244# 0.074434f
C1623 ringtest_0.x4.net4 ringtest_0.x4.counter[1] 3.68e-19
C1624 ringtest_0.x4._16_ a_22164_4362# 0.146025f
C1625 a_13025_23980# VDPWR 0.261817f
C1626 ringtest_0.x4._18_ VDPWR 0.686881f
C1627 ringtest_0.x4.clknet_1_0__leaf_clk a_22350_5878# 3.26e-19
C1628 ringtest_0.x4.net6 a_22775_5878# 5.88e-19
C1629 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[3] 2.42e-19
C1630 a_21845_8816# a_21785_8054# 4.35e-19
C1631 a_21981_8976# a_22399_8976# 3.39e-19
C1632 ringtest_0.x4.clknet_0_clk a_25925_6788# 1.5e-19
C1633 ringtest_0.counter7 VDPWR 2.42695f
C1634 ringtest_0.x4.net6 a_24627_6200# 4.57e-19
C1635 ringtest_0.x4.net9 a_27065_5156# 0.020729f
C1636 muxtest_0.x2.x2.GN4 m3_13302_19985# 7.07e-19
C1637 a_23529_6422# ringtest_0.x4._16_ 1.86e-20
C1638 ringtest_0.x4.net6 ringtest_0.x4.counter[4] 0.003133f
C1639 ringtest_0.x4.net4 a_22390_4566# 0.01239f
C1640 ringtest_0.x4._22_ a_24729_4790# 0.019806f
C1641 a_27191_5712# VDPWR 7.83e-19
C1642 ringtest_0.x4._15_ a_26721_4246# 0.038186f
C1643 ringtest_0.x4.net6 a_23399_3867# 3.58e-19
C1644 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN4 0.141966f
C1645 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._08_ 0.00277f
C1646 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GN3 0.175252f
C1647 ringtest_0.x4._00_ a_21981_9142# 0.005564f
C1648 a_18836_32319# VDPWR 0.001273f
C1649 ringtest_0.x4._24_ a_26555_4790# 3.3e-19
C1650 a_21785_5878# ringtest_0.x4.net5 1.51e-20
C1651 ringtest_0.x4.net7 a_27065_5156# 1.49e-19
C1652 a_22111_10993# ringtest_0.x4._00_ 4.57e-22
C1653 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP2 8.45e-19
C1654 ringtest_0.x4.net1 a_21675_10006# 0.003019f
C1655 a_23949_6654# ringtest_0.x4.net7 0.114197f
C1656 a_24763_6143# VDPWR 0.129866f
C1657 ringtest_0.x4.clknet_1_1__leaf_clk a_25336_4902# 0.046669f
C1658 ringtest_0.x4.net8 a_25225_5334# 0.00311f
C1659 ringtest_0.x4._11_ a_24527_5340# 8.46e-20
C1660 ringtest_0.x4._17_ a_23949_6654# 0.0702f
C1661 ringtest_0.x3.x2.GN1 ua[1] 0.430121f
C1662 a_22295_3867# VDPWR 0.317416f
C1663 a_22139_5878# a_21399_5340# 2.83e-19
C1664 a_16203_12091# ringtest_0.x3.x2.GP1 2.33e-21
C1665 ringtest_0.x4._06_ ringtest_0.x4._16_ 0.064563f
C1666 ringtest_0.x4._08_ a_24800_5334# 1.22e-20
C1667 muxtest_0.x2.x1.nSEL1 a_11845_23906# 0.193944f
C1668 a_16579_11759# ringtest_0.x3.x2.GN3 0.104151f
C1669 a_24070_5852# ringtest_0.x4._16_ 0.035189f
C1670 a_16755_12091# ringtest_0.x3.x2.GN1 3.78e-20
C1671 a_24317_4942# ringtest_0.x4._20_ 0.113204f
C1672 ringtest_0.x4._11_ ringtest_0.x4.clknet_0_clk 0.042991f
C1673 ringtest_0.x4._15_ a_22765_5308# 8.84e-19
C1674 muxtest_0.x1.x3.GP2 a_13501_23906# 6.46e-20
C1675 ringtest_0.x4.net6 a_25393_5308# 0.002597f
C1676 a_21509_4790# a_22541_5058# 0.048748f
C1677 ringtest_0.x4._03_ a_21948_5156# 0.010537f
C1678 ringtest_0.x4.clknet_1_1__leaf_clk VDPWR 3.34801f
C1679 ringtest_0.x4._12_ ringtest_0.x4._11_ 0.214271f
C1680 ringtest_0.x3.x2.GP2 VDPWR 1.81711f
C1681 a_22399_8976# a_22228_8598# 0.001229f
C1682 a_25393_5308# a_24895_4790# 0.002689f
C1683 ringtest_0.x4._22_ ringtest_0.x4.net11 1.96e-19
C1684 a_25225_5334# a_24729_4790# 0.004606f
C1685 muxtest_0.x1.x3.GP3 muxtest_0.R6R7 0.12263f
C1686 a_26569_6422# a_25364_5878# 0.010673f
C1687 ringtest_0.x4._05_ ringtest_0.x4._22_ 0.001519f
C1688 ringtest_0.x4._16_ a_23891_4790# 0.00109f
C1689 ringtest_0.x4.net7 a_24004_6128# 3.79e-19
C1690 a_22765_5308# a_22541_5058# 0.002391f
C1691 a_22097_5334# a_22373_5156# 5.06e-19
C1692 ringtest_0.x4._18_ ringtest_0.x4._21_ 0.005609f
C1693 ringtest_0.x4._23_ ringtest_0.x4._08_ 0.030554f
C1694 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2 3.78674f
C1695 muxtest_0.x2.x1.nSEL0 m2_11882_23495# 3.43e-19
C1696 ringtest_0.x4._16_ a_22373_5156# 6.21e-20
C1697 ringtest_0.x4._17_ a_24004_6128# 0.076419f
C1698 a_26808_5308# a_27233_5308# 1.28e-19
C1699 ringtest_0.x4._08_ a_26367_4790# 0.001269f
C1700 ringtest_0.counter7 ringtest_0.x4.counter[2] 0.003115f
C1701 ringtest_0.counter3 ringtest_0.x4.net5 0.082815f
C1702 a_26367_5340# a_27065_5334# 0.194892f
C1703 ringtest_0.ring_out ringtest_0.x3.x2.GP3 0.080819f
C1704 a_24800_5334# VDPWR 0.255475f
C1705 a_24465_6800# a_24264_6788# 4.67e-20
C1706 a_24336_6544# a_24883_6800# 0.095025f
C1707 a_24536_6699# a_24685_6788# 0.005525f
C1708 ringtest_0.x4.net4 a_22074_4790# 6.57e-19
C1709 muxtest_0.R7R8 ui_in[3] 0.025566f
C1710 a_21425_9686# a_21675_10006# 0.007234f
C1711 a_18662_32213# a_19114_31955# 0.002207f
C1712 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1 1.5157f
C1713 a_12297_23648# a_12425_24040# 0.004764f
C1714 a_12849_23648# a_13025_23980# 0.185422f
C1715 a_23349_6422# ringtest_0.x4._18_ 0.09549f
C1716 a_12297_23648# muxtest_0.x2.x2.GN1 0.012445f
C1717 ringtest_0.x4._21_ a_24763_6143# 1.69e-19
C1718 ringtest_0.x4._17_ a_23381_4818# 6.88e-22
C1719 ringtest_0.x3.x1.nSEL0 ui_in[4] 0.137394f
C1720 muxtest_0.R4R5 muxtest_0.R2R3 7.85e-20
C1721 a_27065_5334# a_27065_5156# 0.01464f
C1722 ringtest_0.x4._23_ VDPWR 1.70159f
C1723 a_21395_6940# ringtest_0.x4._04_ 0.00168f
C1724 a_21951_5878# a_22139_5878# 0.095025f
C1725 a_22817_6146# a_24004_6128# 1.25e-19
C1726 a_22245_8054# ringtest_0.x4._11_ 0.201886f
C1727 a_26367_4790# VDPWR 0.31984f
C1728 a_22295_3867# ringtest_0.x4.counter[2] 0.1107f
C1729 ringtest_0.counter3 a_21007_3867# 2.11e-19
C1730 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C1731 a_16707_12151# VDPWR 0.001127f
C1732 ringtest_0.x4.clknet_1_0__leaf_clk a_21395_6940# 1.67275f
C1733 ringtest_0.x3.x2.GN2 VDPWR 0.602894f
C1734 ringtest_0.x4._22_ ringtest_0.x4._09_ 0.009594f
C1735 muxtest_0.x2.x2.GN4 ua[0] 0.046938f
C1736 ringtest_0.x3.x2.GP1 m3_17036_9140# 5.81e-19
C1737 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._21_ 0.038033f
C1738 ringtest_0.x4._15_ ringtest_0.x4.net8 0.048599f
C1739 ringtest_0.x4.net2 ringtest_0.x4.counter[0] 0.010591f
C1740 ringtest_0.x3.x2.GN3 m3_17032_8096# 0.087318f
C1741 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP3 5.60415f
C1742 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A 0.429865f
C1743 ringtest_0.x4._24_ a_26817_4566# 9.33e-19
C1744 a_23879_6940# a_24763_6143# 1.03e-20
C1745 ringtest_0.x4.net9 ringtest_0.x4._20_ 1.35e-20
C1746 ringtest_0.x4.net3 a_22164_4362# 8.22e-19
C1747 ringtest_0.x4.net7 a_26375_4612# 6.33e-20
C1748 ringtest_0.x4._11_ a_25168_5156# 0.026293f
C1749 a_22021_4220# a_22390_4566# 0.046138f
C1750 ringtest_0.x4._23_ ringtest_0.x4._25_ 0.0063f
C1751 ringtest_0.x4.net5 ringtest_0.x4.counter[4] 0.001223f
C1752 a_27065_5156# a_26627_4246# 2.58e-19
C1753 a_27233_5058# a_27273_4220# 0.005283f
C1754 a_19666_31955# muxtest_0.x1.x3.GN3 0.104183f
C1755 a_21675_9686# a_21561_9116# 1.96e-19
C1756 ringtest_0.counter7 a_21375_3867# 2.81e-20
C1757 ringtest_0.x4.net5 a_23399_3867# 0.233889f
C1758 a_25421_6641# ringtest_0.x4._24_ 1.86e-20
C1759 a_19290_32287# VDPWR 0.194389f
C1760 a_22649_6244# a_22373_5156# 2.6e-20
C1761 a_27065_5156# a_27149_5156# 0.008508f
C1762 ringtest_0.x4._02_ VDPWR 0.325572f
C1763 a_21840_5308# a_22265_5308# 1.28e-19
C1764 a_21399_5340# a_22097_5334# 0.196846f
C1765 muxtest_0.x1.x1.nSEL0 a_18662_32213# 0.081627f
C1766 muxtest_0.x2.x2.GN4 a_13675_24012# 0.001562f
C1767 ringtest_0.x4.net6 a_25083_4790# 0.00565f
C1768 ringtest_0.x4._15_ a_24729_4790# 4.49e-20
C1769 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GN4 0.071281f
C1770 ringtest_0.x4.net8 a_24926_5712# 4.88e-19
C1771 m2_15612_11606# VDPWR 0.14037f
C1772 a_25364_5878# a_26640_5334# 0.01166f
C1773 ringtest_0.x4.net7 ringtest_0.x4._20_ 0.035834f
C1774 ringtest_0.x4._16_ a_21399_5340# 8.97e-20
C1775 muxtest_0.x1.x3.GP1 ui_in[0] 8.18e-19
C1776 VDPWR ui_in[3] 6.025721f
C1777 a_24045_6654# a_24336_6544# 0.192261f
C1778 a_23879_6940# ringtest_0.x4.clknet_1_1__leaf_clk 0.002451f
C1779 muxtest_0.x1.x1.nSEL0 m2_18699_31802# 3.43e-19
C1780 a_24895_4790# a_25083_4790# 0.095025f
C1781 a_25336_4902# a_25593_5156# 0.036838f
C1782 a_24729_4790# a_25263_5156# 0.002698f
C1783 a_20318_32213# ui_in[0] 0.220425f
C1784 ringtest_0.x4._17_ ringtest_0.x4._20_ 1.89e-19
C1785 ringtest_0.x3.nselect2 ringtest_0.x3.x2.GN4 1.53e-20
C1786 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GP1 6.21e-20
C1787 muxtest_0.R3R4 ua[2] 4.52137f
C1788 ui_in[2] ui_in[6] 0.264066f
C1789 ringtest_0.x4.clknet_1_1__leaf_clk a_25309_5334# 0.001538f
C1790 ringtest_0.x4.net6 a_24715_5334# 0.008614f
C1791 muxtest_0.x1.x3.GN4 muxtest_0.R1R2 0.628977f
C1792 a_26895_3867# ringtest_0.x4.counter[9] 2.34e-19
C1793 ringtest_0.x4._14_ a_22765_4478# 0.112679f
C1794 a_26201_5340# a_26201_4790# 0.037572f
C1795 a_21395_6940# ringtest_0.x4.net4 4.87e-19
C1796 uio_in[4] uio_in[3] 0.031023f
C1797 ringtest_0.x4._11_ a_21591_6128# 0.002118f
C1798 a_25593_5156# VDPWR 0.1878f
C1799 a_21375_3867# a_22295_3867# 1.37e-20
C1800 ringtest_0.x4._00_ ui_in[5] 2.67e-19
C1801 a_23879_6940# a_24800_5334# 5.07e-19
C1802 a_24329_6640# a_24545_5878# 2.84e-21
C1803 a_22399_9142# a_22245_8054# 9.03e-20
C1804 muxtest_0.x1.x3.GN2 muxtest_0.R3R4 0.271818f
C1805 muxtest_0.x1.x3.GP2 muxtest_0.x1.x4.A 0.350401f
C1806 a_22116_4902# VDPWR 0.219675f
C1807 ringtest_0.x4.net3 a_21845_8816# 0.008811f
C1808 a_24465_6800# ringtest_0.x4._06_ 4.29e-19
C1809 a_26201_5340# a_26555_5334# 0.062224f
C1810 a_21587_5334# a_21767_5334# 0.001229f
C1811 a_24336_6544# a_24699_6200# 6.47e-19
C1812 a_21845_9116# a_21845_8816# 0.040702f
C1813 ringtest_0.x4._00_ ringtest_0.x4._12_ 4.17e-19
C1814 a_21852_9416# a_21852_8720# 0.027204f
C1815 a_23993_5654# VDPWR 2.25e-21
C1816 ringtest_0.x4._15_ a_22390_4566# 8.81e-20
C1817 a_19666_31955# muxtest_0.x1.x3.GP2 2.46e-19
C1818 ringtest_0.x4._15_ a_26749_6422# 0.001357f
C1819 ringtest_0.x4._19_ a_24287_6422# 1.83e-19
C1820 ringtest_0.x4.net2 a_22201_9142# 1.37e-19
C1821 ringtest_0.x4._15_ ringtest_0.x4.net11 1.7e-19
C1822 ringtest_0.x4.net7 a_26569_6422# 6.19e-19
C1823 ringtest_0.x4.net2 a_21852_9416# 4.89e-19
C1824 ui_in[1] ui_in[2] 2.795f
C1825 ringtest_0.ring_out a_17231_12017# 0.001281f
C1826 ringtest_0.x4._05_ ringtest_0.x4._15_ 9.02e-20
C1827 a_26201_4790# a_27233_5058# 0.048748f
C1828 ringtest_0.x4._09_ a_26640_5156# 0.0221f
C1829 ringtest_0.x4._17_ a_26569_6422# 0.056144f
C1830 ringtest_0.x4.net3 a_22373_5156# 1.53e-21
C1831 ringtest_0.x4._22_ a_24361_5340# 0.016414f
C1832 a_24763_6143# a_24968_5308# 1.06e-19
C1833 a_22541_5058# a_22390_4566# 0.001062f
C1834 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 2.86851f
C1835 muxtest_0.x2.x2.GP1 ua[3] 4.09825f
C1836 ringtest_0.x4._04_ VDPWR 0.27578f
C1837 muxtest_0.x1.x5.GN ui_in[2] 3.98638f
C1838 a_21951_5878# a_22097_5334# 3.42e-19
C1839 a_24699_6200# a_24986_5878# 3.14e-19
C1840 a_22392_5990# a_22265_5308# 0.002135f
C1841 a_24329_6640# a_24317_4942# 8.37e-20
C1842 ringtest_0.x4.clknet_1_0__leaf_clk a_22223_5712# 4.11e-19
C1843 ringtest_0.x4.clknet_0_clk a_24627_6200# 2.68e-20
C1844 a_12297_23648# ua[3] 1.21e-19
C1845 ringtest_0.x4.clknet_1_0__leaf_clk VDPWR 3.74806f
C1846 a_21951_5878# ringtest_0.x4._16_ 1.01e-19
C1847 ringtest_0.x4.net9 a_27489_3702# 0.003439f
C1848 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ui_in[4] 9.08e-20
C1849 a_24045_6654# a_23899_5334# 4.21e-21
C1850 ringtest_0.x4.clknet_1_1__leaf_clk a_24968_5308# 0.01748f
C1851 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.173286f
C1852 ringtest_0.x4.net2 ringtest_0.x4._14_ 0.45134f
C1853 a_21591_6128# a_21785_5878# 5.05e-19
C1854 ringtest_0.x4._18_ a_21233_5340# 3.08e-21
C1855 a_22052_8875# ringtest_0.x4._01_ 0.004715f
C1856 a_26808_5308# a_27149_5334# 9.73e-19
C1857 a_26640_5334# a_26735_5334# 0.007724f
C1858 a_21852_9416# a_22399_8976# 4.5e-20
C1859 ringtest_0.x4._00_ a_22245_8054# 5.19e-20
C1860 a_12849_23648# ui_in[3] 0.086353f
C1861 a_27233_5058# a_27303_4246# 1.25e-19
C1862 a_21803_9508# ringtest_0.x4.clknet_1_0__leaf_clk 7.44e-19
C1863 a_22228_9508# a_22399_9142# 0.001229f
C1864 ringtest_0.drv_out ringtest_0.x4.net6 2.01e-20
C1865 ringtest_0.x4._11_ ringtest_0.x4._18_ 0.035586f
C1866 ringtest_0.x4.net7 a_24287_6422# 6.13e-20
C1867 ringtest_0.x4._11_ ringtest_0.counter7 2.85e-19
C1868 ringtest_0.x4._17_ a_22392_5990# 2.52e-22
C1869 a_24527_5340# a_25393_5308# 0.034054f
C1870 a_24361_5340# a_25225_5334# 0.030894f
C1871 ringtest_0.x4.net1 ringtest_0.x4.clknet_1_0__leaf_clk 0.561165f
C1872 a_21399_5340# a_21587_5334# 0.097818f
C1873 a_24968_5308# a_24800_5334# 0.239923f
C1874 a_18662_32213# muxtest_0.x1.x3.GN2 0.039612f
C1875 ringtest_0.x4._15_ ringtest_0.x4._09_ 0.030214f
C1876 ringtest_0.x4.clknet_1_1__leaf_clk a_25925_6788# 0.001522f
C1877 ringtest_0.x4._17_ a_24287_6422# 0.002375f
C1878 ringtest_0.x4._21_ a_23993_5654# 4.25e-19
C1879 muxtest_0.x1.x3.GN3 ua[0] 0.007815f
C1880 a_24329_6640# ringtest_0.x4._19_ 0.074331f
C1881 ringtest_0.x4.clknet_0_clk a_25393_5308# 0.01296f
C1882 ringtest_0.x4._03_ a_22164_4362# 0.005187f
C1883 ringtest_0.x4.net4 a_22223_5712# 3.33e-19
C1884 a_24317_4942# a_24551_4790# 0.005167f
C1885 ringtest_0.x4._15_ a_26766_5712# 4.15e-19
C1886 a_17377_14114# VDPWR 0.006305f
C1887 ringtest_0.x4.net4 VDPWR 1.18326f
C1888 a_16755_12091# ui_in[4] 0.127717f
C1889 ringtest_0.x4._24_ a_27233_5308# 0.009415f
C1890 ringtest_0.x4._11_ a_24763_6143# 0.004209f
C1891 a_21948_5156# ringtest_0.x4.net5 4.4e-19
C1892 a_22373_5156# a_22457_5156# 0.008508f
C1893 ringtest_0.x4.net3 a_21399_5340# 0.007798f
C1894 a_22765_5308# a_22765_4478# 8.07e-19
C1895 ringtest_0.x4._08_ ringtest_0.x4._22_ 1.19e-20
C1896 ringtest_0.x4.net8 a_25975_3867# 0.2272f
C1897 ringtest_0.x4._18_ a_23899_5654# 9.76e-19
C1898 ringtest_0.x4._11_ a_22295_3867# 3.83e-19
C1899 a_21951_5878# a_22649_6244# 0.194203f
C1900 a_22392_5990# a_22817_6146# 1.28e-19
C1901 ringtest_0.x4._16_ a_23381_4584# 0.039613f
C1902 a_12425_24040# VDPWR 4.32e-19
C1903 muxtest_0.x1.x4.A muxtest_0.R3R4 4.53278f
C1904 a_23899_5334# a_23809_4790# 8.68e-19
C1905 ringtest_0.x4.net9 a_25149_4220# 0.125008f
C1906 muxtest_0.x2.x2.GN1 VDPWR 1.60341f
C1907 ringtest_0.x4._01_ a_21803_8598# 2.39e-19
C1908 a_21852_8720# ringtest_0.x4._10_ 6.77e-19
C1909 ringtest_0.x4.net6 ringtest_0.x4._07_ 0.066033f
C1910 a_23529_6422# a_23770_5308# 6.83e-19
C1911 a_22052_8875# a_21785_8054# 0.0033f
C1912 a_24715_5334# a_24895_5334# 0.001229f
C1913 a_24045_6654# ringtest_0.x4._16_ 1.29e-20
C1914 ringtest_0.x4._07_ a_24895_4790# 0.195848f
C1915 a_24329_6640# ringtest_0.x4.net9 6.06e-20
C1916 ringtest_0.x4._22_ a_25336_4902# 0.001181f
C1917 ringtest_0.x4._19_ a_25364_5878# 6.04e-19
C1918 ringtest_0.x4.net2 ringtest_0.x4._10_ 0.006086f
C1919 ringtest_0.x4.net6 a_25055_3867# 0.013611f
C1920 ringtest_0.x4._11_ ringtest_0.x4.clknet_1_1__leaf_clk 0.367667f
C1921 muxtest_0.R3R4 m3_13302_19985# 0.136776f
C1922 a_24895_4790# a_25055_3867# 1.2e-20
C1923 ringtest_0.x4._00_ a_22228_9508# 8.32e-19
C1924 a_25925_6788# ringtest_0.x4._23_ 0.026998f
C1925 ringtest_0.x4._18_ a_21785_5878# 7.56e-20
C1926 ringtest_0.x4.net6 a_24264_6788# 1.91e-20
C1927 ringtest_0.x4.net7 a_25149_4220# 0.212284f
C1928 a_21425_9686# ringtest_0.x4.clknet_1_0__leaf_clk 3.24e-19
C1929 muxtest_0.x1.x5.GN a_19794_32347# 9.76e-20
C1930 muxtest_0.x1.x1.nSEL1 a_19242_32347# 9.57e-19
C1931 ringtest_0.x4.net7 a_26735_5156# 1.13e-19
C1932 muxtest_0.x1.x3.GP2 ua[0] 1.13e-20
C1933 a_21675_4790# a_22295_3867# 7.04e-21
C1934 a_23837_5878# VDPWR 0.004487f
C1935 a_24329_6640# ringtest_0.x4.net7 0.035144f
C1936 ringtest_0.x4._14_ a_21840_5308# 8.48e-21
C1937 ringtest_0.x4._22_ VDPWR 0.56354f
C1938 ringtest_0.x3.x2.GP1 ua[1] 0.352376f
C1939 ringtest_0.x4._06_ a_23770_5308# 0.002127f
C1940 ringtest_0.x4.clknet_1_1__leaf_clk a_25761_5058# 0.084941f
C1941 muxtest_0.R3R4 muxtest_0.x2.x2.GP2 0.171364f
C1942 ringtest_0.x4.net8 a_26367_5340# 5.19e-19
C1943 ringtest_0.x4._11_ a_24800_5334# 2.99e-20
C1944 ringtest_0.x4.net9 a_24545_5878# 0.063508f
C1945 ringtest_0.x4._19_ a_24317_4942# 4.85e-22
C1946 ringtest_0.x4._17_ a_24329_6640# 0.42661f
C1947 a_24070_5852# a_23770_5308# 8.74e-19
C1948 a_24135_3867# VDPWR 0.287214f
C1949 a_17231_12017# a_17405_12123# 0.006584f
C1950 a_16755_12091# ringtest_0.x3.x2.GP1 2.87e-20
C1951 ringtest_0.x4.net2 a_21509_4790# 5.19e-20
C1952 ringtest_0.x4._08_ a_25225_5334# 7.33e-20
C1953 muxtest_0.x2.x1.nSEL1 a_12473_23980# 0.041068f
C1954 a_15749_12123# ringtest_0.x3.x2.GN2 8.86e-19
C1955 a_17231_12017# ringtest_0.x3.x2.GN3 1.07e-20
C1956 ringtest_0.x3.x2.GN1 a_16155_12151# 1.22e-20
C1957 a_24699_6200# ringtest_0.x4._16_ 0.113309f
C1958 a_25364_5878# ringtest_0.x4.net9 0.111158f
C1959 a_23619_6788# VDPWR 0.002157f
C1960 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ui_in[4] 0.001652f
C1961 ringtest_0.x4.net6 a_26201_5340# 2.14e-19
C1962 a_21509_4790# a_23381_4818# 7.98e-21
C1963 ringtest_0.x4._03_ a_22373_5156# 0.001345f
C1964 ringtest_0.x4._15_ a_24361_5340# 0.034785f
C1965 muxtest_0.x1.x4.A muxtest_0.x2.x1.nSEL0 4.83e-20
C1966 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 5.04e-19
C1967 ringtest_0.x4.net4 ringtest_0.x4.counter[2] 0.006188f
C1968 ringtest_0.x4.net7 a_24545_5878# 2.13e-20
C1969 a_25225_5334# a_25336_4902# 0.001204f
C1970 a_25393_5308# a_25168_5156# 0.003655f
C1971 a_16027_11759# VDPWR 0.161536f
C1972 a_21465_8830# ringtest_0.x4._12_ 0.027335f
C1973 muxtest_0.x1.x3.GN4 muxtest_0.R6R7 0.156481f
C1974 ringtest_0.x4._16_ a_24479_4790# 7.06e-20
C1975 ringtest_0.x4._11_ ringtest_0.x4._23_ 0.090724f
C1976 ringtest_0.x4.net2 a_21867_8054# 6.45e-19
C1977 ringtest_0.x4.net7 a_25364_5878# 0.037674f
C1978 ringtest_0.x4.net6 ringtest_0.x4.counter[5] 0.080069f
C1979 ringtest_0.x4._11_ a_26367_4790# 7.13e-19
C1980 a_19842_32287# muxtest_0.R7R8 7.47e-21
C1981 ringtest_0.x4._16_ a_23809_4790# 0.105405f
C1982 ringtest_0.x4.net2 ringtest_0.x4._13_ 0.197255f
C1983 a_15749_12123# ui_in[3] 9.55e-19
C1984 a_23949_6654# ringtest_0.x4.net8 1.16e-19
C1985 a_24527_5340# a_24715_5334# 0.095025f
C1986 ringtest_0.x4._17_ a_25364_5878# 0.002308f
C1987 ringtest_0.x4.net9 a_24317_4942# 3.24e-20
C1988 ringtest_0.counter3 ringtest_0.counter7 3.44556f
C1989 a_25225_5334# VDPWR 0.182006f
C1990 ui_in[2] ui_in[4] 0.015983f
C1991 muxtest_0.R7R8 m3_13316_18955# 0.131878f
C1992 ringtest_0.x4._16_ a_22795_5334# 0.059496f
C1993 a_24465_6800# a_24883_6800# 3.39e-19
C1994 a_21675_10006# ringtest_0.x4._00_ 0.002065f
C1995 a_19114_31955# a_19290_32287# 0.185422f
C1996 ringtest_0.x4._23_ a_25761_5058# 1.37e-20
C1997 a_21233_5340# ringtest_0.x4._02_ 0.184941f
C1998 a_25761_5058# a_26367_4790# 8.52e-19
C1999 a_23529_6422# ringtest_0.x4.net6 1.5e-19
C2000 a_12473_23980# muxtest_0.x2.x2.GN3 0.048646f
C2001 ringtest_0.x4.net7 a_24317_4942# 0.084753f
C2002 a_12849_23648# muxtest_0.x2.x2.GN1 6.43e-20
C2003 ringtest_0.x4._21_ a_23837_5878# 0.002821f
C2004 ringtest_0.counter7 ua[2] 2.06e-19
C2005 ringtest_0.x4._11_ ringtest_0.x4._02_ 0.012298f
C2006 ringtest_0.x4._21_ ringtest_0.x4._22_ 2.96e-19
C2007 ringtest_0.x4._17_ a_24317_4942# 1.09e-21
C2008 a_26749_6422# a_26367_5340# 6.98e-21
C2009 m2_11882_23495# ui_in[3] 0.130999f
C2010 a_27169_6641# a_26201_5340# 7.7e-20
C2011 a_21509_4790# ringtest_0.x4._20_ 1.9e-21
C2012 ringtest_0.x4._03_ a_22499_4790# 9.96e-20
C2013 a_22021_4220# VDPWR 0.377321f
C2014 ringtest_0.counter7 ringtest_0.x4.net10 5.8e-20
C2015 ringtest_0.x4.net8 a_24004_6128# 0.063158f
C2016 a_21951_5878# a_22733_6244# 4.04e-19
C2017 a_26640_5156# VDPWR 0.248502f
C2018 a_22224_6244# a_22139_5878# 0.037333f
C2019 ringtest_0.counter3 a_22295_3867# 5.4e-19
C2020 ringtest_0.x4._12_ a_21780_8964# 0.001666f
C2021 a_21132_8918# a_21049_8598# 2.42e-19
C2022 ringtest_0.x4.net4 a_21375_3867# 7.77e-19
C2023 ringtest_0.x4.net6 ringtest_0.x4._06_ 0.037389f
C2024 ringtest_0.x4._19_ ringtest_0.x4.net9 4.58e-20
C2025 VDPWR ua[3] 11.3115f
C2026 a_23879_6940# a_23837_5878# 1.78e-20
C2027 ringtest_0.x4._24_ a_27491_4566# 5.3e-19
C2028 ringtest_0.x4.net6 a_24070_5852# 0.016498f
C2029 ringtest_0.x3.x2.GP2 ringtest_0.counter3 0.148166f
C2030 a_21399_5340# ringtest_0.x4._03_ 1.23e-19
C2031 a_21840_5308# a_21509_4790# 0.001425f
C2032 a_26201_4790# a_26895_3867# 4.75e-20
C2033 a_23879_6940# ringtest_0.x4._22_ 7.51e-19
C2034 a_21233_5340# a_22116_4902# 0.001786f
C2035 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP1 0.051787f
C2036 ringtest_0.x4.net8 a_23963_4790# 8.5e-20
C2037 ringtest_0.x4._15_ ringtest_0.x4._08_ 0.030258f
C2038 a_22765_4478# a_22390_4566# 4e-20
C2039 muxtest_0.R3R4 ua[0] 3.1523f
C2040 ringtest_0.x4._11_ a_25593_5156# 0.045045f
C2041 a_20492_32319# VDPWR 8.55e-19
C2042 ringtest_0.counter7 ringtest_0.x4.counter[4] 0.007159f
C2043 ui_in[1] ui_in[6] 0.239552f
C2044 a_21561_9116# a_21780_9142# 0.006169f
C2045 a_20318_32213# muxtest_0.x1.x3.GN3 1.07e-20
C2046 a_21675_9686# a_21845_9116# 5.23e-20
C2047 a_21465_9294# a_21852_9416# 0.034054f
C2048 muxtest_0.x1.x3.GN1 a_19242_32347# 1.22e-20
C2049 ringtest_0.counter7 a_23399_3867# 2.81e-20
C2050 a_18836_32319# muxtest_0.x1.x3.GN2 8.86e-19
C2051 a_19842_32287# VDPWR 0.261767f
C2052 a_27065_5156# ringtest_0.x4.net11 0.003417f
C2053 ringtest_0.x4._11_ a_22116_4902# 0.004479f
C2054 ringtest_0.x4._19_ ringtest_0.x4.net7 0.552257f
C2055 muxtest_0.x1.x1.nSEL0 a_19290_32287# 0.001174f
C2056 ringtest_0.x4._15_ a_25336_4902# 4.59e-21
C2057 a_22649_6244# a_22795_5334# 1.65e-19
C2058 ringtest_0.x4._11_ a_23993_5654# 5.64e-19
C2059 ringtest_0.x4._16_ a_21672_5334# 1.68e-20
C2060 a_24045_6654# a_24465_6800# 0.036838f
C2061 a_24329_6640# a_24536_6699# 0.260055f
C2062 a_23949_6654# ringtest_0.x4._05_ 1.85e-19
C2063 ringtest_0.x4._17_ ringtest_0.x4._19_ 0.214371f
C2064 ringtest_0.x4._24_ a_27149_5334# 8.56e-19
C2065 a_25168_5156# a_25083_4790# 0.037333f
C2066 a_25761_5058# a_25593_5156# 0.310858f
C2067 ua[0] ui_in[5] 0.483363f
C2068 muxtest_0.R3R4 muxtest_0.x2.x2.GN3 3.9625f
C2069 a_21561_8830# VDPWR 0.181976f
C2070 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net10 6.99e-20
C2071 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x1.nSEL1 0.352716f
C2072 ringtest_0.x4._04_ a_21233_5340# 0.001469f
C2073 ringtest_0.drv_out ui_in[5] 0.391919f
C2074 a_27815_3867# ringtest_0.x4.counter[9] 0.039377f
C2075 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ui_in[4] 1.79e-19
C2076 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x3.x2.GN1 2.09e-20
C2077 ringtest_0.x4._15_ VDPWR 1.72333f
C2078 ringtest_0.x4.clknet_1_0__leaf_clk a_21233_5340# 0.318658f
C2079 a_21675_4790# a_22116_4902# 0.127288f
C2080 a_26808_5308# a_26201_4790# 1.99e-20
C2081 ringtest_0.drv_out ringtest_0.x4.clknet_0_clk 0.00889f
C2082 ringtest_0.x4._11_ ringtest_0.x4._04_ 0.257603f
C2083 ui_in[0] ui_in[2] 0.450267f
C2084 a_25263_5156# VDPWR 0.003234f
C2085 a_22295_3867# a_23399_3867# 9e-21
C2086 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.173286f
C2087 a_25364_5878# a_26627_4246# 1.15e-20
C2088 a_24536_6699# a_24545_5878# 1.55e-20
C2089 ringtest_0.x4.net7 ringtest_0.x4.net9 0.742565f
C2090 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._11_ 0.317456f
C2091 a_22541_5058# VDPWR 0.391294f
C2092 ringtest_0.x4.net3 a_22052_8875# 3.02e-19
C2093 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.ring_out 0.083309f
C2094 ringtest_0.x4.net2 ringtest_0.x4.counter[1] 0.015257f
C2095 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP2 0.100463f
C2096 a_25225_5334# a_25309_5334# 0.008508f
C2097 a_26808_5308# a_26555_5334# 3.39e-19
C2098 ringtest_0.x4._17_ ringtest_0.x4.net9 7.02e-19
C2099 a_21845_9116# a_22052_8875# 6.88e-20
C2100 a_22052_9116# a_21852_8720# 1.26e-19
C2101 muxtest_0.x1.x5.GN ui_in[1] 0.141313f
C2102 a_24465_6800# a_24699_6200# 1.61e-19
C2103 a_21981_9142# a_21845_8816# 5.28e-20
C2104 a_24926_5712# VDPWR 0.001185f
C2105 ringtest_0.x3.x2.GN2 ringtest_0.counter3 0.004367f
C2106 ringtest_0.x4._15_ a_23467_4584# 0.001523f
C2107 ringtest_0.x4.net8 ringtest_0.x4._20_ 0.027217f
C2108 ringtest_0.x4._15_ ringtest_0.x4._25_ 0.003323f
C2109 ringtest_0.x4.net1 a_21561_8830# 0.030538f
C2110 ringtest_0.ring_out a_17405_12123# 1.86e-19
C2111 ringtest_0.x4.net2 a_22052_9116# 1.88e-19
C2112 ringtest_0.ring_out ringtest_0.x3.x2.GN3 0.080584f
C2113 a_26201_4790# a_26555_4790# 0.062224f
C2114 a_21951_5878# ringtest_0.x4._03_ 3.92e-19
C2115 ringtest_0.x4._09_ a_27065_5156# 0.024482f
C2116 ringtest_0.x4._07_ a_24527_5340# 0.029939f
C2117 ringtest_0.x4._22_ a_24968_5308# 0.01767f
C2118 ringtest_0.x4.net5 a_22164_4362# 3.95e-20
C2119 ringtest_0.x4._17_ ringtest_0.x4.net7 0.072785f
C2120 ringtest_0.x4.clknet_1_0__leaf_clk a_21675_4790# 0.021572f
C2121 ringtest_0.counter7 a_26808_4902# 1.4e-19
C2122 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN3 4.01e-20
C2123 a_24527_5340# a_25055_3867# 7.09e-22
C2124 ringtest_0.x4._23_ ringtest_0.x4.net10 0.188811f
C2125 ringtest_0.x4.clknet_0_clk ringtest_0.x4._07_ 0.114561f
C2126 a_21049_8598# VDPWR 0.229121f
C2127 ringtest_0.x3.x2.GN4 ringtest_0.counter7 3.94045f
C2128 ringtest_0.counter3 ringtest_0.x4._02_ 0.001266f
C2129 ringtest_0.x4._20_ a_24729_4790# 0.004564f
C2130 a_22224_6244# a_22097_5334# 0.002298f
C2131 ringtest_0.x4.net10 a_26367_4790# 0.003321f
C2132 a_26173_4612# VDPWR 0.001618f
C2133 a_12849_23648# ua[3] 0.001506f
C2134 ringtest_0.x4.net4 a_21233_5340# 0.007432f
C2135 a_22224_6244# ringtest_0.x4._16_ 1.81e-20
C2136 a_26895_3867# ringtest_0.x4.counter[8] 6.92e-19
C2137 muxtest_0.x1.x4.A a_13025_23980# 3.23e-19
C2138 ringtest_0.x4.clknet_1_1__leaf_clk a_25393_5308# 0.005058f
C2139 ringtest_0.x4.net6 a_21399_5340# 1.26e-19
C2140 ringtest_0.x4.clknet_0_clk a_24264_6788# 1.49e-19
C2141 ringtest_0.x4._11_ ringtest_0.x4.net4 0.952686f
C2142 a_21785_5878# ringtest_0.x4._04_ 0.09532f
C2143 ringtest_0.x4._15_ ringtest_0.x4._21_ 0.054317f
C2144 ringtest_0.x4.clknet_1_0__leaf_clk a_21785_5878# 0.245743f
C2145 a_26627_4246# a_26913_4566# 0.010132f
C2146 muxtest_0.x2.x2.GN1 m2_11882_23495# 0.06935f
C2147 a_13501_23906# ui_in[3] 0.220366f
C2148 a_22399_9142# ringtest_0.x4.clknet_1_0__leaf_clk 0.012004f
C2149 ui_in[3] ua[2] 1.63519f
C2150 ringtest_0.x4.net1 a_21049_8598# 0.060735f
C2151 a_21425_9686# a_21561_8830# 6.59e-20
C2152 ringtest_0.x4.net7 a_26095_6788# 0.00717f
C2153 ringtest_0.x4._21_ a_22541_5058# 1.79e-21
C2154 ringtest_0.x4._17_ a_22817_6146# 1.35e-20
C2155 a_21840_5308# a_21798_5712# 4.62e-19
C2156 a_21672_5334# a_21587_5334# 0.037333f
C2157 a_24527_5340# a_26201_5340# 1.33e-19
C2158 a_24968_5308# a_25225_5334# 0.036838f
C2159 a_24361_5340# a_26367_5340# 3.42e-21
C2160 a_19290_32287# muxtest_0.x1.x3.GN2 0.017048f
C2161 ringtest_0.x4.net9 a_27065_5334# 2.45e-19
C2162 ringtest_0.x4.clknet_1_1__leaf_clk a_26808_4902# 2.7e-19
C2163 ringtest_0.x4.net4 a_21675_4790# 0.019846f
C2164 a_13025_23980# muxtest_0.x2.x2.GP2 3.2e-20
C2165 a_24536_6699# ringtest_0.x4._19_ 0.034076f
C2166 muxtest_0.x2.x2.GP3 ui_in[4] 0.00356f
C2167 a_23879_6940# ringtest_0.x4._15_ 2.08e-20
C2168 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP2 8.45e-19
C2169 ringtest_0.x4._03_ a_23381_4584# 2.93e-20
C2170 a_19794_32347# ui_in[0] 0.001558f
C2171 ringtest_0.x4.net4 a_23899_5654# 7.88e-20
C2172 ringtest_0.x3.x2.GN1 ui_in[4] 0.312198f
C2173 ringtest_0.x4._11_ a_23837_5878# 3.73e-19
C2174 a_15575_12017# ringtest_0.x3.x2.GN2 0.039612f
C2175 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN3 0.012418f
C2176 ringtest_0.x4._11_ ringtest_0.x4._22_ 0.420712f
C2177 a_22373_5156# ringtest_0.x4.net5 0.019334f
C2178 ringtest_0.x4.net3 a_21672_5334# 8.21e-19
C2179 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ui_in[4] 1.03e-20
C2180 rst_n clk 0.031023f
C2181 a_22392_5990# ringtest_0.x4.net8 1.22e-20
C2182 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 5.04e-19
C2183 ringtest_0.x4.net9 a_26627_4246# 0.008597f
C2184 muxtest_0.x1.x3.GP1 muxtest_0.R3R4 4.16645f
C2185 ringtest_0.x4._01_ a_21785_8054# 3.94e-19
C2186 a_21981_8976# ringtest_0.x4._10_ 6.67e-19
C2187 a_24045_6654# a_23770_5308# 7.28e-21
C2188 ringtest_0.x4.net9 a_27149_5156# 1.5e-19
C2189 ringtest_0.x4.net4 a_21785_5878# 0.071607f
C2190 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ui_in[3] 1.18e-19
C2191 ringtest_0.x4._11_ a_23619_6788# 1.46e-19
C2192 ringtest_0.x4._07_ a_25168_5156# 0.008539f
C2193 a_24336_6544# ringtest_0.x4._16_ 6.29e-20
C2194 a_24883_6800# a_24712_6422# 0.001229f
C2195 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.ring_out 0.025177f
C2196 a_24536_6699# ringtest_0.x4.net9 4.56e-19
C2197 ringtest_0.x4._22_ a_25761_5058# 3.11e-19
C2198 ui_in[4] ui_in[6] 0.177925f
C2199 ui_in[0] rst_n 0.031023f
C2200 ringtest_0.x4.clknet_0_clk a_23529_6422# 8e-19
C2201 ringtest_0.x4.net6 a_21951_5878# 0.004467f
C2202 ringtest_0.x4._24_ a_27273_4220# 0.003347f
C2203 a_15575_12017# m2_15612_11606# 0.01297f
C2204 a_26569_6422# a_26749_6422# 0.185422f
C2205 a_15575_12017# ui_in[3] 0.048888f
C2206 ringtest_0.x4._24_ a_26766_4790# 6.57e-19
C2207 ringtest_0.x4.net6 a_24883_6800# 9.51e-20
C2208 ringtest_0.x4._00_ ringtest_0.x4.clknet_1_0__leaf_clk 0.144154f
C2209 ringtest_0.x4.net7 a_27149_5156# 3.05e-20
C2210 ringtest_0.x4._23_ a_26808_4902# 0.005759f
C2211 muxtest_0.x1.x1.nSEL1 VDPWR 0.475048f
C2212 a_24763_6143# a_24715_5334# 1.39e-19
C2213 ringtest_0.x4._05_ a_26569_6422# 6.38e-20
C2214 a_26367_4790# a_26808_4902# 0.118966f
C2215 a_24536_6699# ringtest_0.x4.net7 0.026259f
C2216 ringtest_0.x4._14_ a_22265_5308# 1.02e-20
C2217 ringtest_0.x4._06_ a_24527_5340# 0.183131f
C2218 ringtest_0.x4.clknet_1_1__leaf_clk a_25083_4790# 0.011819f
C2219 ringtest_0.x4._16_ a_24986_5878# 3.12e-19
C2220 ringtest_0.x4.net8 a_26640_5334# 2.79e-19
C2221 ringtest_0.x4._11_ a_25225_5334# 7.12e-21
C2222 ringtest_0.x4._17_ a_24536_6699# 0.032936f
C2223 a_24004_6128# a_24361_5340# 4.26e-19
C2224 a_16707_12151# ringtest_0.x3.x2.GN4 3.22e-19
C2225 a_25975_3867# VDPWR 0.309637f
C2226 ringtest_0.x3.x2.GN3 a_17405_12123# 1.07e-20
C2227 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1 1.51569f
C2228 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GN4 8.82e-19
C2229 muxtest_0.x2.x1.nSEL1 a_13025_23980# 1.59e-19
C2230 ringtest_0.x4._08_ a_26367_5340# 0.415957f
C2231 ringtest_0.x4.net5 a_22499_4790# 6.03e-19
C2232 ringtest_0.x4.clknet_0_clk ringtest_0.x4._06_ 2.8e-19
C2233 a_24685_6788# VDPWR 0.002269f
C2234 ringtest_0.x4._04_ a_22775_5878# 6.79e-19
C2235 a_21785_5878# a_23837_5878# 9.88e-21
C2236 ringtest_0.x4.clknet_0_clk a_24070_5852# 7.65e-20
C2237 ringtest_0.x4.clknet_1_1__leaf_clk a_24715_5334# 0.017223f
C2238 ui_in[1] ui_in[4] 4.85e-19
C2239 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x3.nselect2 1.41e-19
C2240 ringtest_0.x4._15_ a_24968_5308# 0.03519f
C2241 a_21233_5340# a_22021_4220# 3.4e-19
C2242 ringtest_0.x4._22_ a_25345_4612# 0.002279f
C2243 ringtest_0.x4._01_ a_22695_8304# 0.012244f
C2244 muxtest_0.x1.x5.A ua[3] 4.51865f
C2245 ringtest_0.counter3 ringtest_0.x4.net4 8.11e-19
C2246 a_25393_5308# a_25593_5156# 4.17e-19
C2247 a_24800_5334# a_25083_4790# 0.001307f
C2248 a_26913_4566# a_26721_4246# 6.96e-20
C2249 muxtest_0.x1.x3.GN3 muxtest_0.R4R5 0.123863f
C2250 a_16579_11759# VDPWR 0.179803f
C2251 ringtest_0.x4.net8 a_25149_4220# 0.1454f
C2252 a_21845_8816# ringtest_0.x4._12_ 0.062549f
C2253 ringtest_0.x4._11_ a_22021_4220# 7.66e-19
C2254 ringtest_0.x4.net9 a_25294_4790# 3.93e-19
C2255 a_23770_5308# a_23809_4790# 2.2e-19
C2256 muxtest_0.x1.x5.GN ui_in[4] 2.49e-19
C2257 ringtest_0.x4.net11 a_27489_3702# 0.250513f
C2258 ringtest_0.x4._11_ a_26640_5156# 5.04e-19
C2259 muxtest_0.x1.x3.GN1 muxtest_0.R7R8 4.45989f
C2260 ringtest_0.x3.x2.GN4 ui_in[3] 0.218716f
C2261 a_24800_5334# a_24715_5334# 0.037333f
C2262 a_24968_5308# a_24926_5712# 4.62e-19
C2263 ringtest_0.x4.net2 a_21132_8918# 0.010623f
C2264 a_22765_5308# a_23151_5334# 0.006406f
C2265 a_24329_6640# ringtest_0.x4.net8 0.001356f
C2266 ringtest_0.x4._08_ a_27065_5156# 3.02e-19
C2267 a_26367_5340# VDPWR 0.31297f
C2268 ringtest_0.x4.net6 a_23381_4584# 1.4e-20
C2269 ringtest_0.x4._16_ a_23899_5334# 0.008193f
C2270 ringtest_0.x4._15_ a_25925_6788# 0.142876f
C2271 ringtest_0.x4._24_ a_26201_4790# 0.03301f
C2272 ringtest_0.drv_out ringtest_0.counter7 2.39e-19
C2273 ringtest_0.x4.net9 a_25351_5712# 3.81e-19
C2274 a_19290_32287# a_19666_31955# 3.02e-19
C2275 muxtest_0.x1.x4.A ui_in[3] 0.00371f
C2276 a_24729_4790# a_25149_4220# 0.009169f
C2277 a_24045_6654# ringtest_0.x4.net6 8.38e-19
C2278 a_13025_23980# muxtest_0.x2.x2.GN3 0.004288f
C2279 a_21675_4790# a_22021_4220# 0.010515f
C2280 a_24329_6640# a_24729_4790# 2.6e-21
C2281 muxtest_0.x2.x2.GN1 ua[2] 0.430038f
C2282 ringtest_0.x4._24_ a_26555_5334# 4.8e-19
C2283 a_27233_5308# a_27273_4220# 1.35e-20
C2284 ringtest_0.x4.net7 a_25351_5712# 1.38e-19
C2285 ringtest_0.x4.net8 a_24545_5878# 0.009814f
C2286 ringtest_0.x4._25_ a_26367_5340# 1.11e-19
C2287 ui_in[0] ui_in[6] 0.281408f
C2288 a_22765_4478# VDPWR 0.201367f
C2289 ringtest_0.x3.nselect2 a_16755_12091# 6.01e-20
C2290 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ui_in[4] 7.73e-20
C2291 a_21507_9686# VDPWR 0.008578f
C2292 ringtest_0.x4.net9 a_26721_4246# 0.003753f
C2293 a_22392_5990# a_22350_5878# 4.62e-19
C2294 a_21951_5878# a_23932_6128# 1.01e-20
C2295 a_27065_5156# VDPWR 0.215619f
C2296 ringtest_0.x4.net8 a_25364_5878# 0.001798f
C2297 ringtest_0.x4._15_ a_21233_5340# 8.17e-21
C2298 a_23949_6654# VDPWR 0.376761f
C2299 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.173286f
C2300 muxtest_0.x1.x3.GP2 muxtest_0.R4R5 0.117653f
C2301 a_21845_8816# a_22245_8054# 4.04e-19
C2302 ringtest_0.x4._12_ a_22201_8964# 0.002771f
C2303 ringtest_0.x4.net4 a_23399_3867# 0.003224f
C2304 muxtest_0.x2.x2.GP2 ui_in[3] 6.63e-19
C2305 muxtest_0.x1.x3.GN1 muxtest_0.R5R6 0.250509f
C2306 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B 0.163894f
C2307 ringtest_0.x4._11_ ringtest_0.x4._15_ 1.40124f
C2308 ringtest_0.x4.net6 a_24699_6200# 0.09145f
C2309 a_21672_5334# ringtest_0.x4._03_ 0.001262f
C2310 a_22265_5308# a_21509_4790# 0.00142f
C2311 ringtest_0.x4.net8 a_24551_4790# 5.79e-19
C2312 a_25364_5878# a_24729_4790# 4.21e-21
C2313 a_24699_6200# a_24895_4790# 8.41e-19
C2314 ringtest_0.drv_out ringtest_0.x4.clknet_1_1__leaf_clk 0.008913f
C2315 ringtest_0.drv_out ringtest_0.x3.x2.GP2 4.09557f
C2316 ringtest_0.counter7 a_25055_3867# 2.81e-20
C2317 a_21561_9116# a_21845_9116# 0.032244f
C2318 ringtest_0.x4._22_ ringtest_0.x4.net10 0.074459f
C2319 a_21951_5878# ringtest_0.x4.net5 3.57e-21
C2320 muxtest_0.x1.x3.GN1 VDPWR 0.915833f
C2321 ringtest_0.x4.net8 a_24317_4942# 0.236033f
C2322 ringtest_0.x4._11_ a_22541_5058# 0.065594f
C2323 ringtest_0.x4.net1 a_21507_9686# 0.010028f
C2324 a_22265_5308# a_22765_5308# 0.016344f
C2325 muxtest_0.x1.x1.nSEL0 a_19842_32287# 1.21e-20
C2326 ui_in[0] ui_in[1] 4.44986f
C2327 ringtest_0.x4.net6 a_24479_4790# 1.78e-19
C2328 ringtest_0.x4._15_ a_25761_5058# 7.77e-19
C2329 ringtest_0.x4._16_ a_22097_5334# 1.35e-19
C2330 a_24329_6640# ringtest_0.x4._05_ 0.196756f
C2331 a_24336_6544# a_24465_6800# 0.110715f
C2332 muxtest_0.x1.x3.GN3 ui_in[2] 0.002225f
C2333 a_24004_6128# VDPWR 0.316019f
C2334 a_24729_4790# a_24551_4790# 1.43e-19
C2335 a_21395_6940# a_21840_5308# 3.17e-20
C2336 a_24763_6143# ringtest_0.x4._07_ 0.001092f
C2337 ringtest_0.x4.net6 a_23809_4790# 0.005791f
C2338 muxtest_0.x1.x5.GN ui_in[0] 0.149831f
C2339 a_21852_8720# VDPWR 0.309635f
C2340 a_24317_4942# a_24729_4790# 0.020429f
C2341 ringtest_0.x4._15_ a_23899_5654# 0.005043f
C2342 ringtest_0.x4.net6 a_22795_5334# 0.007899f
C2343 a_21675_4790# a_22541_5058# 0.034054f
C2344 a_24135_3867# ringtest_0.x4.counter[4] 0.110403f
C2345 a_22116_4902# a_21948_5156# 0.239923f
C2346 ringtest_0.x4.net2 VDPWR 2.41286f
C2347 a_23963_4790# VDPWR 3.08e-19
C2348 a_23399_3867# a_24135_3867# 2.31e-20
C2349 ringtest_0.x4._11_ a_26173_4612# 7.08e-19
C2350 muxtest_0.x1.x3.GP3 muxtest_0.R7R8 0.124327f
C2351 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._07_ 0.44529f
C2352 a_26749_6422# a_25364_5878# 0.006666f
C2353 a_23381_4818# VDPWR 0.254188f
C2354 ringtest_0.x4.net3 ringtest_0.x4._01_ 0.006403f
C2355 a_26640_5334# a_26766_5712# 0.005525f
C2356 ringtest_0.x4._19_ ringtest_0.x4.net8 2.14e-19
C2357 a_21845_9116# ringtest_0.x4._01_ 6.79e-20
C2358 ringtest_0.x4._05_ a_25364_5878# 0.003024f
C2359 a_23949_6654# ringtest_0.x4._21_ 0.001295f
C2360 a_21981_9142# a_22052_8875# 1.77e-19
C2361 a_22052_9116# a_21981_8976# 1.77e-19
C2362 ringtest_0.x4.clknet_1_0__leaf_clk a_21465_8830# 0.01132f
C2363 a_22181_5334# VDPWR 0.007439f
C2364 ringtest_0.x4.clknet_1_1__leaf_clk a_25055_3867# 4.13e-21
C2365 ringtest_0.x4._15_ a_25345_4612# 2.85e-21
C2366 ringtest_0.counter7 ringtest_0.x4.counter[5] 0.007023f
C2367 muxtest_0.x2.x1.nSEL1 ui_in[3] 0.168511f
C2368 ringtest_0.x4.net1 a_21852_8720# 0.00338f
C2369 ringtest_0.drv_out ringtest_0.x3.x2.GN2 3.92936f
C2370 a_26201_4790# a_25977_4220# 2.81e-20
C2371 a_21425_9686# a_21507_9686# 0.006406f
C2372 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP3 3.4436f
C2373 a_21785_5878# a_22541_5058# 3.85e-19
C2374 ringtest_0.x4.net8 a_26735_5334# 7.49e-20
C2375 ringtest_0.x4._04_ a_21948_5156# 3.52e-21
C2376 ringtest_0.x4._07_ a_24800_5334# 0.002926f
C2377 ringtest_0.x4.net1 ringtest_0.x4.net2 0.722672f
C2378 a_25421_6641# ringtest_0.x4.net6 0.019537f
C2379 ringtest_0.x4.net3 a_21863_4790# 7.76e-19
C2380 ringtest_0.x4.net5 a_23381_4584# 0.201023f
C2381 ringtest_0.x4._22_ a_25393_5308# 4.4e-21
C2382 muxtest_0.x1.x3.GP2 ui_in[2] 4.34e-19
C2383 ringtest_0.x4.clknet_1_0__leaf_clk a_21948_5156# 0.003461f
C2384 ringtest_0.x4._18_ a_23529_6422# 0.190808f
C2385 a_24800_5334# a_25055_3867# 3e-19
C2386 a_22399_8976# VDPWR 0.074934f
C2387 ringtest_0.x4._20_ a_25336_4902# 6.25e-20
C2388 a_23879_6940# a_23949_6654# 0.022122f
C2389 a_22817_6146# a_22765_5308# 0.004132f
C2390 muxtest_0.R7R8 muxtest_0.R1R2 0.216753f
C2391 ringtest_0.x4.net10 a_26640_5156# 5.45e-19
C2392 a_26375_4612# VDPWR 1.16e-19
C2393 a_13501_23906# ua[3] 0.003273f
C2394 ua[3] ua[2] 8.93455f
C2395 a_24883_6800# a_24527_5340# 1.11e-20
C2396 a_22649_6244# ringtest_0.x4._16_ 0.003542f
C2397 a_15575_12017# a_16027_11759# 0.002207f
C2398 a_27815_3867# ringtest_0.x4.counter[8] 0.111116f
C2399 ringtest_0.x4.net8 ringtest_0.x4.net9 0.748324f
C2400 a_24004_6128# ringtest_0.x4._21_ 0.128337f
C2401 muxtest_0.R4R5 muxtest_0.R3R4 1.39313f
C2402 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN1 1.38e-21
C2403 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ui_in[4] 1.2e-19
C2404 ringtest_0.x4.clknet_1_1__leaf_clk a_26201_5340# 0.285659f
C2405 ringtest_0.x3.x2.GP3 VDPWR 1.79155f
C2406 ringtest_0.x4._13_ ringtest_0.x4.counter[0] 3.39e-20
C2407 ringtest_0.x4.net6 a_21672_5334# 6.57e-20
C2408 ringtest_0.x4.clknet_0_clk a_24883_6800# 0.004448f
C2409 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 5.04e-19
C2410 muxtest_0.x1.x3.GP3 muxtest_0.R5R6 4.11451f
C2411 ringtest_0.x4._20_ VDPWR 0.175404f
C2412 ringtest_0.x4.net3 a_21785_8054# 0.079675f
C2413 ringtest_0.x4._22_ a_26808_4902# 8.71e-19
C2414 muxtest_0.x1.x3.GN2 ua[3] 0.01442f
C2415 a_22164_4362# a_22295_3867# 0.002548f
C2416 a_26627_4246# a_26721_4246# 0.062574f
C2417 a_27273_4220# a_27491_4566# 0.007234f
C2418 ringtest_0.x4.clknet_1_0__leaf_clk a_21780_8964# 0.001172f
C2419 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B 5.04e-19
C2420 a_13675_24012# ui_in[3] 1.4e-19
C2421 ringtest_0.x4._16_ a_23467_4818# 5.76e-19
C2422 ringtest_0.x4.net7 ringtest_0.x4.net8 1.22349f
C2423 a_25364_5878# ringtest_0.x4._09_ 3.55e-20
C2424 muxtest_0.x2.x2.GN3 ui_in[3] 0.254283f
C2425 ringtest_0.x4.net9 a_24729_4790# 0.006834f
C2426 ringtest_0.x4._18_ ringtest_0.x4._06_ 3.12e-20
C2427 ringtest_0.x4.net1 a_22399_8976# 6.38e-20
C2428 muxtest_0.x1.x3.GP3 VDPWR 3.24635f
C2429 muxtest_0.x1.x3.GN2 a_20492_32319# 8.14e-21
C2430 muxtest_0.x1.x3.GN3 a_19794_32347# 0.001073f
C2431 ringtest_0.x4.net7 a_26839_6788# 1.83e-19
C2432 ringtest_0.x4._18_ a_24070_5852# 7.58e-19
C2433 a_23879_6940# a_24004_6128# 1.01e-19
C2434 ringtest_0.x4._17_ ringtest_0.x4.net8 0.172731f
C2435 a_21840_5308# a_22223_5712# 4.67e-20
C2436 a_25393_5308# a_25225_5334# 0.310858f
C2437 a_19842_32287# muxtest_0.x1.x3.GN2 9.62e-20
C2438 ringtest_0.x4.net6 ringtest_0.x4._24_ 0.002355f
C2439 a_21840_5308# VDPWR 0.200136f
C2440 ringtest_0.x4.net2 a_21425_9686# 0.107098f
C2441 ringtest_0.x4._16_ a_21587_5334# 4.26e-21
C2442 muxtest_0.x1.x1.nSEL1 a_19114_31955# 0.073392f
C2443 ringtest_0.x4.net4 a_21948_5156# 0.004091f
C2444 ringtest_0.x4.clknet_1_1__leaf_clk a_27233_5058# 1.1e-19
C2445 ua[2] ua[6] 0.001584f
C2446 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP2 0.005194f
C2447 ringtest_0.x4._05_ ringtest_0.x4._19_ 0.284135f
C2448 ringtest_0.x4.net7 a_24729_4790# 0.003956f
C2449 a_23529_6422# ringtest_0.x4.clknet_1_1__leaf_clk 1.19e-21
C2450 ringtest_0.x3.x2.GP1 ui_in[4] 8.45e-19
C2451 ringtest_0.x4._17_ a_24729_4790# 1.69e-21
C2452 ringtest_0.x4._15_ ringtest_0.x4.net10 0.289356f
C2453 ringtest_0.x4._06_ a_24763_6143# 9.69e-19
C2454 a_16203_12091# ringtest_0.x3.x2.GN2 0.017071f
C2455 a_23809_4790# ringtest_0.x4.net5 5.06e-20
C2456 ringtest_0.x4._23_ a_26201_5340# 0.029216f
C2457 a_26569_6422# VDPWR 0.206381f
C2458 a_26201_5340# a_26367_4790# 2.64e-19
C2459 muxtest_0.R1R2 VDPWR 1.61319f
C2460 ringtest_0.x4.net3 ringtest_0.x4._16_ 6.72e-19
C2461 ringtest_0.x4._11_ a_25975_3867# 2.18e-19
C2462 a_22817_6146# ringtest_0.x4.net8 5.45e-19
C2463 a_26749_6422# ringtest_0.x4.net9 7.48e-22
C2464 a_24329_6640# a_24361_5340# 0.001493f
C2465 ringtest_0.x4.net9 ringtest_0.x4.net11 0.055197f
C2466 ringtest_0.x4._15_ ringtest_0.x4.counter[4] 9.07e-20
C2467 a_24465_6800# ringtest_0.x4._16_ 2.16e-20
C2468 ringtest_0.x4._07_ a_25593_5156# 5.62e-20
C2469 ringtest_0.x3.x2.GP2 m3_17036_9140# 0.004119f
C2470 ringtest_0.x4._05_ ringtest_0.x4.net9 1.93e-19
C2471 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._06_ 0.005269f
C2472 ringtest_0.x4._22_ a_25083_4790# 0.012798f
C2473 ringtest_0.x4.clknet_0_clk a_24045_6654# 0.00222f
C2474 ringtest_0.x4.net6 a_22224_6244# 3.12e-19
C2475 ringtest_0.x4.net2 a_21375_3867# 0.016821f
C2476 ringtest_0.x4._21_ ringtest_0.x4._20_ 0.296715f
C2477 ringtest_0.x4._14_ a_21509_4790# 0.008544f
C2478 a_25761_5058# a_25975_3867# 2.93e-21
C2479 a_26569_6422# ringtest_0.x4._25_ 0.001476f
C2480 ringtest_0.x4._24_ a_27169_6641# 0.006166f
C2481 a_16203_12091# ui_in[3] 0.143958f
C2482 ringtest_0.x4.net7 a_26749_6422# 5.4e-19
C2483 muxtest_0.R3R4 ui_in[2] 2.94e-19
C2484 ringtest_0.x4._23_ a_27233_5058# 2.3e-19
C2485 ringtest_0.x4.net7 ringtest_0.x4.net11 2.47e-20
C2486 a_26367_4790# a_27233_5058# 0.034054f
C2487 a_26808_4902# a_26640_5156# 0.239923f
C2488 ringtest_0.x4._14_ a_22765_5308# 1.74e-20
C2489 ringtest_0.x4._05_ ringtest_0.x4.net7 0.232588f
C2490 ringtest_0.x4._17_ a_26749_6422# 8.24e-19
C2491 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x1.nSEL1 0.352716f
C2492 ringtest_0.x4._06_ a_24800_5334# 3.32e-19
C2493 ringtest_0.x4.net8 a_27065_5334# 1.1e-19
C2494 ringtest_0.x4._11_ a_26367_5340# 2.03e-20
C2495 a_27489_3702# VDPWR 0.293517f
C2496 ringtest_0.x4._17_ ringtest_0.x4._05_ 0.0576f
C2497 a_24699_6200# a_24527_5340# 1.08e-19
C2498 muxtest_0.x2.x1.nSEL1 a_12425_24040# 9.57e-19
C2499 a_11845_23906# a_12019_24012# 0.006584f
C2500 a_22392_5990# VDPWR 0.177502f
C2501 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN1 0.034862f
C2502 ringtest_0.x4._08_ a_26640_5334# 0.030723f
C2503 ui_in[2] ui_in[5] 0.211146f
C2504 a_24287_6422# VDPWR 0.004852f
C2505 ringtest_0.x4._13_ ringtest_0.x4._14_ 0.074354f
C2506 ringtest_0.x4.clknet_0_clk a_24699_6200# 0.034583f
C2507 a_21509_4790# a_22043_5156# 0.002698f
C2508 ringtest_0.x4._15_ a_25393_5308# 0.031321f
C2509 ringtest_0.x4.counter[0] ringtest_0.x4.counter[1] 0.079742f
C2510 ringtest_0.x4._03_ a_21863_4790# 0.13856f
C2511 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ui_in[4] 1.2e-19
C2512 ringtest_0.x4._22_ a_25547_4612# 0.002069f
C2513 uio_in[3] uio_in[2] 0.031023f
C2514 a_21981_8976# a_21395_6940# 1.29e-20
C2515 muxtest_0.x1.x4.A ua[3] 6.48818f
C2516 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.173286f
C2517 muxtest_0.x2.nselect2 VDPWR 1.22451f
C2518 a_22052_8875# ringtest_0.x4._12_ 0.032034f
C2519 a_17231_12017# VDPWR 0.217593f
C2520 ringtest_0.x4.net8 a_26627_4246# 4.33e-20
C2521 ringtest_0.x4._11_ a_22765_4478# 0.159397f
C2522 a_24361_5340# a_24317_4942# 1.28e-19
C2523 ringtest_0.x4.net9 ringtest_0.x4._09_ 0.571636f
C2524 muxtest_0.x2.x2.GN1 ua[0] 2.35e-19
C2525 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A 0.17253f
C2526 ringtest_0.x4._11_ a_27065_5156# 3.81e-21
C2527 ringtest_0.x3.x2.GN2 m3_17036_9140# 0.099332f
C2528 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A 0.4308f
C2529 a_23770_5308# a_23899_5334# 0.062574f
C2530 ringtest_0.x4._11_ a_23949_6654# 8.65e-19
C2531 a_24536_6699# ringtest_0.x4.net8 5.83e-19
C2532 ringtest_0.x4.clknet_1_1__leaf_clk a_26269_4612# 3.29e-19
C2533 a_26640_5334# VDPWR 0.247111f
C2534 ringtest_0.x4.net6 a_25977_4220# 0.009771f
C2535 a_19114_31955# muxtest_0.x1.x3.GN1 0.012335f
C2536 a_19666_31955# a_19842_32287# 0.185422f
C2537 ringtest_0.x4._15_ a_26808_4902# 0.002208f
C2538 ringtest_0.x4.net7 ringtest_0.x4._09_ 2.46e-19
C2539 a_25336_4902# a_25149_4220# 3.07e-19
C2540 a_24336_6544# ringtest_0.x4.net6 0.001918f
C2541 a_12425_24040# muxtest_0.x2.x2.GN3 5.17e-20
C2542 muxtest_0.x2.x2.GN2 a_12977_24040# 3.11e-20
C2543 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN3 0.002859f
C2544 a_21948_5156# a_22021_4220# 3.53e-19
C2545 a_22116_4902# a_22164_4362# 5.83e-19
C2546 muxtest_0.x2.x2.GP2 ua[3] 0.085048f
C2547 a_18662_32213# ui_in[2] 4.33e-19
C2548 m3_13302_19985# m3_13316_18955# 0.003741f
C2549 ringtest_0.x4.net3 a_21587_5334# 0.003111f
C2550 a_11845_23906# ui_in[4] 0.02803f
C2551 ringtest_0.x4.counter[9] ringtest_0.x4.counter[8] 0.299988f
C2552 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN2 0.154394f
C2553 a_25149_4220# VDPWR 0.405792f
C2554 m2_18699_31802# ui_in[2] 4.4e-19
C2555 ringtest_0.x4._10_ a_21867_8054# 4.63e-20
C2556 a_21785_8054# a_21939_8054# 0.004009f
C2557 a_21465_9294# VDPWR 0.415615f
C2558 ringtest_0.x4._11_ a_24004_6128# 0.043142f
C2559 ringtest_0.x4.net9 a_27659_4246# 3.29e-19
C2560 a_26735_5156# VDPWR 0.002923f
C2561 a_22649_6244# a_22733_6244# 0.008508f
C2562 ringtest_0.x4._19_ a_24361_5340# 9.86e-21
C2563 muxtest_0.R7R8 muxtest_0.R6R7 2.27687f
C2564 a_24287_6422# ringtest_0.x4._21_ 1.26e-19
C2565 ringtest_0.x4._08_ a_25364_5878# 0.011527f
C2566 ringtest_0.x4.net2 a_21233_5340# 3.28e-19
C2567 a_24329_6640# VDPWR 0.438492f
C2568 a_22052_8875# a_22245_8054# 2.48e-20
C2569 ringtest_0.x4._12_ a_21803_8598# 1.13e-19
C2570 a_21852_8720# ringtest_0.x4._11_ 4.06e-19
C2571 ringtest_0.x4.net6 a_24986_5878# 0.001357f
C2572 muxtest_0.x1.x3.GN3 muxtest_0.R2R3 0.27459f
C2573 muxtest_0.x2.x2.GP2 m3_13316_18955# 2.65e-20
C2574 muxtest_0.x1.x3.GN3 ui_in[1] 0.273672f
C2575 ringtest_0.x4.clknet_0_clk a_25421_6641# 0.012442f
C2576 a_21465_8830# a_21561_8830# 0.310858f
C2577 ringtest_0.x4.net6 a_22139_5878# 5.63e-21
C2578 ringtest_0.x4.net2 ringtest_0.x4._11_ 0.001125f
C2579 a_22052_9116# a_22201_9142# 0.005525f
C2580 a_21981_9142# a_21780_9142# 4.67e-20
C2581 ringtest_0.x4._11_ a_23963_4790# 0.001879f
C2582 a_24699_6200# a_25168_5156# 5.18e-21
C2583 a_25364_5878# a_25336_4902# 2.72e-20
C2584 ringtest_0.x4.net11 a_26627_4246# 2.78e-19
C2585 ringtest_0.x4._16_ ringtest_0.x4._03_ 0.005745f
C2586 a_21561_9116# a_21981_9142# 0.036838f
C2587 a_21852_9416# a_22052_9116# 0.074815f
C2588 ringtest_0.x3.x1.nSEL0 m2_15612_11606# 3.43e-19
C2589 ringtest_0.x4._18_ a_21951_5878# 8.49e-20
C2590 ringtest_0.counter7 a_26895_3867# 0.110188f
C2591 ringtest_0.x3.x1.nSEL0 ui_in[3] 0.324822f
C2592 a_22224_6244# ringtest_0.x4.net5 1.47e-19
C2593 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN3 1.7e-19
C2594 ringtest_0.x4._11_ a_23381_4818# 0.163973f
C2595 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN2 0.209954f
C2596 ringtest_0.x4._18_ a_24883_6800# 2.19e-20
C2597 ringtest_0.x4.net1 a_21465_9294# 0.045364f
C2598 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN1 0.002605f
C2599 a_24545_5878# VDPWR 0.011033f
C2600 ringtest_0.x4._06_ a_23993_5654# 6.56e-20
C2601 ringtest_0.x4._15_ a_25083_4790# 7.24e-21
C2602 ringtest_0.x4._13_ a_21509_4790# 6.65e-20
C2603 ringtest_0.x4._11_ a_22181_5334# 7.61e-19
C2604 ringtest_0.x4._16_ a_23770_5308# 0.01721f
C2605 a_24536_6699# ringtest_0.x4._05_ 3.36e-19
C2606 ringtest_0.x4.net9 a_24361_5340# 5.55e-19
C2607 a_24895_4790# a_25677_5156# 3.14e-19
C2608 a_25083_4790# a_25263_5156# 0.001229f
C2609 a_25364_5878# VDPWR 1.3575f
C2610 ringtest_0.counter7 ua[1] 5.26868f
C2611 muxtest_0.x2.x2.GN4 ui_in[4] 0.063283f
C2612 ringtest_0.x4._22_ ringtest_0.x4._07_ 0.503878f
C2613 ringtest_0.x4.net2 a_21675_4790# 3.95e-20
C2614 muxtest_0.x2.nselect2 a_12849_23648# 1.29e-19
C2615 ringtest_0.drv_out a_25225_5334# 2.32e-21
C2616 ringtest_0.x4._14_ ringtest_0.x4.counter[1] 1.03e-21
C2617 a_21981_8976# VDPWR 0.211083f
C2618 ringtest_0.x4.net6 a_23899_5334# 0.044713f
C2619 ringtest_0.x4._15_ a_24715_5334# 0.019231f
C2620 ringtest_0.x4._22_ a_25055_3867# 8.8e-19
C2621 ringtest_0.x4._14_ a_22390_4566# 0.122283f
C2622 a_22116_4902# a_22373_5156# 0.036838f
C2623 a_27065_5334# ringtest_0.x4._09_ 0.001217f
C2624 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ui_in[4] 2.29e-19
C2625 ringtest_0.x4.net7 a_24361_5340# 0.088061f
C2626 a_21785_5878# a_24004_6128# 1.89e-21
C2627 a_22399_8976# ringtest_0.x4._11_ 0.001319f
C2628 ringtest_0.x4._04_ a_24070_5852# 8.65e-21
C2629 muxtest_0.R6R7 muxtest_0.R5R6 2.03637f
C2630 a_24135_3867# a_25055_3867# 1.37e-20
C2631 a_24551_4790# VDPWR 9.47e-20
C2632 muxtest_0.x1.x3.GP2 muxtest_0.R2R3 4.15159f
C2633 ringtest_0.x4.net8 a_26721_4246# 6.89e-20
C2634 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 5.04e-19
C2635 ringtest_0.x4._11_ a_26375_4612# 0.001561f
C2636 ringtest_0.x4._17_ a_24361_5340# 1.12e-20
C2637 muxtest_0.x1.x3.GP2 ui_in[1] 3.1e-20
C2638 a_21465_8830# a_21049_8598# 5.03e-19
C2639 ringtest_0.counter3 a_22765_4478# 8.56e-20
C2640 muxtest_0.x1.x3.GP3 muxtest_0.x1.x5.A 0.358703f
C2641 a_21561_8830# a_21780_8964# 0.006169f
C2642 a_24317_4942# VDPWR 0.226919f
C2643 muxtest_0.x1.x3.GN4 muxtest_0.R7R8 0.13848f
C2644 muxtest_0.R6R7 VDPWR 1.6078f
C2645 a_26808_5308# a_27191_5712# 4.67e-20
C2646 a_26367_5340# ringtest_0.x4.net10 5.04e-19
C2647 a_22399_9142# a_21852_8720# 4.5e-20
C2648 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A 5.04e-19
C2649 a_24329_6640# ringtest_0.x4._21_ 8.19e-20
C2650 ringtest_0.x4.clknet_1_0__leaf_clk a_21845_8816# 0.683552f
C2651 ringtest_0.x4.net4 a_22164_4362# 0.007901f
C2652 ringtest_0.x4.net2 a_21785_5878# 2.26e-20
C2653 a_23151_5334# VDPWR 0.009139f
C2654 ringtest_0.x4._15_ a_25547_4612# 5.62e-21
C2655 ua[3] ua[0] 1.8361f
C2656 ringtest_0.x4.net1 a_21981_8976# 0.001727f
C2657 ringtest_0.x4._11_ ringtest_0.x4._20_ 0.174111f
C2658 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP2 1.7e-20
C2659 ringtest_0.x4.net2 a_22399_9142# 1.04e-19
C2660 ringtest_0.x4.clknet_1_1__leaf_clk a_24883_6800# 3.41e-20
C2661 ringtest_0.x4._09_ a_26627_4246# 0.001692f
C2662 a_21425_9686# a_21465_9294# 1.32e-19
C2663 ringtest_0.x4._00_ a_21507_9686# 6.18e-19
C2664 ringtest_0.x4._09_ a_27149_5156# 6.12e-19
C2665 ringtest_0.x4._04_ a_22373_5156# 0.001409f
C2666 ringtest_0.x4._07_ a_25225_5334# 0.009837f
C2667 ringtest_0.x4._22_ a_26201_5340# 5.82e-21
C2668 ringtest_0.x4._02_ a_21399_5340# 0.275992f
C2669 a_21233_5340# a_21840_5308# 0.141453f
C2670 ringtest_0.x4.clknet_1_0__leaf_clk a_22373_5156# 6.12e-19
C2671 ringtest_0.x3.x2.GP2 ua[1] 0.349381f
C2672 ringtest_0.counter7 a_26555_4790# 2.77e-20
C2673 muxtest_0.R3R4 muxtest_0.x2.x2.GP3 4.09931f
C2674 ringtest_0.x4._18_ a_24045_6654# 2.33e-19
C2675 a_23349_6422# a_24329_6640# 6.46e-21
C2676 a_22228_8598# VDPWR 0.004407f
C2677 ringtest_0.x4._21_ a_24545_5878# 0.053333f
C2678 a_16755_12091# ringtest_0.x3.x2.GP2 3.2e-20
C2679 a_23879_6940# a_24329_6640# 0.022305f
C2680 ringtest_0.x4.clknet_1_0__leaf_clk a_21767_5334# 0.001355f
C2681 ringtest_0.x4._11_ a_21840_5308# 0.005658f
C2682 a_13675_24012# ua[3] 3.17e-19
C2683 ringtest_0.x4._20_ a_25761_5058# 3.47e-20
C2684 a_26913_4566# VDPWR 4.51e-19
C2685 ringtest_0.x4.net10 a_27065_5156# 0.003817f
C2686 muxtest_0.x2.x2.GN3 ua[3] 0.087947f
C2687 ringtest_0.ring_out VDPWR 4.36398f
C2688 ringtest_0.counter3 m3_17032_8096# 0.119717f
C2689 a_25364_5878# ringtest_0.x4._21_ 3.33e-20
C2690 a_16027_11759# a_16203_12091# 0.185422f
C2691 a_22116_4902# a_22499_4790# 4.67e-20
C2692 a_24135_3867# ringtest_0.x4.counter[5] 4.98e-19
C2693 ringtest_0.x4.clknet_1_1__leaf_clk a_26808_5308# 5.16e-19
C2694 ringtest_0.x4._08_ ringtest_0.x4.net9 0.003243f
C2695 ringtest_0.x4._19_ VDPWR 0.197759f
C2696 ringtest_0.x4.net6 a_22097_5334# 5.09e-19
C2697 ringtest_0.x4.clknet_0_clk a_26007_6788# 5.18e-20
C2698 ringtest_0.x4.net6 ringtest_0.x4._16_ 0.291584f
C2699 muxtest_0.x1.x3.GN4 muxtest_0.R5R6 0.304696f
C2700 ringtest_0.x4.clknet_1_0__leaf_clk a_22201_8964# 4.64e-19
C2701 muxtest_0.x2.x2.GN3 m3_13316_18955# 0.016026f
C2702 ringtest_0.x4._23_ a_26895_3867# 7.52e-20
C2703 a_27273_4220# a_27303_4246# 0.025037f
C2704 ringtest_0.x4.net2 ringtest_0.counter3 0.003151f
C2705 a_23879_6940# a_24545_5878# 2.81e-20
C2706 ringtest_0.x4._16_ a_24895_4790# 4.88e-21
C2707 a_26735_5334# VDPWR 0.002923f
C2708 ringtest_0.x4.net9 a_25336_4902# 0.007121f
C2709 a_21840_5308# a_21675_4790# 3.46e-19
C2710 a_21399_5340# a_22116_4902# 0.001879f
C2711 ringtest_0.counter7 m3_17046_7066# 0.117708f
C2712 ringtest_0.drv_out ringtest_0.x4._15_ 0.005511f
C2713 ringtest_0.x4.net7 ringtest_0.x4._08_ 1.97e-19
C2714 ringtest_0.x4._00_ a_21852_8720# 4.06e-19
C2715 ringtest_0.counter7 ringtest_0.x4.counter[6] 0.087745f
C2716 muxtest_0.x1.x3.GN4 VDPWR 1.35388f
C2717 ringtest_0.x4._21_ a_24317_4942# 0.011629f
C2718 a_22265_5308# a_22223_5712# 7.84e-20
C2719 a_25393_5308# a_26367_5340# 2.73e-19
C2720 a_25225_5334# a_26201_5340# 1.07e-19
C2721 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN2 0.142718f
C2722 ringtest_0.x4._19_ ringtest_0.x4._25_ 9.05e-21
C2723 a_22265_5308# VDPWR 0.421579f
C2724 ringtest_0.x4.net2 ringtest_0.x4._00_ 0.002662f
C2725 a_23529_6422# a_23619_6788# 0.004764f
C2726 ringtest_0.x4.clknet_1_1__leaf_clk a_26555_4790# 6.27e-19
C2727 muxtest_0.x1.x1.nSEL1 a_19666_31955# 7.84e-19
C2728 ringtest_0.x4.net4 a_22373_5156# 0.022715f
C2729 ringtest_0.x4.net7 a_25336_4902# 0.005145f
C2730 ringtest_0.x4.net3 ringtest_0.x4._03_ 0.019455f
C2731 ringtest_0.x4.net9 VDPWR 0.964697f
C2732 a_24045_6654# ringtest_0.x4.clknet_1_1__leaf_clk 1.54e-20
C2733 ui_in[6] ui_in[5] 6.50488f
C2734 a_21509_4790# a_22390_4566# 3.11e-19
C2735 ringtest_0.x3.x2.GN2 ua[1] 0.42933f
C2736 ringtest_0.x4._06_ a_23837_5878# 4.79e-19
C2737 ringtest_0.x4._06_ ringtest_0.x4._22_ 0.004416f
C2738 a_16579_11759# ringtest_0.x3.x2.GN4 6.84e-19
C2739 ringtest_0.x4._04_ a_21399_5340# 0.011144f
C2740 a_24070_5852# a_23837_5878# 0.005961f
C2741 a_16755_12091# ringtest_0.x3.x2.GN2 5.62e-20
C2742 a_21785_5878# a_21840_5308# 0.002941f
C2743 a_24699_6200# a_24763_6143# 0.266837f
C2744 a_21863_4790# ringtest_0.x4.net5 2.02e-19
C2745 ringtest_0.x4._23_ a_26808_5308# 0.006211f
C2746 muxtest_0.R3R4 muxtest_0.R2R3 2.48395f
C2747 ringtest_0.x4.clknet_1_0__leaf_clk a_21399_5340# 0.158653f
C2748 ringtest_0.x4._18_ a_22795_5334# 4.57e-20
C2749 a_26808_5308# a_26367_4790# 2.96e-21
C2750 ringtest_0.x4.net7 VDPWR 1.83862f
C2751 a_26367_5340# a_26808_4902# 2.96e-21
C2752 a_26201_5340# a_26640_5156# 1.73e-19
C2753 ringtest_0.x4._11_ a_22392_5990# 0.032361f
C2754 a_21561_9116# ui_in[5] 2.06e-20
C2755 a_24336_6544# a_24527_5340# 6.46e-19
C2756 ringtest_0.x4.net3 a_21939_8054# 8.45e-20
C2757 a_24329_6640# a_24968_5308# 2.9e-20
C2758 ringtest_0.x4._15_ ringtest_0.x4._07_ 0.022092f
C2759 a_24536_6699# a_24361_5340# 2.08e-22
C2760 a_27273_4220# ringtest_0.x4.counter[8] 0.001844f
C2761 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.173286f
C2762 muxtest_0.x1.x3.GN3 ui_in[4] 7.93e-20
C2763 ringtest_0.x4._17_ VDPWR 2.38225f
C2764 ringtest_0.x4._07_ a_25263_5156# 2.91e-19
C2765 ringtest_0.x3.x2.GP2 m3_17046_7066# 2.65e-20
C2766 ringtest_0.x3.x1.nSEL1 VDPWR 0.646724f
C2767 ringtest_0.x4._19_ ringtest_0.x4._21_ 7.87e-20
C2768 ringtest_0.x4.clknet_0_clk a_24336_6544# 0.025079f
C2769 ringtest_0.x4.net6 a_22649_6244# 0.021756f
C2770 ui_in[3] ua[1] 4.1e-22
C2771 ringtest_0.x3.x2.GP3 ringtest_0.counter3 4.0653f
C2772 ringtest_0.x4.clknet_1_1__leaf_clk a_24699_6200# 7.2e-19
C2773 ringtest_0.x4._00_ a_22399_8976# 0.001531f
C2774 a_21561_9116# ringtest_0.x4._12_ 1.23e-19
C2775 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y 0.17253f
C2776 a_23963_4790# ringtest_0.x4.counter[4] 4.17e-20
C2777 ui_in[1] ui_in[5] 0.187526f
C2778 ringtest_0.x4._09_ a_26721_4246# 2.04e-21
C2779 ringtest_0.x4.net8 a_24729_4790# 0.009204f
C2780 a_16755_12091# ui_in[3] 0.279858f
C2781 a_22021_4220# a_22164_4362# 0.221119f
C2782 ringtest_0.x4.net7 ringtest_0.x4._25_ 3.01e-19
C2783 ringtest_0.x4._23_ a_26555_4790# 0.012973f
C2784 a_27065_5156# a_27191_4790# 0.006169f
C2785 ringtest_0.x4.net4 a_22499_4790# 0.00133f
C2786 a_26367_4790# a_26555_4790# 0.097994f
C2787 a_26808_4902# a_27065_5156# 0.036838f
C2788 a_24329_6640# a_25925_6788# 2.69e-21
C2789 ringtest_0.x4._17_ ringtest_0.x4._25_ 1.89e-19
C2790 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP1 2.55932f
C2791 ringtest_0.x4._06_ a_25225_5334# 9.38e-20
C2792 a_23349_6422# ringtest_0.x4._19_ 0.001413f
C2793 ringtest_0.x4._11_ a_26640_5334# 6.96e-20
C2794 a_24699_6200# a_24800_5334# 0.001605f
C2795 a_23879_6940# ringtest_0.x4._19_ 5.98e-19
C2796 ringtest_0.x4.counter[0] VDPWR 0.661077f
C2797 a_12297_23648# muxtest_0.x2.x2.GN2 0.106178f
C2798 a_22817_6146# VDPWR 0.386139f
C2799 ringtest_0.x4.clknet_1_1__leaf_clk a_23809_4790# 2.42e-19
C2800 ringtest_0.x4._08_ a_27065_5334# 0.013878f
C2801 ringtest_0.x4._21_ ringtest_0.x4.net9 0.170283f
C2802 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR 0.787508f
C2803 a_26095_6788# VDPWR 0.002069f
C2804 ringtest_0.x4.net4 a_21399_5340# 0.002039f
C2805 ringtest_0.x3.nselect2 ui_in[4] 0.001177f
C2806 ringtest_0.x4.clknet_1_1__leaf_clk a_22795_5334# 7.11e-20
C2807 ringtest_0.x4._15_ a_26201_5340# 0.069151f
C2808 ringtest_0.x4.net6 a_21587_5334# 1.35e-20
C2809 ringtest_0.x3.x1.nSEL0 a_16027_11759# 0.03096f
C2810 ringtest_0.x4._22_ a_26269_4612# 6.12e-20
C2811 ringtest_0.x4._13_ a_22350_5878# 2.65e-20
C2812 a_17405_12123# VDPWR 7.45e-19
C2813 ua[2] ua[5] 0.002786f
C2814 ringtest_0.x4._04_ a_21951_5878# 0.215918f
C2815 a_21785_5878# a_22392_5990# 0.136461f
C2816 ringtest_0.x3.x2.GN3 VDPWR 0.649844f
C2817 muxtest_0.x1.x3.GP1 ua[3] 0.0076f
C2818 ringtest_0.x4._01_ ringtest_0.x4._12_ 0.353697f
C2819 ringtest_0.x4._11_ a_25149_4220# 2.67e-19
C2820 a_25925_6788# a_25364_5878# 0.010774f
C2821 ringtest_0.x4.net7 ringtest_0.x4._21_ 0.326643f
C2822 ringtest_0.x4.clknet_1_0__leaf_clk a_21951_5878# 0.020113f
C2823 ringtest_0.x3.x2.GN4 m3_17032_8096# 7.07e-19
C2824 a_26749_6422# a_26839_6788# 0.004764f
C2825 a_18662_32213# ui_in[1] 0.02803f
C2826 ringtest_0.x4._16_ ringtest_0.x4.net5 0.096932f
C2827 ringtest_0.x4._08_ a_27149_5156# 1.22e-19
C2828 ringtest_0.x4._17_ ringtest_0.x4._21_ 0.019243f
C2829 a_23879_6940# ringtest_0.x4.net9 1.97e-19
C2830 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A 0.428132f
C2831 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP3 0.060268f
C2832 ringtest_0.x4._11_ a_24329_6640# 2.33e-19
C2833 a_20318_32213# a_20492_32319# 0.006584f
C2834 a_27065_5334# VDPWR 0.233266f
C2835 ringtest_0.x4._15_ a_22164_4362# 4.86e-20
C2836 ringtest_0.x4.net6 a_27273_4220# 4.97e-21
C2837 m2_18699_31802# ui_in[1] 0.183786f
C2838 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ui_in[3] 1.1e-22
C2839 a_19666_31955# muxtest_0.x1.x3.GN1 7.37e-20
C2840 muxtest_0.x1.x5.GN a_18662_32213# 0.001336f
C2841 a_24465_6800# ringtest_0.x4.net6 0.001158f
C2842 ringtest_0.x4.clknet_1_1__leaf_clk a_25421_6641# 0.035969f
C2843 a_23529_6422# ringtest_0.x4._15_ 2e-21
C2844 a_13501_23906# muxtest_0.R1R2 5.05e-21
C2845 a_23349_6422# ringtest_0.x4.net7 2.88e-19
C2846 a_23879_6940# ringtest_0.x4.net7 0.002812f
C2847 muxtest_0.x1.x5.GN m2_18699_31802# 4e-19
C2848 muxtest_0.x1.x3.GN3 ui_in[0] 0.254198f
C2849 a_19290_32287# ui_in[2] 1.22e-19
C2850 ringtest_0.x4._17_ a_23349_6422# 0.250762f
C2851 a_23879_6940# ringtest_0.x4._17_ 7.15e-19
C2852 a_12473_23980# ui_in[4] 0.254026f
C2853 ringtest_0.x4.net7 a_25309_5334# 0.001255f
C2854 ringtest_0.x4._11_ a_24545_5878# 1.22e-19
C2855 a_22201_9142# VDPWR 0.003202f
C2856 a_26627_4246# VDPWR 0.152186f
C2857 a_21852_9416# VDPWR 0.335402f
C2858 a_22817_6146# ringtest_0.x4._21_ 1.76e-19
C2859 a_27149_5156# VDPWR 0.005629f
C2860 ui_in[2] ui_in[3] 0.170107f
C2861 ringtest_0.x4._11_ a_25364_5878# 0.049204f
C2862 muxtest_0.x1.x3.GN2 muxtest_0.R1R2 0.006936f
C2863 a_24536_6699# VDPWR 0.266088f
C2864 muxtest_0.x1.x5.A muxtest_0.R6R7 4.52052f
C2865 ringtest_0.x4._01_ a_22245_8054# 0.014882f
C2866 ringtest_0.x4._12_ a_21785_8054# 0.001375f
C2867 ringtest_0.x4.net4 a_21951_5878# 0.34974f
C2868 ringtest_0.x4._15_ ringtest_0.x4._06_ 0.139237f
C2869 a_21561_8830# a_21845_8816# 0.030894f
C2870 ringtest_0.x4._15_ a_24070_5852# 6.77e-20
C2871 a_21465_8830# a_21852_8720# 0.034054f
C2872 ringtest_0.x4.net8 ringtest_0.x4._09_ 2.1e-20
C2873 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y 5.04e-19
C2874 ringtest_0.x4._23_ a_26817_4566# 4.18e-19
C2875 a_25149_4220# a_25345_4612# 0.00119f
C2876 ringtest_0.x4._11_ a_24551_4790# 0.001398f
C2877 a_25593_5156# ringtest_0.x4.counter[6] 2e-19
C2878 a_25364_5878# a_25761_5058# 0.001883f
C2879 a_21845_9116# a_21981_9142# 0.141453f
C2880 a_21233_5340# a_23151_5334# 4.04e-20
C2881 a_21852_9416# a_21803_9508# 6.32e-19
C2882 a_21675_9686# ringtest_0.x4.clknet_1_0__leaf_clk 2.59e-19
C2883 ringtest_0.x4.net2 a_21465_8830# 0.004306f
C2884 ringtest_0.x4._18_ a_22224_6244# 5.13e-20
C2885 a_22649_6244# ringtest_0.x4.net5 4.89e-20
C2886 ringtest_0.x4._11_ a_24317_4942# 0.046716f
C2887 a_25421_6641# ringtest_0.x4._23_ 1.03e-19
C2888 ringtest_0.x4._05_ a_26749_6422# 4.21e-20
C2889 ringtest_0.x4.net1 a_21852_9416# 0.006588f
C2890 a_22111_10993# a_21845_9116# 6.9e-23
C2891 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._24_ 0.041474f
C2892 ringtest_0.x4.net10 a_27489_3702# 1.3e-21
C2893 ringtest_0.x4._14_ VDPWR 0.685574f
C2894 ringtest_0.x4.net6 a_26201_4790# 5.6e-22
C2895 ringtest_0.x4._15_ a_23891_4790# 1.25e-19
C2896 ringtest_0.x4._11_ a_23151_5334# 0.00137f
C2897 ringtest_0.x4._16_ a_24527_5340# 9.89e-20
C2898 a_13025_23980# muxtest_0.x2.x2.GP3 5.21e-19
C2899 ringtest_0.x4.net9 a_24968_5308# 2.05e-20
C2900 muxtest_0.x1.x3.GP2 ui_in[0] 4.71e-19
C2901 a_22319_6244# VDPWR 0.003961f
C2902 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP3 3.4436f
C2903 a_25336_4902# a_25294_4790# 4.62e-19
C2904 a_24895_4790# a_26201_4790# 3.23e-19
C2905 ringtest_0.x4._15_ a_22373_5156# 1.6e-20
C2906 muxtest_0.x2.nselect2 a_13501_23906# 9.77e-20
C2907 ringtest_0.x4.clknet_0_clk ringtest_0.x4._16_ 0.019509f
C2908 ringtest_0.x4.net5 a_23467_4818# 2.72e-19
C2909 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR 0.639974f
C2910 ringtest_0.x4.net6 a_26555_5334# 3.93e-20
C2911 muxtest_0.R7R8 muxtest_0.x2.x2.GN2 1.22e-19
C2912 ringtest_0.x4._22_ a_26895_3867# 1.85e-19
C2913 a_22392_5990# a_22775_5878# 4.67e-20
C2914 muxtest_0.R3R4 ui_in[4] 3.8e-21
C2915 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x2.GN2 3.88e-22
C2916 a_22541_5058# a_22373_5156# 0.310858f
C2917 clk ena 0.031023f
C2918 ringtest_0.x4.net7 a_24968_5308# 0.040813f
C2919 a_24883_6800# ringtest_0.x4._22_ 0.001069f
C2920 a_21785_8054# a_22245_8054# 0.001479f
C2921 ringtest_0.x4._12_ a_22695_8304# 0.001754f
C2922 a_25055_3867# a_25975_3867# 1.37e-20
C2923 a_25294_4790# VDPWR 1.42e-19
C2924 ringtest_0.x4._17_ a_24968_5308# 1.03e-20
C2925 a_22043_5156# VDPWR 0.005794f
C2926 muxtest_0.x1.x3.GP3 muxtest_0.x1.x4.A 0.358376f
C2927 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A 0.446595f
C2928 a_26640_5334# ringtest_0.x4.net10 3.33e-19
C2929 a_27233_5308# a_27191_5712# 7.84e-20
C2930 ringtest_0.x4.clknet_1_0__leaf_clk a_22052_8875# 0.037641f
C2931 ringtest_0.x4.net4 a_23381_4584# 0.083888f
C2932 a_24536_6699# ringtest_0.x4._21_ 0.0043f
C2933 ui_in[4] ui_in[5] 0.278355f
C2934 ringtest_0.x4._11_ ringtest_0.x4._19_ 0.032711f
C2935 ringtest_0.x4._15_ a_26269_4612# 0.00403f
C2936 a_19666_31955# muxtest_0.x1.x3.GP3 0.001353f
C2937 ringtest_0.x4._23_ ringtest_0.x4._24_ 0.206353f
C2938 ringtest_0.x4.net7 a_25925_6788# 0.168744f
C2939 ringtest_0.x4._24_ a_26367_4790# 0.03707f
C2940 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ui_in[3] 0.001551f
C2941 ringtest_0.x4._00_ a_21465_9294# 0.001095f
C2942 a_21425_9686# a_21852_9416# 0.00324f
C2943 a_26749_6422# ringtest_0.x4._09_ 2.51e-21
C2944 ringtest_0.x4._09_ ringtest_0.x4.net11 0.071633f
C2945 ringtest_0.x4.net3 ringtest_0.x4.net5 9.15e-21
C2946 ringtest_0.x4._02_ a_21672_5334# 8.22e-19
C2947 a_21233_5340# a_22265_5308# 0.048748f
C2948 ringtest_0.x4._22_ a_26808_5308# 9.3e-20
C2949 ringtest_0.x4._17_ a_25925_6788# 0.139841f
C2950 ringtest_0.x4._04_ a_22795_5334# 0.072162f
C2951 ringtest_0.x4._18_ a_24336_6544# 1.59e-19
C2952 ringtest_0.x4._10_ VDPWR 0.249351f
C2953 ringtest_0.x4._20_ a_25083_4790# 5.09e-20
C2954 ringtest_0.x4.net8 a_24361_5340# 0.036074f
C2955 a_23879_6940# a_24536_6699# 0.007109f
C2956 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP2 0.005192f
C2957 ringtest_0.x4._11_ a_22265_5308# 0.033019f
C2958 a_26721_4246# VDPWR 0.191262f
C2959 muxtest_0.x1.x4.A muxtest_0.R1R2 4.5214f
C2960 muxtest_0.x2.x1.nSEL0 ui_in[4] 0.13767f
C2961 a_16203_12091# a_16579_11759# 3.02e-19
C2962 ringtest_0.x3.x1.nSEL1 a_15749_12123# 0.00175f
C2963 a_22541_5058# a_22499_4790# 7.84e-20
C2964 ringtest_0.x4._11_ ringtest_0.x4.net9 0.233741f
C2965 ringtest_0.x4.clknet_1_1__leaf_clk a_27233_5308# 9.45e-20
C2966 muxtest_0.x1.x3.GN3 muxtest_0.x2.x2.GN4 8.02e-21
C2967 a_12977_24040# VDPWR 0.001496f
C2968 ringtest_0.x4.net6 a_23770_5308# 0.050235f
C2969 ringtest_0.x4.clknet_0_clk a_26201_6788# 6.75e-20
C2970 muxtest_0.x2.x2.GN2 VDPWR 0.601936f
C2971 a_24361_5340# a_24729_4790# 0.012779f
C2972 ringtest_0.x4.net3 a_21007_3867# 0.006292f
C2973 ringtest_0.x4.clknet_1_0__leaf_clk a_21803_8598# 0.002574f
C2974 a_24045_6654# a_23837_5878# 9.42e-20
C2975 ringtest_0.x4._16_ a_25168_5156# 7.37e-22
C2976 a_24336_6544# a_24763_6143# 0.003687f
C2977 a_21509_4790# VDPWR 0.741952f
C2978 ringtest_0.x4._11_ ringtest_0.x4.net7 0.966176f
C2979 a_26640_5156# a_26895_3867# 6.36e-19
C2980 ringtest_0.x4.net9 a_25761_5058# 0.115737f
C2981 ringtest_0.x4.net11 a_27659_4246# 0.004987f
C2982 a_22265_5308# a_21675_4790# 0.00183f
C2983 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A 0.17253f
C2984 ringtest_0.x4.net1 ringtest_0.x4._10_ 0.033245f
C2985 a_25925_6788# a_26095_6788# 0.001675f
C2986 ringtest_0.x4._11_ ringtest_0.x4._17_ 0.113734f
C2987 a_26201_5340# a_26367_5340# 0.970499f
C2988 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GP1 1.17e-19
C2989 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN4 2.26e-20
C2990 a_22765_5308# VDPWR 0.252112f
C2991 ringtest_0.x4.clknet_1_1__leaf_clk a_25977_4220# 3.39e-19
C2992 a_23949_6654# a_24264_6788# 7.84e-20
C2993 ringtest_0.x4._16_ a_22983_5654# 3.98e-19
C2994 a_25364_5878# ringtest_0.x4.net10 3.58e-19
C2995 muxtest_0.x1.x5.GN a_18836_32319# 1.95e-19
C2996 ringtest_0.x4.net7 a_25761_5058# 0.064911f
C2997 ringtest_0.x4._03_ a_22939_4584# 1.17e-19
C2998 a_24336_6544# ringtest_0.x4.clknet_1_1__leaf_clk 0.013843f
C2999 a_12297_23648# muxtest_0.x2.x2.GP1 9.92e-19
C3000 a_21867_8054# VDPWR 2.01e-19
C3001 ringtest_0.x4.net4 a_22795_5334# 0.005199f
C3002 a_24627_6200# a_24545_5878# 2.78e-19
C3003 a_24763_6143# a_24986_5878# 3.74e-19
C3004 ringtest_0.x4._13_ VDPWR 0.524973f
C3005 a_17231_12017# ringtest_0.x3.x2.GN4 0.134079f
C3006 ringtest_0.x3.x2.GN2 a_16155_12151# 0.002418f
C3007 ua[3] ua[1] 0.003505f
C3008 a_21785_5878# a_22265_5308# 4.12e-19
C3009 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN2 0.065153f
C3010 ringtest_0.x4._04_ a_21672_5334# 3.3e-20
C3011 ringtest_0.x4._22_ ringtest_0.x4.counter[6] 9.35e-22
C3012 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR 0.636657f
C3013 a_24699_6200# ringtest_0.x4._22_ 0.019192f
C3014 ui_in[0] ui_in[5] 0.21609f
C3015 ringtest_0.x4._23_ a_27233_5308# 1.75e-20
C3016 ringtest_0.x4.clknet_1_0__leaf_clk a_21672_5334# 0.032164f
C3017 a_26201_5340# a_27065_5156# 1.29e-19
C3018 a_26640_5334# a_26808_4902# 3.15e-19
C3019 a_26808_5308# a_26640_5156# 3.15e-19
C3020 ringtest_0.x4._18_ a_23899_5334# 3.94e-20
C3021 ringtest_0.x4._16_ a_22486_4246# 0.00427f
C3022 muxtest_0.x1.x4.A muxtest_0.x2.nselect2 0.01287f
C3023 ringtest_0.x4._11_ a_22817_6146# 0.052724f
C3024 a_21845_9116# ui_in[5] 1.25e-19
C3025 ringtest_0.x4.net9 a_25345_4612# 0.001755f
C3026 a_24336_6544# a_24800_5334# 9.47e-20
C3027 ringtest_0.x4._08_ ringtest_0.x4.net8 2.38e-19
C3028 ringtest_0.x4._11_ a_26095_6788# 0.001703f
C3029 muxtest_0.x2.x2.GP3 ui_in[3] 4.18e-19
C3030 ringtest_0.x4.net3 ringtest_0.x4._12_ 0.271994f
C3031 ringtest_0.x4._15_ a_26895_3867# 0.006207f
C3032 muxtest_0.x1.x3.GN2 muxtest_0.R6R7 4.03742f
C3033 ringtest_0.x4.net1 a_21867_8054# 0.00162f
C3034 ringtest_0.x4.clknet_0_clk a_24465_6800# 0.003343f
C3035 a_21845_9116# ringtest_0.x4._12_ 2.52e-19
C3036 ringtest_0.x4._07_ a_23381_4818# 2.73e-21
C3037 ringtest_0.x3.x2.GN1 m2_15612_11606# 0.06935f
C3038 ringtest_0.x4._09_ a_27659_4246# 2.25e-19
C3039 ringtest_0.counter7 ringtest_0.x4.counter[9] 2.14e-19
C3040 ringtest_0.x4._23_ a_25977_4220# 0.130093f
C3041 ringtest_0.x3.x2.GN1 ui_in[3] 0.021168f
C3042 ringtest_0.x4.net8 a_25336_4902# 0.00264f
C3043 ringtest_0.drv_out ringtest_0.x3.x2.GP3 0.077808f
C3044 ringtest_0.x4._17_ a_21785_5878# 1.5e-21
C3045 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ui_in[3] 1.61e-19
C3046 muxtest_0.x1.x3.GP3 ua[0] 0.17111f
C3047 a_26640_5156# a_26555_4790# 0.037333f
C3048 a_21951_5878# a_22541_5058# 8.13e-20
C3049 a_27233_5058# a_27065_5156# 0.310858f
C3050 ringtest_0.x4.net10 a_26913_4566# 0.002966f
C3051 ringtest_0.x4.clknet_1_1__leaf_clk a_25677_5156# 1.62e-19
C3052 ringtest_0.x4.net6 a_24895_4790# 0.045685f
C3053 a_12849_23648# a_12977_24040# 0.004764f
C3054 a_25364_5878# a_25393_5308# 0.009572f
C3055 a_23529_6422# a_23949_6654# 0.017007f
C3056 ringtest_0.x4.net8 VDPWR 1.78891f
C3057 a_12849_23648# muxtest_0.x2.x2.GN2 1.63e-19
C3058 a_24729_4790# a_25336_4902# 0.141453f
C3059 ui_in[3] ui_in[6] 0.153563f
C3060 a_18662_32213# ui_in[0] 0.048888f
C3061 a_26839_6788# VDPWR 6.35e-19
C3062 ringtest_0.x4.net4 a_21672_5334# 4.27e-19
C3063 ringtest_0.x4.clknet_1_1__leaf_clk a_23899_5334# 0.001857f
C3064 ringtest_0.x4._03_ ringtest_0.x4.net5 3.86e-19
C3065 ringtest_0.x3.x1.nSEL0 a_16579_11759# 1.91e-20
C3066 ringtest_0.x4._15_ a_26808_5308# 4.57e-19
C3067 m2_18699_31802# ui_in[0] 0.130999f
C3068 ringtest_0.x4._22_ a_26817_4566# 1.37e-20
C3069 ringtest_0.x4.net10 a_26735_5334# 8.52e-20
C3070 a_21785_5878# a_22817_6146# 0.048608f
C3071 ringtest_0.x4._04_ a_22224_6244# 0.01404f
C3072 a_24729_4790# VDPWR 0.727748f
C3073 ringtest_0.x4.net3 a_22245_8054# 0.001478f
C3074 ringtest_0.x4._11_ a_26627_4246# 0.054652f
C3075 muxtest_0.R1R2 ua[0] 2.31469f
C3076 ringtest_0.x4.clknet_1_0__leaf_clk a_22224_6244# 0.002436f
C3077 a_21845_9116# a_22245_8054# 4.52e-21
C3078 ringtest_0.x4._18_ ringtest_0.x4._16_ 0.283975f
C3079 ringtest_0.x4._07_ ringtest_0.x4._20_ 1.72e-19
C3080 a_25364_5878# a_26808_4902# 7.13e-20
C3081 a_26749_6422# ringtest_0.x4._08_ 0.001905f
C3082 a_19290_32287# ui_in[1] 0.254026f
C3083 ringtest_0.x4._25_ a_26839_6788# 8.17e-20
C3084 a_24968_5308# a_25351_5712# 4.67e-20
C3085 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A 5.04e-19
C3086 ringtest_0.x4._11_ a_24536_6699# 3.53e-20
C3087 a_23949_6654# a_24070_5852# 0.002561f
C3088 a_21465_9294# a_21465_8830# 0.025128f
C3089 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GN4 0.057602f
C3090 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1 2.99928f
C3091 a_21798_5712# VDPWR 4.21e-19
C3092 a_19242_32347# VDPWR 5.13e-19
C3093 ringtest_0.x4._15_ a_23381_4584# 0.110742f
C3094 ringtest_0.x4.net9 ringtest_0.x4.net10 0.022804f
C3095 ringtest_0.x4.net6 a_27169_6641# 1.17e-21
C3096 ui_in[1] ui_in[3] 0.006066f
C3097 ui_in[2] ua[3] 0.781024f
C3098 ringtest_0.x4._15_ a_26555_4790# 0.005742f
C3099 a_25593_5156# a_25977_4220# 0.009905f
C3100 muxtest_0.x1.x5.GN a_19290_32287# 3.26e-19
C3101 a_25593_5156# a_25719_4790# 0.006169f
C3102 a_24045_6654# ringtest_0.x4._15_ 1.09e-20
C3103 ringtest_0.x4._14_ a_21233_5340# 0.001276f
C3104 a_22373_5156# a_22765_4478# 0.001309f
C3105 ringtest_0.x4.counter[1] VDPWR 0.349593f
C3106 a_24763_6143# ringtest_0.x4._16_ 0.060109f
C3107 m3_17036_9140# m3_17032_8096# 0.003764f
C3108 muxtest_0.R3R4 muxtest_0.x2.x2.GN4 0.269437f
C3109 ringtest_0.x4.net9 a_24627_6200# 0.004319f
C3110 ringtest_0.x4.net7 ringtest_0.x4.net10 6.54e-19
C3111 a_13025_23980# ui_in[4] 0.127717f
C3112 ringtest_0.x4._11_ ringtest_0.x4._14_ 0.007676f
C3113 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.nselect2 0.047548f
C3114 muxtest_0.x2.x1.nSEL0 a_11845_23906# 0.081627f
C3115 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR 0.636415f
C3116 a_22390_4566# VDPWR 0.007674f
C3117 ringtest_0.x4._16_ a_22295_3867# 4.24e-19
C3118 a_24004_6128# ringtest_0.x4._06_ 0.111795f
C3119 a_26749_6422# VDPWR 0.178246f
C3120 a_22052_9116# VDPWR 0.286747f
C3121 ringtest_0.x4.net11 VDPWR 0.794015f
C3122 ringtest_0.x4.net8 ringtest_0.x4._21_ 0.333812f
C3123 ringtest_0.x4._11_ a_22319_6244# 0.00121f
C3124 ringtest_0.counter3 ringtest_0.x4.counter[0] 0.117902f
C3125 a_24070_5852# a_24004_6128# 0.221119f
C3126 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A a_16027_11759# 2.51e-19
C3127 a_24329_6640# a_24715_5334# 6.17e-21
C3128 ringtest_0.x4._05_ VDPWR 0.240335f
C3129 ringtest_0.x4._24_ ringtest_0.x4._22_ 0.01067f
C3130 ringtest_0.x4.net4 a_22224_6244# 0.034877f
C3131 ringtest_0.x4._23_ ringtest_0.x4.counter[9] 7.62e-19
C3132 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._16_ 0.001692f
C3133 ringtest_0.x4.net3 a_21591_6128# 0.001185f
C3134 a_21465_8830# a_21981_8976# 1.28e-19
C3135 ringtest_0.x4._15_ a_24699_6200# 2.91e-20
C3136 a_21845_8816# a_21852_8720# 0.969092f
C3137 ringtest_0.x4.net6 a_23932_6128# 0.002624f
C3138 ringtest_0.x4.net3 a_22486_4246# 1.66e-19
C3139 ringtest_0.x4._17_ a_24627_6200# 4.44e-20
C3140 ringtest_0.x4._23_ a_27491_4566# 3.52e-19
C3141 a_25149_4220# a_25547_4612# 0.005781f
C3142 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP2 4.55678f
C3143 ringtest_0.x4._11_ a_25294_4790# 0.002651f
C3144 ringtest_0.x4._14_ a_21675_4790# 5.98e-19
C3145 ringtest_0.x4._21_ a_24729_4790# 5.62e-21
C3146 ringtest_0.x4.clknet_1_0__leaf_clk a_21780_9142# 0.001704f
C3147 a_26749_6422# ringtest_0.x4._25_ 0.082413f
C3148 ringtest_0.x3.x2.GN3 ringtest_0.counter3 3.89796f
C3149 ringtest_0.x4.counter[0] ua[2] 1.11e-19
C3150 a_21852_9416# a_22399_9142# 0.095025f
C3151 ringtest_0.x4._08_ ringtest_0.x4._09_ 0.013938f
C3152 a_21561_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.038899f
C3153 ringtest_0.x4.net2 a_21845_8816# 3.07e-19
C3154 a_21845_9116# a_22228_9508# 0.002698f
C3155 ringtest_0.x4._18_ a_22649_6244# 3.43e-19
C3156 a_23879_6940# ringtest_0.x4.net8 0.001938f
C3157 ringtest_0.x4._11_ a_22043_5156# 6.67e-19
C3158 ringtest_0.ring_out ringtest_0.x3.x2.GN4 0.080391f
C3159 ringtest_0.x4._05_ ringtest_0.x4._25_ 4.6e-21
C3160 ringtest_0.x4.net1 a_22052_9116# 0.002893f
C3161 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ui_in[3] 5.64e-20
C3162 ringtest_0.drv_out a_17231_12017# 3.86e-20
C3163 ringtest_0.x4.net8 a_25309_5334# 9.28e-20
C3164 ua[2] ua[4] 0.002786f
C3165 ringtest_0.x4._16_ a_24800_5334# 0.00213f
C3166 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP3 0.002439f
C3167 ringtest_0.x4.net9 a_25393_5308# 0.007609f
C3168 ringtest_0.x4._08_ a_26766_5712# 0.001882f
C3169 a_22350_5878# VDPWR 3.37e-19
C3170 a_25593_5156# a_25677_5156# 0.008508f
C3171 ringtest_0.x4.clknet_0_clk a_23770_5308# 8.98e-21
C3172 ringtest_0.x4.net6 ringtest_0.x4.net5 0.003368f
C3173 ringtest_0.x4._15_ a_23809_4790# 0.080244f
C3174 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN4 2.26e-20
C3175 muxtest_0.x2.nselect2 muxtest_0.x2.x2.GN3 7.39e-21
C3176 ringtest_0.x3.x2.GP2 ui_in[4] 1.37e-19
C3177 ringtest_0.x4.net6 a_24895_5334# 0.001259f
C3178 a_22817_6146# a_22775_5878# 7.84e-20
C3179 a_17377_14114# ui_in[6] 0.040112f
C3180 ringtest_0.x4.counter[1] ringtest_0.x4.counter[2] 0.070133f
C3181 a_22116_4902# a_21863_4790# 3.39e-19
C3182 a_22541_5058# a_23809_4790# 3.71e-21
C3183 ringtest_0.x3.x1.nSEL1 a_15575_12017# 0.193944f
C3184 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A a_16579_11759# 2.51e-19
C3185 ringtest_0.x4.net7 a_25393_5308# 0.08513f
C3186 muxtest_0.x2.x2.GP1 VDPWR 1.85798f
C3187 a_25975_3867# a_26895_3867# 1.37e-20
C3188 a_21785_5878# a_22319_6244# 0.002698f
C3189 ringtest_0.x4._09_ VDPWR 0.262387f
C3190 ringtest_0.x4._04_ a_22139_5878# 0.126198f
C3191 ringtest_0.x4._10_ ringtest_0.x4._11_ 0.033565f
C3192 ringtest_0.x4._11_ a_26721_4246# 0.039972f
C3193 a_22795_5334# a_22541_5058# 0.001352f
C3194 ringtest_0.x4._23_ ringtest_0.x4._16_ 3.32e-22
C3195 ringtest_0.x4.net9 a_27191_4790# 6.87e-19
C3196 a_12297_23648# VDPWR 0.161892f
C3197 ringtest_0.x4._17_ a_25393_5308# 4.35e-22
C3198 ringtest_0.x4.clknet_1_0__leaf_clk a_22139_5878# 0.003123f
C3199 a_21852_8720# a_22201_8964# 2.36e-19
C3200 a_21981_8976# a_21780_8964# 4.67e-20
C3201 a_21845_8816# a_22399_8976# 0.057611f
C3202 a_21561_8830# a_21803_8598# 0.008508f
C3203 a_22074_4790# VDPWR 0.003212f
C3204 ringtest_0.x4.net9 a_26808_4902# 0.022365f
C3205 ringtest_0.x3.x2.GP3 m3_17036_9140# 9.67e-19
C3206 a_27065_5334# ringtest_0.x4.net10 0.00375f
C3207 a_23993_5654# a_23899_5334# 1.26e-19
C3208 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A 0.446529f
C3209 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP3 0.061475f
C3210 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._01_ 0.05158f
C3211 a_12019_24012# ui_in[3] 9.55e-19
C3212 a_21233_5340# a_21509_4790# 0.001876f
C3213 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A 0.17253f
C3214 ringtest_0.x4._15_ a_26817_4566# 0.004129f
C3215 a_19666_31955# muxtest_0.x1.x3.GN4 6.84e-19
C3216 ringtest_0.drv_out a_24329_6640# 4.16e-19
C3217 ringtest_0.x4._24_ a_26640_5156# 0.010089f
C3218 ringtest_0.x4._00_ a_21852_9416# 0.208988f
C3219 ringtest_0.x4._11_ a_21509_4790# 0.005486f
C3220 ringtest_0.x4.net7 a_26808_4902# 1.23e-19
C3221 ringtest_0.x4.net3 ringtest_0.counter7 4.2e-20
C3222 a_21233_5340# a_22765_5308# 1.05e-19
C3223 ringtest_0.x4._02_ a_22097_5334# 3.18e-19
C3224 ringtest_0.x4.net5 a_22939_4584# 0.002311f
C3225 ringtest_0.x4.clknet_1_0__leaf_clk a_21863_4790# 0.003207f
C3226 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP2 0.043302f
C3227 ringtest_0.x4._16_ ringtest_0.x4._02_ 3.22e-20
C3228 ringtest_0.x4._18_ a_24465_6800# 7.52e-20
C3229 ringtest_0.x4.net10 a_26627_4246# 0.27342f
C3230 a_23349_6422# ringtest_0.x4._05_ 4.45e-20
C3231 a_23879_6940# ringtest_0.x4._05_ 0.005813f
C3232 ringtest_0.x4.net8 a_24968_5308# 0.001066f
C3233 a_18836_32319# ui_in[0] 9.55e-19
C3234 ringtest_0.x4._11_ a_22765_5308# 0.001227f
C3235 a_27659_4246# VDPWR 0.009314f
C3236 ringtest_0.x4.net10 a_27149_5156# 3.08e-19
C3237 ringtest_0.x3.x2.GN2 ui_in[4] 0.108649f
C3238 a_16027_11759# a_16155_12151# 0.004764f
C3239 ringtest_0.x4._08_ a_24361_5340# 3.42e-20
C3240 a_16027_11759# ringtest_0.x3.x2.GN1 0.012445f
C3241 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR 0.636415f
C3242 a_16579_11759# a_16755_12091# 0.185422f
C3243 ringtest_0.x4._13_ a_21233_5340# 3.88e-19
C3244 muxtest_0.x1.x3.GP1 muxtest_0.R1R2 2.46e-21
C3245 ringtest_0.x4._11_ a_21867_8054# 1.17e-19
C3246 ringtest_0.x4._07_ a_25149_4220# 9.24e-19
C3247 uio_in[2] uio_in[1] 0.031023f
C3248 a_21509_4790# a_21675_4790# 0.970278f
C3249 ringtest_0.x4.net6 a_24527_5340# 0.048602f
C3250 a_21375_3867# ringtest_0.x4.counter[1] 0.1107f
C3251 ringtest_0.x4.clknet_0_clk a_24712_6422# 4.01e-19
C3252 ringtest_0.drv_out a_25364_5878# 1.27e-19
C3253 ringtest_0.x4._22_ a_25977_4220# 0.191159f
C3254 ringtest_0.x4.net4 a_22139_5878# 0.011292f
C3255 ringtest_0.x4._11_ ringtest_0.x4._13_ 0.217373f
C3256 a_24361_5340# a_25336_4902# 3.92e-19
C3257 ringtest_0.x4._22_ a_25719_4790# 7.63e-20
C3258 a_24968_5308# a_24729_4790# 1.62e-19
C3259 a_24527_5340# a_24895_4790# 1.17e-19
C3260 muxtest_0.x1.x3.GN3 muxtest_0.R3R4 0.377005f
C3261 ringtest_0.x4.net3 a_22295_3867# 0.001252f
C3262 ringtest_0.x4.clknet_1_0__leaf_clk a_21785_8054# 0.024338f
C3263 a_25149_4220# a_25055_3867# 3.27e-19
C3264 a_24329_6640# ringtest_0.x4._07_ 5.99e-19
C3265 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net6 0.087511f
C3266 a_24336_6544# ringtest_0.x4._22_ 8.56e-19
C3267 ringtest_0.x4.net9 a_25083_4790# 1.61e-19
C3268 a_27233_5058# a_27489_3702# 3.35e-20
C3269 a_22265_5308# a_21948_5156# 0.005602f
C3270 a_22097_5334# a_22116_4902# 3.73e-19
C3271 ringtest_0.x4.clknet_0_clk a_24895_4790# 3.43e-21
C3272 ringtest_0.x4._18_ a_22733_6244# 1.72e-19
C3273 m2_15612_11606# ui_in[4] 0.183786f
C3274 ringtest_0.x4._16_ a_22116_4902# 0.005579f
C3275 a_26367_5340# a_26808_5308# 0.118966f
C3276 a_26201_5340# a_26640_5334# 0.273138f
C3277 a_21399_5340# a_22181_5334# 6.32e-19
C3278 ui_in[3] ui_in[4] 13.523f
C3279 ringtest_0.x4._15_ ringtest_0.x4._24_ 0.032103f
C3280 a_24361_5340# VDPWR 0.421866f
C3281 ringtest_0.x4._16_ a_23993_5654# 3.31e-19
C3282 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ui_in[3] 9.57e-20
C3283 ringtest_0.x4.net4 a_21863_4790# 4.45e-19
C3284 ringtest_0.x4.net9 a_24715_5334# 1.41e-19
C3285 a_21785_5878# a_21509_4790# 2.82e-20
C3286 ringtest_0.x4.net7 a_25083_4790# 4.68e-19
C3287 a_12849_23648# muxtest_0.x2.x2.GP1 1.21e-20
C3288 a_24465_6800# ringtest_0.x4.clknet_1_1__leaf_clk 1.17e-20
C3289 a_21395_6940# VDPWR 1.52032f
C3290 ringtest_0.counter7 a_26201_4790# 2.09e-20
C3291 ringtest_0.x3.x2.GN4 a_17405_12123# 0.001562f
C3292 ringtest_0.x4._22_ a_24986_5878# 0.006962f
C3293 muxtest_0.x2.x2.GP3 ua[3] 0.084041f
C3294 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP1 2.56189f
C3295 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GN4 0.071282f
C3296 a_21132_8918# VDPWR 4.93e-19
C3297 muxtest_0.x1.x1.nSEL1 ui_in[2] 0.164995f
C3298 ringtest_0.x4._04_ a_22097_5334# 0.001211f
C3299 a_21785_5878# a_22765_5308# 0.002539f
C3300 a_25364_5878# ringtest_0.x4._07_ 0.022424f
C3301 ringtest_0.x4.net7 a_24715_5334# 0.014734f
C3302 ringtest_0.x4._04_ ringtest_0.x4._16_ 0.025302f
C3303 ringtest_0.x4.clknet_1_0__leaf_clk a_22097_5334# 0.004501f
C3304 a_25975_3867# ringtest_0.x4.counter[6] 0.1107f
C3305 a_26367_5340# a_26555_4790# 1.41e-20
C3306 ringtest_0.x4._11_ ringtest_0.x4.net8 0.418201f
C3307 ringtest_0.x4.net9 a_25547_4612# 6.77e-19
C3308 a_21951_5878# a_24004_6128# 1.23e-20
C3309 a_21981_9142# ui_in[5] 2.79e-20
C3310 muxtest_0.R7R8 muxtest_0.R5R6 0.318606f
C3311 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._16_ 4.14e-20
C3312 ringtest_0.x4._05_ a_24968_5308# 8.7e-19
C3313 muxtest_0.x1.x3.GP2 muxtest_0.R3R4 0.170487f
C3314 ringtest_0.x4._13_ a_21785_5878# 0.002226f
C3315 muxtest_0.x2.x2.GP3 m3_13316_18955# 0.006132f
C3316 a_22111_10993# ui_in[5] 0.231636f
C3317 ringtest_0.ring_out ringtest_0.drv_out 2.13841f
C3318 muxtest_0.x1.x3.GN1 muxtest_0.R4R5 0.334962f
C3319 ringtest_0.x4.net1 a_21395_6940# 0.001584f
C3320 muxtest_0.R7R8 VDPWR 3.21675f
C3321 a_21981_9142# ringtest_0.x4._12_ 7.61e-20
C3322 ringtest_0.x4._07_ a_24317_4942# 1.81e-19
C3323 ringtest_0.x3.x2.GP1 ui_in[3] 8.3e-19
C3324 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A 5.04e-19
C3325 ringtest_0.x4._23_ a_27273_4220# 0.220841f
C3326 ringtest_0.x4.net1 a_21132_8918# 0.001512f
C3327 ringtest_0.x4.net7 a_25547_4612# 0.001525f
C3328 a_22765_4478# a_23381_4584# 0.013543f
C3329 ringtest_0.drv_out ringtest_0.x4._19_ 0.013619f
C3330 ringtest_0.x4.net8 a_25761_5058# 0.020836f
C3331 ringtest_0.x4._11_ a_24729_4790# 0.029022f
C3332 a_26808_4902# a_26627_4246# 3.15e-19
C3333 ringtest_0.x4._23_ a_26766_4790# 6.82e-19
C3334 a_19114_31955# a_19242_32347# 0.004764f
C3335 ringtest_0.x4._02_ a_21587_5334# 0.114994f
C3336 a_26808_4902# a_27149_5156# 9.73e-19
C3337 a_22224_6244# a_22541_5058# 2.18e-19
C3338 ringtest_0.x4._05_ a_25925_6788# 1.27e-19
C3339 muxtest_0.x1.x3.GN4 ua[0] 4.10932f
C3340 a_21399_5340# a_21840_5308# 0.127288f
C3341 ringtest_0.x4.clknet_1_1__leaf_clk a_26201_4790# 0.306202f
C3342 ringtest_0.x4.net10 a_26721_4246# 0.007482f
C3343 ringtest_0.x4.net6 a_25168_5156# 6.05e-21
C3344 a_13025_23980# muxtest_0.x2.x2.GN4 0.003699f
C3345 ringtest_0.x4._11_ a_21798_5712# 4.01e-19
C3346 ringtest_0.x4._21_ a_24361_5340# 0.016583f
C3347 a_25364_5878# a_26201_5340# 0.016172f
C3348 a_13501_23906# muxtest_0.x2.x2.GN2 7.58e-21
C3349 muxtest_0.x2.x2.GN1 a_12019_24012# 0.001144f
C3350 a_23949_6654# a_24045_6654# 0.310858f
C3351 a_23529_6422# a_24329_6640# 2.3e-20
C3352 muxtest_0.x2.x2.GN2 ua[2] 0.429379f
C3353 a_24895_4790# a_25168_5156# 0.074022f
C3354 a_24729_4790# a_25761_5058# 0.048748f
C3355 a_19290_32287# ui_in[0] 0.143958f
C3356 ringtest_0.x4._08_ VDPWR 0.467036f
C3357 ringtest_0.x4.net4 a_22097_5334# 0.006897f
C3358 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR 0.636362f
C3359 ringtest_0.x4.clknet_1_1__leaf_clk a_26555_5334# 3.58e-19
C3360 muxtest_0.R2R3 ua[3] 0.017699f
C3361 ringtest_0.x4._15_ a_27233_5308# 1.61e-19
C3362 ringtest_0.x4.net6 a_22983_5654# 0.001315f
C3363 ringtest_0.x4.net3 ringtest_0.x4._02_ 0.031079f
C3364 ringtest_0.x4._22_ a_27491_4566# 3.34e-21
C3365 ringtest_0.x4.net4 ringtest_0.x4._16_ 0.442589f
C3366 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GN3 1.1e-19
C3367 ringtest_0.drv_out ringtest_0.x4.net9 4.05e-20
C3368 ui_in[0] ui_in[3] 0.001641f
C3369 ringtest_0.counter3 ringtest_0.x4._13_ 0.003357f
C3370 ringtest_0.x4._04_ a_22649_6244# 0.006456f
C3371 a_21785_5878# ringtest_0.x4.net8 9.67e-20
C3372 a_25336_4902# VDPWR 0.183641f
C3373 ringtest_0.x4.net8 a_25345_4612# 0.005557f
C3374 ringtest_0.x4._18_ a_23770_5308# 0.079699f
C3375 ringtest_0.x4._11_ a_22390_4566# 9.44e-19
C3376 a_23879_6940# a_24361_5340# 3.84e-19
C3377 a_20492_32319# ui_in[1] 8.84e-19
C3378 ringtest_0.x4.clknet_1_0__leaf_clk a_22649_6244# 6.75e-21
C3379 ringtest_0.x4._11_ ringtest_0.x4.net11 2.31e-19
C3380 muxtest_0.R5R6 VDPWR 1.61253f
C3381 muxtest_0.x1.x5.GN ua[3] 0.820663f
C3382 a_24329_6640# ringtest_0.x4._06_ 0.002324f
C3383 ringtest_0.x4._25_ ringtest_0.x4._08_ 0.208467f
C3384 a_19842_32287# ui_in[1] 0.127717f
C3385 a_25393_5308# a_25351_5712# 7.84e-20
C3386 ringtest_0.x4._11_ ringtest_0.x4._05_ 0.023537f
C3387 a_24045_6654# a_24004_6128# 0.001715f
C3388 ringtest_0.x4.net6 a_21591_6128# 4.71e-21
C3389 a_21561_9116# a_21561_8830# 0.015931f
C3390 ringtest_0.counter7 ringtest_0.x4.counter[8] 0.068429f
C3391 ringtest_0.drv_out ringtest_0.x4.net7 6.87e-19
C3392 a_22223_5712# VDPWR 0.002609f
C3393 ringtest_0.x4._15_ a_25977_4220# 0.086673f
C3394 ringtest_0.x4._19_ a_24264_6788# 1.38e-19
C3395 muxtest_0.x1.x1.nSEL1 a_19794_32347# 4.08e-19
C3396 ringtest_0.drv_out ringtest_0.x4._17_ 1.68e-19
C3397 muxtest_0.x1.x1.nSEL0 a_19242_32347# 2.51e-19
C3398 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ui_in[3] 9.57e-20
C3399 ringtest_0.x4.net2 a_21675_9686# 0.008042f
C3400 ringtest_0.x4._23_ a_26201_4790# 0.029061f
C3401 muxtest_0.x1.x5.GN a_19842_32287# 2.26e-19
C3402 a_26201_4790# a_26367_4790# 0.970499f
C3403 a_24336_6544# ringtest_0.x4._15_ 1.53e-20
C3404 ringtest_0.x4.net3 a_22116_4902# 3.22e-20
C3405 ringtest_0.x3.x2.GP3 ua[1] 0.357364f
C3406 a_21675_4790# a_22390_4566# 4.63e-19
C3407 a_23381_4818# a_23381_4584# 0.012876f
C3408 ringtest_0.x4._16_ a_23837_5878# 0.061172f
C3409 ringtest_0.x4._04_ a_21587_5334# 3.27e-21
C3410 a_16755_12091# ringtest_0.x3.x2.GP3 5.21e-19
C3411 muxtest_0.x1.x3.GN1 ui_in[2] 0.054229f
C3412 m3_17032_8096# m3_17046_7066# 0.003741f
C3413 ringtest_0.x4._06_ a_24545_5878# 0.046896f
C3414 ringtest_0.x4.net9 ringtest_0.x4._07_ 0.03749f
C3415 ringtest_0.x4._22_ ringtest_0.x4._16_ 0.135659f
C3416 muxtest_0.x2.x2.GN1 ui_in[4] 0.312374f
C3417 ringtest_0.x4._23_ a_26555_5334# 0.014354f
C3418 a_22795_5334# a_22765_4478# 6.77e-20
C3419 muxtest_0.x2.x1.nSEL0 a_12473_23980# 0.001174f
C3420 ringtest_0.x4.clknet_1_0__leaf_clk a_21587_5334# 0.03291f
C3421 a_23467_4584# VDPWR 0.002731f
C3422 a_26555_5334# a_26367_4790# 1.41e-20
C3423 ringtest_0.x4._25_ VDPWR 0.22908f
C3424 a_21803_9508# VDPWR 0.005315f
C3425 ringtest_0.x4._11_ a_22350_5878# 0.003523f
C3426 a_24004_6128# a_24699_6200# 5.89e-19
C3427 ringtest_0.x4.net1 VDPWR 1.47718f
C3428 ringtest_0.x4.clknet_1_1__leaf_clk a_23770_5308# 0.048773f
C3429 muxtest_0.x1.x3.GP3 muxtest_0.R4R5 0.346864f
C3430 ringtest_0.x4.net4 a_22649_6244# 0.002624f
C3431 ringtest_0.x4.net7 ringtest_0.x4._07_ 0.047771f
C3432 muxtest_0.x1.x3.GP1 muxtest_0.R6R7 0.271251f
C3433 ringtest_0.x4.net3 ringtest_0.x4._04_ 5.28e-22
C3434 a_21852_8720# a_22052_8875# 0.080195f
C3435 a_21785_5878# a_22390_4566# 4.07e-21
C3436 a_21561_8830# ringtest_0.x4._01_ 8.93e-19
C3437 a_21845_8816# a_21981_8976# 0.136009f
C3438 a_26201_5340# a_26735_5334# 0.002698f
C3439 ringtest_0.x4._17_ ringtest_0.x4._07_ 3.97e-20
C3440 ringtest_0.x4._23_ a_27303_4246# 0.113094f
C3441 ringtest_0.x4.net7 a_25055_3867# 0.201574f
C3442 a_25977_4220# a_26173_4612# 0.00119f
C3443 ringtest_0.x4._11_ ringtest_0.x4._09_ 0.004259f
C3444 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net3 0.373279f
C3445 ringtest_0.x4._14_ a_21948_5156# 9.43e-20
C3446 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A 0.17253f
C3447 a_26808_4902# a_26721_4246# 5.71e-20
C3448 a_11845_23906# ui_in[3] 0.048888f
C3449 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.308902f
C3450 ringtest_0.x4.net2 a_22052_8875# 3.35e-21
C3451 a_22052_9116# a_22399_9142# 0.037333f
C3452 ringtest_0.x4._06_ a_24317_4942# 2.49e-19
C3453 ringtest_0.x4.net7 a_24264_6788# 0.001683f
C3454 ringtest_0.drv_out ringtest_0.x3.x2.GN3 0.243642f
C3455 a_24004_6128# a_23809_4790# 5.65e-20
C3456 ringtest_0.x4.net1 a_21803_9508# 8.57e-19
C3457 a_24361_5340# a_24968_5308# 0.136009f
C3458 ringtest_0.x4.net8 ringtest_0.x4.net10 1.02e-19
C3459 ringtest_0.x4.net9 a_26201_5340# 8.34e-19
C3460 a_25593_5156# a_26201_4790# 3.54e-19
C3461 a_23529_6422# ringtest_0.x4._19_ 0.082191f
C3462 ringtest_0.x4._18_ ringtest_0.x4.net6 0.081404f
C3463 a_25761_5058# ringtest_0.x4._09_ 0.001669f
C3464 ringtest_0.x4._21_ VDPWR 0.492491f
C3465 ringtest_0.x4.clknet_0_clk a_24527_5340# 5.94e-19
C3466 ringtest_0.x4.counter[2] VDPWR 0.494938f
C3467 ringtest_0.counter7 ringtest_0.x4.net6 6.88e-20
C3468 a_24045_6654# ringtest_0.x4._20_ 1.76e-19
C3469 ringtest_0.x4.net4 a_21587_5334# 1.97e-19
C3470 a_23809_4790# a_23963_4790# 0.004009f
C3471 ringtest_0.x4._15_ a_23899_5334# 0.046541f
C3472 a_16027_11759# ui_in[4] 0.03417f
C3473 muxtest_0.x1.x4.A a_12977_24040# 3.86e-20
C3474 ringtest_0.x4._24_ a_26367_5340# 0.035946f
C3475 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR 0.636314f
C3476 ringtest_0.x3.x1.nSEL1 a_16203_12091# 0.041068f
C3477 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN2 1.03e-20
C3478 a_21675_4790# a_22074_4790# 0.001351f
C3479 a_22116_4902# a_22457_5156# 9.73e-19
C3480 a_23381_4818# a_23809_4790# 0.00155f
C3481 a_21948_5156# a_22043_5156# 0.007724f
C3482 ringtest_0.counter3 ringtest_0.x4.counter[1] 0.099026f
C3483 ringtest_0.x4.net7 a_26201_5340# 8.61e-20
C3484 a_22265_5308# a_22164_4362# 6.81e-19
C3485 a_21425_9686# VDPWR 0.260172f
C3486 ringtest_0.x4._16_ a_22021_4220# 0.184103f
C3487 a_21951_5878# a_22392_5990# 0.111047f
C3488 a_23349_6422# VDPWR 0.252612f
C3489 a_12849_23648# VDPWR 0.180589f
C3490 a_21845_8816# a_22228_8598# 0.001632f
C3491 a_21852_8720# a_21803_8598# 4.04e-19
C3492 a_22052_8875# a_22399_8976# 0.037333f
C3493 a_21981_8976# a_22201_8964# 4.62e-19
C3494 ringtest_0.x4._23_ ringtest_0.x4.counter[8] 9.18e-19
C3495 a_23879_6940# VDPWR 1.29479f
C3496 ringtest_0.x4.net6 a_24763_6143# 0.027058f
C3497 ringtest_0.x4.net9 a_27233_5058# 0.001937f
C3498 ringtest_0.x3.x2.GP3 m3_17046_7066# 0.006132f
C3499 ringtest_0.x4._19_ ringtest_0.x4._06_ 7.42e-21
C3500 ringtest_0.x4.net7 ringtest_0.x4.counter[5] 0.002945f
C3501 ringtest_0.x4.net3 ringtest_0.x4.net4 0.0313f
C3502 muxtest_0.x2.x2.GN2 m3_13302_19985# 0.016745f
C3503 muxtest_0.x2.x2.GN4 ui_in[3] 0.218988f
C3504 a_25309_5334# VDPWR 0.004428f
C3505 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP1 0.062377f
C3506 ringtest_0.x4.counter[1] ua[2] 1.11e-19
C3507 a_20318_32213# muxtest_0.x1.x3.GN4 0.134079f
C3508 muxtest_0.x1.x3.GN2 a_19242_32347# 0.002395f
C3509 ringtest_0.x4._00_ a_22052_9116# 0.00938f
C3510 ringtest_0.x4._24_ a_27065_5156# 0.012283f
C3511 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ui_in[3] 9.57e-20
C3512 ringtest_0.x4.net7 a_27233_5058# 8.32e-20
C3513 ringtest_0.x4.net1 a_21425_9686# 0.224922f
C3514 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2 2.14737f
C3515 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net6 0.323735f
C3516 ringtest_0.ring_out ringtest_0.x3.x1.nSEL0 1.86e-21
C3517 muxtest_0.x1.x3.GP3 ui_in[2] 1.6e-19
C3518 a_23529_6422# ringtest_0.x4.net7 0.002934f
C3519 ringtest_0.x4.clknet_1_1__leaf_clk a_24895_4790# 0.486375f
C3520 ringtest_0.x4.net8 a_25393_5308# 0.084103f
C3521 ringtest_0.x4._17_ a_23529_6422# 0.043588f
C3522 ringtest_0.x4._11_ a_24361_5340# 1.58e-19
C3523 a_21375_3867# VDPWR 0.272145f
C3524 ringtest_0.x4.net10 ringtest_0.x4.net11 0.310558f
C3525 a_16027_11759# ringtest_0.x3.x2.GP1 9.92e-19
C3526 a_16203_12091# ringtest_0.x3.x2.GN3 0.048646f
C3527 ringtest_0.x4._08_ a_24968_5308# 9.82e-20
C3528 ringtest_0.x4._06_ ringtest_0.x4.net9 0.017291f
C3529 a_16579_11759# ringtest_0.x3.x2.GN1 6.43e-20
C3530 a_23809_4790# ringtest_0.x4._20_ 0.237238f
C3531 ua[3] ui_in[4] 1.14709f
C3532 ringtest_0.x4._11_ a_21395_6940# 0.055744f
C3533 a_21509_4790# a_21948_5156# 0.273138f
C3534 ringtest_0.x4._15_ a_22097_5334# 7.5e-20
C3535 ringtest_0.x4.net6 a_24800_5334# 0.019975f
C3536 ringtest_0.x4._03_ a_22116_4902# 0.006259f
C3537 ringtest_0.x4._22_ a_27273_4220# 4.31e-19
C3538 ringtest_0.x4._12_ a_22245_8054# 0.026119f
C3539 muxtest_0.x1.x5.A muxtest_0.R7R8 4.52065f
C3540 a_24527_5340# a_25168_5156# 7.62e-19
C3541 a_24800_5334# a_24895_4790# 8.92e-19
C3542 ringtest_0.x4._15_ ringtest_0.x4._16_ 0.656968f
C3543 a_25393_5308# a_24729_4790# 0.002274f
C3544 a_25977_4220# a_25975_3867# 0.01226f
C3545 ringtest_0.x4.net7 ringtest_0.x4._06_ 0.141876f
C3546 ringtest_0.x4.net7 a_24070_5852# 0.003377f
C3547 ringtest_0.x4.clknet_0_clk a_25168_5156# 4.63e-19
C3548 ringtest_0.x4._18_ a_23932_6128# 0.00112f
C3549 ringtest_0.x4._17_ ringtest_0.x4._06_ 0.001225f
C3550 muxtest_0.x1.x1.nSEL1 ui_in[1] 0.275603f
C3551 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A 5.04e-19
C3552 a_23879_6940# ringtest_0.x4._21_ 0.001038f
C3553 ringtest_0.x4._16_ a_22541_5058# 1.37e-19
C3554 a_26808_5308# a_26640_5334# 0.239923f
C3555 a_26201_5340# a_27065_5334# 0.032244f
C3556 a_23770_5308# a_23993_5654# 0.011458f
C3557 a_26367_5340# a_27233_5308# 0.034054f
C3558 ringtest_0.x4._17_ a_24070_5852# 0.062168f
C3559 a_24968_5308# VDPWR 0.185172f
C3560 ringtest_0.x4.net6 ringtest_0.x4._23_ 0.023006f
C3561 a_24329_6640# a_24883_6800# 0.057611f
C3562 a_24045_6654# a_24287_6422# 0.008508f
C3563 ringtest_0.x4.net4 a_22457_5156# 8.77e-19
C3564 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x5.GN 0.10521f
C3565 muxtest_0.x2.x2.GP1 ua[2] 0.352897f
C3566 a_24895_4790# a_26367_4790# 0.002814f
C3567 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._03_ 0.00668f
C3568 a_18662_32213# m2_18699_31802# 0.01297f
C3569 muxtest_0.x2.x1.nSEL1 a_12977_24040# 4.08e-19
C3570 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN2 0.209956f
C3571 a_11845_23906# muxtest_0.x2.x2.GN1 0.12869f
C3572 ringtest_0.x4.net10 ringtest_0.x4._09_ 0.081678f
C3573 ringtest_0.counter7 ringtest_0.x4.net5 6.88e-20
C3574 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR 0.636314f
C3575 a_27233_5308# a_27065_5156# 7.04e-19
C3576 a_22817_6146# ringtest_0.x4._06_ 1.81e-20
C3577 a_25925_6788# VDPWR 0.455589f
C3578 a_27065_5334# a_27233_5058# 7.04e-19
C3579 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x1.nSEL1 0.352716f
C3580 a_21395_6940# a_21785_5878# 5.49e-20
C3581 a_21375_3867# ringtest_0.x4.counter[2] 4.98e-19
C3582 a_22817_6146# a_24070_5852# 2.22e-20
C3583 muxtest_0.x1.x5.A muxtest_0.R5R6 4.5214f
C3584 uio_in[7] uio_in[6] 0.031023f
C3585 ringtest_0.x4.net6 ringtest_0.x4._02_ 0.001309f
C3586 ringtest_0.x4._11_ ringtest_0.x4._08_ 1.44e-20
C3587 ringtest_0.x4.clknet_1_0__leaf_clk a_21939_8054# 3.8e-19
C3588 a_15749_12123# VDPWR 9.25e-19
C3589 ringtest_0.x4._22_ a_26201_4790# 4.68e-20
C3590 muxtest_0.x2.x2.GN2 ua[0] 4.0283f
C3591 muxtest_0.x1.x5.A VDPWR 14.1646f
C3592 a_19794_32347# muxtest_0.x1.x3.GP3 4.39e-19
C3593 ringtest_0.x3.x2.GN3 m3_17036_9140# 0.001446f
C3594 ringtest_0.x4.net3 a_22021_4220# 0.002183f
C3595 ringtest_0.x4._15_ a_26201_6788# 0.001194f
C3596 ringtest_0.x4.net7 a_26269_4612# 5.42e-19
C3597 a_25925_6788# ringtest_0.x4._25_ 1.87e-19
C3598 ringtest_0.x4._11_ a_25336_4902# 0.039242f
C3599 ringtest_0.x4._23_ a_27169_6641# 6.47e-19
C3600 ringtest_0.x4.net11 a_27191_4790# 3e-19
C3601 ringtest_0.x4._07_ a_25351_5712# 5.27e-19
C3602 a_21675_9686# a_21465_9294# 3.08e-19
C3603 a_19290_32287# muxtest_0.x1.x3.GN3 0.048646f
C3604 ringtest_0.x4._02_ a_21055_5334# 0.01416f
C3605 ringtest_0.counter7 a_21007_3867# 2.81e-20
C3606 a_26749_6422# a_26808_4902# 1.02e-20
C3607 a_19114_31955# VDPWR 0.164569f
C3608 a_26640_5156# a_26766_4790# 0.005525f
C3609 a_26555_4790# a_26735_5156# 0.001229f
C3610 a_21233_5340# VDPWR 0.684183f
C3611 a_21399_5340# a_22265_5308# 0.034054f
C3612 a_21840_5308# a_21672_5334# 0.239923f
C3613 ringtest_0.x4.net4 ringtest_0.x4._03_ 0.031989f
C3614 ringtest_0.x4.net10 a_27659_4246# 0.003077f
C3615 ringtest_0.ring_out ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.167117f
C3616 muxtest_0.x2.x2.GN3 a_12977_24040# 0.001073f
C3617 muxtest_0.x2.x2.GN2 a_13675_24012# 8.14e-21
C3618 m2_11882_23495# VDPWR 0.139985f
C3619 ringtest_0.x4.net8 a_24715_5334# 0.005878f
C3620 ringtest_0.x4._11_ a_22223_5712# 6.78e-19
C3621 ringtest_0.x4.net6 a_25593_5156# 4.38e-19
C3622 ringtest_0.x4._15_ a_23467_4818# 7.85e-19
C3623 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GN3 0.067465f
C3624 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN4 0.001074f
C3625 a_25364_5878# a_26808_5308# 0.006157f
C3626 a_24045_6654# a_24329_6640# 0.030894f
C3627 a_23949_6654# a_24336_6544# 0.034054f
C3628 a_20492_32319# ui_in[0] 1.77e-19
C3629 ringtest_0.x4._11_ VDPWR 5.18499f
C3630 a_25336_4902# a_25761_5058# 1.28e-19
C3631 a_24729_4790# a_25083_4790# 0.062224f
C3632 a_24895_4790# a_25593_5156# 0.193199f
C3633 a_19842_32287# ui_in[0] 0.279876f
C3634 ringtest_0.x4.net4 a_23770_5308# 1.34e-19
C3635 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN3 4.01e-20
C3636 ringtest_0.x4.clknet_1_1__leaf_clk a_24895_5334# 0.002214f
C3637 ringtest_0.x4._22_ a_27303_4246# 6.52e-20
C3638 a_25975_3867# ringtest_0.x4.counter[9] 2.37e-20
C3639 muxtest_0.R6R7 muxtest_0.R4R5 2.49e-19
C3640 ringtest_0.x4._14_ a_22164_4362# 0.089653f
C3641 a_25761_5058# VDPWR 0.400861f
C3642 ringtest_0.x4.net8 a_25547_4612# 1.72e-20
C3643 a_23879_6940# a_24968_5308# 8.05e-21
C3644 ringtest_0.x4._11_ a_23467_4584# 6.46e-19
C3645 ringtest_0.x4._11_ ringtest_0.x4._25_ 2.54e-20
C3646 muxtest_0.x1.x3.GN1 muxtest_0.R2R3 2.55e-19
C3647 a_25364_5878# a_26555_4790# 1.26e-19
C3648 a_21675_4790# VDPWR 0.342267f
C3649 ringtest_0.x4.net3 a_21561_8830# 0.006429f
C3650 a_24536_6699# ringtest_0.x4._06_ 2.41e-19
C3651 muxtest_0.x1.x3.GN1 ui_in[1] 0.312176f
C3652 ringtest_0.x4.net1 ringtest_0.x4._11_ 0.002334f
C3653 ringtest_0.x4.clknet_0_clk ringtest_0.x4._18_ 0.002702f
C3654 a_24968_5308# a_25309_5334# 9.73e-19
C3655 a_24800_5334# a_24895_5334# 0.007724f
C3656 a_21561_9116# a_21852_8720# 1.53e-19
C3657 a_21845_9116# a_21561_8830# 9.64e-20
C3658 a_24336_6544# a_24004_6128# 0.002652f
C3659 a_24329_6640# a_24699_6200# 0.007926f
C3660 ringtest_0.x4.net6 ringtest_0.x4._04_ 0.050232f
C3661 a_21852_9416# a_21845_8816# 3.36e-19
C3662 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A 0.17253f
C3663 a_23899_5654# VDPWR 5.6e-19
C3664 a_26569_6422# ringtest_0.x4._24_ 0.095435f
C3665 ringtest_0.x4.net2 a_21780_9142# 2.28e-19
C3666 ringtest_0.x4._19_ a_24883_6800# 0.014678f
C3667 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net6 6.56e-20
C3668 ringtest_0.x3.nselect2 ui_in[3] 1.88e-19
C3669 ringtest_0.ring_out ua[1] 4.51997f
C3670 ringtest_0.x4.net2 a_21561_9116# 0.019416f
C3671 ringtest_0.x4._09_ a_27191_4790# 0.001794f
C3672 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN1 0.645006f
C3673 muxtest_0.x1.x1.nSEL0 VDPWR 0.389106f
C3674 ringtest_0.ring_out a_16755_12091# 2.55e-19
C3675 a_24465_6800# ringtest_0.x4._15_ 2.35e-21
C3676 ringtest_0.x4._09_ a_26808_4902# 0.039926f
C3677 a_26201_4790# a_26640_5156# 0.273138f
C3678 a_24763_6143# a_24527_5340# 0.003413f
C3679 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP3 0.002437f
C3680 a_21785_5878# VDPWR 0.6434f
C3681 a_24045_6654# a_24317_4942# 5.98e-21
C3682 a_21951_5878# a_22265_5308# 0.003783f
C3683 muxtest_0.x2.x1.nSEL0 a_13025_23980# 1.21e-20
C3684 a_24699_6200# a_24545_5878# 0.049785f
C3685 ringtest_0.x4.clknet_0_clk a_24763_6143# 7.62e-19
C3686 ringtest_0.x4.clknet_1_0__leaf_clk a_21055_5334# 1.21e-20
C3687 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP1 1.16e-20
C3688 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR 0.63819f
C3689 a_22399_9142# VDPWR 0.080219f
C3690 ringtest_0.x4.net9 a_26895_3867# 0.202772f
C3691 ringtest_0.x4._11_ ringtest_0.x4._21_ 0.059807f
C3692 muxtest_0.R7R8 ua[2] 4.51509f
C3693 a_23949_6654# a_23899_5334# 2.76e-21
C3694 ringtest_0.x4.clknet_1_1__leaf_clk a_24527_5340# 0.079788f
C3695 muxtest_0.x1.x3.GN4 muxtest_0.R4R5 4.23588f
C3696 muxtest_0.x2.x2.GP1 m3_13302_19985# 3.25e-21
C3697 a_21852_8720# ringtest_0.x4._01_ 0.239739f
C3698 ringtest_0.x4.net3 a_21049_8598# 0.042192f
C3699 a_22052_8875# a_21981_8976# 0.239923f
C3700 a_26367_5340# a_27149_5334# 6.32e-19
C3701 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_1_1__leaf_clk 0.335671f
C3702 muxtest_0.x1.x3.GN2 muxtest_0.R7R8 0.260757f
C3703 a_25977_4220# a_26375_4612# 0.005781f
C3704 ringtest_0.x4._14_ a_22373_5156# 0.002114f
C3705 ringtest_0.x4.net6 ringtest_0.x4.net4 0.008308f
C3706 a_21981_9142# ringtest_0.x4.clknet_1_0__leaf_clk 0.050329f
C3707 a_12473_23980# ui_in[3] 0.143958f
C3708 ringtest_0.x4.net2 ringtest_0.x4._01_ 9.85e-20
C3709 ringtest_0.x4._11_ a_23349_6422# 0.001422f
C3710 ringtest_0.x4.net7 a_24883_6800# 0.019182f
C3711 ringtest_0.x4._11_ a_23879_6940# 4.59e-19
C3712 ringtest_0.x4._17_ a_21951_5878# 9.29e-21
C3713 a_24361_5340# a_25393_5308# 0.048748f
C3714 a_24527_5340# a_24800_5334# 0.074815f
C3715 ringtest_0.x4.net1 a_22399_9142# 5.53e-20
C3716 a_18662_32213# a_18836_32319# 0.006584f
C3717 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP2 0.043402f
C3718 ringtest_0.x4._17_ a_24883_6800# 0.016586f
C3719 ringtest_0.x4._15_ a_26201_4790# 0.02569f
C3720 ringtest_0.x4._21_ a_23899_5654# 2.03e-19
C3721 ringtest_0.x4.net9 a_26808_5308# 2.66e-21
C3722 ringtest_0.ring_out ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C3723 a_24045_6654# ringtest_0.x4._19_ 0.046625f
C3724 ringtest_0.x4._08_ ringtest_0.x4.net10 0.001321f
C3725 a_24329_6640# a_25421_6641# 5.23e-20
C3726 ringtest_0.x4.clknet_0_clk a_24800_5334# 4.59e-20
C3727 ringtest_0.counter3 VDPWR 2.51653f
C3728 ringtest_0.x4._03_ a_22021_4220# 0.112166f
C3729 a_21509_4790# a_22164_4362# 0.00127f
C3730 a_24317_4942# a_24479_4790# 0.004009f
C3731 muxtest_0.x2.x2.GN4 ua[3] 0.085877f
C3732 ringtest_0.x4._15_ a_26555_5334# 0.007874f
C3733 ringtest_0.x4.net8 ringtest_0.x4._07_ 0.001136f
C3734 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x3.x2.GN3 7.01e-21
C3735 ringtest_0.x4._24_ a_26640_5334# 0.010979f
C3736 a_16579_11759# ui_in[4] 0.261734f
C3737 ringtest_0.x3.x1.nSEL1 a_16755_12091# 1.59e-19
C3738 a_23809_4790# a_24317_4942# 0.017774f
C3739 a_22116_4902# ringtest_0.x4.net5 0.001073f
C3740 a_21948_5156# a_22074_4790# 0.005525f
C3741 ringtest_0.x4._00_ VDPWR 0.655201f
C3742 a_27489_3702# a_27815_3867# 0.024477f
C3743 ringtest_0.x4.net8 a_25055_3867# 3.76e-19
C3744 muxtest_0.x1.x3.GP3 muxtest_0.R2R3 0.115101f
C3745 a_22392_5990# a_22224_6244# 0.239923f
C3746 a_21951_5878# a_22817_6146# 0.034054f
C3747 ringtest_0.x4._16_ a_22765_4478# 0.01632f
C3748 a_13501_23906# VDPWR 0.218058f
C3749 VDPWR ua[2] 13.246901f
C3750 a_21852_8720# a_21785_8054# 1.58e-19
C3751 a_21981_8976# a_21803_8598# 9.73e-19
C3752 a_22052_8875# a_22228_8598# 0.007724f
C3753 muxtest_0.x1.x3.GP3 ui_in[1] 0.003199f
C3754 ringtest_0.x4.net6 a_23837_5878# 4.02e-19
C3755 a_21845_8816# ringtest_0.x4._10_ 0.011255f
C3756 ringtest_0.x4._01_ a_22399_8976# 0.121379f
C3757 ringtest_0.x4.clknet_0_clk ringtest_0.x4._23_ 2.29e-20
C3758 ringtest_0.x4.net6 ringtest_0.x4._22_ 0.641715f
C3759 ringtest_0.x4.net9 a_26555_4790# 0.016338f
C3760 muxtest_0.x2.x2.GN4 m3_13316_18955# 0.084813f
C3761 muxtest_0.x1.x3.GN2 muxtest_0.R5R6 0.122627f
C3762 ringtest_0.x4._07_ a_24729_4790# 0.112051f
C3763 a_23949_6654# ringtest_0.x4._16_ 3.45e-20
C3764 ringtest_0.x4._19_ a_24699_6200# 1.87e-20
C3765 ringtest_0.x4._22_ a_24895_4790# 0.02378f
C3766 ringtest_0.x4.net10 VDPWR 1.28398f
C3767 ringtest_0.x4.net6 a_24135_3867# 0.195979f
C3768 ringtest_0.x4.net2 a_21785_8054# 0.165774f
C3769 ringtest_0.x4.counter[0] ua[1] 3.21e-19
C3770 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A 5.04e-19
C3771 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP3 3.82e-20
C3772 ringtest_0.drv_out ringtest_0.x4._05_ 0.0016f
C3773 a_24729_4790# a_25055_3867# 1.63e-21
C3774 ringtest_0.x4._24_ a_26735_5156# 7.21e-19
C3775 muxtest_0.x1.x3.GN2 VDPWR 0.701394f
C3776 ringtest_0.x4._00_ a_21803_9508# 3.7e-19
C3777 ringtest_0.x4.net7 a_23381_4584# 2.04e-20
C3778 ringtest_0.x4._04_ ringtest_0.x4.net5 0.003846f
C3779 ringtest_0.x4.net7 a_26555_4790# 2.26e-19
C3780 ua[1] ua[4] 0.001128f
C3781 ringtest_0.x4.net1 ringtest_0.x4._00_ 0.056053f
C3782 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net5 6.12e-20
C3783 ringtest_0.x4._14_ a_21399_5340# 4.89e-20
C3784 a_24045_6654# ringtest_0.x4.net7 0.037726f
C3785 a_24627_6200# VDPWR 0.001301f
C3786 muxtest_0.x1.x3.GN4 ui_in[2] 5.71e-20
C3787 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GP1 1.21e-19
C3788 ringtest_0.x4.clknet_1_1__leaf_clk a_25168_5156# 0.042872f
C3789 ringtest_0.x4._06_ a_22765_5308# 1.6e-20
C3790 ringtest_0.x4.counter[4] VDPWR 0.454642f
C3791 ringtest_0.x4.net8 a_26201_5340# 0.001229f
C3792 muxtest_0.R2R3 muxtest_0.R1R2 1.9897f
C3793 ringtest_0.x3.x2.GN3 ua[1] 0.429944f
C3794 ringtest_0.x4._11_ a_24968_5308# 7.26e-20
C3795 ringtest_0.x4._17_ a_24045_6654# 0.036473f
C3796 a_23399_3867# VDPWR 0.316408f
C3797 a_16579_11759# ringtest_0.x3.x2.GP1 1.21e-20
C3798 ui_in[3] ui_in[5] 0.13854f
C3799 ringtest_0.x4._08_ a_25393_5308# 9.54e-19
C3800 muxtest_0.x2.x1.nSEL1 a_12297_23648# 0.073392f
C3801 a_16755_12091# ringtest_0.x3.x2.GN3 0.004288f
C3802 muxtest_0.x1.x1.nSEL1 ui_in[0] 0.169954f
C3803 a_24004_6128# ringtest_0.x4._16_ 0.029136f
C3804 ringtest_0.x4.net9 ringtest_0.x4.counter[6] 3.69e-19
C3805 a_24699_6200# ringtest_0.x4.net9 0.170073f
C3806 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR 0.92605f
C3807 ringtest_0.counter3 ringtest_0.x4.counter[2] 0.16993f
C3808 a_21509_4790# a_22373_5156# 0.032244f
C3809 a_23899_5334# ringtest_0.x4._20_ 1.05e-19
C3810 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x3.x1.nSEL1 1.23e-19
C3811 ringtest_0.x4.net6 a_25225_5334# 8.63e-19
C3812 ringtest_0.x4._03_ a_22541_5058# 3.08e-19
C3813 ringtest_0.x4._15_ a_23770_5308# 0.229149f
C3814 a_25225_5334# a_24895_4790# 1.5e-19
C3815 a_25393_5308# a_25336_4902# 6.84e-19
C3816 ringtest_0.x4.net2 ringtest_0.x4._16_ 5.41e-20
C3817 muxtest_0.x2.x2.GP1 ua[0] 0.128232f
C3818 ringtest_0.x4._24_ a_25364_5878# 0.025563f
C3819 a_26627_4246# a_26895_3867# 1.23e-19
C3820 a_15575_12017# VDPWR 0.211635f
C3821 ringtest_0.x4.net7 ringtest_0.x4.counter[6] 1.8e-19
C3822 ringtest_0.x4._16_ a_23963_4790# 5.12e-19
C3823 a_22649_6244# a_22765_4478# 3.06e-22
C3824 ringtest_0.x4._11_ a_25925_6788# 0.087773f
C3825 a_21840_5308# a_21863_4790# 6.87e-19
C3826 ringtest_0.x4.net9 a_24479_4790# 8.5e-21
C3827 ringtest_0.x4.net7 a_24699_6200# 6.37e-20
C3828 a_22765_5308# a_22373_5156# 0.006202f
C3829 a_19666_31955# muxtest_0.R7R8 7.47e-21
C3830 ringtest_0.x4._16_ a_23381_4818# 0.113241f
C3831 ringtest_0.x4.counter[2] ua[2] 1.11e-19
C3832 a_26808_5308# a_27065_5334# 0.036838f
C3833 a_22265_5308# a_22795_5334# 2.84e-19
C3834 a_24361_5340# a_24715_5334# 0.057611f
C3835 a_22097_5334# a_22181_5334# 0.008508f
C3836 ringtest_0.x4._17_ a_24699_6200# 7.49e-19
C3837 muxtest_0.x2.x1.nSEL0 ui_in[3] 0.32698f
C3838 muxtest_0.R7R8 m3_13302_19985# 0.001045f
C3839 a_25393_5308# VDPWR 0.406789f
C3840 a_24336_6544# a_24287_6422# 4.04e-19
C3841 a_24536_6699# a_24883_6800# 0.037333f
C3842 a_24465_6800# a_24685_6788# 4.62e-19
C3843 a_21425_9686# ringtest_0.x4._00_ 0.167554f
C3844 ringtest_0.x4.net4 ringtest_0.x4.net5 0.483177f
C3845 ringtest_0.x4.net7 a_24479_4790# 1.98e-19
C3846 a_25421_6641# ringtest_0.x4._19_ 0.214472f
C3847 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP1 0.001426f
C3848 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.001676f
C3849 a_12297_23648# muxtest_0.x2.x2.GN3 6.68e-19
C3850 ringtest_0.x4.net7 a_23809_4790# 0.003261f
C3851 a_12473_23980# muxtest_0.x2.x2.GN1 1.46e-19
C3852 muxtest_0.R7R8 muxtest_0.x2.x2.GP2 1.13e-20
C3853 a_23932_6128# a_23837_5878# 0.002032f
C3854 ringtest_0.x4._11_ a_21233_5340# 0.00462f
C3855 ringtest_0.x4._17_ a_23809_4790# 1e-20
C3856 a_21951_5878# ringtest_0.x4._14_ 3.24e-22
C3857 a_26749_6422# a_26201_5340# 6.06e-21
C3858 ringtest_0.x4.net8 ringtest_0.x4._06_ 0.209874f
C3859 a_27191_4790# VDPWR 4.71e-19
C3860 ringtest_0.x4.net8 a_24070_5852# 0.028641f
C3861 a_22392_5990# a_22139_5878# 3.39e-19
C3862 a_26808_4902# VDPWR 0.186041f
C3863 ringtest_0.counter3 a_21375_3867# 4.27e-20
C3864 ringtest_0.x3.x2.GN4 VDPWR 1.23317f
C3865 muxtest_0.x1.x4.A muxtest_0.R5R6 1.64e-20
C3866 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_0_clk 0.004956f
C3867 muxtest_0.x1.x3.GN3 ua[3] 0.014498f
C3868 muxtest_0.x1.x5.GN muxtest_0.x2.nselect2 4.76e-21
C3869 a_25421_6641# ringtest_0.x4.net9 3.61e-20
C3870 ringtest_0.x3.x2.GP1 m3_17032_8096# 3.25e-21
C3871 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._12_ 0.075464f
C3872 ringtest_0.x3.x2.GN3 m3_17046_7066# 0.016026f
C3873 ringtest_0.x4._24_ a_26913_4566# 0.002926f
C3874 ringtest_0.x4._16_ ringtest_0.x4._20_ 0.011071f
C3875 muxtest_0.x1.x4.A VDPWR 15.014299f
C3876 a_21233_5340# a_21675_4790# 2.24e-19
C3877 ringtest_0.x4._22_ ringtest_0.x4.net5 4.26e-20
C3878 a_21399_5340# a_21509_4790# 0.010101f
C3879 a_19794_32347# muxtest_0.x1.x3.GN4 3.22e-19
C3880 ringtest_0.x4.net8 a_23891_4790# 4.38e-20
C3881 muxtest_0.x1.x3.GN3 a_20492_32319# 1.07e-20
C3882 a_22164_4362# a_22390_4566# 0.005961f
C3883 ringtest_0.x4._11_ a_25761_5058# 0.028602f
C3884 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A 0.17253f
C3885 a_21465_9294# a_21780_9142# 7.84e-20
C3886 a_27065_5156# a_27273_4220# 0.003595f
C3887 a_19842_32287# muxtest_0.x1.x3.GN3 0.004289f
C3888 a_21675_9686# a_21852_9416# 0.001655f
C3889 a_21465_9294# a_21561_9116# 0.310858f
C3890 ringtest_0.x4.net5 a_24135_3867# 0.001724f
C3891 ringtest_0.counter7 a_22295_3867# 2.81e-20
C3892 a_27233_5058# ringtest_0.x4.net11 0.092457f
C3893 ringtest_0.x4._19_ ringtest_0.x4._24_ 8.27e-21
C3894 a_19666_31955# VDPWR 0.171399f
C3895 ringtest_0.x4._11_ a_21675_4790# 0.03376f
C3896 ringtest_0.x4.net6 ringtest_0.x4._15_ 0.117386f
C3897 a_21840_5308# a_22097_5334# 0.036838f
C3898 a_25421_6641# ringtest_0.x4.net7 0.030401f
C3899 muxtest_0.x1.x1.nSEL0 a_19114_31955# 0.03096f
C3900 ringtest_0.x4._15_ a_24895_4790# 2.57e-20
C3901 ringtest_0.x4._16_ a_21840_5308# 1.76e-20
C3902 ringtest_0.x4._17_ a_25421_6641# 0.019971f
C3903 a_23529_6422# ringtest_0.x4._05_ 4.91e-20
C3904 a_23949_6654# a_24465_6800# 1.28e-19
C3905 ringtest_0.x4._18_ ringtest_0.x4.clknet_1_1__leaf_clk 3.06e-19
C3906 a_24329_6640# a_24336_6544# 0.961627f
C3907 ringtest_0.x4._24_ a_26735_5334# 7.21e-19
C3908 a_25336_4902# a_25083_4790# 3.39e-19
C3909 ringtest_0.x3.x2.GP2 ringtest_0.counter7 1.13e-20
C3910 ringtest_0.x3.x2.GP3 ui_in[4] 0.003259f
C3911 muxtest_0.x1.x3.GN1 ui_in[0] 0.023343f
C3912 a_21465_8830# VDPWR 0.399249f
C3913 a_23381_4818# a_23467_4818# 0.006584f
C3914 a_21785_5878# a_21233_5340# 0.002682f
C3915 ringtest_0.x4._13_ a_21399_5340# 1.58e-19
C3916 ringtest_0.x4.net6 a_24926_5712# 0.001426f
C3917 a_27489_3702# ringtest_0.x4.counter[9] 0.109832f
C3918 muxtest_0.x2.x2.GP2 VDPWR 1.81003f
C3919 a_26201_5340# ringtest_0.x4._09_ 1.11e-19
C3920 a_26367_5340# a_26201_4790# 2.64e-19
C3921 ringtest_0.x4._14_ a_23381_4584# 9.06e-21
C3922 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x1.nSEL1 2.53e-21
C3923 ringtest_0.x4._11_ a_21785_5878# 0.205946f
C3924 a_26721_4246# a_26895_3867# 2.21e-19
C3925 a_25083_4790# VDPWR 0.079731f
C3926 ringtest_0.x4._24_ ringtest_0.x4.net9 0.165357f
C3927 muxtest_0.x1.x3.GP2 ua[3] 0.023177f
C3928 a_25364_5878# a_25977_4220# 4.57e-20
C3929 a_22399_9142# ringtest_0.x4._11_ 2.48e-19
C3930 ringtest_0.x4.clknet_1_0__leaf_clk a_22245_8054# 0.00537f
C3931 a_21948_5156# VDPWR 0.286549f
C3932 ringtest_0.x4.net3 a_21852_8720# 0.005586f
C3933 a_26367_5340# a_26555_5334# 0.097994f
C3934 a_21852_9416# a_22052_8875# 1.26e-19
C3935 a_21845_9116# a_21852_8720# 3.36e-19
C3936 a_22052_9116# a_21845_8816# 6.88e-20
C3937 a_24715_5334# VDPWR 0.084103f
C3938 ringtest_0.x4._15_ a_22939_4584# 1.81e-19
C3939 a_19842_32287# muxtest_0.x1.x3.GP2 2.95e-20
C3940 ringtest_0.x4.net1 a_21465_8830# 0.081622f
C3941 ringtest_0.x4.net2 ringtest_0.x4.net3 1.28152f
C3942 ringtest_0.x4._15_ a_27169_6641# 8.98e-20
C3943 muxtest_0.R7R8 ua[0] 2.33155f
C3944 ringtest_0.x4.net7 ringtest_0.x4._24_ 2.68e-19
C3945 ringtest_0.x4.net2 a_21845_9116# 4.59e-19
C3946 ringtest_0.ring_out ringtest_0.x3.x2.GN1 4.6809f
C3947 a_21951_5878# a_21509_4790# 1.21e-19
C3948 a_21785_5878# a_21675_4790# 3.23e-21
C3949 ringtest_0.x4._09_ a_27233_5058# 0.010518f
C3950 a_26201_4790# a_27065_5156# 0.032244f
C3951 ringtest_0.x4._07_ a_24361_5340# 0.022853f
C3952 ringtest_0.x4._17_ ringtest_0.x4._24_ 0.004444f
C3953 ringtest_0.counter7 ringtest_0.x4._23_ 0.004833f
C3954 a_24763_6143# a_24800_5334# 1.41e-19
C3955 ringtest_0.x4.net5 a_22021_4220# 0.006016f
C3956 ringtest_0.x4._22_ a_24527_5340# 0.015364f
C3957 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.025028f
C3958 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP3 0.001226f
C3959 ringtest_0.counter7 a_26367_4790# 5.88e-20
C3960 muxtest_0.R1R2 ui_in[4] 8.73e-20
C3961 ringtest_0.x4._04_ a_22983_5654# 0.002919f
C3962 muxtest_0.x2.x1.nSEL0 a_12425_24040# 2.51e-19
C3963 a_24361_5340# a_25055_3867# 1.7e-21
C3964 a_21780_8964# VDPWR 3.44e-19
C3965 a_22224_6244# a_22265_5308# 0.004197f
C3966 a_22392_5990# a_22097_5334# 0.004484f
C3967 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN1 0.004375f
C3968 a_24336_6544# a_24317_4942# 2.42e-19
C3969 ringtest_0.x4.clknet_1_0__leaf_clk a_22983_5654# 1.8e-20
C3970 ringtest_0.x4.clknet_0_clk ringtest_0.x4._22_ 0.003156f
C3971 ua[4] VSS 0.139799f
C3972 ua[5] VSS 0.141076f
C3973 ua[6] VSS 0.141964f
C3974 ua[7] VSS 0.146962f
C3975 ena VSS 0.072324f
C3976 clk VSS 0.044814f
C3977 rst_n VSS 0.044814f
C3978 ui_in[7] VSS 0.044814f
C3979 uio_in[0] VSS 0.047326f
C3980 uio_in[1] VSS 0.048926f
C3981 uio_in[2] VSS 0.044814f
C3982 uio_in[3] VSS 0.044814f
C3983 uio_in[4] VSS 0.044814f
C3984 uio_in[5] VSS 0.044814f
C3985 uio_in[6] VSS 0.044814f
C3986 uio_in[7] VSS 0.075838f
C3987 ua[1] VSS 28.486887f
C3988 ui_in[5] VSS 17.64489f
C3989 ui_in[6] VSS 24.291725f
C3990 ua[2] VSS 34.46381f
C3991 ua[0] VSS 51.530293f
C3992 ui_in[4] VSS 31.64427f
C3993 ui_in[3] VSS 32.74676f
C3994 ua[3] VSS 54.146942f
C3995 ui_in[2] VSS 26.529623f
C3996 ui_in[1] VSS 10.570298f
C3997 ui_in[0] VSS 10.700917f
C3998 VDPWR VSS 0.699931p
C3999 m3_17046_7066# VSS 0.075151f $ **FLOATING
C4000 m3_17032_8096# VSS 0.073094f $ **FLOATING
C4001 m3_17036_9140# VSS 0.148749f $ **FLOATING
C4002 m3_13316_18955# VSS 0.066786f $ **FLOATING
C4003 m3_13302_19985# VSS 0.064102f $ **FLOATING
C4004 m2_15612_11606# VSS 0.070212f $ **FLOATING
C4005 m2_11882_23495# VSS 0.065655f $ **FLOATING
C4006 m2_18699_31802# VSS 0.065655f $ **FLOATING
C4007 ringtest_0.x4.counter[8] VSS 0.58641f
C4008 ringtest_0.x4.counter[9] VSS 0.88818f
C4009 ringtest_0.x4.counter[6] VSS 0.659827f
C4010 ringtest_0.x4.counter[5] VSS 0.636589f
C4011 ringtest_0.x4.counter[4] VSS 0.791173f
C4012 ringtest_0.x4.counter[2] VSS 0.606277f
C4013 ringtest_0.x4.counter[1] VSS 0.591348f
C4014 ringtest_0.x4.counter[0] VSS 0.938564f
C4015 a_27815_3867# VSS 0.270206f
C4016 a_27489_3702# VSS 0.257101f
C4017 a_26895_3867# VSS 0.296141f
C4018 a_25975_3867# VSS 0.269288f
C4019 a_25055_3867# VSS 0.278393f
C4020 a_24135_3867# VSS 0.327843f
C4021 a_23399_3867# VSS 0.269041f
C4022 a_22295_3867# VSS 0.276333f
C4023 a_21375_3867# VSS 0.316834f
C4024 a_21007_3867# VSS 0.25238f
C4025 a_27659_4246# VSS 8.84e-19
C4026 a_27303_4246# VSS 0.004608f
C4027 a_26721_4246# VSS 0.01879f
C4028 a_27491_4566# VSS 0.00589f
C4029 a_26913_4566# VSS 0.010025f
C4030 a_26817_4566# VSS 0.006433f
C4031 a_26375_4612# VSS 0.001566f
C4032 a_26269_4612# VSS 0.003693f
C4033 a_26173_4612# VSS 0.003656f
C4034 a_25547_4612# VSS 0.003203f
C4035 a_25441_4612# VSS 0.005457f
C4036 a_25345_4612# VSS 0.005167f
C4037 a_22486_4246# VSS 0.001114f
C4038 a_23467_4584# VSS 0.004685f
C4039 a_22939_4584# VSS 0.007506f
C4040 a_22390_4566# VSS 0.183329f
C4041 a_27273_4220# VSS 0.369297f
C4042 a_26627_4246# VSS 0.344415f
C4043 a_25977_4220# VSS 0.261046f
C4044 a_25149_4220# VSS 0.294745f
C4045 a_23381_4584# VSS 0.255389f
C4046 a_22765_4478# VSS 0.284107f
C4047 a_22164_4362# VSS 0.207092f
C4048 a_22021_4220# VSS 0.20644f
C4049 a_27191_4790# VSS 0.004938f
C4050 ringtest_0.x4.net11 VSS 0.763831f
C4051 a_26766_4790# VSS 0.009249f
C4052 a_27149_5156# VSS 3.75e-19
C4053 a_25719_4790# VSS 0.004164f
C4054 a_26735_5156# VSS 0.002645f
C4055 a_26555_4790# VSS 0.063923f
C4056 a_27065_5156# VSS 0.26998f
C4057 a_27233_5058# VSS 0.379784f
C4058 a_26640_5156# VSS 0.228155f
C4059 a_26808_4902# VSS 0.258239f
C4060 a_26367_4790# VSS 0.335157f
C4061 ringtest_0.x4._09_ VSS 0.545207f
C4062 a_26201_4790# VSS 0.497148f
C4063 a_25294_4790# VSS 0.008691f
C4064 a_25677_5156# VSS 2.5e-19
C4065 a_24551_4790# VSS 7.68e-19
C4066 a_24479_4790# VSS 0.002515f
C4067 a_23963_4790# VSS 0.002664f
C4068 a_23891_4790# VSS 7.95e-19
C4069 a_25263_5156# VSS 7.5e-19
C4070 a_25083_4790# VSS 0.062716f
C4071 a_25593_5156# VSS 0.275541f
C4072 a_25761_5058# VSS 0.356576f
C4073 a_25168_5156# VSS 0.218254f
C4074 a_25336_4902# VSS 0.278138f
C4075 a_24895_4790# VSS 0.323857f
C4076 a_24729_4790# VSS 0.485385f
C4077 a_23467_4818# VSS 0.004685f
C4078 ringtest_0.x4._20_ VSS 0.296302f
C4079 a_22499_4790# VSS 0.004794f
C4080 ringtest_0.x4.net5 VSS 1.52232f
C4081 a_22074_4790# VSS 0.007478f
C4082 a_22457_5156# VSS 3.28e-19
C4083 a_21863_4790# VSS 0.069011f
C4084 a_24317_4942# VSS 0.233023f
C4085 a_23809_4790# VSS 0.25233f
C4086 a_23381_4818# VSS 0.250617f
C4087 a_22373_5156# VSS 0.29125f
C4088 a_22541_5058# VSS 0.405228f
C4089 a_21948_5156# VSS 0.210325f
C4090 a_22116_4902# VSS 0.255348f
C4091 a_21675_4790# VSS 0.417108f
C4092 ringtest_0.x4._03_ VSS 0.578555f
C4093 a_21509_4790# VSS 0.557931f
C4094 a_27149_5334# VSS 0.001033f
C4095 a_26735_5334# VSS 0.002645f
C4096 ringtest_0.x4.net10 VSS 1.58326f
C4097 a_27191_5712# VSS 0.005282f
C4098 a_25309_5334# VSS 0.002002f
C4099 a_26766_5712# VSS 0.010952f
C4100 a_26555_5334# VSS 0.070151f
C4101 a_25351_5712# VSS 0.005844f
C4102 a_23899_5334# VSS 0.014804f
C4103 a_23151_5334# VSS 0.001519f
C4104 a_22795_5334# VSS 0.026188f
C4105 a_22181_5334# VSS 4.07e-19
C4106 a_21767_5334# VSS 6.93e-19
C4107 a_24926_5712# VSS 0.006941f
C4108 a_24715_5334# VSS 0.060618f
C4109 a_23993_5654# VSS 0.006538f
C4110 a_23899_5654# VSS 0.008165f
C4111 a_22983_5654# VSS 0.007253f
C4112 a_22223_5712# VSS 0.004473f
C4113 a_21055_5334# VSS 4.64e-19
C4114 a_21798_5712# VSS 0.008558f
C4115 a_21587_5334# VSS 0.080622f
C4116 a_27065_5334# VSS 0.275172f
C4117 a_27233_5308# VSS 0.371259f
C4118 a_26640_5334# VSS 0.237292f
C4119 a_26808_5308# VSS 0.266551f
C4120 a_26367_5340# VSS 0.344626f
C4121 a_26201_5340# VSS 0.532322f
C4122 a_25225_5334# VSS 0.288597f
C4123 a_25393_5308# VSS 0.391747f
C4124 a_24800_5334# VSS 0.200127f
C4125 a_24968_5308# VSS 0.247676f
C4126 a_24527_5340# VSS 0.312142f
C4127 a_24361_5340# VSS 0.480598f
C4128 a_23770_5308# VSS 0.352433f
C4129 a_22765_5308# VSS 0.430766f
C4130 a_22097_5334# VSS 0.280567f
C4131 a_22265_5308# VSS 0.367396f
C4132 a_21672_5334# VSS 0.214988f
C4133 a_21840_5308# VSS 0.263107f
C4134 a_21399_5340# VSS 0.41156f
C4135 ringtest_0.x4._02_ VSS 0.384112f
C4136 a_21233_5340# VSS 0.551857f
C4137 ringtest_0.x4._14_ VSS 1.2474f
C4138 a_24986_5878# VSS 0.004249f
C4139 a_24545_5878# VSS 0.154917f
C4140 ringtest_0.x4._07_ VSS 0.467795f
C4141 a_23837_5878# VSS 0.204157f
C4142 a_22775_5878# VSS 0.00681f
C4143 ringtest_0.x4._16_ VSS 2.102403f
C4144 ringtest_0.x4._22_ VSS 1.57042f
C4145 a_24627_6200# VSS 8.25e-20
C4146 a_24763_6143# VSS 0.189132f
C4147 ringtest_0.x4.net9 VSS 1.9761f
C4148 ringtest_0.x4._06_ VSS 0.355082f
C4149 ringtest_0.x4._21_ VSS 0.491639f
C4150 a_23932_6128# VSS 9.9e-19
C4151 a_22350_5878# VSS 0.007439f
C4152 a_22733_6244# VSS 0.002478f
C4153 a_22319_6244# VSS 5.31e-19
C4154 a_22139_5878# VSS 0.062654f
C4155 a_25364_5878# VSS 2.07482f
C4156 a_24699_6200# VSS 0.166512f
C4157 a_24004_6128# VSS 0.208373f
C4158 a_24070_5852# VSS 0.228425f
C4159 ringtest_0.x4.net8 VSS 1.78641f
C4160 a_22649_6244# VSS 0.331871f
C4161 a_22817_6146# VSS 0.427232f
C4162 a_22224_6244# VSS 0.220057f
C4163 a_22392_5990# VSS 0.267836f
C4164 a_21951_5878# VSS 0.384412f
C4165 ringtest_0.x4._04_ VSS 0.647447f
C4166 a_21785_5878# VSS 0.561386f
C4167 a_21591_6128# VSS 0.005123f
C4168 ringtest_0.x4._13_ VSS 1.13412f
C4169 ringtest_0.x4.net4 VSS 1.31635f
C4170 ringtest_0.x4._08_ VSS 0.728198f
C4171 a_26839_6788# VSS 0.008414f
C4172 a_26201_6788# VSS 0.003851f
C4173 a_26095_6788# VSS 0.003674f
C4174 a_26007_6788# VSS 0.001688f
C4175 a_24287_6422# VSS 7.93e-19
C4176 a_24883_6800# VSS 0.060853f
C4177 a_24685_6788# VSS 0.006624f
C4178 a_24264_6788# VSS 0.005539f
C4179 a_23619_6788# VSS 0.005238f
C4180 ringtest_0.x4._25_ VSS 0.368024f
C4181 a_27169_6641# VSS 0.273817f
C4182 a_26749_6422# VSS 0.263282f
C4183 ringtest_0.x4._24_ VSS 0.69832f
C4184 a_26569_6422# VSS 0.271803f
C4185 ringtest_0.x4._23_ VSS 0.976575f
C4186 a_25925_6788# VSS 0.264561f
C4187 ringtest_0.x4._15_ VSS 3.54948f
C4188 ringtest_0.x4.net7 VSS 2.72071f
C4189 ringtest_0.x4.net6 VSS 3.218643f
C4190 ringtest_0.x4._19_ VSS 0.32708f
C4191 a_25421_6641# VSS 0.252712f
C4192 ringtest_0.x4.clknet_1_1__leaf_clk VSS 3.414301f
C4193 ringtest_0.x4._05_ VSS 0.318608f
C4194 a_24465_6800# VSS 0.241882f
C4195 a_24536_6699# VSS 0.198121f
C4196 a_24336_6544# VSS 0.303545f
C4197 a_24329_6640# VSS 0.46613f
C4198 a_24045_6654# VSS 0.281525f
C4199 a_23949_6654# VSS 0.378965f
C4200 a_23529_6422# VSS 0.234926f
C4201 ringtest_0.x4._18_ VSS 0.468402f
C4202 a_23349_6422# VSS 0.254342f
C4203 ringtest_0.x4._17_ VSS 0.622485f
C4204 ringtest_0.counter7 VSS 17.349024f
C4205 a_23879_6940# VSS 2.29287f
C4206 ringtest_0.x4.clknet_0_clk VSS 4.193551f
C4207 a_21395_6940# VSS 2.29289f
C4208 a_21939_8054# VSS 0.002457f
C4209 a_21867_8054# VSS 0.001303f
C4210 a_22695_8304# VSS 0.005104f
C4211 ringtest_0.counter3 VSS 14.338387f
C4212 ringtest_0.x4._11_ VSS 5.669866f
C4213 a_22245_8054# VSS 0.298451f
C4214 ringtest_0.x4._10_ VSS 0.339714f
C4215 a_21785_8054# VSS 0.252154f
C4216 a_21803_8598# VSS 6.89e-19
C4217 a_22399_8976# VSS 0.064411f
C4218 a_22201_8964# VSS 0.006624f
C4219 a_21049_8598# VSS 0.017559f
C4220 a_21780_8964# VSS 0.004183f
C4221 ringtest_0.x4._12_ VSS 1.2616f
C4222 a_21132_8918# VSS 0.004429f
C4223 ringtest_0.x4._01_ VSS 0.405148f
C4224 a_21981_8976# VSS 0.238144f
C4225 a_22052_8875# VSS 0.195482f
C4226 a_21852_8720# VSS 0.31379f
C4227 a_21845_8816# VSS 0.552106f
C4228 a_21561_8830# VSS 0.279727f
C4229 a_21465_8830# VSS 0.390267f
C4230 ringtest_0.x4.net3 VSS 2.298238f
C4231 a_22201_9142# VSS 0.007478f
C4232 a_21780_9142# VSS 0.004654f
C4233 ringtest_0.x4.clknet_1_0__leaf_clk VSS 4.010709f
C4234 a_22399_9142# VSS 0.069779f
C4235 a_21803_9508# VSS 6.84e-19
C4236 a_21981_9142# VSS 0.264386f
C4237 a_22052_9116# VSS 0.210923f
C4238 a_21845_9116# VSS 0.580201f
C4239 a_21852_9416# VSS 0.340144f
C4240 a_21561_9116# VSS 0.287469f
C4241 a_21465_9294# VSS 0.412387f
C4242 a_21675_9686# VSS 0.013142f
C4243 a_21507_9686# VSS 0.006974f
C4244 ringtest_0.x4._00_ VSS 0.757573f
C4245 a_21675_10006# VSS 0.006222f
C4246 a_21425_9686# VSS 0.393994f
C4247 ringtest_0.x4.net2 VSS 3.500251f
C4248 ringtest_0.x4.net1 VSS 1.81106f
C4249 a_22111_10993# VSS 0.293097f
C4250 ringtest_0.x3.x2.GP3 VSS 1.64575f
C4251 ringtest_0.x3.x2.GP2 VSS 5.54164f
C4252 ringtest_0.x3.x2.GP1 VSS 4.63625f
C4253 a_17405_12123# VSS 0.006782f
C4254 ringtest_0.x3.x2.GN4 VSS 3.79271f
C4255 a_16707_12151# VSS 0.007327f
C4256 ringtest_0.x3.x2.GN3 VSS 3.64172f
C4257 a_16155_12151# VSS 0.004704f
C4258 ringtest_0.x3.x2.GN2 VSS 3.91967f
C4259 a_15749_12123# VSS 0.006793f
C4260 ringtest_0.x3.x2.GN1 VSS 4.84443f
C4261 a_17231_12017# VSS 0.3167f
C4262 a_16755_12091# VSS 0.251626f
C4263 a_16579_11759# VSS 0.236732f
C4264 a_16203_12091# VSS 0.236633f
C4265 a_16027_11759# VSS 0.222621f
C4266 a_15575_12017# VSS 0.270062f
C4267 ringtest_0.x3.nselect2 VSS 0.455447f
C4268 ringtest_0.x3.x1.nSEL1 VSS 0.740163f
C4269 ringtest_0.x3.x1.nSEL0 VSS 0.685116f
C4270 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VSS 0.505562f
C4271 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VSS 0.498424f
C4272 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VSS 0.498285f
C4273 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VSS 0.499488f
C4274 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VSS 0.500758f
C4275 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VSS 0.50136f
C4276 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VSS 0.501617f
C4277 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VSS 0.52312f
C4278 ringtest_0.drv_out VSS 29.368195f
C4279 a_17377_14114# VSS 0.332619f
C4280 ringtest_0.ring_out VSS 16.289782f
C4281 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VSS 0.632983f
C4282 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VSS 0.508122f
C4283 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VSS 0.498331f
C4284 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VSS 0.498331f
C4285 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VSS 0.498339f
C4286 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VSS 0.498632f
C4287 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VSS 0.498682f
C4288 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VSS 0.498707f
C4289 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VSS 0.507755f
C4290 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VSS 0.971227f
C4291 muxtest_0.x2.x2.GP3 VSS 1.68554f
C4292 muxtest_0.x2.x2.GP2 VSS 5.5641f
C4293 muxtest_0.x2.x2.GP1 VSS 4.625069f
C4294 muxtest_0.R1R2 VSS 6.645505f
C4295 a_13675_24012# VSS 0.006439f
C4296 muxtest_0.x2.x2.GN4 VSS 3.796f
C4297 a_12977_24040# VSS 0.006801f
C4298 muxtest_0.x2.x2.GN3 VSS 3.65554f
C4299 a_12425_24040# VSS 0.004461f
C4300 muxtest_0.x2.x2.GN2 VSS 3.88834f
C4301 a_12019_24012# VSS 0.006505f
C4302 muxtest_0.x2.x2.GN1 VSS 4.79625f
C4303 a_13501_23906# VSS 0.306555f
C4304 a_13025_23980# VSS 0.249538f
C4305 a_12849_23648# VSS 0.232764f
C4306 a_12473_23980# VSS 0.23458f
C4307 a_12297_23648# VSS 0.220868f
C4308 a_11845_23906# VSS 0.267622f
C4309 muxtest_0.x2.nselect2 VSS 0.451665f
C4310 muxtest_0.x2.x1.nSEL1 VSS 0.686441f
C4311 muxtest_0.x2.x1.nSEL0 VSS 0.647345f
C4312 muxtest_0.R2R3 VSS 7.982832f
C4313 muxtest_0.R3R4 VSS 15.859409f
C4314 muxtest_0.R4R5 VSS 7.656276f
C4315 muxtest_0.R5R6 VSS 7.957228f
C4316 muxtest_0.R6R7 VSS 7.795067f
C4317 muxtest_0.R7R8 VSS 29.82938f
C4318 muxtest_0.x1.x5.A VSS 13.867701f
C4319 muxtest_0.x1.x4.A VSS 16.1317f
C4320 muxtest_0.x1.x3.GP3 VSS 3.18231f
C4321 muxtest_0.x1.x3.GP2 VSS 10.304811f
C4322 muxtest_0.x1.x3.GP1 VSS 10.781407f
C4323 a_20492_32319# VSS 0.006616f
C4324 muxtest_0.x1.x3.GN4 VSS 7.04004f
C4325 a_19794_32347# VSS 0.006984f
C4326 muxtest_0.x1.x3.GN3 VSS 6.77674f
C4327 a_19242_32347# VSS 0.004523f
C4328 muxtest_0.x1.x3.GN2 VSS 7.175951f
C4329 a_18836_32319# VSS 0.006515f
C4330 muxtest_0.x1.x3.GN1 VSS 8.91731f
C4331 a_20318_32213# VSS 0.311491f
C4332 a_19842_32287# VSS 0.24978f
C4333 a_19666_31955# VSS 0.233122f
C4334 a_19290_32287# VSS 0.234813f
C4335 a_19114_31955# VSS 0.221018f
C4336 a_18662_32213# VSS 0.267639f
C4337 muxtest_0.x1.x5.GN VSS 5.73587f
C4338 muxtest_0.x1.x1.nSEL1 VSS 0.683011f
C4339 muxtest_0.x1.x1.nSEL0 VSS 0.650421f
C4340 ui_in[5].t1 VSS 0.0025f
C4341 ui_in[5].t0 VSS 0.004008f
C4342 ui_in[5].n0 VSS 0.008077f
C4343 ui_in[5].n1 VSS 0.003407f
C4344 ui_in[5].n2 VSS 0.33124f
C4345 ui_in[5].n3 VSS 3.27797f
C4346 ui_in[6].t0 VSS 0.00254f
C4347 ui_in[6].t2 VSS 0.001497f
C4348 ui_in[6].n0 VSS 0.003424f
C4349 ui_in[6].t1 VSS 0.00254f
C4350 ui_in[6].t3 VSS 0.001497f
C4351 ui_in[6].n1 VSS 0.003424f
C4352 ui_in[6].n2 VSS 0.001687f
C4353 ui_in[6].n3 VSS 0.224459f
C4354 muxtest_0.R2R3.t0 VSS 0.626391f
C4355 muxtest_0.R2R3.t1 VSS 0.443113f
C4356 muxtest_0.R2R3.n0 VSS 3.43546f
C4357 muxtest_0.R2R3.t2 VSS 0.347912f
C4358 muxtest_0.R2R3.t3 VSS 0.638083f
C4359 muxtest_0.R2R3.n1 VSS 3.5698f
C4360 muxtest_0.R2R3.n2 VSS 0.568983f
C4361 muxtest_0.R2R3.n3 VSS 0.116677f
C4362 muxtest_0.R2R3.t4 VSS 0.210663f
C4363 muxtest_0.R2R3.t5 VSS 0.170342f
C4364 muxtest_0.R2R3.n4 VSS 3.38019f
C4365 muxtest_0.R4R5.t1 VSS 0.627578f
C4366 muxtest_0.R4R5.t2 VSS 0.443953f
C4367 muxtest_0.R4R5.n0 VSS 3.44197f
C4368 muxtest_0.R4R5.t4 VSS 0.348571f
C4369 muxtest_0.R4R5.t5 VSS 0.639293f
C4370 muxtest_0.R4R5.n1 VSS 3.57657f
C4371 muxtest_0.R4R5.n2 VSS 0.570061f
C4372 muxtest_0.R4R5.n3 VSS 0.119407f
C4373 muxtest_0.R4R5.t0 VSS 0.212944f
C4374 muxtest_0.R4R5.t3 VSS 0.170665f
C4375 muxtest_0.R4R5.n4 VSS 3.47489f
C4376 muxtest_0.x2.x2.x4.GP VSS 2.57727f
C4377 muxtest_0.x2.x1.gpo3 VSS 1.20603f
C4378 muxtest_0.x2.x2.GP4.t1 VSS 0.012374f
C4379 muxtest_0.x2.x2.GP4.t0 VSS 0.012374f
C4380 muxtest_0.x2.x2.GP4.n0 VSS 0.027184f
C4381 muxtest_0.x2.x1.x14.Y VSS 0.076955f
C4382 muxtest_0.x2.x2.GP4.n1 VSS 0.01052f
C4383 muxtest_0.x2.x2.GP4.t5 VSS 0.626223f
C4384 muxtest_0.x2.x2.GP4.t4 VSS 0.643686f
C4385 muxtest_0.x2.x2.GP4.n2 VSS 2.28835f
C4386 muxtest_0.x2.x2.GP4.n3 VSS 0.048401f
C4387 muxtest_0.x2.x2.GP4.t3 VSS 0.019037f
C4388 muxtest_0.x2.x2.GP4.t2 VSS 0.019037f
C4389 muxtest_0.x2.x2.GP4.n4 VSS 0.043773f
C4390 muxtest_0.x2.x2.GP4.n5 VSS 0.088779f
C4391 ringtest_0.x3.x2.GP2.t1 VSS 0.016198f
C4392 ringtest_0.x3.x2.GP2.t0 VSS 0.016198f
C4393 ringtest_0.x3.x2.GP2.n0 VSS 0.035585f
C4394 ringtest_0.x3.x2.GP2.n1 VSS 0.023f
C4395 ringtest_0.x3.x2.GP2.t5 VSS 0.819754f
C4396 ringtest_0.x3.x2.GP2.t4 VSS 0.842614f
C4397 ringtest_0.x3.x2.GP2.n2 VSS 2.98946f
C4398 ringtest_0.x3.x2.GP2.t3 VSS 0.02492f
C4399 ringtest_0.x3.x2.GP2.t2 VSS 0.02492f
C4400 ringtest_0.x3.x2.GP2.n3 VSS 0.051391f
C4401 ringtest_0.x3.x2.GP2.n4 VSS 0.120168f
C4402 ringtest_0.x3.x2.GP2.n5 VSS 0.027176f
C4403 ringtest_0.ring_out.t13 VSS 0.143976f
C4404 ringtest_0.ring_out.t12 VSS 0.066482f
C4405 ringtest_0.ring_out.n0 VSS 1.43742f
C4406 ringtest_0.ring_out.t2 VSS 0.011895f
C4407 ringtest_0.ring_out.t1 VSS 0.011895f
C4408 ringtest_0.ring_out.n1 VSS 0.036116f
C4409 ringtest_0.ring_out.t7 VSS 0.011895f
C4410 ringtest_0.ring_out.t8 VSS 0.011895f
C4411 ringtest_0.ring_out.n2 VSS 0.026441f
C4412 ringtest_0.ring_out.n3 VSS 0.119642f
C4413 ringtest_0.ring_out.t9 VSS 0.007732f
C4414 ringtest_0.ring_out.t0 VSS 0.007732f
C4415 ringtest_0.ring_out.n4 VSS 0.017154f
C4416 ringtest_0.ring_out.n5 VSS 0.032249f
C4417 ringtest_0.ring_out.n6 VSS 0.009203f
C4418 ringtest_0.ring_out.t14 VSS 0.010903f
C4419 ringtest_0.ring_out.t10 VSS 0.018503f
C4420 ringtest_0.ring_out.t15 VSS 0.010903f
C4421 ringtest_0.ring_out.t11 VSS 0.018503f
C4422 ringtest_0.ring_out.n7 VSS 0.031045f
C4423 ringtest_0.ring_out.n8 VSS 0.04596f
C4424 ringtest_0.ring_out.n9 VSS 0.181049f
C4425 ringtest_0.ring_out.n10 VSS 0.421446f
C4426 ringtest_0.ring_out.t5 VSS 0.673389f
C4427 ringtest_0.ring_out.t6 VSS 0.47636f
C4428 ringtest_0.ring_out.n11 VSS 3.69323f
C4429 ringtest_0.ring_out.t3 VSS 0.374016f
C4430 ringtest_0.ring_out.t4 VSS 0.685959f
C4431 ringtest_0.ring_out.n12 VSS 3.83764f
C4432 ringtest_0.ring_out.n13 VSS 0.611674f
C4433 ringtest_0.x3.x2.GP1.t1 VSS 0.012908f
C4434 ringtest_0.x3.x2.GP1.t0 VSS 0.012908f
C4435 ringtest_0.x3.x2.GP1.n0 VSS 0.028358f
C4436 ringtest_0.x3.x2.GP1.n1 VSS 0.018329f
C4437 ringtest_0.x3.x2.GP1.t4 VSS 0.653268f
C4438 ringtest_0.x3.x2.GP1.t5 VSS 0.671486f
C4439 ringtest_0.x3.x2.GP1.n2 VSS 2.37213f
C4440 ringtest_0.x3.x2.GP1.t3 VSS 0.019859f
C4441 ringtest_0.x3.x2.GP1.t2 VSS 0.019859f
C4442 ringtest_0.x3.x2.GP1.n3 VSS 0.04092f
C4443 ringtest_0.x3.x2.GP1.n4 VSS 0.100085f
C4444 ringtest_0.x3.x2.GP1.n5 VSS 0.021877f
C4445 ui_in[3].t3 VSS 0.007332f
C4446 ui_in[3].t12 VSS 0.00432f
C4447 ui_in[3].t18 VSS 0.007332f
C4448 ui_in[3].t2 VSS 0.00432f
C4449 ui_in[3].n0 VSS 0.012301f
C4450 ui_in[3].n1 VSS 0.018181f
C4451 ui_in[3].n2 VSS 0.005713f
C4452 ui_in[3].t6 VSS 0.003611f
C4453 ui_in[3].t10 VSS 0.005245f
C4454 ui_in[3].n3 VSS 0.012493f
C4455 ui_in[3].n4 VSS 0.006939f
C4456 ui_in[3].t9 VSS 0.004276f
C4457 ui_in[3].t19 VSS 0.006297f
C4458 ui_in[3].n5 VSS 0.014878f
C4459 ui_in[3].n6 VSS 0.00309f
C4460 ui_in[3].n7 VSS 0.001204f
C4461 ui_in[3].n8 VSS 0.110032f
C4462 ui_in[3].t17 VSS 0.007155f
C4463 ui_in[3].t15 VSS 0.003393f
C4464 ui_in[3].n9 VSS 0.025691f
C4465 ui_in[3].n10 VSS 0.004978f
C4466 ui_in[3].n11 VSS 0.126236f
C4467 ui_in[3].n12 VSS 0.082029f
C4468 ui_in[3].t8 VSS 0.007332f
C4469 ui_in[3].t16 VSS 0.00432f
C4470 ui_in[3].t5 VSS 0.007332f
C4471 ui_in[3].t13 VSS 0.00432f
C4472 ui_in[3].n13 VSS 0.012301f
C4473 ui_in[3].n14 VSS 0.018181f
C4474 ui_in[3].n15 VSS 0.005713f
C4475 ui_in[3].t7 VSS 0.003611f
C4476 ui_in[3].t11 VSS 0.005245f
C4477 ui_in[3].n16 VSS 0.012493f
C4478 ui_in[3].n17 VSS 0.006939f
C4479 ui_in[3].t14 VSS 0.004276f
C4480 ui_in[3].t0 VSS 0.006297f
C4481 ui_in[3].n18 VSS 0.014878f
C4482 ui_in[3].n19 VSS 0.00309f
C4483 ui_in[3].n20 VSS 0.001204f
C4484 ui_in[3].n21 VSS 0.110032f
C4485 ui_in[3].t4 VSS 0.007155f
C4486 ui_in[3].t1 VSS 0.003393f
C4487 ui_in[3].n22 VSS 0.025691f
C4488 ui_in[3].n23 VSS 0.004978f
C4489 ui_in[3].n24 VSS 0.126236f
C4490 ui_in[3].n25 VSS 0.082029f
C4491 ui_in[3].n26 VSS 10.0315f
C4492 muxtest_0.R7R8.t4 VSS 0.570638f
C4493 muxtest_0.R7R8.t3 VSS 0.403673f
C4494 muxtest_0.R7R8.n0 VSS 3.12968f
C4495 muxtest_0.R7R8.t0 VSS 0.316945f
C4496 muxtest_0.R7R8.t1 VSS 0.58129f
C4497 muxtest_0.R7R8.n1 VSS 3.25206f
C4498 muxtest_0.R7R8.n2 VSS 0.51834f
C4499 muxtest_0.R7R8.n3 VSS 0.107649f
C4500 muxtest_0.R7R8.t9 VSS 0.157299f
C4501 muxtest_0.R7R8.t2 VSS 0.858788f
C4502 muxtest_0.R7R8.n4 VSS 1.55412f
C4503 muxtest_0.R7R8.t5 VSS 0.570638f
C4504 muxtest_0.R7R8.t6 VSS 0.403673f
C4505 muxtest_0.R7R8.n5 VSS 3.12968f
C4506 muxtest_0.R7R8.t7 VSS 0.316945f
C4507 muxtest_0.R7R8.t8 VSS 0.58129f
C4508 muxtest_0.R7R8.n6 VSS 3.25206f
C4509 muxtest_0.R7R8.n7 VSS 0.51834f
C4510 muxtest_0.R7R8.n8 VSS 0.108573f
C4511 muxtest_0.R7R8.n9 VSS 9.50513f
C4512 ua[0].t5 VSS 0.319126f
C4513 ua[0].t6 VSS 0.225752f
C4514 ua[0].n0 VSS 1.75026f
C4515 ua[0].t8 VSS 0.17725f
C4516 ua[0].t7 VSS 0.325083f
C4517 ua[0].n1 VSS 1.8187f
C4518 ua[0].n2 VSS 0.289879f
C4519 ua[0].n3 VSS 0.060719f
C4520 ua[0].t4 VSS 0.086784f
C4521 ua[0].n4 VSS 1.50131f
C4522 ua[0].n5 VSS 11.5833f
C4523 ua[0].t3 VSS 0.319126f
C4524 ua[0].t2 VSS 0.225752f
C4525 ua[0].n6 VSS 1.75026f
C4526 ua[0].t1 VSS 0.17725f
C4527 ua[0].t0 VSS 0.325083f
C4528 ua[0].n7 VSS 1.8187f
C4529 ua[0].n8 VSS 0.289879f
C4530 ua[0].n9 VSS 0.059443f
C4531 muxtest_0.R6R7.t1 VSS 0.693927f
C4532 muxtest_0.R6R7.t0 VSS 0.490889f
C4533 muxtest_0.R6R7.n0 VSS 3.80587f
C4534 muxtest_0.R6R7.t2 VSS 0.385423f
C4535 muxtest_0.R6R7.t3 VSS 0.706881f
C4536 muxtest_0.R6R7.n1 VSS 3.95469f
C4537 muxtest_0.R6R7.n2 VSS 0.63033f
C4538 muxtest_0.R6R7.n3 VSS 0.129257f
C4539 muxtest_0.R6R7.t4 VSS 0.920517f
C4540 muxtest_0.R6R7.t5 VSS 0.188708f
C4541 muxtest_0.R6R7.n4 VSS 2.80582f
C4542 muxtest_0.R6R7.n5 VSS 1.24461f
C4543 muxtest_0.x2.x2.GP2.t0 VSS 0.016198f
C4544 muxtest_0.x2.x2.GP2.t1 VSS 0.016198f
C4545 muxtest_0.x2.x2.GP2.n0 VSS 0.035585f
C4546 muxtest_0.x2.x2.GP2.n1 VSS 0.023f
C4547 muxtest_0.x2.x2.GP2.t5 VSS 0.819754f
C4548 muxtest_0.x2.x2.GP2.t4 VSS 0.842614f
C4549 muxtest_0.x2.x2.GP2.n2 VSS 2.98946f
C4550 muxtest_0.x2.x2.GP2.t3 VSS 0.02492f
C4551 muxtest_0.x2.x2.GP2.t2 VSS 0.02492f
C4552 muxtest_0.x2.x2.GP2.n3 VSS 0.051391f
C4553 muxtest_0.x2.x2.GP2.n4 VSS 0.120168f
C4554 muxtest_0.x2.x2.GP2.n5 VSS 0.027176f
C4555 ringtest_0.x4._16_.t0 VSS 0.046376f
C4556 ringtest_0.x4._16_.n0 VSS 0.026397f
C4557 ringtest_0.x4._16_.t7 VSS 0.021164f
C4558 ringtest_0.x4._16_.t2 VSS 0.017507f
C4559 ringtest_0.x4._16_.n1 VSS 0.047954f
C4560 ringtest_0.x4._16_.n2 VSS 0.154756f
C4561 ringtest_0.x4._16_.t9 VSS 0.020065f
C4562 ringtest_0.x4._16_.t3 VSS 0.031953f
C4563 ringtest_0.x4._16_.n3 VSS 0.045672f
C4564 ringtest_0.x4._16_.n4 VSS 0.0375f
C4565 ringtest_0.x4._16_.t4 VSS 0.020065f
C4566 ringtest_0.x4._16_.t8 VSS 0.031953f
C4567 ringtest_0.x4._16_.n5 VSS 0.058943f
C4568 ringtest_0.x4._16_.n6 VSS 0.063595f
C4569 ringtest_0.x4._16_.n7 VSS 0.426096f
C4570 ringtest_0.x4._16_.t5 VSS 0.012893f
C4571 ringtest_0.x4._16_.t6 VSS 0.013824f
C4572 ringtest_0.x4._16_.n8 VSS 0.03796f
C4573 ringtest_0.x4._16_.n9 VSS 0.022428f
C4574 ringtest_0.x4._16_.n10 VSS 0.327394f
C4575 ringtest_0.x4._16_.n11 VSS 0.020414f
C4576 ringtest_0.x4._16_.t1 VSS 0.119992f
C4577 ringtest_0.x4._16_.n12 VSS 0.021583f
C4578 ringtest_0.x4._16_.n13 VSS 0.021194f
C4579 muxtest_0.R5R6.t0 VSS 0.695132f
C4580 muxtest_0.R5R6.t1 VSS 0.491742f
C4581 muxtest_0.R5R6.n0 VSS 3.81248f
C4582 muxtest_0.R5R6.t5 VSS 0.386092f
C4583 muxtest_0.R5R6.t4 VSS 0.708108f
C4584 muxtest_0.R5R6.n1 VSS 3.96156f
C4585 muxtest_0.R5R6.n2 VSS 0.631424f
C4586 muxtest_0.R5R6.n3 VSS 0.129973f
C4587 muxtest_0.R5R6.t3 VSS 0.191095f
C4588 muxtest_0.R5R6.t2 VSS 1.13104f
C4589 muxtest_0.R5R6.n4 VSS 2.8297f
C4590 muxtest_0.x1.x3.GP2.t0 VSS 0.018287f
C4591 muxtest_0.x1.x3.GP2.t1 VSS 0.018287f
C4592 muxtest_0.x1.x3.GP2.n0 VSS 0.040174f
C4593 muxtest_0.x1.x3.GP2.n1 VSS 0.025967f
C4594 muxtest_0.x1.x3.GP2.t6 VSS 0.925483f
C4595 muxtest_0.x1.x3.GP2.t7 VSS 0.951291f
C4596 muxtest_0.x1.x3.GP2.n2 VSS 3.37503f
C4597 muxtest_0.x1.x3.GP2.t5 VSS 0.925483f
C4598 muxtest_0.x1.x3.GP2.t4 VSS 0.951291f
C4599 muxtest_0.x1.x3.GP2.n3 VSS 3.37503f
C4600 muxtest_0.x1.x3.GP2.n4 VSS 1.97357f
C4601 muxtest_0.x1.x3.GP2.t2 VSS 0.028134f
C4602 muxtest_0.x1.x3.GP2.t3 VSS 0.028134f
C4603 muxtest_0.x1.x3.GP2.n5 VSS 0.058019f
C4604 muxtest_0.x1.x3.GP2.n6 VSS 0.132927f
C4605 muxtest_0.x1.x3.GP2.n7 VSS 0.030681f
C4606 ringtest_0.counter3.t3 VSS 0.033829f
C4607 ringtest_0.counter3.n0 VSS 0.005886f
C4608 ringtest_0.counter3.t2 VSS 0.023398f
C4609 ringtest_0.counter3.n1 VSS 0.028682f
C4610 ringtest_0.counter3.n2 VSS 0.036901f
C4611 ringtest_0.counter3.n3 VSS 0.371589f
C4612 ringtest_0.counter3.t1 VSS 0.740343f
C4613 ringtest_0.counter3.t0 VSS 0.523724f
C4614 ringtest_0.counter3.n4 VSS 4.06044f
C4615 ringtest_0.counter3.t4 VSS 0.410954f
C4616 ringtest_0.counter3.t5 VSS 0.761665f
C4617 ringtest_0.counter3.n5 VSS 4.29752f
C4618 ringtest_0.counter3.n6 VSS 0.672491f
C4619 ringtest_0.x4.clknet_1_0__leaf_clk.t38 VSS 0.022262f
C4620 ringtest_0.x4.clknet_1_0__leaf_clk.t41 VSS 0.014894f
C4621 ringtest_0.x4.clknet_1_0__leaf_clk.n0 VSS 0.04068f
C4622 ringtest_0.x4.clknet_1_0__leaf_clk.n1 VSS 0.107083f
C4623 ringtest_0.x4.clknet_1_0__leaf_clk.t37 VSS 0.014894f
C4624 ringtest_0.x4.clknet_1_0__leaf_clk.t32 VSS 0.022262f
C4625 ringtest_0.x4.clknet_1_0__leaf_clk.n2 VSS 0.041145f
C4626 ringtest_0.x4.clknet_1_0__leaf_clk.n3 VSS 0.437523f
C4627 ringtest_0.x4.clknet_1_0__leaf_clk.t30 VSS 0.014222f
C4628 ringtest_0.x4.clknet_1_0__leaf_clk.t16 VSS 0.014222f
C4629 ringtest_0.x4.clknet_1_0__leaf_clk.n4 VSS 0.029978f
C4630 ringtest_0.x4.clknet_1_0__leaf_clk.t27 VSS 0.014222f
C4631 ringtest_0.x4.clknet_1_0__leaf_clk.t29 VSS 0.014222f
C4632 ringtest_0.x4.clknet_1_0__leaf_clk.n5 VSS 0.029589f
C4633 ringtest_0.x4.clknet_1_0__leaf_clk.t8 VSS 0.005973f
C4634 ringtest_0.x4.clknet_1_0__leaf_clk.t11 VSS 0.005973f
C4635 ringtest_0.x4.clknet_1_0__leaf_clk.n6 VSS 0.021211f
C4636 ringtest_0.x4.clknet_1_0__leaf_clk.t13 VSS 0.005973f
C4637 ringtest_0.x4.clknet_1_0__leaf_clk.t15 VSS 0.005973f
C4638 ringtest_0.x4.clknet_1_0__leaf_clk.n7 VSS 0.013636f
C4639 ringtest_0.x4.clknet_1_0__leaf_clk.n8 VSS 0.086164f
C4640 ringtest_0.x4.clknet_1_0__leaf_clk.t10 VSS 0.005973f
C4641 ringtest_0.x4.clknet_1_0__leaf_clk.t12 VSS 0.005973f
C4642 ringtest_0.x4.clknet_1_0__leaf_clk.n9 VSS 0.013636f
C4643 ringtest_0.x4.clknet_1_0__leaf_clk.n10 VSS 0.051791f
C4644 ringtest_0.x4.clknet_1_0__leaf_clk.t14 VSS 0.005973f
C4645 ringtest_0.x4.clknet_1_0__leaf_clk.t9 VSS 0.005973f
C4646 ringtest_0.x4.clknet_1_0__leaf_clk.n11 VSS 0.013644f
C4647 ringtest_0.x4.clknet_1_0__leaf_clk.n12 VSS 0.053424f
C4648 ringtest_0.x4.clknet_1_0__leaf_clk.t1 VSS 0.005973f
C4649 ringtest_0.x4.clknet_1_0__leaf_clk.t4 VSS 0.005973f
C4650 ringtest_0.x4.clknet_1_0__leaf_clk.n13 VSS 0.013636f
C4651 ringtest_0.x4.clknet_1_0__leaf_clk.n14 VSS 0.051791f
C4652 ringtest_0.x4.clknet_1_0__leaf_clk.t6 VSS 0.005973f
C4653 ringtest_0.x4.clknet_1_0__leaf_clk.t7 VSS 0.005973f
C4654 ringtest_0.x4.clknet_1_0__leaf_clk.n15 VSS 0.013636f
C4655 ringtest_0.x4.clknet_1_0__leaf_clk.n16 VSS 0.05205f
C4656 ringtest_0.x4.clknet_1_0__leaf_clk.t3 VSS 0.005973f
C4657 ringtest_0.x4.clknet_1_0__leaf_clk.t5 VSS 0.005973f
C4658 ringtest_0.x4.clknet_1_0__leaf_clk.n17 VSS 0.013636f
C4659 ringtest_0.x4.clknet_1_0__leaf_clk.n18 VSS 0.04471f
C4660 ringtest_0.x4.clknet_1_0__leaf_clk.t0 VSS 0.005973f
C4661 ringtest_0.x4.clknet_1_0__leaf_clk.t2 VSS 0.005973f
C4662 ringtest_0.x4.clknet_1_0__leaf_clk.n19 VSS 0.013163f
C4663 ringtest_0.x4.clknet_1_0__leaf_clk.n20 VSS 0.043256f
C4664 ringtest_0.x4.clknet_1_0__leaf_clk.n21 VSS 0.09308f
C4665 ringtest_0.x4.clknet_1_0__leaf_clk.n22 VSS 0.067594f
C4666 ringtest_0.x4.clknet_1_0__leaf_clk.t19 VSS 0.014222f
C4667 ringtest_0.x4.clknet_1_0__leaf_clk.t22 VSS 0.014222f
C4668 ringtest_0.x4.clknet_1_0__leaf_clk.n23 VSS 0.036128f
C4669 ringtest_0.x4.clknet_1_0__leaf_clk.t24 VSS 0.014222f
C4670 ringtest_0.x4.clknet_1_0__leaf_clk.t26 VSS 0.014222f
C4671 ringtest_0.x4.clknet_1_0__leaf_clk.n24 VSS 0.029978f
C4672 ringtest_0.x4.clknet_1_0__leaf_clk.n25 VSS 0.136621f
C4673 ringtest_0.x4.clknet_1_0__leaf_clk.t21 VSS 0.014222f
C4674 ringtest_0.x4.clknet_1_0__leaf_clk.t23 VSS 0.014222f
C4675 ringtest_0.x4.clknet_1_0__leaf_clk.n26 VSS 0.029978f
C4676 ringtest_0.x4.clknet_1_0__leaf_clk.n27 VSS 0.0787f
C4677 ringtest_0.x4.clknet_1_0__leaf_clk.t25 VSS 0.014222f
C4678 ringtest_0.x4.clknet_1_0__leaf_clk.t20 VSS 0.014222f
C4679 ringtest_0.x4.clknet_1_0__leaf_clk.n28 VSS 0.029978f
C4680 ringtest_0.x4.clknet_1_0__leaf_clk.n29 VSS 0.078334f
C4681 ringtest_0.x4.clknet_1_0__leaf_clk.t28 VSS 0.014222f
C4682 ringtest_0.x4.clknet_1_0__leaf_clk.t31 VSS 0.014222f
C4683 ringtest_0.x4.clknet_1_0__leaf_clk.n30 VSS 0.029978f
C4684 ringtest_0.x4.clknet_1_0__leaf_clk.n31 VSS 0.078334f
C4685 ringtest_0.x4.clknet_1_0__leaf_clk.n32 VSS 0.04742f
C4686 ringtest_0.x4.clknet_1_0__leaf_clk.t17 VSS 0.014222f
C4687 ringtest_0.x4.clknet_1_0__leaf_clk.t18 VSS 0.014222f
C4688 ringtest_0.x4.clknet_1_0__leaf_clk.n33 VSS 0.028445f
C4689 ringtest_0.x4.clknet_1_0__leaf_clk.n34 VSS 0.022411f
C4690 ringtest_0.x4.clknet_1_0__leaf_clk.n35 VSS 0.171468f
C4691 ringtest_0.x4.clknet_1_0__leaf_clk.t39 VSS 0.014894f
C4692 ringtest_0.x4.clknet_1_0__leaf_clk.t36 VSS 0.022262f
C4693 ringtest_0.x4.clknet_1_0__leaf_clk.n36 VSS 0.040782f
C4694 ringtest_0.x4.clknet_1_0__leaf_clk.n37 VSS 0.024896f
C4695 ringtest_0.x4.clknet_1_0__leaf_clk.t33 VSS 0.022262f
C4696 ringtest_0.x4.clknet_1_0__leaf_clk.t40 VSS 0.014894f
C4697 ringtest_0.x4.clknet_1_0__leaf_clk.n38 VSS 0.040732f
C4698 ringtest_0.x4.clknet_1_0__leaf_clk.n39 VSS 0.086433f
C4699 ringtest_0.x4.clknet_1_0__leaf_clk.n40 VSS 0.225449f
C4700 ringtest_0.x4.clknet_1_0__leaf_clk.t35 VSS 0.022262f
C4701 ringtest_0.x4.clknet_1_0__leaf_clk.t34 VSS 0.014894f
C4702 ringtest_0.x4.clknet_1_0__leaf_clk.n41 VSS 0.04068f
C4703 ringtest_0.x4.clknet_1_0__leaf_clk.n42 VSS 0.027948f
C4704 ringtest_0.x4.clknet_1_0__leaf_clk.n43 VSS 0.145937f
C4705 ua[1].t0 VSS 0.322568f
C4706 ua[1].n0 VSS 0.401178f
C4707 ua[1].t5 VSS 0.24977f
C4708 ua[1].t1 VSS 0.33145f
C4709 ua[1].n1 VSS 1.6726f
C4710 ua[1].n2 VSS 0.565936f
C4711 ua[1].t6 VSS 0.244855f
C4712 ua[1].n3 VSS 0.365612f
C4713 ua[1].n4 VSS 0.509787f
C4714 ua[1].t4 VSS 0.322568f
C4715 ua[1].n5 VSS 0.401178f
C4716 ua[1].t8 VSS 0.24977f
C4717 ua[1].t12 VSS 0.33145f
C4718 ua[1].n6 VSS 1.6726f
C4719 ua[1].n7 VSS 0.565936f
C4720 ua[1].t9 VSS 0.244855f
C4721 ua[1].n8 VSS 0.365612f
C4722 ua[1].n9 VSS 0.495416f
C4723 ua[1].n10 VSS 0.270615f
C4724 ua[1].t13 VSS 0.322568f
C4725 ua[1].n11 VSS 0.401178f
C4726 ua[1].t11 VSS 0.24977f
C4727 ua[1].t7 VSS 0.33145f
C4728 ua[1].n12 VSS 1.6726f
C4729 ua[1].n13 VSS 0.565936f
C4730 ua[1].t10 VSS 0.244855f
C4731 ua[1].n14 VSS 0.365612f
C4732 ua[1].n15 VSS 0.495991f
C4733 ua[1].n16 VSS 0.268745f
C4734 ua[1].n17 VSS 0.801201f
C4735 ua[1].t3 VSS 0.322568f
C4736 ua[1].n18 VSS 0.401178f
C4737 ua[1].t15 VSS 0.24977f
C4738 ua[1].t2 VSS 0.33145f
C4739 ua[1].n19 VSS 1.6726f
C4740 ua[1].n20 VSS 0.565936f
C4741 ua[1].t14 VSS 0.244855f
C4742 ua[1].n21 VSS 0.365612f
C4743 ua[1].n22 VSS 0.500412f
C4744 ua[1].n23 VSS 0.264233f
C4745 ua[1].n24 VSS 0.382993f
C4746 ua[1].n25 VSS 7.827061f
C4747 ringtest_0.counter7.t5 VSS 0.031678f
C4748 ringtest_0.counter7.n0 VSS 0.005512f
C4749 ringtest_0.counter7.t4 VSS 0.021911f
C4750 ringtest_0.counter7.n1 VSS 0.026858f
C4751 ringtest_0.counter7.n2 VSS 0.039564f
C4752 ringtest_0.counter7.n3 VSS 0.38767f
C4753 ringtest_0.counter7.t0 VSS 0.693272f
C4754 ringtest_0.counter7.t1 VSS 0.490426f
C4755 ringtest_0.counter7.n4 VSS 3.80227f
C4756 ringtest_0.counter7.t2 VSS 0.385059f
C4757 ringtest_0.counter7.t3 VSS 0.706213f
C4758 ringtest_0.counter7.n5 VSS 3.95096f
C4759 ringtest_0.counter7.n6 VSS 0.629734f
C4760 ringtest_0.x3.x2.x4.GP VSS 2.5438f
C4761 ringtest_0.x3.x1.gpo3 VSS 1.19037f
C4762 ringtest_0.x3.x2.GP4.t1 VSS 0.012213f
C4763 ringtest_0.x3.x2.GP4.t0 VSS 0.012213f
C4764 ringtest_0.x3.x2.GP4.n0 VSS 0.026831f
C4765 ringtest_0.x3.x1.x14.Y VSS 0.075955f
C4766 ringtest_0.x3.x2.GP4.n1 VSS 0.010383f
C4767 ringtest_0.x3.x2.GP4.t4 VSS 0.618091f
C4768 ringtest_0.x3.x2.GP4.t5 VSS 0.635327f
C4769 ringtest_0.x3.x2.GP4.n2 VSS 2.25863f
C4770 ringtest_0.x3.x2.GP4.n3 VSS 0.047772f
C4771 ringtest_0.x3.x2.GP4.t3 VSS 0.01879f
C4772 ringtest_0.x3.x2.GP4.t2 VSS 0.01879f
C4773 ringtest_0.x3.x2.GP4.n4 VSS 0.043205f
C4774 ringtest_0.x3.x2.GP4.n5 VSS 0.087626f
C4775 ui_in[2].t7 VSS 0.320078f
C4776 ui_in[2].t1 VSS 0.312355f
C4777 ui_in[2].n0 VSS 1.40142f
C4778 ui_in[2].n1 VSS 0.46615f
C4779 ui_in[2].t6 VSS 0.375993f
C4780 ui_in[2].t0 VSS 0.386477f
C4781 ui_in[2].n2 VSS 1.40813f
C4782 ui_in[2].n3 VSS 0.945344f
C4783 ui_in[2].n4 VSS 2.4766f
C4784 ui_in[2].t3 VSS 0.01778f
C4785 ui_in[2].t5 VSS 0.010478f
C4786 ui_in[2].t2 VSS 0.01778f
C4787 ui_in[2].t4 VSS 0.010478f
C4788 ui_in[2].n5 VSS 0.029832f
C4789 ui_in[2].n6 VSS 0.044104f
C4790 ui_in[2].n7 VSS 0.043804f
C4791 ui_in[2].n8 VSS 0.708274f
C4792 ringtest_0.x4.net3.t1 VSS 0.067779f
C4793 ringtest_0.x4.net3.t2 VSS 0.019614f
C4794 ringtest_0.x4.net3.t7 VSS 0.031428f
C4795 ringtest_0.x4.net3.n0 VSS 0.061838f
C4796 ringtest_0.x4.net3.n1 VSS 0.008618f
C4797 ringtest_0.x4.net3.n2 VSS 0.005246f
C4798 ringtest_0.x4.net3.t6 VSS 0.029572f
C4799 ringtest_0.x4.net3.t5 VSS 0.018443f
C4800 ringtest_0.x4.net3.n3 VSS 0.059457f
C4801 ringtest_0.x4.net3.n4 VSS 0.019056f
C4802 ringtest_0.x4.net3.t4 VSS 0.030361f
C4803 ringtest_0.x4.net3.t3 VSS 0.055573f
C4804 ringtest_0.x4.net3.n5 VSS 0.744487f
C4805 ringtest_0.x4.net3.n6 VSS 0.124162f
C4806 ringtest_0.x4.net3.n7 VSS 0.092279f
C4807 ringtest_0.x4.net3.t0 VSS 0.037792f
C4808 ringtest_0.x4.net3.n8 VSS 0.040884f
C4809 ringtest_0.drv_out.t19 VSS 0.591341f
C4810 ringtest_0.drv_out.t0 VSS 0.418319f
C4811 ringtest_0.drv_out.n0 VSS 3.24323f
C4812 ringtest_0.drv_out.t2 VSS 0.328444f
C4813 ringtest_0.drv_out.t1 VSS 0.602379f
C4814 ringtest_0.drv_out.n1 VSS 3.37005f
C4815 ringtest_0.drv_out.n2 VSS 0.537145f
C4816 ringtest_0.drv_out.n3 VSS 0.110148f
C4817 ringtest_0.drv_out.t21 VSS 0.015262f
C4818 ringtest_0.drv_out.t25 VSS 0.007138f
C4819 ringtest_0.drv_out.t20 VSS 0.015262f
C4820 ringtest_0.drv_out.t24 VSS 0.007138f
C4821 ringtest_0.drv_out.t23 VSS 0.015262f
C4822 ringtest_0.drv_out.t27 VSS 0.007138f
C4823 ringtest_0.drv_out.t22 VSS 0.015262f
C4824 ringtest_0.drv_out.t26 VSS 0.007138f
C4825 ringtest_0.drv_out.n4 VSS 0.034841f
C4826 ringtest_0.drv_out.n5 VSS 0.04589f
C4827 ringtest_0.drv_out.n6 VSS 0.04589f
C4828 ringtest_0.drv_out.n7 VSS 0.055736f
C4829 ringtest_0.drv_out.n8 VSS 0.015444f
C4830 ringtest_0.drv_out.n9 VSS 0.346765f
C4831 ringtest_0.drv_out.n10 VSS 0.764086f
C4832 ringtest_0.drv_out.n11 VSS 5.53733f
C4833 ringtest_0.drv_out.t17 VSS 0.1149f
C4834 ringtest_0.drv_out.t12 VSS 0.1149f
C4835 ringtest_0.drv_out.n12 VSS 0.273611f
C4836 ringtest_0.drv_out.t14 VSS 0.1149f
C4837 ringtest_0.drv_out.t16 VSS 0.1149f
C4838 ringtest_0.drv_out.n13 VSS 0.273611f
C4839 ringtest_0.drv_out.t13 VSS 0.1149f
C4840 ringtest_0.drv_out.t15 VSS 0.1149f
C4841 ringtest_0.drv_out.n14 VSS 0.273611f
C4842 ringtest_0.drv_out.t18 VSS 0.1149f
C4843 ringtest_0.drv_out.t11 VSS 0.1149f
C4844 ringtest_0.drv_out.n15 VSS 0.273611f
C4845 ringtest_0.drv_out.n16 VSS 4.32f
C4846 ringtest_0.drv_out.t6 VSS 0.0383f
C4847 ringtest_0.drv_out.t8 VSS 0.0383f
C4848 ringtest_0.drv_out.n17 VSS 0.093269f
C4849 ringtest_0.drv_out.t7 VSS 0.0383f
C4850 ringtest_0.drv_out.t9 VSS 0.0383f
C4851 ringtest_0.drv_out.n18 VSS 0.093269f
C4852 ringtest_0.drv_out.t3 VSS 0.0383f
C4853 ringtest_0.drv_out.t4 VSS 0.0383f
C4854 ringtest_0.drv_out.n19 VSS 0.093269f
C4855 ringtest_0.drv_out.t10 VSS 0.0383f
C4856 ringtest_0.drv_out.t5 VSS 0.0383f
C4857 ringtest_0.drv_out.n20 VSS 0.093269f
C4858 ringtest_0.drv_out.n21 VSS 1.9949f
C4859 ringtest_0.drv_out.n22 VSS 2.14485f
C4860 a_19289_13081.t12 VSS 0.136375f
C4861 a_19289_13081.t2 VSS 0.13635f
C4862 a_19289_13081.n0 VSS 0.157675f
C4863 a_19289_13081.t13 VSS 0.13635f
C4864 a_19289_13081.n1 VSS 0.086028f
C4865 a_19289_13081.t7 VSS 0.13635f
C4866 a_19289_13081.n2 VSS 0.160734f
C4867 a_19289_13081.t4 VSS 0.049796f
C4868 a_19289_13081.t15 VSS 0.049764f
C4869 a_19289_13081.n3 VSS 0.09498f
C4870 a_19289_13081.t5 VSS 0.049764f
C4871 a_19289_13081.n4 VSS 0.055718f
C4872 a_19289_13081.t11 VSS 0.049764f
C4873 a_19289_13081.n5 VSS 0.086134f
C4874 a_19289_13081.t0 VSS 0.098833f
C4875 a_19289_13081.n6 VSS 0.831842f
C4876 a_19289_13081.t6 VSS 0.049771f
C4877 a_19289_13081.t9 VSS 0.13635f
C4878 a_19289_13081.n7 VSS 0.503671f
C4879 a_19289_13081.t16 VSS 0.049764f
C4880 a_19289_13081.n8 VSS 0.212248f
C4881 a_19289_13081.t17 VSS 0.13635f
C4882 a_19289_13081.n9 VSS 0.242932f
C4883 a_19289_13081.t8 VSS 0.049764f
C4884 a_19289_13081.n10 VSS 0.212248f
C4885 a_19289_13081.t10 VSS 0.13635f
C4886 a_19289_13081.n11 VSS 0.242932f
C4887 a_19289_13081.t3 VSS 0.049764f
C4888 a_19289_13081.n12 VSS 0.212248f
C4889 a_19289_13081.t14 VSS 0.13635f
C4890 a_19289_13081.n13 VSS 0.494157f
C4891 a_19289_13081.n14 VSS 1.47337f
C4892 a_19289_13081.n15 VSS 2.33573f
C4893 a_19289_13081.t1 VSS 0.309542f
C4894 muxtest_0.R1R2.t1 VSS 0.625209f
C4895 muxtest_0.R1R2.t0 VSS 0.442278f
C4896 muxtest_0.R1R2.n0 VSS 3.42898f
C4897 muxtest_0.R1R2.t4 VSS 0.347255f
C4898 muxtest_0.R1R2.t5 VSS 0.63688f
C4899 muxtest_0.R1R2.n1 VSS 3.56307f
C4900 muxtest_0.R1R2.n2 VSS 0.56791f
C4901 muxtest_0.R1R2.n3 VSS 0.116899f
C4902 muxtest_0.R1R2.t3 VSS 0.207548f
C4903 muxtest_0.R1R2.t2 VSS 0.169702f
C4904 muxtest_0.R1R2.n4 VSS 3.13805f
C4905 muxtest_0.R1R2.n5 VSS 1.09366f
C4906 ui_in[4].t4 VSS 0.008207f
C4907 ui_in[4].t10 VSS 0.004836f
C4908 ui_in[4].t6 VSS 0.008207f
C4909 ui_in[4].t16 VSS 0.004836f
C4910 ui_in[4].n0 VSS 0.01377f
C4911 ui_in[4].n1 VSS 0.020344f
C4912 ui_in[4].n2 VSS 0.012412f
C4913 ui_in[4].t19 VSS 0.008009f
C4914 ui_in[4].t13 VSS 0.003797f
C4915 ui_in[4].n3 VSS 0.028758f
C4916 ui_in[4].n4 VSS 0.005576f
C4917 ui_in[4].n5 VSS 0.00476f
C4918 ui_in[4].t7 VSS 0.003976f
C4919 ui_in[4].t12 VSS 0.005786f
C4920 ui_in[4].n6 VSS 0.016813f
C4921 ui_in[4].n7 VSS 0.003873f
C4922 ui_in[4].n8 VSS 0.027736f
C4923 ui_in[4].n9 VSS 0.100485f
C4924 ui_in[4].t5 VSS 0.004786f
C4925 ui_in[4].t0 VSS 0.007049f
C4926 ui_in[4].n10 VSS 0.016654f
C4927 ui_in[4].n11 VSS 0.002169f
C4928 ui_in[4].n12 VSS 0.024508f
C4929 ui_in[4].n13 VSS 0.115979f
C4930 ui_in[4].n14 VSS 0.151491f
C4931 ui_in[4].n15 VSS 0.034981f
C4932 ui_in[4].t15 VSS 0.008207f
C4933 ui_in[4].t2 VSS 0.004836f
C4934 ui_in[4].t9 VSS 0.008207f
C4935 ui_in[4].t18 VSS 0.004836f
C4936 ui_in[4].n16 VSS 0.01377f
C4937 ui_in[4].n17 VSS 0.020344f
C4938 ui_in[4].n18 VSS 0.012412f
C4939 ui_in[4].t1 VSS 0.008009f
C4940 ui_in[4].t17 VSS 0.003797f
C4941 ui_in[4].n19 VSS 0.028758f
C4942 ui_in[4].n20 VSS 0.005576f
C4943 ui_in[4].n21 VSS 0.00476f
C4944 ui_in[4].t11 VSS 0.003976f
C4945 ui_in[4].t14 VSS 0.005786f
C4946 ui_in[4].n22 VSS 0.016813f
C4947 ui_in[4].n23 VSS 0.003873f
C4948 ui_in[4].n24 VSS 0.027736f
C4949 ui_in[4].n25 VSS 0.100485f
C4950 ui_in[4].t8 VSS 0.004786f
C4951 ui_in[4].t3 VSS 0.007049f
C4952 ui_in[4].n26 VSS 0.016654f
C4953 ui_in[4].n27 VSS 0.002169f
C4954 ui_in[4].n28 VSS 0.024508f
C4955 ui_in[4].n29 VSS 0.115979f
C4956 ui_in[4].n30 VSS 0.151491f
C4957 ui_in[4].n31 VSS 12.0273f
C4958 muxtest_0.R3R4.t6 VSS 0.65338f
C4959 muxtest_0.R3R4.t5 VSS 0.462206f
C4960 muxtest_0.R3R4.n0 VSS 3.58348f
C4961 muxtest_0.R3R4.t1 VSS 0.362902f
C4962 muxtest_0.R3R4.t0 VSS 0.665576f
C4963 muxtest_0.R3R4.n1 VSS 3.72361f
C4964 muxtest_0.R3R4.n2 VSS 0.593498f
C4965 muxtest_0.R3R4.n3 VSS 0.123258f
C4966 muxtest_0.R3R4.t4 VSS 1.02738f
C4967 muxtest_0.R3R4.t7 VSS 0.177328f
C4968 muxtest_0.R3R4.n4 VSS 2.29699f
C4969 muxtest_0.R3R4.t3 VSS 0.65338f
C4970 muxtest_0.R3R4.t2 VSS 0.462206f
C4971 muxtest_0.R3R4.n5 VSS 3.58348f
C4972 muxtest_0.R3R4.t8 VSS 0.362902f
C4973 muxtest_0.R3R4.t9 VSS 0.665576f
C4974 muxtest_0.R3R4.n6 VSS 3.72361f
C4975 muxtest_0.R3R4.n7 VSS 0.593498f
C4976 muxtest_0.R3R4.n8 VSS 0.122166f
C4977 muxtest_0.R3R4.n9 VSS 0.05979f
C4978 muxtest_0.R3R4.n10 VSS 6.98972f
C4979 muxtest_0.R3R4.n11 VSS 7.31123f
C4980 muxtest_0.R3R4.n12 VSS 1.03011f
C4981 ui_in[0].t6 VSS 0.006125f
C4982 ui_in[0].t0 VSS 0.003609f
C4983 ui_in[0].t8 VSS 0.006125f
C4984 ui_in[0].t3 VSS 0.003609f
C4985 ui_in[0].n0 VSS 0.010276f
C4986 ui_in[0].n1 VSS 0.015187f
C4987 ui_in[0].n2 VSS 0.004773f
C4988 ui_in[0].t9 VSS 0.003016f
C4989 ui_in[0].t5 VSS 0.004381f
C4990 ui_in[0].n3 VSS 0.010436f
C4991 ui_in[0].n4 VSS 0.005796f
C4992 ui_in[0].t1 VSS 0.003572f
C4993 ui_in[0].t7 VSS 0.00526f
C4994 ui_in[0].n5 VSS 0.012428f
C4995 ui_in[0].n6 VSS 0.002581f
C4996 ui_in[0].n7 VSS 0.001006f
C4997 ui_in[0].n8 VSS 0.091917f
C4998 ui_in[0].t4 VSS 0.005977f
C4999 ui_in[0].t2 VSS 0.002834f
C5000 ui_in[0].n9 VSS 0.021461f
C5001 ui_in[0].n10 VSS 0.004159f
C5002 ui_in[0].n11 VSS 0.105454f
C5003 ui_in[0].n12 VSS 0.068524f
C5004 ui_in[0].n13 VSS 2.54475f
C5005 ringtest_0.x4._11_.t3 VSS 0.02558f
C5006 ringtest_0.x4._11_.t2 VSS 0.02558f
C5007 ringtest_0.x4._11_.n0 VSS 0.053419f
C5008 ringtest_0.x4._11_.t12 VSS 0.042601f
C5009 ringtest_0.x4._11_.t9 VSS 0.026392f
C5010 ringtest_0.x4._11_.n1 VSS 0.086305f
C5011 ringtest_0.x4._11_.n2 VSS 0.024278f
C5012 ringtest_0.x4._11_.t7 VSS 0.027069f
C5013 ringtest_0.x4._11_.t13 VSS 0.043108f
C5014 ringtest_0.x4._11_.n3 VSS 0.058737f
C5015 ringtest_0.x4._11_.n4 VSS 0.032841f
C5016 ringtest_0.x4._11_.t17 VSS 0.023619f
C5017 ringtest_0.x4._11_.t5 VSS 0.034667f
C5018 ringtest_0.x4._11_.n5 VSS 0.06984f
C5019 ringtest_0.x4._11_.n6 VSS 0.034707f
C5020 ringtest_0.x4._11_.n7 VSS 0.494881f
C5021 ringtest_0.x4._11_.t21 VSS 0.027069f
C5022 ringtest_0.x4._11_.t10 VSS 0.043108f
C5023 ringtest_0.x4._11_.n8 VSS 0.058739f
C5024 ringtest_0.x4._11_.n9 VSS 0.133927f
C5025 ringtest_0.x4._11_.n10 VSS 0.765831f
C5026 ringtest_0.x4._11_.t11 VSS 0.021102f
C5027 ringtest_0.x4._11_.t18 VSS 0.017461f
C5028 ringtest_0.x4._11_.n11 VSS 0.092223f
C5029 ringtest_0.x4._11_.n12 VSS 0.043963f
C5030 ringtest_0.x4._11_.n13 VSS 0.150035f
C5031 ringtest_0.x4._11_.t14 VSS 0.028052f
C5032 ringtest_0.x4._11_.t4 VSS 0.019277f
C5033 ringtest_0.x4._11_.n14 VSS 0.081517f
C5034 ringtest_0.x4._11_.n15 VSS 0.011369f
C5035 ringtest_0.x4._11_.n16 VSS 0.03744f
C5036 ringtest_0.x4._11_.n17 VSS 0.156255f
C5037 ringtest_0.x4._11_.t15 VSS 0.019598f
C5038 ringtest_0.x4._11_.t19 VSS 0.028465f
C5039 ringtest_0.x4._11_.n18 VSS 0.067767f
C5040 ringtest_0.x4._11_.n19 VSS 0.143997f
C5041 ringtest_0.x4._11_.n20 VSS 0.492685f
C5042 ringtest_0.x4._11_.t8 VSS 0.042359f
C5043 ringtest_0.x4._11_.t16 VSS 0.026451f
C5044 ringtest_0.x4._11_.n21 VSS 0.080165f
C5045 ringtest_0.x4._11_.n22 VSS 0.023455f
C5046 ringtest_0.x4._11_.n23 VSS 0.356691f
C5047 ringtest_0.x4._11_.t20 VSS 0.023619f
C5048 ringtest_0.x4._11_.t6 VSS 0.034667f
C5049 ringtest_0.x4._11_.n24 VSS 0.06984f
C5050 ringtest_0.x4._11_.n25 VSS 0.014495f
C5051 ringtest_0.x4._11_.n26 VSS 0.490885f
C5052 ringtest_0.x4._11_.n27 VSS 1.19049f
C5053 ringtest_0.x4._11_.n28 VSS 0.353781f
C5054 ringtest_0.x4._11_.n29 VSS 0.021904f
C5055 ringtest_0.x4._11_.t0 VSS 0.010743f
C5056 ringtest_0.x4._11_.t1 VSS 0.010743f
C5057 ringtest_0.x4._11_.n30 VSS 0.02648f
C5058 muxtest_0.x1.x3.x4.GP VSS 2.932f
C5059 muxtest_0.x1.x2.x4.GP VSS 2.29581f
C5060 muxtest_0.x1.x1.gpo3 VSS 1.43031f
C5061 muxtest_0.x1.x3.GP4.t1 VSS 0.01297f
C5062 muxtest_0.x1.x3.GP4.t0 VSS 0.01297f
C5063 muxtest_0.x1.x3.GP4.n0 VSS 0.028494f
C5064 muxtest_0.x1.x1.x14.Y VSS 0.080663f
C5065 muxtest_0.x1.x3.GP4.n1 VSS 0.011026f
C5066 muxtest_0.x1.x3.GP4.t6 VSS 0.656398f
C5067 muxtest_0.x1.x3.GP4.t7 VSS 0.674702f
C5068 muxtest_0.x1.x3.GP4.n2 VSS 2.39862f
C5069 muxtest_0.x1.x3.GP4.t4 VSS 0.656398f
C5070 muxtest_0.x1.x3.GP4.t5 VSS 0.674702f
C5071 muxtest_0.x1.x3.GP4.n3 VSS 2.39862f
C5072 muxtest_0.x1.x3.GP4.n4 VSS 2.8073f
C5073 muxtest_0.x1.x3.GP4.n5 VSS 0.050183f
C5074 muxtest_0.x1.x3.GP4.t2 VSS 0.019954f
C5075 muxtest_0.x1.x3.GP4.t3 VSS 0.019954f
C5076 muxtest_0.x1.x3.GP4.n6 VSS 0.045883f
C5077 muxtest_0.x1.x3.GP4.n7 VSS 0.093057f
C5078 muxtest_0.x1.x3.GP1.t1 VSS 0.018021f
C5079 muxtest_0.x1.x3.GP1.t0 VSS 0.018021f
C5080 muxtest_0.x1.x3.GP1.n0 VSS 0.039591f
C5081 muxtest_0.x1.x3.GP1.n1 VSS 0.02559f
C5082 muxtest_0.x1.x3.GP1.t7 VSS 0.912037f
C5083 muxtest_0.x1.x3.GP1.t6 VSS 0.937471f
C5084 muxtest_0.x1.x3.GP1.n2 VSS 3.31176f
C5085 muxtest_0.x1.x3.GP1.t5 VSS 0.912037f
C5086 muxtest_0.x1.x3.GP1.t4 VSS 0.937471f
C5087 muxtest_0.x1.x3.GP1.n3 VSS 3.31176f
C5088 muxtest_0.x1.x3.GP1.n4 VSS 1.73806f
C5089 muxtest_0.x1.x3.GP1.t2 VSS 0.027725f
C5090 muxtest_0.x1.x3.GP1.t3 VSS 0.027725f
C5091 muxtest_0.x1.x3.GP1.n5 VSS 0.057129f
C5092 muxtest_0.x1.x3.GP1.n6 VSS 0.132634f
C5093 muxtest_0.x1.x3.GP1.n7 VSS 0.030542f
C5094 ui_in[1].t2 VSS 0.013664f
C5095 ui_in[1].t6 VSS 0.008052f
C5096 ui_in[1].t0 VSS 0.013664f
C5097 ui_in[1].t5 VSS 0.008052f
C5098 ui_in[1].n0 VSS 0.022926f
C5099 ui_in[1].n1 VSS 0.033873f
C5100 ui_in[1].n2 VSS 0.020666f
C5101 ui_in[1].t1 VSS 0.013334f
C5102 ui_in[1].t4 VSS 0.006323f
C5103 ui_in[1].n3 VSS 0.047881f
C5104 ui_in[1].n4 VSS 0.009284f
C5105 ui_in[1].n5 VSS 0.007925f
C5106 ui_in[1].t3 VSS 0.00662f
C5107 ui_in[1].t7 VSS 0.009633f
C5108 ui_in[1].n6 VSS 0.027992f
C5109 ui_in[1].n7 VSS 0.006448f
C5110 ui_in[1].n8 VSS 0.04618f
C5111 ui_in[1].n9 VSS 0.167305f
C5112 ui_in[1].t9 VSS 0.007969f
C5113 ui_in[1].t8 VSS 0.011736f
C5114 ui_in[1].n10 VSS 0.027728f
C5115 ui_in[1].n11 VSS 0.003611f
C5116 ui_in[1].n12 VSS 0.040805f
C5117 ui_in[1].n13 VSS 0.193102f
C5118 ui_in[1].n14 VSS 0.252228f
C5119 ui_in[1].n15 VSS 0.051098f
C5120 ui_in[1].n16 VSS 5.24829f
C5121 ringtest_0.x4.clknet_1_1__leaf_clk.t13 VSS 0.005541f
C5122 ringtest_0.x4.clknet_1_1__leaf_clk.t14 VSS 0.005541f
C5123 ringtest_0.x4.clknet_1_1__leaf_clk.n0 VSS 0.019676f
C5124 ringtest_0.x4.clknet_1_1__leaf_clk.t15 VSS 0.005541f
C5125 ringtest_0.x4.clknet_1_1__leaf_clk.t12 VSS 0.005541f
C5126 ringtest_0.x4.clknet_1_1__leaf_clk.n1 VSS 0.01265f
C5127 ringtest_0.x4.clknet_1_1__leaf_clk.n2 VSS 0.07993f
C5128 ringtest_0.x4.clknet_1_1__leaf_clk.t11 VSS 0.005541f
C5129 ringtest_0.x4.clknet_1_1__leaf_clk.t10 VSS 0.005541f
C5130 ringtest_0.x4.clknet_1_1__leaf_clk.n3 VSS 0.01265f
C5131 ringtest_0.x4.clknet_1_1__leaf_clk.n4 VSS 0.048044f
C5132 ringtest_0.x4.clknet_1_1__leaf_clk.t6 VSS 0.005541f
C5133 ringtest_0.x4.clknet_1_1__leaf_clk.t8 VSS 0.005541f
C5134 ringtest_0.x4.clknet_1_1__leaf_clk.n5 VSS 0.012657f
C5135 ringtest_0.x4.clknet_1_1__leaf_clk.n6 VSS 0.049559f
C5136 ringtest_0.x4.clknet_1_1__leaf_clk.t2 VSS 0.005541f
C5137 ringtest_0.x4.clknet_1_1__leaf_clk.t4 VSS 0.005541f
C5138 ringtest_0.x4.clknet_1_1__leaf_clk.n7 VSS 0.01265f
C5139 ringtest_0.x4.clknet_1_1__leaf_clk.n8 VSS 0.048044f
C5140 ringtest_0.x4.clknet_1_1__leaf_clk.t5 VSS 0.005541f
C5141 ringtest_0.x4.clknet_1_1__leaf_clk.t7 VSS 0.005541f
C5142 ringtest_0.x4.clknet_1_1__leaf_clk.n9 VSS 0.011247f
C5143 ringtest_0.x4.clknet_1_1__leaf_clk.t37 VSS 0.013817f
C5144 ringtest_0.x4.clknet_1_1__leaf_clk.t32 VSS 0.020651f
C5145 ringtest_0.x4.clknet_1_1__leaf_clk.n10 VSS 0.038168f
C5146 ringtest_0.x4.clknet_1_1__leaf_clk.t41 VSS 0.020651f
C5147 ringtest_0.x4.clknet_1_1__leaf_clk.t35 VSS 0.013817f
C5148 ringtest_0.x4.clknet_1_1__leaf_clk.n11 VSS 0.037785f
C5149 ringtest_0.x4.clknet_1_1__leaf_clk.n12 VSS 0.039947f
C5150 ringtest_0.x4.clknet_1_1__leaf_clk.t38 VSS 0.013817f
C5151 ringtest_0.x4.clknet_1_1__leaf_clk.t34 VSS 0.020651f
C5152 ringtest_0.x4.clknet_1_1__leaf_clk.n13 VSS 0.038168f
C5153 ringtest_0.x4.clknet_1_1__leaf_clk.n14 VSS 0.30833f
C5154 ringtest_0.x4.clknet_1_1__leaf_clk.t33 VSS 0.020651f
C5155 ringtest_0.x4.clknet_1_1__leaf_clk.t40 VSS 0.013817f
C5156 ringtest_0.x4.clknet_1_1__leaf_clk.n15 VSS 0.037785f
C5157 ringtest_0.x4.clknet_1_1__leaf_clk.n16 VSS 0.030886f
C5158 ringtest_0.x4.clknet_1_1__leaf_clk.n17 VSS 0.118422f
C5159 ringtest_0.x4.clknet_1_1__leaf_clk.t39 VSS 0.013817f
C5160 ringtest_0.x4.clknet_1_1__leaf_clk.t36 VSS 0.020651f
C5161 ringtest_0.x4.clknet_1_1__leaf_clk.n18 VSS 0.037832f
C5162 ringtest_0.x4.clknet_1_1__leaf_clk.n19 VSS 0.022005f
C5163 ringtest_0.x4.clknet_1_1__leaf_clk.n20 VSS 0.128874f
C5164 ringtest_0.x4.clknet_1_1__leaf_clk.n21 VSS 0.280206f
C5165 ringtest_0.x4.clknet_1_1__leaf_clk.n22 VSS 0.023331f
C5166 ringtest_0.x4.clknet_1_1__leaf_clk.n23 VSS 0.030986f
C5167 ringtest_0.x4.clknet_1_1__leaf_clk.t1 VSS 0.005541f
C5168 ringtest_0.x4.clknet_1_1__leaf_clk.t9 VSS 0.005541f
C5169 ringtest_0.x4.clknet_1_1__leaf_clk.n24 VSS 0.01265f
C5170 ringtest_0.x4.clknet_1_1__leaf_clk.n25 VSS 0.041476f
C5171 ringtest_0.x4.clknet_1_1__leaf_clk.t25 VSS 0.013193f
C5172 ringtest_0.x4.clknet_1_1__leaf_clk.t22 VSS 0.013193f
C5173 ringtest_0.x4.clknet_1_1__leaf_clk.n26 VSS 0.027449f
C5174 ringtest_0.x4.clknet_1_1__leaf_clk.t19 VSS 0.013193f
C5175 ringtest_0.x4.clknet_1_1__leaf_clk.t20 VSS 0.013193f
C5176 ringtest_0.x4.clknet_1_1__leaf_clk.n27 VSS 0.033515f
C5177 ringtest_0.x4.clknet_1_1__leaf_clk.t21 VSS 0.013193f
C5178 ringtest_0.x4.clknet_1_1__leaf_clk.t18 VSS 0.013193f
C5179 ringtest_0.x4.clknet_1_1__leaf_clk.n28 VSS 0.02781f
C5180 ringtest_0.x4.clknet_1_1__leaf_clk.n29 VSS 0.126738f
C5181 ringtest_0.x4.clknet_1_1__leaf_clk.t17 VSS 0.013193f
C5182 ringtest_0.x4.clknet_1_1__leaf_clk.t16 VSS 0.013193f
C5183 ringtest_0.x4.clknet_1_1__leaf_clk.n30 VSS 0.02781f
C5184 ringtest_0.x4.clknet_1_1__leaf_clk.n31 VSS 0.073006f
C5185 ringtest_0.x4.clknet_1_1__leaf_clk.t28 VSS 0.013193f
C5186 ringtest_0.x4.clknet_1_1__leaf_clk.t30 VSS 0.013193f
C5187 ringtest_0.x4.clknet_1_1__leaf_clk.n32 VSS 0.02781f
C5188 ringtest_0.x4.clknet_1_1__leaf_clk.n33 VSS 0.072667f
C5189 ringtest_0.x4.clknet_1_1__leaf_clk.t24 VSS 0.013193f
C5190 ringtest_0.x4.clknet_1_1__leaf_clk.t26 VSS 0.013193f
C5191 ringtest_0.x4.clknet_1_1__leaf_clk.n34 VSS 0.02781f
C5192 ringtest_0.x4.clknet_1_1__leaf_clk.n35 VSS 0.072667f
C5193 ringtest_0.x4.clknet_1_1__leaf_clk.t27 VSS 0.013193f
C5194 ringtest_0.x4.clknet_1_1__leaf_clk.t29 VSS 0.013193f
C5195 ringtest_0.x4.clknet_1_1__leaf_clk.n36 VSS 0.02781f
C5196 ringtest_0.x4.clknet_1_1__leaf_clk.n37 VSS 0.073006f
C5197 ringtest_0.x4.clknet_1_1__leaf_clk.t23 VSS 0.013193f
C5198 ringtest_0.x4.clknet_1_1__leaf_clk.t31 VSS 0.013193f
C5199 ringtest_0.x4.clknet_1_1__leaf_clk.n38 VSS 0.02781f
C5200 ringtest_0.x4.clknet_1_1__leaf_clk.n39 VSS 0.062704f
C5201 ringtest_0.x4.clknet_1_1__leaf_clk.n40 VSS 0.086346f
C5202 ringtest_0.x4.clknet_1_1__leaf_clk.n41 VSS 0.040127f
C5203 ringtest_0.x4.clknet_1_1__leaf_clk.t3 VSS 0.005541f
C5204 ringtest_0.x4.clknet_1_1__leaf_clk.t0 VSS 0.005541f
C5205 ringtest_0.x4.clknet_1_1__leaf_clk.n42 VSS 0.012211f
C5206 ringtest_0.x4.net6.t8 VSS 0.023291f
C5207 ringtest_0.x4.net6.t4 VSS 0.034395f
C5208 ringtest_0.x4.net6.n0 VSS 0.095831f
C5209 ringtest_0.x4.net6.t2 VSS 0.040459f
C5210 ringtest_0.x4.net6.t12 VSS 0.025233f
C5211 ringtest_0.x4.net6.n1 VSS 0.081347f
C5212 ringtest_0.x4.net6.n2 VSS 0.124436f
C5213 ringtest_0.x4.net6.t6 VSS 0.023291f
C5214 ringtest_0.x4.net6.t13 VSS 0.034395f
C5215 ringtest_0.x4.net6.n3 VSS 0.095831f
C5216 ringtest_0.x4.net6.n4 VSS 0.41789f
C5217 ringtest_0.x4.net6.t10 VSS 0.021456f
C5218 ringtest_0.x4.net6.t3 VSS 0.017754f
C5219 ringtest_0.x4.net6.n5 VSS 0.093771f
C5220 ringtest_0.x4.net6.n6 VSS 0.080526f
C5221 ringtest_0.x4.net6.n7 VSS 0.286209f
C5222 ringtest_0.x4.net6.t11 VSS 0.027524f
C5223 ringtest_0.x4.net6.t5 VSS 0.043832f
C5224 ringtest_0.x4.net6.n8 VSS 0.059723f
C5225 ringtest_0.x4.net6.n9 VSS 0.146037f
C5226 ringtest_0.x4.net6.n10 VSS 0.772479f
C5227 ringtest_0.x4.net6.n11 VSS 0.732404f
C5228 ringtest_0.x4.net6.t9 VSS 0.023842f
C5229 ringtest_0.x4.net6.t14 VSS 0.040459f
C5230 ringtest_0.x4.net6.n12 VSS 0.051672f
C5231 ringtest_0.x4.net6.t15 VSS 0.023842f
C5232 ringtest_0.x4.net6.t7 VSS 0.040459f
C5233 ringtest_0.x4.net6.n13 VSS 0.057394f
C5234 ringtest_0.x4.net6.n14 VSS 0.027196f
C5235 ringtest_0.x4.net6.n15 VSS 0.1061f
C5236 ringtest_0.x4.net6.n16 VSS 0.491563f
C5237 ringtest_0.x4.net6.t1 VSS 0.092732f
C5238 ringtest_0.x4.net6.n17 VSS 0.127274f
C5239 ringtest_0.x4.net6.t0 VSS 0.050895f
C5240 ringtest_0.x4.net6.n18 VSS 0.064268f
C5241 ringtest_0.x4.clknet_0_clk.t2 VSS 0.004717f
C5242 ringtest_0.x4.clknet_0_clk.t15 VSS 0.004717f
C5243 ringtest_0.x4.clknet_0_clk.n0 VSS 0.016749f
C5244 ringtest_0.x4.clknet_0_clk.t4 VSS 0.004717f
C5245 ringtest_0.x4.clknet_0_clk.t6 VSS 0.004717f
C5246 ringtest_0.x4.clknet_0_clk.n1 VSS 0.010767f
C5247 ringtest_0.x4.clknet_0_clk.n2 VSS 0.068037f
C5248 ringtest_0.x4.clknet_0_clk.t8 VSS 0.004717f
C5249 ringtest_0.x4.clknet_0_clk.t10 VSS 0.004717f
C5250 ringtest_0.x4.clknet_0_clk.n3 VSS 0.010767f
C5251 ringtest_0.x4.clknet_0_clk.n4 VSS 0.040895f
C5252 ringtest_0.x4.clknet_0_clk.t5 VSS 0.004717f
C5253 ringtest_0.x4.clknet_0_clk.t7 VSS 0.004717f
C5254 ringtest_0.x4.clknet_0_clk.n5 VSS 0.010774f
C5255 ringtest_0.x4.clknet_0_clk.n6 VSS 0.042184f
C5256 ringtest_0.x4.clknet_0_clk.t9 VSS 0.004717f
C5257 ringtest_0.x4.clknet_0_clk.t11 VSS 0.004717f
C5258 ringtest_0.x4.clknet_0_clk.n7 VSS 0.010767f
C5259 ringtest_0.x4.clknet_0_clk.n8 VSS 0.040895f
C5260 ringtest_0.x4.clknet_0_clk.t0 VSS 0.004717f
C5261 ringtest_0.x4.clknet_0_clk.t13 VSS 0.004717f
C5262 ringtest_0.x4.clknet_0_clk.n9 VSS 0.009573f
C5263 ringtest_0.x4.clknet_0_clk.t39 VSS 0.015823f
C5264 ringtest_0.x4.clknet_0_clk.t47 VSS 0.0074f
C5265 ringtest_0.x4.clknet_0_clk.t40 VSS 0.015823f
C5266 ringtest_0.x4.clknet_0_clk.t32 VSS 0.0074f
C5267 ringtest_0.x4.clknet_0_clk.t37 VSS 0.015823f
C5268 ringtest_0.x4.clknet_0_clk.t44 VSS 0.0074f
C5269 ringtest_0.x4.clknet_0_clk.t41 VSS 0.015823f
C5270 ringtest_0.x4.clknet_0_clk.t33 VSS 0.0074f
C5271 ringtest_0.x4.clknet_0_clk.n10 VSS 0.036121f
C5272 ringtest_0.x4.clknet_0_clk.n11 VSS 0.047576f
C5273 ringtest_0.x4.clknet_0_clk.n12 VSS 0.047576f
C5274 ringtest_0.x4.clknet_0_clk.n13 VSS 0.057784f
C5275 ringtest_0.x4.clknet_0_clk.n14 VSS 0.075138f
C5276 ringtest_0.x4.clknet_0_clk.t46 VSS 0.015823f
C5277 ringtest_0.x4.clknet_0_clk.t38 VSS 0.0074f
C5278 ringtest_0.x4.clknet_0_clk.t43 VSS 0.015823f
C5279 ringtest_0.x4.clknet_0_clk.t35 VSS 0.0074f
C5280 ringtest_0.x4.clknet_0_clk.t42 VSS 0.015823f
C5281 ringtest_0.x4.clknet_0_clk.t34 VSS 0.0074f
C5282 ringtest_0.x4.clknet_0_clk.t45 VSS 0.015823f
C5283 ringtest_0.x4.clknet_0_clk.t36 VSS 0.0074f
C5284 ringtest_0.x4.clknet_0_clk.n15 VSS 0.036121f
C5285 ringtest_0.x4.clknet_0_clk.n16 VSS 0.047576f
C5286 ringtest_0.x4.clknet_0_clk.n17 VSS 0.047576f
C5287 ringtest_0.x4.clknet_0_clk.n18 VSS 0.057941f
C5288 ringtest_0.x4.clknet_0_clk.n19 VSS 0.038186f
C5289 ringtest_0.x4.clknet_0_clk.n20 VSS 0.145873f
C5290 ringtest_0.x4.clknet_0_clk.n21 VSS 0.015919f
C5291 ringtest_0.x4.clknet_0_clk.n22 VSS 0.026375f
C5292 ringtest_0.x4.clknet_0_clk.t14 VSS 0.004717f
C5293 ringtest_0.x4.clknet_0_clk.t12 VSS 0.004717f
C5294 ringtest_0.x4.clknet_0_clk.n23 VSS 0.010767f
C5295 ringtest_0.x4.clknet_0_clk.n24 VSS 0.035304f
C5296 ringtest_0.x4.clknet_0_clk.t26 VSS 0.01123f
C5297 ringtest_0.x4.clknet_0_clk.t28 VSS 0.01123f
C5298 ringtest_0.x4.clknet_0_clk.n25 VSS 0.023364f
C5299 ringtest_0.x4.clknet_0_clk.t23 VSS 0.01123f
C5300 ringtest_0.x4.clknet_0_clk.t21 VSS 0.01123f
C5301 ringtest_0.x4.clknet_0_clk.n26 VSS 0.023672f
C5302 ringtest_0.x4.clknet_0_clk.t25 VSS 0.01123f
C5303 ringtest_0.x4.clknet_0_clk.t22 VSS 0.01123f
C5304 ringtest_0.x4.clknet_0_clk.n27 VSS 0.023672f
C5305 ringtest_0.x4.clknet_0_clk.t18 VSS 0.01123f
C5306 ringtest_0.x4.clknet_0_clk.t20 VSS 0.01123f
C5307 ringtest_0.x4.clknet_0_clk.n28 VSS 0.023672f
C5308 ringtest_0.x4.clknet_0_clk.t30 VSS 0.01123f
C5309 ringtest_0.x4.clknet_0_clk.t16 VSS 0.01123f
C5310 ringtest_0.x4.clknet_0_clk.n29 VSS 0.023672f
C5311 ringtest_0.x4.clknet_0_clk.t17 VSS 0.01123f
C5312 ringtest_0.x4.clknet_0_clk.t19 VSS 0.01123f
C5313 ringtest_0.x4.clknet_0_clk.n30 VSS 0.023672f
C5314 ringtest_0.x4.clknet_0_clk.t27 VSS 0.01123f
C5315 ringtest_0.x4.clknet_0_clk.t24 VSS 0.01123f
C5316 ringtest_0.x4.clknet_0_clk.n31 VSS 0.028528f
C5317 ringtest_0.x4.clknet_0_clk.t29 VSS 0.01123f
C5318 ringtest_0.x4.clknet_0_clk.t31 VSS 0.01123f
C5319 ringtest_0.x4.clknet_0_clk.n32 VSS 0.023672f
C5320 ringtest_0.x4.clknet_0_clk.n33 VSS 0.107879f
C5321 ringtest_0.x4.clknet_0_clk.n34 VSS 0.062143f
C5322 ringtest_0.x4.clknet_0_clk.n35 VSS 0.061854f
C5323 ringtest_0.x4.clknet_0_clk.n36 VSS 0.061854f
C5324 ringtest_0.x4.clknet_0_clk.n37 VSS 0.062143f
C5325 ringtest_0.x4.clknet_0_clk.n38 VSS 0.053374f
C5326 ringtest_0.x4.clknet_0_clk.n39 VSS 0.073498f
C5327 ringtest_0.x4.clknet_0_clk.n40 VSS 0.034156f
C5328 ringtest_0.x4.clknet_0_clk.t1 VSS 0.004717f
C5329 ringtest_0.x4.clknet_0_clk.t3 VSS 0.004717f
C5330 ringtest_0.x4.clknet_0_clk.n41 VSS 0.010394f
C5331 ua[2].t8 VSS 0.247385f
C5332 ua[2].n0 VSS 0.307673f
C5333 ua[2].t12 VSS 0.191554f
C5334 ua[2].t9 VSS 0.254197f
C5335 ua[2].n1 VSS 1.28275f
C5336 ua[2].n2 VSS 0.434029f
C5337 ua[2].t13 VSS 0.187785f
C5338 ua[2].n3 VSS 0.280396f
C5339 ua[2].n4 VSS 0.390968f
C5340 ua[2].t3 VSS 0.247385f
C5341 ua[2].n5 VSS 0.307673f
C5342 ua[2].t15 VSS 0.191554f
C5343 ua[2].t2 VSS 0.254197f
C5344 ua[2].n6 VSS 1.28275f
C5345 ua[2].n7 VSS 0.434029f
C5346 ua[2].t14 VSS 0.187785f
C5347 ua[2].n8 VSS 0.280396f
C5348 ua[2].n9 VSS 0.385643f
C5349 ua[2].n10 VSS 0.201153f
C5350 ua[2].n11 VSS 0.0295f
C5351 ua[2].n12 VSS 0.068599f
C5352 ua[2].n13 VSS 0.274656f
C5353 ua[2].t7 VSS 0.247385f
C5354 ua[2].n14 VSS 0.307673f
C5355 ua[2].t1 VSS 0.191554f
C5356 ua[2].t6 VSS 0.254197f
C5357 ua[2].n15 VSS 1.28275f
C5358 ua[2].n16 VSS 0.434029f
C5359 ua[2].t0 VSS 0.187785f
C5360 ua[2].n17 VSS 0.280396f
C5361 ua[2].n18 VSS 0.380387f
C5362 ua[2].n19 VSS 0.206106f
C5363 ua[2].n20 VSS 0.522334f
C5364 ua[2].t5 VSS 0.247385f
C5365 ua[2].n21 VSS 0.307673f
C5366 ua[2].t10 VSS 0.191554f
C5367 ua[2].t4 VSS 0.254197f
C5368 ua[2].n22 VSS 1.28275f
C5369 ua[2].n23 VSS 0.434029f
C5370 ua[2].t11 VSS 0.187785f
C5371 ua[2].n24 VSS 0.280396f
C5372 ua[2].n25 VSS 0.383777f
C5373 ua[2].n26 VSS 0.202647f
C5374 ua[2].n27 VSS 0.509311f
C5375 ua[2].n28 VSS 9.99833f
C5376 ua[3].t7 VSS 0.195583f
C5377 ua[3].n0 VSS 0.292041f
C5378 ua[3].t9 VSS 0.199509f
C5379 ua[3].t3 VSS 0.264753f
C5380 ua[3].n1 VSS 1.33602f
C5381 ua[3].n2 VSS 0.452054f
C5382 ua[3].t2 VSS 0.257658f
C5383 ua[3].n3 VSS 0.32045f
C5384 ua[3].n4 VSS 0.405279f
C5385 ua[3].t0 VSS 0.195583f
C5386 ua[3].n5 VSS 0.292041f
C5387 ua[3].t1 VSS 0.199509f
C5388 ua[3].t6 VSS 0.264753f
C5389 ua[3].n6 VSS 1.33602f
C5390 ua[3].n7 VSS 0.452054f
C5391 ua[3].t8 VSS 0.257658f
C5392 ua[3].n8 VSS 0.32045f
C5393 ua[3].n9 VSS 0.407204f
C5394 ua[3].t4 VSS 0.370241f
C5395 ua[3].t5 VSS 0.261912f
C5396 ua[3].n10 VSS 2.0306f
C5397 ua[3].t11 VSS 0.205641f
C5398 ua[3].t10 VSS 0.377153f
C5399 ua[3].n11 VSS 2.11001f
C5400 ua[3].n12 VSS 0.336309f
C5401 ua[3].n13 VSS 0.069845f
C5402 ua[3].n14 VSS 0.028001f
C5403 ua[3].n15 VSS 1.71586f
C5404 ua[3].n16 VSS 0.514233f
C5405 ua[3].n17 VSS 0.337655f
C5406 muxtest_0.x2.x2.GP1.t1 VSS 0.012908f
C5407 muxtest_0.x2.x2.GP1.t0 VSS 0.012908f
C5408 muxtest_0.x2.x2.GP1.n0 VSS 0.028358f
C5409 muxtest_0.x2.x2.GP1.n1 VSS 0.018329f
C5410 muxtest_0.x2.x2.GP1.t5 VSS 0.653268f
C5411 muxtest_0.x2.x2.GP1.t4 VSS 0.671486f
C5412 muxtest_0.x2.x2.GP1.n2 VSS 2.37213f
C5413 muxtest_0.x2.x2.GP1.t3 VSS 0.019859f
C5414 muxtest_0.x2.x2.GP1.t2 VSS 0.019859f
C5415 muxtest_0.x2.x2.GP1.n3 VSS 0.04092f
C5416 muxtest_0.x2.x2.GP1.n4 VSS 0.100085f
C5417 muxtest_0.x2.x2.GP1.n5 VSS 0.021877f
C5418 VDPWR.n0 VSS 0.003488f
C5419 VDPWR.t881 VSS 0.007172f
C5420 VDPWR.n1 VSS 0.007983f
C5421 VDPWR.t113 VSS 7.56e-19
C5422 VDPWR.t197 VSS 0.001148f
C5423 VDPWR.n2 VSS 0.001983f
C5424 VDPWR.t879 VSS 0.007175f
C5425 VDPWR.t307 VSS 0.00704f
C5426 VDPWR.n3 VSS 0.006705f
C5427 VDPWR.n4 VSS 0.003488f
C5428 VDPWR.n5 VSS 0.003158f
C5429 VDPWR.t56 VSS 0.001036f
C5430 VDPWR.n6 VSS 0.00294f
C5431 VDPWR.t217 VSS 0.004259f
C5432 VDPWR.n7 VSS 0.00392f
C5433 VDPWR.n8 VSS 0.003499f
C5434 VDPWR.t305 VSS 0.007175f
C5435 VDPWR.n9 VSS 5.76e-19
C5436 VDPWR.t988 VSS 0.003015f
C5437 VDPWR.t662 VSS 0.004984f
C5438 VDPWR.n10 VSS 0.004913f
C5439 VDPWR.n11 VSS 0.005888f
C5440 VDPWR.t1217 VSS 0.020799f
C5441 VDPWR.n12 VSS 0.018812f
C5442 VDPWR.t261 VSS 5.64e-19
C5443 VDPWR.t793 VSS 0.001513f
C5444 VDPWR.n13 VSS 0.006904f
C5445 VDPWR.n14 VSS 0.003647f
C5446 VDPWR.t663 VSS 0.004984f
C5447 VDPWR.n15 VSS 0.01361f
C5448 VDPWR.n16 VSS 0.010753f
C5449 VDPWR.n17 VSS 0.013967f
C5450 VDPWR.n18 VSS 0.008065f
C5451 VDPWR.n19 VSS 0.005888f
C5452 VDPWR.n20 VSS 0.004416f
C5453 VDPWR.n21 VSS 0.005354f
C5454 VDPWR.n22 VSS 0.006068f
C5455 VDPWR.n23 VSS 0.013691f
C5456 VDPWR.t1038 VSS 0.014151f
C5457 VDPWR.n24 VSS 7.37e-19
C5458 VDPWR.n25 VSS 0.004416f
C5459 VDPWR.n26 VSS 0.00136f
C5460 VDPWR.t131 VSS 7.56e-19
C5461 VDPWR.t961 VSS 0.001148f
C5462 VDPWR.n27 VSS 0.001983f
C5463 VDPWR.n28 VSS 0.005856f
C5464 VDPWR.n29 VSS 0.003488f
C5465 VDPWR.t1282 VSS 0.020799f
C5466 VDPWR.n30 VSS 0.005184f
C5467 VDPWR.n31 VSS 0.003488f
C5468 VDPWR.t207 VSS 5.64e-19
C5469 VDPWR.t909 VSS 0.001513f
C5470 VDPWR.n32 VSS 0.006904f
C5471 VDPWR.t1268 VSS 0.020799f
C5472 VDPWR.t927 VSS 0.003047f
C5473 VDPWR.n33 VSS 0.009651f
C5474 VDPWR.n34 VSS 0.005344f
C5475 VDPWR.n35 VSS 0.002933f
C5476 VDPWR.t529 VSS 0.004984f
C5477 VDPWR.n36 VSS 0.004913f
C5478 VDPWR.n37 VSS 0.018812f
C5479 VDPWR.n38 VSS 0.008065f
C5480 VDPWR.n39 VSS 0.013967f
C5481 VDPWR.t926 VSS 0.02849f
C5482 VDPWR.t908 VSS 0.027547f
C5483 VDPWR.t528 VSS 0.020377f
C5484 VDPWR.t206 VSS 0.029245f
C5485 VDPWR.t1136 VSS 0.02849f
C5486 VDPWR.t930 VSS 0.032453f
C5487 VDPWR.t960 VSS 0.023585f
C5488 VDPWR.t130 VSS 0.012641f
C5489 VDPWR.t208 VSS 0.005849f
C5490 VDPWR.t210 VSS 0.020566f
C5491 VDPWR.n40 VSS 0.026837f
C5492 VDPWR.t211 VSS 0.007137f
C5493 VDPWR.n41 VSS 0.002016f
C5494 VDPWR.n42 VSS 0.0024f
C5495 VDPWR.n43 VSS 0.018611f
C5496 VDPWR.n44 VSS 0.005471f
C5497 VDPWR.t530 VSS 0.004984f
C5498 VDPWR.n45 VSS 0.008777f
C5499 VDPWR.n46 VSS 0.010753f
C5500 VDPWR.n47 VSS 0.003648f
C5501 VDPWR.n48 VSS 0.02906f
C5502 VDPWR.n49 VSS 0.039529f
C5503 VDPWR.t712 VSS 0.004984f
C5504 VDPWR.n50 VSS 0.009746f
C5505 VDPWR.n51 VSS 0.018812f
C5506 VDPWR.n52 VSS 0.011593f
C5507 VDPWR.t950 VSS 0.007172f
C5508 VDPWR.n53 VSS 0.00838f
C5509 VDPWR.n54 VSS 0.003488f
C5510 VDPWR.n55 VSS 0.001519f
C5511 VDPWR.n56 VSS 0.001519f
C5512 VDPWR.n57 VSS 0.1025f
C5513 VDPWR.t569 VSS 0.004984f
C5514 VDPWR.n58 VSS 0.004913f
C5515 VDPWR.n59 VSS 0.005888f
C5516 VDPWR.t1215 VSS 0.020799f
C5517 VDPWR.n60 VSS 0.018812f
C5518 VDPWR.n61 VSS 0.003647f
C5519 VDPWR.t570 VSS 0.004984f
C5520 VDPWR.n62 VSS 0.01361f
C5521 VDPWR.n63 VSS 0.014953f
C5522 VDPWR.n64 VSS 0.011593f
C5523 VDPWR.n65 VSS 0.005888f
C5524 VDPWR.n66 VSS 0.004416f
C5525 VDPWR.n67 VSS 0.005604f
C5526 VDPWR.t1032 VSS 0.007175f
C5527 VDPWR.n68 VSS 0.009278f
C5528 VDPWR.n69 VSS 0.003488f
C5529 VDPWR.n70 VSS 0.005888f
C5530 VDPWR.n71 VSS 0.004416f
C5531 VDPWR.t60 VSS 0.007172f
C5532 VDPWR.n72 VSS 0.00847f
C5533 VDPWR.t929 VSS 0.007175f
C5534 VDPWR.n73 VSS 0.009165f
C5535 VDPWR.n74 VSS 0.003488f
C5536 VDPWR.n75 VSS 0.005888f
C5537 VDPWR.n76 VSS 0.004416f
C5538 VDPWR.t1022 VSS 0.007172f
C5539 VDPWR.n77 VSS 0.00847f
C5540 VDPWR.t947 VSS 0.007175f
C5541 VDPWR.n78 VSS 0.009165f
C5542 VDPWR.n79 VSS 0.001519f
C5543 VDPWR.n80 VSS 0.005888f
C5544 VDPWR.n81 VSS 0.004416f
C5545 VDPWR.n82 VSS 0.00224f
C5546 VDPWR.t711 VSS 0.064097f
C5547 VDPWR.t568 VSS 0.039378f
C5548 VDPWR.t1031 VSS 0.016158f
C5549 VDPWR.t59 VSS 0.022364f
C5550 VDPWR.t928 VSS 0.016158f
C5551 VDPWR.t1021 VSS 0.022364f
C5552 VDPWR.t946 VSS 0.016158f
C5553 VDPWR.t949 VSS 0.024184f
C5554 VDPWR.n83 VSS 0.026472f
C5555 VDPWR.n84 VSS 0.012237f
C5556 VDPWR.n85 VSS 0.005471f
C5557 VDPWR.t713 VSS 0.004984f
C5558 VDPWR.n86 VSS 0.008777f
C5559 VDPWR.n87 VSS 0.014953f
C5560 VDPWR.n88 VSS 0.002976f
C5561 VDPWR.n89 VSS 0.027044f
C5562 VDPWR.n90 VSS 0.026223f
C5563 VDPWR.n91 VSS 6.08e-19
C5564 VDPWR.t209 VSS 0.007136f
C5565 VDPWR.n92 VSS 0.013312f
C5566 VDPWR.t1138 VSS 0.007172f
C5567 VDPWR.n93 VSS 0.008357f
C5568 VDPWR.t931 VSS 0.002363f
C5569 VDPWR.t1039 VSS 0.006281f
C5570 VDPWR.n94 VSS 0.003563f
C5571 VDPWR.t1137 VSS 0.007041f
C5572 VDPWR.n95 VSS 0.007429f
C5573 VDPWR.n96 VSS 0.009555f
C5574 VDPWR.n97 VSS 0.001258f
C5575 VDPWR.n98 VSS 0.005888f
C5576 VDPWR.n99 VSS 0.003488f
C5577 VDPWR.n100 VSS 0.002016f
C5578 VDPWR.n101 VSS 0.00224f
C5579 VDPWR.n102 VSS 0.012275f
C5580 VDPWR.n103 VSS 0.032875f
C5581 VDPWR.t112 VSS 0.006226f
C5582 VDPWR.t880 VSS 0.016226f
C5583 VDPWR.t878 VSS 0.018113f
C5584 VDPWR.t196 VSS 0.012641f
C5585 VDPWR.t55 VSS 0.023585f
C5586 VDPWR.t306 VSS 0.033207f
C5587 VDPWR.t304 VSS 0.016226f
C5588 VDPWR.t216 VSS 0.012641f
C5589 VDPWR.t260 VSS 0.029245f
C5590 VDPWR.t661 VSS 0.020377f
C5591 VDPWR.t792 VSS 0.027547f
C5592 VDPWR.t987 VSS 0.02849f
C5593 VDPWR.n104 VSS 0.019402f
C5594 VDPWR.n105 VSS 0.005637f
C5595 VDPWR.n106 VSS 0.003862f
C5596 VDPWR.n107 VSS 0.009272f
C5597 VDPWR.n108 VSS 0.002696f
C5598 VDPWR.n109 VSS 0.005888f
C5599 VDPWR.n110 VSS 0.004416f
C5600 VDPWR.n111 VSS 0.002625f
C5601 VDPWR.n112 VSS 0.008924f
C5602 VDPWR.n113 VSS 0.006148f
C5603 VDPWR.n114 VSS 0.004064f
C5604 VDPWR.n115 VSS 0.011493f
C5605 VDPWR.n116 VSS 0.0731f
C5606 VDPWR.n117 VSS 7.840919f
C5607 VDPWR.n118 VSS 0.489074f
C5608 VDPWR.t893 VSS 0.007172f
C5609 VDPWR.n119 VSS 0.00838f
C5610 VDPWR.t369 VSS 0.007175f
C5611 VDPWR.n120 VSS 0.009029f
C5612 VDPWR.n121 VSS 0.023921f
C5613 VDPWR.t371 VSS 0.007172f
C5614 VDPWR.t75 VSS 0.007175f
C5615 VDPWR.n122 VSS 0.010921f
C5616 VDPWR.t77 VSS 0.007172f
C5617 VDPWR.n123 VSS 0.00847f
C5618 VDPWR.t245 VSS 0.007175f
C5619 VDPWR.t247 VSS 0.007172f
C5620 VDPWR.n124 VSS 0.00847f
C5621 VDPWR.t87 VSS 0.007175f
C5622 VDPWR.t85 VSS 0.007172f
C5623 VDPWR.n125 VSS 0.00847f
C5624 VDPWR.t89 VSS 0.007175f
C5625 VDPWR.t91 VSS 0.007172f
C5626 VDPWR.n126 VSS 0.00847f
C5627 VDPWR.n127 VSS 0.014476f
C5628 VDPWR.n128 VSS 0.013372f
C5629 VDPWR.t885 VSS 0.007172f
C5630 VDPWR.n129 VSS 0.00847f
C5631 VDPWR.n130 VSS 0.001519f
C5632 VDPWR.n131 VSS 0.001519f
C5633 VDPWR.n132 VSS 0.001519f
C5634 VDPWR.n133 VSS 0.001519f
C5635 VDPWR.n134 VSS 0.022941f
C5636 VDPWR.t905 VSS 0.007172f
C5637 VDPWR.n135 VSS 0.00838f
C5638 VDPWR.n136 VSS 0.01181f
C5639 VDPWR.n137 VSS 0.008587f
C5640 VDPWR.n138 VSS 0.013249f
C5641 VDPWR.t241 VSS 0.007179f
C5642 VDPWR.t861 VSS 0.0018f
C5643 VDPWR.t243 VSS 0.0018f
C5644 VDPWR.n139 VSS 0.003864f
C5645 VDPWR.n140 VSS 0.005287f
C5646 VDPWR.t859 VSS 0.006979f
C5647 VDPWR.n141 VSS 0.009924f
C5648 VDPWR.n142 VSS 0.04768f
C5649 VDPWR.n143 VSS 0.001711f
C5650 VDPWR.n144 VSS 0.010005f
C5651 VDPWR.n145 VSS 0.01181f
C5652 VDPWR.t858 VSS 0.041519f
C5653 VDPWR.t860 VSS 0.017977f
C5654 VDPWR.t242 VSS 0.017977f
C5655 VDPWR.t240 VSS 0.015837f
C5656 VDPWR.n146 VSS 0.021229f
C5657 VDPWR.n147 VSS 0.022941f
C5658 VDPWR.n148 VSS 0.01181f
C5659 VDPWR.n149 VSS 0.008587f
C5660 VDPWR.n150 VSS 0.008587f
C5661 VDPWR.n151 VSS 0.013372f
C5662 VDPWR.n152 VSS 0.001519f
C5663 VDPWR.n153 VSS 0.001519f
C5664 VDPWR.n154 VSS 0.001519f
C5665 VDPWR.t887 VSS 0.007175f
C5666 VDPWR.n155 VSS 0.009165f
C5667 VDPWR.n156 VSS 0.013372f
C5668 VDPWR.n157 VSS 0.022572f
C5669 VDPWR.n158 VSS 0.016929f
C5670 VDPWR.t889 VSS 0.007172f
C5671 VDPWR.n159 VSS 0.00847f
C5672 VDPWR.t181 VSS 0.007175f
C5673 VDPWR.n160 VSS 0.009165f
C5674 VDPWR.n161 VSS 0.013372f
C5675 VDPWR.n162 VSS 0.022572f
C5676 VDPWR.n163 VSS 0.016929f
C5677 VDPWR.t183 VSS 0.007172f
C5678 VDPWR.n164 VSS 0.00847f
C5679 VDPWR.t171 VSS 0.007175f
C5680 VDPWR.n165 VSS 0.009165f
C5681 VDPWR.n166 VSS 0.013372f
C5682 VDPWR.n167 VSS 0.022572f
C5683 VDPWR.n168 VSS 0.016929f
C5684 VDPWR.t173 VSS 0.007172f
C5685 VDPWR.n169 VSS 0.00847f
C5686 VDPWR.t903 VSS 0.007175f
C5687 VDPWR.n170 VSS 0.009165f
C5688 VDPWR.n171 VSS 0.001519f
C5689 VDPWR.n172 VSS 0.022572f
C5690 VDPWR.n173 VSS 0.016929f
C5691 VDPWR.n174 VSS 0.008587f
C5692 VDPWR.n175 VSS 0.011946f
C5693 VDPWR.n176 VSS 0.028292f
C5694 VDPWR.t904 VSS 0.024184f
C5695 VDPWR.t902 VSS 0.015813f
C5696 VDPWR.t172 VSS 0.022364f
C5697 VDPWR.t170 VSS 0.016158f
C5698 VDPWR.t182 VSS 0.022364f
C5699 VDPWR.t180 VSS 0.016158f
C5700 VDPWR.t888 VSS 0.022364f
C5701 VDPWR.t886 VSS 0.016158f
C5702 VDPWR.t884 VSS 0.022364f
C5703 VDPWR.t882 VSS 0.016158f
C5704 VDPWR.t291 VSS 0.022364f
C5705 VDPWR.t289 VSS 0.016158f
C5706 VDPWR.t842 VSS 0.022364f
C5707 VDPWR.t844 VSS 0.016158f
C5708 VDPWR.t840 VSS 0.022364f
C5709 VDPWR.t838 VSS 0.016158f
C5710 VDPWR.t898 VSS 0.022364f
C5711 VDPWR.t896 VSS 0.016158f
C5712 VDPWR.n177 VSS 0.008587f
C5713 VDPWR.n178 VSS 0.026055f
C5714 VDPWR.t897 VSS 0.007175f
C5715 VDPWR.n179 VSS 0.009029f
C5716 VDPWR.n180 VSS 0.013372f
C5717 VDPWR.n181 VSS 0.022572f
C5718 VDPWR.n182 VSS 0.016929f
C5719 VDPWR.t899 VSS 0.007172f
C5720 VDPWR.n183 VSS 0.00847f
C5721 VDPWR.t839 VSS 0.007175f
C5722 VDPWR.n184 VSS 0.009165f
C5723 VDPWR.n185 VSS 0.013372f
C5724 VDPWR.n186 VSS 0.022572f
C5725 VDPWR.n187 VSS 0.016929f
C5726 VDPWR.t841 VSS 0.007172f
C5727 VDPWR.n188 VSS 0.00847f
C5728 VDPWR.t845 VSS 0.007175f
C5729 VDPWR.n189 VSS 0.009165f
C5730 VDPWR.n190 VSS 0.013372f
C5731 VDPWR.n191 VSS 0.022572f
C5732 VDPWR.n192 VSS 0.016929f
C5733 VDPWR.t843 VSS 0.007172f
C5734 VDPWR.n193 VSS 0.00847f
C5735 VDPWR.t290 VSS 0.007175f
C5736 VDPWR.n194 VSS 0.009165f
C5737 VDPWR.n195 VSS 0.013372f
C5738 VDPWR.n196 VSS 0.022572f
C5739 VDPWR.n197 VSS 0.016929f
C5740 VDPWR.t292 VSS 0.007172f
C5741 VDPWR.n198 VSS 0.00847f
C5742 VDPWR.t883 VSS 0.007175f
C5743 VDPWR.n199 VSS 0.009165f
C5744 VDPWR.n200 VSS 0.001519f
C5745 VDPWR.n201 VSS 0.01374f
C5746 VDPWR.n202 VSS 1.62819f
C5747 VDPWR.n203 VSS 1.62991f
C5748 VDPWR.t313 VSS 0.007175f
C5749 VDPWR.t311 VSS 0.007172f
C5750 VDPWR.n204 VSS 0.00847f
C5751 VDPWR.t276 VSS 0.007175f
C5752 VDPWR.t274 VSS 0.007172f
C5753 VDPWR.n205 VSS 0.00847f
C5754 VDPWR.t278 VSS 0.007175f
C5755 VDPWR.t280 VSS 0.007172f
C5756 VDPWR.n206 VSS 0.00847f
C5757 VDPWR.t895 VSS 0.007175f
C5758 VDPWR.n207 VSS 0.023921f
C5759 VDPWR.n208 VSS 0.028948f
C5760 VDPWR.n209 VSS 0.001519f
C5761 VDPWR.n210 VSS 0.009165f
C5762 VDPWR.n211 VSS 0.010921f
C5763 VDPWR.n212 VSS 0.023921f
C5764 VDPWR.n213 VSS 0.028948f
C5765 VDPWR.n214 VSS 0.001519f
C5766 VDPWR.n215 VSS 0.009165f
C5767 VDPWR.n216 VSS 0.010921f
C5768 VDPWR.n217 VSS 0.023921f
C5769 VDPWR.n218 VSS 0.028948f
C5770 VDPWR.n219 VSS 0.001519f
C5771 VDPWR.n220 VSS 0.009165f
C5772 VDPWR.n221 VSS 0.010921f
C5773 VDPWR.n222 VSS 0.023921f
C5774 VDPWR.n223 VSS 0.028948f
C5775 VDPWR.n224 VSS 0.001519f
C5776 VDPWR.n225 VSS 0.009165f
C5777 VDPWR.n226 VSS 0.010921f
C5778 VDPWR.n227 VSS 0.023921f
C5779 VDPWR.n228 VSS 0.019415f
C5780 VDPWR.n229 VSS 0.001519f
C5781 VDPWR.n230 VSS 0.009165f
C5782 VDPWR.n231 VSS 0.010921f
C5783 VDPWR.n232 VSS 0.023921f
C5784 VDPWR.n233 VSS 0.028948f
C5785 VDPWR.n234 VSS 0.001519f
C5786 VDPWR.n235 VSS 0.009165f
C5787 VDPWR.n236 VSS 0.010921f
C5788 VDPWR.n237 VSS 0.023921f
C5789 VDPWR.n238 VSS 0.028948f
C5790 VDPWR.n239 VSS 0.001519f
C5791 VDPWR.n240 VSS 0.009165f
C5792 VDPWR.n241 VSS 0.010921f
C5793 VDPWR.n242 VSS 0.023921f
C5794 VDPWR.n243 VSS 0.028948f
C5795 VDPWR.n244 VSS 0.001519f
C5796 VDPWR.n245 VSS 0.009165f
C5797 VDPWR.n246 VSS 0.00847f
C5798 VDPWR.n247 VSS 0.001519f
C5799 VDPWR.n248 VSS 0.028948f
C5800 VDPWR.n249 VSS 0.010921f
C5801 VDPWR.n250 VSS 0.031124f
C5802 VDPWR.t368 VSS 0.01252f
C5803 VDPWR.t370 VSS 0.026002f
C5804 VDPWR.t74 VSS 0.01252f
C5805 VDPWR.t76 VSS 0.026002f
C5806 VDPWR.t244 VSS 0.01252f
C5807 VDPWR.t246 VSS 0.026002f
C5808 VDPWR.t86 VSS 0.01252f
C5809 VDPWR.t84 VSS 0.026002f
C5810 VDPWR.t88 VSS 0.01252f
C5811 VDPWR.t90 VSS 0.026002f
C5812 VDPWR.t312 VSS 0.01252f
C5813 VDPWR.t310 VSS 0.026002f
C5814 VDPWR.t275 VSS 0.01252f
C5815 VDPWR.t273 VSS 0.026002f
C5816 VDPWR.t277 VSS 0.01252f
C5817 VDPWR.t279 VSS 0.026002f
C5818 VDPWR.t894 VSS 0.01252f
C5819 VDPWR.t892 VSS 0.03644f
C5820 VDPWR.n251 VSS 0.035343f
C5821 VDPWR.n252 VSS 0.012134f
C5822 VDPWR.n253 VSS 3.92216f
C5823 VDPWR.n254 VSS 0.058044f
C5824 VDPWR.n255 VSS 0.105387f
C5825 VDPWR.n256 VSS 4.47053f
C5826 VDPWR.n257 VSS 2.12953f
C5827 VDPWR.n258 VSS 0.003488f
C5828 VDPWR.t177 VSS 0.007172f
C5829 VDPWR.n259 VSS 0.007983f
C5830 VDPWR.t109 VSS 7.56e-19
C5831 VDPWR.t990 VSS 0.001148f
C5832 VDPWR.n260 VSS 0.001983f
C5833 VDPWR.t179 VSS 0.007175f
C5834 VDPWR.t71 VSS 0.00704f
C5835 VDPWR.n261 VSS 0.006705f
C5836 VDPWR.n262 VSS 0.003488f
C5837 VDPWR.n263 VSS 0.003158f
C5838 VDPWR.t1090 VSS 0.001036f
C5839 VDPWR.n264 VSS 0.00294f
C5840 VDPWR.t189 VSS 0.004259f
C5841 VDPWR.n265 VSS 0.00392f
C5842 VDPWR.n266 VSS 0.003499f
C5843 VDPWR.t73 VSS 0.007175f
C5844 VDPWR.n267 VSS 5.76e-19
C5845 VDPWR.t765 VSS 0.003015f
C5846 VDPWR.t540 VSS 0.004984f
C5847 VDPWR.n268 VSS 0.004913f
C5848 VDPWR.n269 VSS 0.005888f
C5849 VDPWR.t1228 VSS 0.020799f
C5850 VDPWR.n270 VSS 0.018812f
C5851 VDPWR.t286 VSS 5.64e-19
C5852 VDPWR.t62 VSS 0.001513f
C5853 VDPWR.n271 VSS 0.006904f
C5854 VDPWR.n272 VSS 0.003647f
C5855 VDPWR.t541 VSS 0.004984f
C5856 VDPWR.n273 VSS 0.01361f
C5857 VDPWR.n274 VSS 0.010753f
C5858 VDPWR.n275 VSS 0.013967f
C5859 VDPWR.n276 VSS 0.008065f
C5860 VDPWR.n277 VSS 0.005888f
C5861 VDPWR.n278 VSS 0.004416f
C5862 VDPWR.n279 VSS 0.005354f
C5863 VDPWR.n280 VSS 0.006068f
C5864 VDPWR.n281 VSS 0.013691f
C5865 VDPWR.t110 VSS 0.014151f
C5866 VDPWR.n282 VSS 7.37e-19
C5867 VDPWR.n283 VSS 0.004416f
C5868 VDPWR.n284 VSS 0.00136f
C5869 VDPWR.t236 VSS 7.56e-19
C5870 VDPWR.t849 VSS 0.001148f
C5871 VDPWR.n285 VSS 0.001983f
C5872 VDPWR.n286 VSS 0.005856f
C5873 VDPWR.n287 VSS 0.003488f
C5874 VDPWR.t1201 VSS 0.020799f
C5875 VDPWR.n288 VSS 0.005184f
C5876 VDPWR.n289 VSS 0.003488f
C5877 VDPWR.t303 VSS 5.64e-19
C5878 VDPWR.t1092 VSS 0.001513f
C5879 VDPWR.n290 VSS 0.006904f
C5880 VDPWR.t1200 VSS 0.020799f
C5881 VDPWR.t107 VSS 0.003047f
C5882 VDPWR.n291 VSS 0.009651f
C5883 VDPWR.n292 VSS 0.005344f
C5884 VDPWR.n293 VSS 0.002933f
C5885 VDPWR.t600 VSS 0.004984f
C5886 VDPWR.n294 VSS 0.004913f
C5887 VDPWR.n295 VSS 0.018812f
C5888 VDPWR.n296 VSS 0.008065f
C5889 VDPWR.n297 VSS 0.013967f
C5890 VDPWR.t106 VSS 0.02849f
C5891 VDPWR.t1091 VSS 0.027547f
C5892 VDPWR.t599 VSS 0.020377f
C5893 VDPWR.t302 VSS 0.029245f
C5894 VDPWR.t851 VSS 0.02849f
C5895 VDPWR.t104 VSS 0.032453f
C5896 VDPWR.t848 VSS 0.023585f
C5897 VDPWR.t235 VSS 0.012641f
C5898 VDPWR.t1010 VSS 0.005849f
C5899 VDPWR.t1008 VSS 0.020566f
C5900 VDPWR.n298 VSS 0.026837f
C5901 VDPWR.t1009 VSS 0.007137f
C5902 VDPWR.n299 VSS 0.002016f
C5903 VDPWR.n300 VSS 0.0024f
C5904 VDPWR.n301 VSS 0.018611f
C5905 VDPWR.n302 VSS 0.005471f
C5906 VDPWR.t601 VSS 0.004984f
C5907 VDPWR.n303 VSS 0.008777f
C5908 VDPWR.n304 VSS 0.010753f
C5909 VDPWR.n305 VSS 0.003648f
C5910 VDPWR.n306 VSS 0.02906f
C5911 VDPWR.n307 VSS 0.039529f
C5912 VDPWR.t597 VSS 0.004984f
C5913 VDPWR.n308 VSS 0.009746f
C5914 VDPWR.n309 VSS 0.018812f
C5915 VDPWR.n310 VSS 0.011593f
C5916 VDPWR.t1097 VSS 0.007172f
C5917 VDPWR.n311 VSS 0.00838f
C5918 VDPWR.n312 VSS 0.003488f
C5919 VDPWR.n313 VSS 0.001519f
C5920 VDPWR.n314 VSS 0.001519f
C5921 VDPWR.n315 VSS 0.1025f
C5922 VDPWR.t436 VSS 0.004984f
C5923 VDPWR.n316 VSS 0.004913f
C5924 VDPWR.n317 VSS 0.005888f
C5925 VDPWR.t1263 VSS 0.020799f
C5926 VDPWR.n318 VSS 0.018812f
C5927 VDPWR.t437 VSS 0.004984f
C5928 VDPWR.n319 VSS 0.003647f
C5929 VDPWR.n320 VSS 0.01361f
C5930 VDPWR.n321 VSS 0.014953f
C5931 VDPWR.n322 VSS 0.011593f
C5932 VDPWR.n323 VSS 0.005888f
C5933 VDPWR.n324 VSS 0.004416f
C5934 VDPWR.n325 VSS 0.005604f
C5935 VDPWR.t234 VSS 0.007175f
C5936 VDPWR.n326 VSS 0.009278f
C5937 VDPWR.n327 VSS 0.003488f
C5938 VDPWR.n328 VSS 0.005888f
C5939 VDPWR.n329 VSS 0.004416f
C5940 VDPWR.t238 VSS 0.007172f
C5941 VDPWR.n330 VSS 0.00847f
C5942 VDPWR.t815 VSS 0.007175f
C5943 VDPWR.n331 VSS 0.009165f
C5944 VDPWR.n332 VSS 0.003488f
C5945 VDPWR.n333 VSS 0.005888f
C5946 VDPWR.n334 VSS 0.004416f
C5947 VDPWR.t1046 VSS 0.007172f
C5948 VDPWR.n335 VSS 0.00847f
C5949 VDPWR.t1099 VSS 0.007175f
C5950 VDPWR.n336 VSS 0.009165f
C5951 VDPWR.n337 VSS 0.001519f
C5952 VDPWR.n338 VSS 0.005888f
C5953 VDPWR.n339 VSS 0.004416f
C5954 VDPWR.n340 VSS 0.00224f
C5955 VDPWR.t596 VSS 0.064097f
C5956 VDPWR.t435 VSS 0.039378f
C5957 VDPWR.t233 VSS 0.016158f
C5958 VDPWR.t237 VSS 0.022364f
C5959 VDPWR.t814 VSS 0.016158f
C5960 VDPWR.t1045 VSS 0.022364f
C5961 VDPWR.t1098 VSS 0.016158f
C5962 VDPWR.t1096 VSS 0.024184f
C5963 VDPWR.n341 VSS 0.026472f
C5964 VDPWR.n342 VSS 0.012237f
C5965 VDPWR.n343 VSS 0.005471f
C5966 VDPWR.t598 VSS 0.004984f
C5967 VDPWR.n344 VSS 0.008777f
C5968 VDPWR.n345 VSS 0.014953f
C5969 VDPWR.n346 VSS 0.002976f
C5970 VDPWR.n347 VSS 0.027044f
C5971 VDPWR.n348 VSS 0.026223f
C5972 VDPWR.n349 VSS 6.08e-19
C5973 VDPWR.t1011 VSS 0.007136f
C5974 VDPWR.n350 VSS 0.013312f
C5975 VDPWR.t850 VSS 0.007172f
C5976 VDPWR.n351 VSS 0.008357f
C5977 VDPWR.t105 VSS 0.002363f
C5978 VDPWR.t111 VSS 0.006281f
C5979 VDPWR.n352 VSS 0.003563f
C5980 VDPWR.t852 VSS 0.007041f
C5981 VDPWR.n353 VSS 0.007429f
C5982 VDPWR.n354 VSS 0.009555f
C5983 VDPWR.n355 VSS 0.001258f
C5984 VDPWR.n356 VSS 0.005888f
C5985 VDPWR.n357 VSS 0.003488f
C5986 VDPWR.n358 VSS 0.002016f
C5987 VDPWR.n359 VSS 0.00224f
C5988 VDPWR.n360 VSS 0.012275f
C5989 VDPWR.n361 VSS 0.032875f
C5990 VDPWR.t108 VSS 0.006226f
C5991 VDPWR.t176 VSS 0.016226f
C5992 VDPWR.t178 VSS 0.018113f
C5993 VDPWR.t989 VSS 0.012641f
C5994 VDPWR.t1089 VSS 0.023585f
C5995 VDPWR.t70 VSS 0.033207f
C5996 VDPWR.t72 VSS 0.016226f
C5997 VDPWR.t188 VSS 0.012641f
C5998 VDPWR.t285 VSS 0.029245f
C5999 VDPWR.t539 VSS 0.020377f
C6000 VDPWR.t61 VSS 0.027547f
C6001 VDPWR.t764 VSS 0.02849f
C6002 VDPWR.n362 VSS 0.019402f
C6003 VDPWR.n363 VSS 0.005637f
C6004 VDPWR.n364 VSS 0.003862f
C6005 VDPWR.n365 VSS 0.009272f
C6006 VDPWR.n366 VSS 0.002696f
C6007 VDPWR.n367 VSS 0.005888f
C6008 VDPWR.n368 VSS 0.004416f
C6009 VDPWR.n369 VSS 0.002625f
C6010 VDPWR.n370 VSS 0.008924f
C6011 VDPWR.n371 VSS 0.006148f
C6012 VDPWR.n372 VSS 0.004064f
C6013 VDPWR.n373 VSS 0.011493f
C6014 VDPWR.n374 VSS 0.089674f
C6015 VDPWR.n375 VSS 0.05908f
C6016 VDPWR.n376 VSS 0.114583f
C6017 VDPWR.n377 VSS 0.318185f
C6018 VDPWR.n378 VSS 0.114492f
C6019 VDPWR.n379 VSS 0.056224f
C6020 VDPWR.n380 VSS 0.076648f
C6021 VDPWR.n381 VSS 0.056138f
C6022 VDPWR.n382 VSS 0.465708f
C6023 VDPWR.t772 VSS 0.619228f
C6024 VDPWR.n385 VSS 0.465708f
C6025 VDPWR.n386 VSS 0.055408f
C6026 VDPWR.n387 VSS 0.036337f
C6027 VDPWR.n388 VSS 0.073206f
C6028 VDPWR.n389 VSS 0.038046f
C6029 VDPWR.n390 VSS 0.114492f
C6030 VDPWR.n391 VSS 0.056224f
C6031 VDPWR.n392 VSS 0.076648f
C6032 VDPWR.n393 VSS 0.056138f
C6033 VDPWR.n394 VSS 0.465708f
C6034 VDPWR.t119 VSS 0.619228f
C6035 VDPWR.n397 VSS 0.465708f
C6036 VDPWR.n398 VSS 0.055408f
C6037 VDPWR.n399 VSS 0.036337f
C6038 VDPWR.n400 VSS 0.073206f
C6039 VDPWR.n401 VSS 0.071425f
C6040 VDPWR.n402 VSS 0.171041f
C6041 VDPWR.n403 VSS 0.073588f
C6042 VDPWR.n404 VSS 0.035269f
C6043 VDPWR.n405 VSS 0.114487f
C6044 VDPWR.n406 VSS 0.055474f
C6045 VDPWR.n407 VSS 0.055474f
C6046 VDPWR.n408 VSS 0.055293f
C6047 VDPWR.n409 VSS 0.076656f
C6048 VDPWR.n410 VSS 0.247132f
C6049 VDPWR.t345 VSS 0.356671f
C6050 VDPWR.n411 VSS 0.344366f
C6051 VDPWR.t1037 VSS 0.356671f
C6052 VDPWR.n412 VSS 0.247132f
C6053 VDPWR.n413 VSS 2.15e-19
C6054 VDPWR.n414 VSS 0.025894f
C6055 VDPWR.n415 VSS 0.035269f
C6056 VDPWR.n416 VSS 0.076656f
C6057 VDPWR.n417 VSS 0.247132f
C6058 VDPWR.n418 VSS 2.38e-19
C6059 VDPWR.n419 VSS 0.247132f
C6060 VDPWR.t958 VSS 0.356671f
C6061 VDPWR.t959 VSS 0.356671f
C6062 VDPWR.n420 VSS 0.055293f
C6063 VDPWR.n421 VSS 0.055474f
C6064 VDPWR.n422 VSS 0.344366f
C6065 VDPWR.n423 VSS 0.055474f
C6066 VDPWR.n424 VSS 0.114487f
C6067 VDPWR.n425 VSS 0.060635f
C6068 VDPWR.n426 VSS 0.018181f
C6069 VDPWR.n427 VSS 0.029454f
C6070 VDPWR.n428 VSS 0.073168f
C6071 VDPWR.n429 VSS 0.084539f
C6072 VDPWR.n430 VSS 0.035235f
C6073 VDPWR.n431 VSS 0.114487f
C6074 VDPWR.n432 VSS 0.00445f
C6075 VDPWR.n433 VSS 0.055474f
C6076 VDPWR.n434 VSS 0.055474f
C6077 VDPWR.n435 VSS 0.055293f
C6078 VDPWR.n436 VSS 0.076656f
C6079 VDPWR.n437 VSS 0.247132f
C6080 VDPWR.t120 VSS 0.356671f
C6081 VDPWR.n438 VSS 0.344366f
C6082 VDPWR.t123 VSS 0.356671f
C6083 VDPWR.n439 VSS 0.247132f
C6084 VDPWR.n440 VSS 0.002025f
C6085 VDPWR.n441 VSS 0.060694f
C6086 VDPWR.n442 VSS 0.018181f
C6087 VDPWR.n443 VSS 0.029169f
C6088 VDPWR.n444 VSS 0.067579f
C6089 VDPWR.n445 VSS 0.082325f
C6090 VDPWR.n446 VSS 0.035121f
C6091 VDPWR.n447 VSS 0.114487f
C6092 VDPWR.n448 VSS 0.004458f
C6093 VDPWR.n449 VSS 0.055474f
C6094 VDPWR.n450 VSS 0.055474f
C6095 VDPWR.n451 VSS 0.055293f
C6096 VDPWR.n452 VSS 0.076656f
C6097 VDPWR.n453 VSS 0.247132f
C6098 VDPWR.t68 VSS 0.356671f
C6099 VDPWR.n454 VSS 0.344366f
C6100 VDPWR.t69 VSS 0.356671f
C6101 VDPWR.n455 VSS 0.247132f
C6102 VDPWR.n456 VSS 0.002138f
C6103 VDPWR.n457 VSS 0.060694f
C6104 VDPWR.n458 VSS 0.018181f
C6105 VDPWR.n459 VSS 0.029169f
C6106 VDPWR.n460 VSS 0.065201f
C6107 VDPWR.n461 VSS 0.075229f
C6108 VDPWR.n462 VSS 0.006257f
C6109 VDPWR.n463 VSS 0.060659f
C6110 VDPWR.n464 VSS 0.018181f
C6111 VDPWR.n465 VSS 0.029431f
C6112 VDPWR.n466 VSS 0.064503f
C6113 VDPWR.n467 VSS 0.08621f
C6114 VDPWR.n468 VSS 0.035269f
C6115 VDPWR.n469 VSS 0.114487f
C6116 VDPWR.n470 VSS 0.055474f
C6117 VDPWR.n471 VSS 0.055474f
C6118 VDPWR.n472 VSS 0.055293f
C6119 VDPWR.n473 VSS 0.076656f
C6120 VDPWR.n474 VSS 0.247132f
C6121 VDPWR.t956 VSS 0.356671f
C6122 VDPWR.n475 VSS 0.344366f
C6123 VDPWR.t957 VSS 0.356671f
C6124 VDPWR.n476 VSS 0.247132f
C6125 VDPWR.n477 VSS 2.38e-19
C6126 VDPWR.n478 VSS 0.006274f
C6127 VDPWR.n479 VSS 0.060635f
C6128 VDPWR.n480 VSS 0.018181f
C6129 VDPWR.n481 VSS 0.029454f
C6130 VDPWR.n482 VSS 0.043811f
C6131 VDPWR.n483 VSS 0.106582f
C6132 VDPWR.n484 VSS 0.035235f
C6133 VDPWR.n485 VSS 0.114487f
C6134 VDPWR.n486 VSS 0.00445f
C6135 VDPWR.n487 VSS 0.055474f
C6136 VDPWR.n488 VSS 0.055474f
C6137 VDPWR.n489 VSS 0.055293f
C6138 VDPWR.n490 VSS 0.076656f
C6139 VDPWR.n491 VSS 0.247132f
C6140 VDPWR.t122 VSS 0.356671f
C6141 VDPWR.n492 VSS 0.344366f
C6142 VDPWR.t121 VSS 0.356671f
C6143 VDPWR.n493 VSS 0.247132f
C6144 VDPWR.n494 VSS 0.002025f
C6145 VDPWR.n495 VSS 0.060694f
C6146 VDPWR.n496 VSS 0.018181f
C6147 VDPWR.n497 VSS 0.029169f
C6148 VDPWR.n498 VSS 0.067579f
C6149 VDPWR.n499 VSS 0.082325f
C6150 VDPWR.n500 VSS 0.035121f
C6151 VDPWR.n501 VSS 0.114487f
C6152 VDPWR.n502 VSS 0.004458f
C6153 VDPWR.n503 VSS 0.055474f
C6154 VDPWR.n504 VSS 0.055474f
C6155 VDPWR.n505 VSS 0.055293f
C6156 VDPWR.n506 VSS 0.076656f
C6157 VDPWR.n507 VSS 0.247132f
C6158 VDPWR.t67 VSS 0.356671f
C6159 VDPWR.n508 VSS 0.344366f
C6160 VDPWR.t13 VSS 0.356671f
C6161 VDPWR.n509 VSS 0.247132f
C6162 VDPWR.n510 VSS 0.002138f
C6163 VDPWR.n511 VSS 0.060694f
C6164 VDPWR.n512 VSS 0.018181f
C6165 VDPWR.n513 VSS 0.029169f
C6166 VDPWR.n514 VSS 0.064853f
C6167 VDPWR.n515 VSS 0.086126f
C6168 VDPWR.n516 VSS 0.035269f
C6169 VDPWR.n517 VSS 0.114487f
C6170 VDPWR.n518 VSS 0.055474f
C6171 VDPWR.n519 VSS 0.055474f
C6172 VDPWR.n520 VSS 0.055293f
C6173 VDPWR.n521 VSS 0.076656f
C6174 VDPWR.n522 VSS 0.247132f
C6175 VDPWR.t1036 VSS 0.356671f
C6176 VDPWR.n523 VSS 0.344366f
C6177 VDPWR.t1035 VSS 0.356671f
C6178 VDPWR.n524 VSS 0.247132f
C6179 VDPWR.n525 VSS 2.15e-19
C6180 VDPWR.n526 VSS 0.006257f
C6181 VDPWR.n527 VSS 0.060659f
C6182 VDPWR.n528 VSS 0.018181f
C6183 VDPWR.n529 VSS 0.029432f
C6184 VDPWR.n530 VSS 0.108553f
C6185 VDPWR.n531 VSS 0.406145f
C6186 VDPWR.n532 VSS 1.02472f
C6187 VDPWR.t951 VSS 0.0028f
C6188 VDPWR.t1202 VSS 0.00165f
C6189 VDPWR.t942 VSS 0.0028f
C6190 VDPWR.t1193 VSS 0.00165f
C6191 VDPWR.n533 VSS 0.004698f
C6192 VDPWR.n534 VSS 0.006946f
C6193 VDPWR.n535 VSS 0.006899f
C6194 VDPWR.n536 VSS 0.002816f
C6195 VDPWR.n537 VSS 0.366828f
C6196 VDPWR.n538 VSS 0.003488f
C6197 VDPWR.t187 VSS 0.007172f
C6198 VDPWR.n539 VSS 0.007983f
C6199 VDPWR.t789 VSS 7.56e-19
C6200 VDPWR.t19 VSS 0.001148f
C6201 VDPWR.n540 VSS 0.001983f
C6202 VDPWR.t185 VSS 0.007175f
C6203 VDPWR.t1165 VSS 0.00704f
C6204 VDPWR.n541 VSS 0.006705f
C6205 VDPWR.n542 VSS 0.003488f
C6206 VDPWR.n543 VSS 0.003158f
C6207 VDPWR.t911 VSS 0.001036f
C6208 VDPWR.n544 VSS 0.00294f
C6209 VDPWR.t965 VSS 0.004259f
C6210 VDPWR.n545 VSS 0.00392f
C6211 VDPWR.n546 VSS 0.003499f
C6212 VDPWR.t1163 VSS 0.007175f
C6213 VDPWR.n547 VSS 5.76e-19
C6214 VDPWR.t146 VSS 0.003015f
C6215 VDPWR.t682 VSS 0.004984f
C6216 VDPWR.n548 VSS 0.004913f
C6217 VDPWR.n549 VSS 0.005888f
C6218 VDPWR.t1207 VSS 0.020799f
C6219 VDPWR.n550 VSS 0.018812f
C6220 VDPWR.t288 VSS 5.64e-19
C6221 VDPWR.t329 VSS 0.001513f
C6222 VDPWR.n551 VSS 0.006904f
C6223 VDPWR.n552 VSS 0.003647f
C6224 VDPWR.t683 VSS 0.004984f
C6225 VDPWR.n553 VSS 0.01361f
C6226 VDPWR.n554 VSS 0.010753f
C6227 VDPWR.n555 VSS 0.013967f
C6228 VDPWR.n556 VSS 0.008065f
C6229 VDPWR.n557 VSS 0.005888f
C6230 VDPWR.n558 VSS 0.004416f
C6231 VDPWR.n559 VSS 0.005354f
C6232 VDPWR.n560 VSS 0.006068f
C6233 VDPWR.n561 VSS 0.013691f
C6234 VDPWR.t28 VSS 0.014151f
C6235 VDPWR.n562 VSS 7.37e-19
C6236 VDPWR.n563 VSS 0.004416f
C6237 VDPWR.n564 VSS 0.00136f
C6238 VDPWR.t856 VSS 7.56e-19
C6239 VDPWR.t31 VSS 0.001148f
C6240 VDPWR.n565 VSS 0.001983f
C6241 VDPWR.n566 VSS 0.005856f
C6242 VDPWR.n567 VSS 0.003488f
C6243 VDPWR.t1261 VSS 0.020799f
C6244 VDPWR.n568 VSS 0.005184f
C6245 VDPWR.n569 VSS 0.003488f
C6246 VDPWR.t5 VSS 5.64e-19
C6247 VDPWR.t1034 VSS 0.001513f
C6248 VDPWR.n570 VSS 0.006904f
C6249 VDPWR.t1214 VSS 0.020799f
C6250 VDPWR.t1024 VSS 0.003047f
C6251 VDPWR.n571 VSS 0.009651f
C6252 VDPWR.n572 VSS 0.005344f
C6253 VDPWR.n573 VSS 0.002933f
C6254 VDPWR.t668 VSS 0.004984f
C6255 VDPWR.n574 VSS 0.004913f
C6256 VDPWR.n575 VSS 0.018812f
C6257 VDPWR.n576 VSS 0.008065f
C6258 VDPWR.n577 VSS 0.013967f
C6259 VDPWR.t1023 VSS 0.02849f
C6260 VDPWR.t1033 VSS 0.027547f
C6261 VDPWR.t667 VSS 0.020377f
C6262 VDPWR.t4 VSS 0.029245f
C6263 VDPWR.t971 VSS 0.02849f
C6264 VDPWR.t924 VSS 0.032453f
C6265 VDPWR.t30 VSS 0.023585f
C6266 VDPWR.t855 VSS 0.012641f
C6267 VDPWR.t979 VSS 0.005849f
C6268 VDPWR.t981 VSS 0.020566f
C6269 VDPWR.n578 VSS 0.026837f
C6270 VDPWR.t982 VSS 0.007137f
C6271 VDPWR.n579 VSS 0.002016f
C6272 VDPWR.n580 VSS 0.0024f
C6273 VDPWR.n581 VSS 0.018611f
C6274 VDPWR.n582 VSS 0.005471f
C6275 VDPWR.t669 VSS 0.004984f
C6276 VDPWR.n583 VSS 0.008777f
C6277 VDPWR.n584 VSS 0.010753f
C6278 VDPWR.n585 VSS 0.003648f
C6279 VDPWR.n586 VSS 0.02906f
C6280 VDPWR.n587 VSS 0.039529f
C6281 VDPWR.t700 VSS 0.004984f
C6282 VDPWR.n588 VSS 0.009746f
C6283 VDPWR.n589 VSS 0.018812f
C6284 VDPWR.n590 VSS 0.011593f
C6285 VDPWR.t944 VSS 0.007172f
C6286 VDPWR.n591 VSS 0.00838f
C6287 VDPWR.n592 VSS 0.003488f
C6288 VDPWR.n593 VSS 0.001519f
C6289 VDPWR.n594 VSS 0.001519f
C6290 VDPWR.n595 VSS 0.1025f
C6291 VDPWR.t517 VSS 0.004984f
C6292 VDPWR.n596 VSS 0.004913f
C6293 VDPWR.n597 VSS 0.005888f
C6294 VDPWR.t1205 VSS 0.020799f
C6295 VDPWR.n598 VSS 0.018812f
C6296 VDPWR.n599 VSS 0.003647f
C6297 VDPWR.t518 VSS 0.004984f
C6298 VDPWR.n600 VSS 0.01361f
C6299 VDPWR.n601 VSS 0.014953f
C6300 VDPWR.n602 VSS 0.011593f
C6301 VDPWR.n603 VSS 0.005888f
C6302 VDPWR.n604 VSS 0.004416f
C6303 VDPWR.n605 VSS 0.005604f
C6304 VDPWR.t58 VSS 0.007175f
C6305 VDPWR.n606 VSS 0.009278f
C6306 VDPWR.n607 VSS 0.003488f
C6307 VDPWR.n608 VSS 0.005888f
C6308 VDPWR.n609 VSS 0.004416f
C6309 VDPWR.t854 VSS 0.007172f
C6310 VDPWR.n610 VSS 0.00847f
C6311 VDPWR.t115 VSS 0.007175f
C6312 VDPWR.n611 VSS 0.009165f
C6313 VDPWR.n612 VSS 0.003488f
C6314 VDPWR.n613 VSS 0.005888f
C6315 VDPWR.n614 VSS 0.004416f
C6316 VDPWR.t117 VSS 0.007172f
C6317 VDPWR.n615 VSS 0.00847f
C6318 VDPWR.t953 VSS 0.007175f
C6319 VDPWR.n616 VSS 0.009165f
C6320 VDPWR.n617 VSS 0.001519f
C6321 VDPWR.n618 VSS 0.005888f
C6322 VDPWR.n619 VSS 0.004416f
C6323 VDPWR.n620 VSS 0.00224f
C6324 VDPWR.t699 VSS 0.064097f
C6325 VDPWR.t516 VSS 0.039378f
C6326 VDPWR.t57 VSS 0.016158f
C6327 VDPWR.t853 VSS 0.022364f
C6328 VDPWR.t114 VSS 0.016158f
C6329 VDPWR.t116 VSS 0.022364f
C6330 VDPWR.t952 VSS 0.016158f
C6331 VDPWR.t943 VSS 0.024184f
C6332 VDPWR.n621 VSS 0.026472f
C6333 VDPWR.n622 VSS 0.012237f
C6334 VDPWR.n623 VSS 0.005471f
C6335 VDPWR.t701 VSS 0.004984f
C6336 VDPWR.n624 VSS 0.008777f
C6337 VDPWR.n625 VSS 0.014953f
C6338 VDPWR.n626 VSS 0.002976f
C6339 VDPWR.n627 VSS 0.027044f
C6340 VDPWR.n628 VSS 0.026223f
C6341 VDPWR.n629 VSS 6.08e-19
C6342 VDPWR.t980 VSS 0.007136f
C6343 VDPWR.n630 VSS 0.013312f
C6344 VDPWR.t970 VSS 0.007172f
C6345 VDPWR.n631 VSS 0.008357f
C6346 VDPWR.t925 VSS 0.002363f
C6347 VDPWR.t29 VSS 0.006281f
C6348 VDPWR.n632 VSS 0.003563f
C6349 VDPWR.t972 VSS 0.007041f
C6350 VDPWR.n633 VSS 0.007429f
C6351 VDPWR.n634 VSS 0.009555f
C6352 VDPWR.n635 VSS 0.001258f
C6353 VDPWR.n636 VSS 0.005888f
C6354 VDPWR.n637 VSS 0.003488f
C6355 VDPWR.n638 VSS 0.002016f
C6356 VDPWR.n639 VSS 0.00224f
C6357 VDPWR.n640 VSS 0.012275f
C6358 VDPWR.n641 VSS 0.032875f
C6359 VDPWR.t788 VSS 0.006226f
C6360 VDPWR.t186 VSS 0.016226f
C6361 VDPWR.t184 VSS 0.018113f
C6362 VDPWR.t18 VSS 0.012641f
C6363 VDPWR.t910 VSS 0.023585f
C6364 VDPWR.t1164 VSS 0.033207f
C6365 VDPWR.t1162 VSS 0.016226f
C6366 VDPWR.t964 VSS 0.012641f
C6367 VDPWR.t287 VSS 0.029245f
C6368 VDPWR.t681 VSS 0.020377f
C6369 VDPWR.t328 VSS 0.027547f
C6370 VDPWR.t145 VSS 0.02849f
C6371 VDPWR.n642 VSS 0.019402f
C6372 VDPWR.n643 VSS 0.005637f
C6373 VDPWR.n644 VSS 0.003862f
C6374 VDPWR.n645 VSS 0.009272f
C6375 VDPWR.n646 VSS 0.002696f
C6376 VDPWR.n647 VSS 0.005888f
C6377 VDPWR.n648 VSS 0.004416f
C6378 VDPWR.n649 VSS 0.002625f
C6379 VDPWR.n650 VSS 0.008924f
C6380 VDPWR.n651 VSS 0.006148f
C6381 VDPWR.n652 VSS 0.004064f
C6382 VDPWR.n653 VSS 0.011493f
C6383 VDPWR.n654 VSS 0.0731f
C6384 VDPWR.n655 VSS 0.037381f
C6385 VDPWR.n656 VSS 0.117598f
C6386 VDPWR.n657 VSS 0.025894f
C6387 VDPWR.n658 VSS 0.035269f
C6388 VDPWR.n659 VSS 0.076656f
C6389 VDPWR.n660 VSS 0.247132f
C6390 VDPWR.n661 VSS 2.38e-19
C6391 VDPWR.n662 VSS 0.247132f
C6392 VDPWR.t763 VSS 0.356671f
C6393 VDPWR.t762 VSS 0.356671f
C6394 VDPWR.n663 VSS 0.055293f
C6395 VDPWR.n664 VSS 0.055474f
C6396 VDPWR.n665 VSS 0.344366f
C6397 VDPWR.n666 VSS 0.055474f
C6398 VDPWR.n667 VSS 0.114487f
C6399 VDPWR.n668 VSS 0.060635f
C6400 VDPWR.n669 VSS 0.018181f
C6401 VDPWR.n670 VSS 0.029454f
C6402 VDPWR.n671 VSS 0.073168f
C6403 VDPWR.n672 VSS 0.084539f
C6404 VDPWR.n673 VSS 0.035235f
C6405 VDPWR.n674 VSS 0.114487f
C6406 VDPWR.n675 VSS 0.00445f
C6407 VDPWR.n676 VSS 0.055474f
C6408 VDPWR.n677 VSS 0.055474f
C6409 VDPWR.n678 VSS 0.055293f
C6410 VDPWR.n679 VSS 0.076656f
C6411 VDPWR.n680 VSS 0.247132f
C6412 VDPWR.t281 VSS 0.356671f
C6413 VDPWR.n681 VSS 0.344366f
C6414 VDPWR.t282 VSS 0.356671f
C6415 VDPWR.n682 VSS 0.247132f
C6416 VDPWR.n683 VSS 0.002025f
C6417 VDPWR.n684 VSS 0.060694f
C6418 VDPWR.n685 VSS 0.018181f
C6419 VDPWR.n686 VSS 0.029169f
C6420 VDPWR.n687 VSS 0.067579f
C6421 VDPWR.n688 VSS 0.082325f
C6422 VDPWR.n689 VSS 0.035121f
C6423 VDPWR.n690 VSS 0.114487f
C6424 VDPWR.n691 VSS 0.004458f
C6425 VDPWR.n692 VSS 0.055474f
C6426 VDPWR.n693 VSS 0.055474f
C6427 VDPWR.n694 VSS 0.055293f
C6428 VDPWR.n695 VSS 0.076656f
C6429 VDPWR.n696 VSS 0.247132f
C6430 VDPWR.t760 VSS 0.356671f
C6431 VDPWR.n697 VSS 0.344366f
C6432 VDPWR.t761 VSS 0.356671f
C6433 VDPWR.n698 VSS 0.247132f
C6434 VDPWR.n699 VSS 0.002138f
C6435 VDPWR.n700 VSS 0.060694f
C6436 VDPWR.n701 VSS 0.018181f
C6437 VDPWR.n702 VSS 0.029169f
C6438 VDPWR.n703 VSS 0.064853f
C6439 VDPWR.n704 VSS 0.086053f
C6440 VDPWR.n705 VSS 0.035269f
C6441 VDPWR.n706 VSS 0.114487f
C6442 VDPWR.n707 VSS 0.055474f
C6443 VDPWR.n708 VSS 0.055474f
C6444 VDPWR.n709 VSS 0.055293f
C6445 VDPWR.n710 VSS 0.076656f
C6446 VDPWR.n711 VSS 0.247132f
C6447 VDPWR.t315 VSS 0.356671f
C6448 VDPWR.n712 VSS 0.344366f
C6449 VDPWR.t314 VSS 0.356671f
C6450 VDPWR.n713 VSS 0.247132f
C6451 VDPWR.n714 VSS 2.15e-19
C6452 VDPWR.n715 VSS 0.006257f
C6453 VDPWR.n716 VSS 0.060659f
C6454 VDPWR.n717 VSS 0.018181f
C6455 VDPWR.n718 VSS 0.029432f
C6456 VDPWR.n719 VSS 0.059483f
C6457 VDPWR.n720 VSS 0.358402f
C6458 VDPWR.n721 VSS 5.33642f
C6459 VDPWR.t373 VSS 0.120007f
C6460 VDPWR.t340 VSS 0.074568f
C6461 VDPWR.t822 VSS 0.019801f
C6462 VDPWR.t219 VSS 0.019801f
C6463 VDPWR.n722 VSS 0.047461f
C6464 VDPWR.n723 VSS 0.423604f
C6465 VDPWR.t344 VSS 0.07455f
C6466 VDPWR.t824 VSS 0.019801f
C6467 VDPWR.t820 VSS 0.019801f
C6468 VDPWR.n724 VSS 0.047461f
C6469 VDPWR.n725 VSS 0.413821f
C6470 VDPWR.t253 VSS 0.019801f
C6471 VDPWR.t342 VSS 0.019801f
C6472 VDPWR.n726 VSS 0.047461f
C6473 VDPWR.n727 VSS 0.158951f
C6474 VDPWR.n728 VSS 0.064745f
C6475 VDPWR.n729 VSS 0.023069f
C6476 VDPWR.n730 VSS 0.03559f
C6477 VDPWR.n731 VSS 0.03559f
C6478 VDPWR.n732 VSS 0.03559f
C6479 VDPWR.n733 VSS 0.034528f
C6480 VDPWR.n734 VSS 0.218283f
C6481 VDPWR.t339 VSS 0.209454f
C6482 VDPWR.t821 VSS 0.143241f
C6483 VDPWR.t218 VSS 0.143241f
C6484 VDPWR.t252 VSS 0.107431f
C6485 VDPWR.n735 VSS 0.071621f
C6486 VDPWR.t341 VSS 0.107431f
C6487 VDPWR.t823 VSS 0.143241f
C6488 VDPWR.t819 VSS 0.143241f
C6489 VDPWR.t343 VSS 0.209454f
C6490 VDPWR.n736 VSS 0.218283f
C6491 VDPWR.n737 VSS 0.034517f
C6492 VDPWR.n738 VSS 0.023068f
C6493 VDPWR.n739 VSS 0.302545f
C6494 VDPWR.n740 VSS 0.014605f
C6495 VDPWR.n741 VSS 0.02803f
C6496 VDPWR.n742 VSS 0.02803f
C6497 VDPWR.t372 VSS 0.269964f
C6498 VDPWR.n743 VSS 0.027307f
C6499 VDPWR.n745 VSS 0.207311f
C6500 VDPWR.n746 VSS 0.02803f
C6501 VDPWR.n748 VSS 0.207311f
C6502 VDPWR.n749 VSS 0.027294f
C6503 VDPWR.n750 VSS 0.014601f
C6504 VDPWR.n751 VSS 0.170811f
C6505 VDPWR.n752 VSS 0.317852f
C6506 VDPWR.n753 VSS 0.465132f
C6507 VDPWR.n754 VSS 0.951569f
C6508 VDPWR.n755 VSS 1.09773f
C6509 VDPWR.n756 VSS 4.26152f
C6510 VDPWR.n757 VSS 3.16295f
C6511 VDPWR.n758 VSS 1.27886f
C6512 VDPWR.n759 VSS 0.16157f
C6513 VDPWR.n760 VSS 0.035269f
C6514 VDPWR.n761 VSS 0.114487f
C6515 VDPWR.n762 VSS 0.055474f
C6516 VDPWR.n763 VSS 0.055474f
C6517 VDPWR.n764 VSS 0.055293f
C6518 VDPWR.n765 VSS 0.076656f
C6519 VDPWR.n766 VSS 0.247132f
C6520 VDPWR.t1012 VSS 0.356671f
C6521 VDPWR.n767 VSS 0.344366f
C6522 VDPWR.t118 VSS 0.356671f
C6523 VDPWR.n768 VSS 0.247132f
C6524 VDPWR.n769 VSS 2.15e-19
C6525 VDPWR.n770 VSS 0.348256f
C6526 VDPWR.n771 VSS 0.012843f
C6527 VDPWR.n772 VSS 0.003054f
C6528 VDPWR.n773 VSS 0.001579f
C6529 VDPWR.n774 VSS 0.001579f
C6530 VDPWR.n775 VSS 0.116061f
C6531 VDPWR.n776 VSS 0.281618f
C6532 VDPWR.n777 VSS 0.096641f
C6533 VDPWR.n778 VSS 0.219213f
C6534 VDPWR.n779 VSS 0.281574f
C6535 VDPWR.n780 VSS 0.060111f
C6536 VDPWR.n781 VSS 0.096641f
C6537 VDPWR.n782 VSS 0.107527f
C6538 VDPWR.n783 VSS 0.001579f
C6539 VDPWR.n784 VSS 0.003054f
C6540 VDPWR.n785 VSS 0.003054f
C6541 VDPWR.n786 VSS 0.001973f
C6542 VDPWR.n787 VSS 0.002048f
C6543 VDPWR.n788 VSS 5.48e-19
C6544 VDPWR.t871 VSS 0.003019f
C6545 VDPWR.n789 VSS 0.006163f
C6546 VDPWR.n790 VSS 0.00224f
C6547 VDPWR.t531 VSS 0.052075f
C6548 VDPWR.t78 VSS 0.028868f
C6549 VDPWR.t938 VSS 0.022453f
C6550 VDPWR.t542 VSS 0.029245f
C6551 VDPWR.t962 VSS 0.03434f
C6552 VDPWR.t757 VSS 0.022453f
C6553 VDPWR.t507 VSS 0.029245f
C6554 VDPWR.t471 VSS 0.031509f
C6555 VDPWR.t248 VSS 0.033585f
C6556 VDPWR.t1146 VSS 0.02283f
C6557 VDPWR.t38 VSS 0.041132f
C6558 VDPWR.t265 VSS 0.016604f
C6559 VDPWR.t874 VSS 0.010566f
C6560 VDPWR.t966 VSS 0.017358f
C6561 VDPWR.t128 VSS 0.055283f
C6562 VDPWR.t998 VSS 0.060189f
C6563 VDPWR.t627 VSS 0.020377f
C6564 VDPWR.t916 VSS 0.027547f
C6565 VDPWR.t868 VSS 0.02849f
C6566 VDPWR.n791 VSS 0.038158f
C6567 VDPWR.t628 VSS 0.004984f
C6568 VDPWR.n792 VSS 0.008777f
C6569 VDPWR.t869 VSS 0.003019f
C6570 VDPWR.t1198 VSS 0.036876f
C6571 VDPWR.n793 VSS 0.011929f
C6572 VDPWR.n794 VSS 0.004416f
C6573 VDPWR.t999 VSS 5.64e-19
C6574 VDPWR.t917 VSS 0.001513f
C6575 VDPWR.n795 VSS 0.006904f
C6576 VDPWR.n796 VSS 0.013967f
C6577 VDPWR.t129 VSS 0.007511f
C6578 VDPWR.n797 VSS 0.016861f
C6579 VDPWR.t629 VSS 0.004984f
C6580 VDPWR.n798 VSS 0.004829f
C6581 VDPWR.t875 VSS 0.001527f
C6582 VDPWR.t39 VSS 0.001527f
C6583 VDPWR.n799 VSS 0.003322f
C6584 VDPWR.n800 VSS 0.007816f
C6585 VDPWR.n801 VSS 0.002048f
C6586 VDPWR.n802 VSS 0.001973f
C6587 VDPWR.n803 VSS 0.001579f
C6588 VDPWR.n804 VSS 0.003054f
C6589 VDPWR.n805 VSS 0.001973f
C6590 VDPWR.n806 VSS 0.002949f
C6591 VDPWR.t266 VSS 0.007332f
C6592 VDPWR.n807 VSS 0.005407f
C6593 VDPWR.n808 VSS 0.001734f
C6594 VDPWR.n809 VSS 0.001472f
C6595 VDPWR.n810 VSS 0.001472f
C6596 VDPWR.n811 VSS 8.32e-19
C6597 VDPWR.n812 VSS 0.001599f
C6598 VDPWR.t1147 VSS 0.001372f
C6599 VDPWR.t249 VSS 0.002267f
C6600 VDPWR.n813 VSS 0.006267f
C6601 VDPWR.n814 VSS 0.008122f
C6602 VDPWR.t1259 VSS 0.029301f
C6603 VDPWR.n815 VSS 0.015457f
C6604 VDPWR.n816 VSS 0.003488f
C6605 VDPWR.t508 VSS 0.005024f
C6606 VDPWR.t1265 VSS 0.010664f
C6607 VDPWR.n818 VSS 0.027341f
C6608 VDPWR.t509 VSS 0.005024f
C6609 VDPWR.n819 VSS 0.013522f
C6610 VDPWR.t543 VSS 0.005019f
C6611 VDPWR.n820 VSS 0.002332f
C6612 VDPWR.t758 VSS 0.001527f
C6613 VDPWR.t963 VSS 0.001527f
C6614 VDPWR.n821 VSS 0.003322f
C6615 VDPWR.n822 VSS 0.011761f
C6616 VDPWR.t1245 VSS 0.03788f
C6617 VDPWR.n823 VSS 0.06464f
C6618 VDPWR.n824 VSS 0.019984f
C6619 VDPWR.t939 VSS 0.001527f
C6620 VDPWR.t79 VSS 0.001527f
C6621 VDPWR.n825 VSS 0.003322f
C6622 VDPWR.n826 VSS 0.021375f
C6623 VDPWR.n827 VSS 7.36e-19
C6624 VDPWR.n828 VSS 0.001973f
C6625 VDPWR.n829 VSS 0.002944f
C6626 VDPWR.t544 VSS 0.004984f
C6627 VDPWR.n830 VSS 0.008777f
C6628 VDPWR.n831 VSS 0.005471f
C6629 VDPWR.t532 VSS 0.005024f
C6630 VDPWR.t1248 VSS 0.010664f
C6631 VDPWR.n833 VSS 0.027341f
C6632 VDPWR.t533 VSS 0.005024f
C6633 VDPWR.n834 VSS 0.014893f
C6634 VDPWR.n835 VSS 0.002048f
C6635 VDPWR.t656 VSS 0.005024f
C6636 VDPWR.t1185 VSS 0.010664f
C6637 VDPWR.n837 VSS 0.027341f
C6638 VDPWR.t657 VSS 0.005024f
C6639 VDPWR.n838 VSS 0.014893f
C6640 VDPWR.n839 VSS 0.001973f
C6641 VDPWR.n840 VSS 0.002112f
C6642 VDPWR.n841 VSS 0.002885f
C6643 VDPWR.n842 VSS 0.001376f
C6644 VDPWR.n843 VSS 0.012553f
C6645 VDPWR.n844 VSS 0.002048f
C6646 VDPWR.n845 VSS 0.001472f
C6647 VDPWR.n846 VSS 0.001973f
C6648 VDPWR.n847 VSS 0.003054f
C6649 VDPWR.n848 VSS 0.002949f
C6650 VDPWR.n849 VSS 0.005152f
C6651 VDPWR.n850 VSS 0.002016f
C6652 VDPWR.n851 VSS 0.015457f
C6653 VDPWR.n852 VSS 0.012685f
C6654 VDPWR.n853 VSS 0.00224f
C6655 VDPWR.n854 VSS 0.006234f
C6656 VDPWR.n855 VSS 0.002016f
C6657 VDPWR.n856 VSS 0.00475f
C6658 VDPWR.t473 VSS 0.005064f
C6659 VDPWR.n857 VSS 0.007505f
C6660 VDPWR.n858 VSS 0.018913f
C6661 VDPWR.n859 VSS 0.020217f
C6662 VDPWR.n860 VSS 0.005888f
C6663 VDPWR.n861 VSS 0.004416f
C6664 VDPWR.n862 VSS 0.0024f
C6665 VDPWR.n863 VSS 0.039775f
C6666 VDPWR.t472 VSS 0.004984f
C6667 VDPWR.n864 VSS 0.008777f
C6668 VDPWR.n865 VSS 0.002829f
C6669 VDPWR.n866 VSS 0.002048f
C6670 VDPWR.n867 VSS 0.001472f
C6671 VDPWR.n868 VSS 0.001973f
C6672 VDPWR.n869 VSS 0.001579f
C6673 VDPWR.n870 VSS 0.128008f
C6674 VDPWR.n871 VSS 0.281618f
C6675 VDPWR.n872 VSS 0.128862f
C6676 VDPWR.n873 VSS 0.003404f
C6677 VDPWR.n874 VSS 0.00352f
C6678 VDPWR.n875 VSS 0.002757f
C6679 VDPWR.n876 VSS 0.001579f
C6680 VDPWR.n877 VSS 0.002944f
C6681 VDPWR.t1270 VSS 0.020799f
C6682 VDPWR.n878 VSS 0.015788f
C6683 VDPWR.t915 VSS 0.003019f
C6684 VDPWR.n879 VSS 0.012345f
C6685 VDPWR.n880 VSS 0.002048f
C6686 VDPWR.n881 VSS 0.001973f
C6687 VDPWR.n882 VSS 0.00352f
C6688 VDPWR.n883 VSS 0.001579f
C6689 VDPWR.t485 VSS 0.004984f
C6690 VDPWR.n884 VSS 0.004325f
C6691 VDPWR.n885 VSS 0.005471f
C6692 VDPWR.t426 VSS 0.052075f
C6693 VDPWR.t876 VSS 0.028868f
C6694 VDPWR.t967 VSS 0.019245f
C6695 VDPWR.t553 VSS 0.017547f
C6696 VDPWR.t392 VSS 0.024906f
C6697 VDPWR.t974 VSS 0.039811f
C6698 VDPWR.t9 VSS 0.009057f
C6699 VDPWR.t1015 VSS 0.016038f
C6700 VDPWR.t294 VSS 0.015849f
C6701 VDPWR.t334 VSS 0.017924f
C6702 VDPWR.t973 VSS 0.035472f
C6703 VDPWR.t250 VSS 0.019434f
C6704 VDPWR.t890 VSS 0.016038f
C6705 VDPWR.t338 VSS 0.024906f
C6706 VDPWR.t271 VSS 0.017924f
C6707 VDPWR.t333 VSS 0.017924f
C6708 VDPWR.t976 VSS 0.019434f
C6709 VDPWR.t864 VSS 0.015849f
C6710 VDPWR.t293 VSS 0.024906f
C6711 VDPWR.t862 VSS 0.021509f
C6712 VDPWR.t212 VSS 0.017924f
C6713 VDPWR.t336 VSS 0.030566f
C6714 VDPWR.t337 VSS 0.024906f
C6715 VDPWR.t36 VSS 0.021509f
C6716 VDPWR.t204 VSS 0.015849f
C6717 VDPWR.t214 VSS 0.039623f
C6718 VDPWR.t269 VSS 0.038868f
C6719 VDPWR.t991 VSS 0.015849f
C6720 VDPWR.t202 VSS 0.035472f
C6721 VDPWR.t1150 VSS 0.025094f
C6722 VDPWR.t1027 VSS 0.020566f
C6723 VDPWR.t730 VSS 0.015849f
C6724 VDPWR.t326 VSS 0.024151f
C6725 VDPWR.t771 VSS 0.023208f
C6726 VDPWR.n886 VSS 0.020611f
C6727 VDPWR.t327 VSS 0.0018f
C6728 VDPWR.t1028 VSS 0.0018f
C6729 VDPWR.n887 VSS 0.003918f
C6730 VDPWR.n888 VSS 0.004957f
C6731 VDPWR.t731 VSS 0.005024f
C6732 VDPWR.t1180 VSS 0.010664f
C6733 VDPWR.n890 VSS 0.027341f
C6734 VDPWR.t732 VSS 0.005024f
C6735 VDPWR.n891 VSS 0.014893f
C6736 VDPWR.t1151 VSS 0.00632f
C6737 VDPWR.n892 VSS 0.001133f
C6738 VDPWR.t203 VSS 0.0018f
C6739 VDPWR.t270 VSS 0.0018f
C6740 VDPWR.n893 VSS 0.004032f
C6741 VDPWR.n894 VSS 0.00519f
C6742 VDPWR.n895 VSS 0.004416f
C6743 VDPWR.t205 VSS 0.002834f
C6744 VDPWR.t215 VSS 0.0018f
C6745 VDPWR.t37 VSS 0.0018f
C6746 VDPWR.n896 VSS 0.004032f
C6747 VDPWR.n897 VSS 0.00519f
C6748 VDPWR.n898 VSS 0.004672f
C6749 VDPWR.t213 VSS 0.002834f
C6750 VDPWR.t863 VSS 0.00135f
C6751 VDPWR.t865 VSS 0.002785f
C6752 VDPWR.n899 VSS 0.00567f
C6753 VDPWR.n900 VSS 0.004406f
C6754 VDPWR.n901 VSS 0.002949f
C6755 VDPWR.n902 VSS 0.002112f
C6756 VDPWR.n903 VSS 0.003083f
C6757 VDPWR.n904 VSS 0.001973f
C6758 VDPWR.n905 VSS 0.001579f
C6759 VDPWR.n906 VSS 0.001973f
C6760 VDPWR.n907 VSS 0.002048f
C6761 VDPWR.n908 VSS 0.005888f
C6762 VDPWR.n909 VSS 0.002944f
C6763 VDPWR.n910 VSS 0.002048f
C6764 VDPWR.n911 VSS 0.001598f
C6765 VDPWR.n912 VSS 0.002085f
C6766 VDPWR.t272 VSS 0.00135f
C6767 VDPWR.t891 VSS 0.002785f
C6768 VDPWR.n913 VSS 0.00567f
C6769 VDPWR.n914 VSS 0.005888f
C6770 VDPWR.t251 VSS 0.002776f
C6771 VDPWR.t335 VSS 0.001152f
C6772 VDPWR.t1016 VSS 0.001152f
C6773 VDPWR.n915 VSS 0.002399f
C6774 VDPWR.n916 VSS 0.006924f
C6775 VDPWR.t10 VSS 0.002776f
C6776 VDPWR.t554 VSS 0.004984f
C6777 VDPWR.n917 VSS 0.008777f
C6778 VDPWR.n918 VSS 0.003488f
C6779 VDPWR.t1250 VSS 0.029301f
C6780 VDPWR.t975 VSS 0.001152f
C6781 VDPWR.t393 VSS 0.001152f
C6782 VDPWR.n919 VSS 0.002373f
C6783 VDPWR.n920 VSS 0.014953f
C6784 VDPWR.n921 VSS 7.36e-19
C6785 VDPWR.n922 VSS 0.001973f
C6786 VDPWR.n923 VSS 0.116061f
C6787 VDPWR.n924 VSS 0.003404f
C6788 VDPWR.n925 VSS 0.003083f
C6789 VDPWR.n926 VSS 0.00352f
C6790 VDPWR.n927 VSS 0.001973f
C6791 VDPWR.n928 VSS 0.002048f
C6792 VDPWR.n929 VSS 0.007329f
C6793 VDPWR.t676 VSS 0.005024f
C6794 VDPWR.t1190 VSS 0.010664f
C6795 VDPWR.n931 VSS 0.027341f
C6796 VDPWR.t677 VSS 0.005024f
C6797 VDPWR.n932 VSS 0.014893f
C6798 VDPWR.n933 VSS 0.005888f
C6799 VDPWR.t1247 VSS 0.029301f
C6800 VDPWR.n934 VSS 0.044937f
C6801 VDPWR.n935 VSS 0.005445f
C6802 VDPWR.t154 VSS 0.001152f
C6803 VDPWR.t391 VSS 0.001152f
C6804 VDPWR.n936 VSS 0.002373f
C6805 VDPWR.n937 VSS 0.008042f
C6806 VDPWR.n938 VSS 0.0048f
C6807 VDPWR.t978 VSS 0.002755f
C6808 VDPWR.t716 VSS 0.005483f
C6809 VDPWR.n939 VSS 0.00426f
C6810 VDPWR.n940 VSS 0.002944f
C6811 VDPWR.n941 VSS 0.001973f
C6812 VDPWR.n942 VSS 0.00352f
C6813 VDPWR.n943 VSS 0.116061f
C6814 VDPWR.n944 VSS 0.00352f
C6815 VDPWR.n945 VSS 0.002949f
C6816 VDPWR.n946 VSS 0.001579f
C6817 VDPWR.n947 VSS 0.002048f
C6818 VDPWR.n948 VSS 0.005687f
C6819 VDPWR.n949 VSS 0.005888f
C6820 VDPWR.t1178 VSS 0.072626f
C6821 VDPWR.n950 VSS 0.033923f
C6822 VDPWR.n951 VSS 0.005888f
C6823 VDPWR.t813 VSS 0.00281f
C6824 VDPWR.t811 VSS 0.0018f
C6825 VDPWR.t158 VSS 0.0018f
C6826 VDPWR.n952 VSS 0.004032f
C6827 VDPWR.n953 VSS 0.007616f
C6828 VDPWR.n954 VSS 0.01243f
C6829 VDPWR.n955 VSS 0.002048f
C6830 VDPWR.n956 VSS 0.001973f
C6831 VDPWR.n957 VSS 0.00352f
C6832 VDPWR.n958 VSS 0.001579f
C6833 VDPWR.n959 VSS 0.002048f
C6834 VDPWR.n960 VSS 0.002944f
C6835 VDPWR.t1236 VSS 0.020799f
C6836 VDPWR.n961 VSS 0.007141f
C6837 VDPWR.t796 VSS 0.007646f
C6838 VDPWR.n962 VSS 0.011292f
C6839 VDPWR.n963 VSS 0.005888f
C6840 VDPWR.t54 VSS 0.0018f
C6841 VDPWR.t378 VSS 0.0018f
C6842 VDPWR.n964 VSS 0.004032f
C6843 VDPWR.t380 VSS 0.002834f
C6844 VDPWR.n965 VSS 0.006409f
C6845 VDPWR.n966 VSS 0.005344f
C6846 VDPWR.n967 VSS 0.001099f
C6847 VDPWR.n968 VSS 0.002949f
C6848 VDPWR.n969 VSS 0.002763f
C6849 VDPWR.n970 VSS 0.00288f
C6850 VDPWR.n971 VSS 0.001579f
C6851 VDPWR.n972 VSS 0.00352f
C6852 VDPWR.n973 VSS 0.116061f
C6853 VDPWR.n974 VSS 0.128008f
C6854 VDPWR.n975 VSS 0.00352f
C6855 VDPWR.n976 VSS 0.002949f
C6856 VDPWR.n977 VSS 0.001973f
C6857 VDPWR.n978 VSS 0.001579f
C6858 VDPWR.t1149 VSS 0.001148f
C6859 VDPWR.t367 VSS -7.28e-19
C6860 VDPWR.n979 VSS 0.007328f
C6861 VDPWR.n980 VSS 0.005643f
C6862 VDPWR.t1135 VSS 0.002776f
C6863 VDPWR.n981 VSS 0.001349f
C6864 VDPWR.n982 VSS 0.001151f
C6865 VDPWR.t1105 VSS 0.001867f
C6866 VDPWR.t1107 VSS 0.001867f
C6867 VDPWR.n983 VSS 0.003854f
C6868 VDPWR.n984 VSS 0.001131f
C6869 VDPWR.n985 VSS 0.002048f
C6870 VDPWR.n986 VSS 0.001973f
C6871 VDPWR.n987 VSS 0.00352f
C6872 VDPWR.n988 VSS 0.116061f
C6873 VDPWR.n989 VSS 0.128008f
C6874 VDPWR.n990 VSS 0.00352f
C6875 VDPWR.n991 VSS 0.002949f
C6876 VDPWR.n992 VSS 0.001579f
C6877 VDPWR.n993 VSS 0.002048f
C6878 VDPWR.n994 VSS 0.002944f
C6879 VDPWR.t1043 VSS 0.001036f
C6880 VDPWR.t226 VSS 0.001036f
C6881 VDPWR.n995 VSS 0.002169f
C6882 VDPWR.t1129 VSS 0.001867f
C6883 VDPWR.t1103 VSS 0.001867f
C6884 VDPWR.n996 VSS 0.003854f
C6885 VDPWR.t1121 VSS 0.0018f
C6886 VDPWR.t1125 VSS 0.001867f
C6887 VDPWR.n997 VSS 0.003787f
C6888 VDPWR.n998 VSS 0.005527f
C6889 VDPWR.n999 VSS 0.004432f
C6890 VDPWR.t1131 VSS 0.001867f
C6891 VDPWR.t1123 VSS 0.001867f
C6892 VDPWR.n1000 VSS 0.003881f
C6893 VDPWR.n1001 VSS 0.006736f
C6894 VDPWR.n1002 VSS 0.005888f
C6895 VDPWR.t1119 VSS 0.00659f
C6896 VDPWR.n1003 VSS 0.008378f
C6897 VDPWR.n1004 VSS 0.005344f
C6898 VDPWR.t901 VSS 0.001527f
C6899 VDPWR.t955 VSS 0.001527f
C6900 VDPWR.n1005 VSS 0.003322f
C6901 VDPWR.n1006 VSS 0.019777f
C6902 VDPWR.n1007 VSS 0.001973f
C6903 VDPWR.n1008 VSS 0.00352f
C6904 VDPWR.n1009 VSS 0.140809f
C6905 VDPWR.n1010 VSS 0.167264f
C6906 VDPWR.n1011 VSS 0.281618f
C6907 VDPWR.n1012 VSS 0.116061f
C6908 VDPWR.n1013 VSS 0.003404f
C6909 VDPWR.n1014 VSS 0.00352f
C6910 VDPWR.n1015 VSS 0.002757f
C6911 VDPWR.n1016 VSS 0.001579f
C6912 VDPWR.n1017 VSS 0.002944f
C6913 VDPWR.t1273 VSS 0.020799f
C6914 VDPWR.n1018 VSS 0.021306f
C6915 VDPWR.t729 VSS 0.004984f
C6916 VDPWR.n1019 VSS 0.011445f
C6917 VDPWR.n1020 VSS 0.002048f
C6918 VDPWR.n1021 VSS 0.001973f
C6919 VDPWR.n1022 VSS 0.00352f
C6920 VDPWR.n1023 VSS 0.001579f
C6921 VDPWR.t583 VSS 0.052075f
C6922 VDPWR.t696 VSS 0.085094f
C6923 VDPWR.t1081 VSS 0.069434f
C6924 VDPWR.t589 VSS 0.016226f
C6925 VDPWR.t1077 VSS 0.018868f
C6926 VDPWR.t1055 VSS 0.032453f
C6927 VDPWR.t1083 VSS 0.032453f
C6928 VDPWR.t1059 VSS 0.032453f
C6929 VDPWR.t1057 VSS 0.032453f
C6930 VDPWR.t1085 VSS 0.032453f
C6931 VDPWR.t1079 VSS 0.025849f
C6932 VDPWR.t1063 VSS 0.022642f
C6933 VDPWR.t1073 VSS 0.032453f
C6934 VDPWR.t1069 VSS 0.032453f
C6935 VDPWR.t1065 VSS 0.032453f
C6936 VDPWR.t1075 VSS 0.032453f
C6937 VDPWR.t1071 VSS 0.027358f
C6938 VDPWR.t630 VSS 0.016226f
C6939 VDPWR.t1067 VSS 0.021321f
C6940 VDPWR.t1061 VSS 0.032453f
C6941 VDPWR.t1154 VSS 0.032453f
C6942 VDPWR.t779 VSS 0.032453f
C6943 VDPWR.t1152 VSS 0.032453f
C6944 VDPWR.t1156 VSS 0.022264f
C6945 VDPWR.n1024 VSS 0.037412f
C6946 VDPWR.n1025 VSS 0.008952f
C6947 VDPWR.n1026 VSS 0.002791f
C6948 VDPWR.n1027 VSS 0.005888f
C6949 VDPWR.t1157 VSS 0.006898f
C6950 VDPWR.n1028 VSS 0.006782f
C6951 VDPWR.t631 VSS 0.005483f
C6952 VDPWR.n1029 VSS 0.004139f
C6953 VDPWR.t1153 VSS 0.001867f
C6954 VDPWR.t780 VSS 0.001867f
C6955 VDPWR.n1030 VSS 0.004011f
C6956 VDPWR.t1216 VSS 0.073477f
C6957 VDPWR.n1031 VSS 0.030131f
C6958 VDPWR.n1032 VSS 0.005888f
C6959 VDPWR.t1155 VSS 0.001867f
C6960 VDPWR.t1062 VSS 0.001867f
C6961 VDPWR.n1033 VSS 0.004002f
C6962 VDPWR.n1034 VSS 0.008485f
C6963 VDPWR.t1068 VSS 0.001867f
C6964 VDPWR.t1072 VSS 0.001867f
C6965 VDPWR.n1035 VSS 0.003854f
C6966 VDPWR.n1036 VSS 0.005775f
C6967 VDPWR.n1037 VSS 0.002949f
C6968 VDPWR.t1076 VSS 0.001867f
C6969 VDPWR.t1066 VSS 0.001867f
C6970 VDPWR.n1038 VSS 0.003854f
C6971 VDPWR.n1039 VSS 0.008648f
C6972 VDPWR.t1070 VSS 0.001867f
C6973 VDPWR.t1074 VSS 0.001867f
C6974 VDPWR.n1040 VSS 0.003854f
C6975 VDPWR.n1041 VSS 0.008648f
C6976 VDPWR.n1042 VSS 0.002112f
C6977 VDPWR.n1043 VSS 0.003083f
C6978 VDPWR.n1044 VSS 0.001973f
C6979 VDPWR.n1045 VSS 0.00352f
C6980 VDPWR.n1046 VSS 0.116061f
C6981 VDPWR.n1047 VSS 0.001579f
C6982 VDPWR.n1048 VSS 0.001973f
C6983 VDPWR.n1049 VSS 0.005888f
C6984 VDPWR.t1064 VSS 0.001867f
C6985 VDPWR.t1080 VSS 0.0018f
C6986 VDPWR.n1050 VSS 0.003797f
C6987 VDPWR.t632 VSS 0.005483f
C6988 VDPWR.n1051 VSS 0.004291f
C6989 VDPWR.n1052 VSS 0.005694f
C6990 VDPWR.n1053 VSS 0.002048f
C6991 VDPWR.n1054 VSS 0.002944f
C6992 VDPWR.n1055 VSS 0.001504f
C6993 VDPWR.n1056 VSS 0.001321f
C6994 VDPWR.n1057 VSS 0.006783f
C6995 VDPWR.t1086 VSS 0.001867f
C6996 VDPWR.t1058 VSS 0.001867f
C6997 VDPWR.n1058 VSS 0.003854f
C6998 VDPWR.n1059 VSS 0.003782f
C6999 VDPWR.n1060 VSS 0.005888f
C7000 VDPWR.t1230 VSS 0.072626f
C7001 VDPWR.t1060 VSS 0.001867f
C7002 VDPWR.t1084 VSS 0.001867f
C7003 VDPWR.n1061 VSS 0.003854f
C7004 VDPWR.n1062 VSS 0.00661f
C7005 VDPWR.n1063 VSS 0.033913f
C7006 VDPWR.t1056 VSS 0.001867f
C7007 VDPWR.t1078 VSS 0.001867f
C7008 VDPWR.n1064 VSS 0.003854f
C7009 VDPWR.t1082 VSS 0.006558f
C7010 VDPWR.n1065 VSS 0.009583f
C7011 VDPWR.t697 VSS 0.004984f
C7012 VDPWR.n1066 VSS 0.006247f
C7013 VDPWR.n1067 VSS 0.005696f
C7014 VDPWR.t1284 VSS 0.020799f
C7015 VDPWR.n1068 VSS 0.021306f
C7016 VDPWR.t698 VSS 0.004984f
C7017 VDPWR.t584 VSS 0.005024f
C7018 VDPWR.t1234 VSS 0.010664f
C7019 VDPWR.n1070 VSS 0.027341f
C7020 VDPWR.t585 VSS 0.005024f
C7021 VDPWR.n1071 VSS 0.014893f
C7022 VDPWR.t692 VSS 0.005024f
C7023 VDPWR.t1167 VSS 0.010664f
C7024 VDPWR.n1073 VSS 0.027341f
C7025 VDPWR.t693 VSS 0.005024f
C7026 VDPWR.n1074 VSS 0.014893f
C7027 VDPWR.n1075 VSS 0.012551f
C7028 VDPWR.n1076 VSS 0.002949f
C7029 VDPWR.n1077 VSS 0.002048f
C7030 VDPWR.n1078 VSS 0.003083f
C7031 VDPWR.n1079 VSS 0.001973f
C7032 VDPWR.n1080 VSS 0.003404f
C7033 VDPWR.n1081 VSS 0.001579f
C7034 VDPWR.n1082 VSS 0.001973f
C7035 VDPWR.n1083 VSS 0.002944f
C7036 VDPWR.n1084 VSS 0.002048f
C7037 VDPWR.n1085 VSS 0.002112f
C7038 VDPWR.n1086 VSS 0.001376f
C7039 VDPWR.n1087 VSS 0.002885f
C7040 VDPWR.n1088 VSS 0.003083f
C7041 VDPWR.n1089 VSS 0.140809f
C7042 VDPWR.n1090 VSS 0.532156f
C7043 VDPWR.n1091 VSS 0.140809f
C7044 VDPWR.n1092 VSS 0.003404f
C7045 VDPWR.n1093 VSS 0.00352f
C7046 VDPWR.n1094 VSS 0.002949f
C7047 VDPWR.n1095 VSS 0.001579f
C7048 VDPWR.n1096 VSS 0.002048f
C7049 VDPWR.n1097 VSS 0.00288f
C7050 VDPWR.t425 VSS 0.001867f
C7051 VDPWR.t397 VSS 0.001867f
C7052 VDPWR.n1098 VSS 0.003854f
C7053 VDPWR.t1283 VSS 0.072626f
C7054 VDPWR.t411 VSS 0.001867f
C7055 VDPWR.t421 VSS 0.001867f
C7056 VDPWR.n1099 VSS 0.003854f
C7057 VDPWR.n1100 VSS 0.008648f
C7058 VDPWR.n1101 VSS 0.005888f
C7059 VDPWR.t257 VSS 0.001867f
C7060 VDPWR.t417 VSS 0.001867f
C7061 VDPWR.n1102 VSS 0.004002f
C7062 VDPWR.n1103 VSS 0.005793f
C7063 VDPWR.t255 VSS 0.006898f
C7064 VDPWR.n1104 VSS 0.006887f
C7065 VDPWR.n1105 VSS 0.005836f
C7066 VDPWR.t1240 VSS 0.020636f
C7067 VDPWR.n1106 VSS 0.010252f
C7068 VDPWR.n1107 VSS 0.003941f
C7069 VDPWR.t563 VSS 0.004984f
C7070 VDPWR.n1108 VSS 0.002657f
C7071 VDPWR.t525 VSS 0.066226f
C7072 VDPWR.t678 VSS 0.055472f
C7073 VDPWR.t556 VSS 0.092264f
C7074 VDPWR.t492 VSS 0.063962f
C7075 VDPWR.t640 VSS 0.109622f
C7076 VDPWR.t704 VSS 0.098679f
C7077 VDPWR.t727 VSS 0.063962f
C7078 VDPWR.t736 VSS 0.040566f
C7079 VDPWR.t418 VSS 0.048868f
C7080 VDPWR.t414 VSS 0.032453f
C7081 VDPWR.t404 VSS 0.032453f
C7082 VDPWR.t408 VSS 0.032453f
C7083 VDPWR.t406 VSS 0.022453f
C7084 VDPWR.t412 VSS 0.026226f
C7085 VDPWR.t402 VSS 0.032453f
C7086 VDPWR.t398 VSS 0.032264f
C7087 VDPWR.t394 VSS 0.032264f
C7088 VDPWR.t422 VSS 0.032453f
C7089 VDPWR.t400 VSS 0.023962f
C7090 VDPWR.t432 VSS 0.016226f
C7091 VDPWR.t396 VSS 0.024717f
C7092 VDPWR.t424 VSS 0.032453f
C7093 VDPWR.t420 VSS 0.032453f
C7094 VDPWR.t410 VSS 0.032453f
C7095 VDPWR.t416 VSS 0.032453f
C7096 VDPWR.t256 VSS 0.032453f
C7097 VDPWR.t258 VSS 0.02f
C7098 VDPWR.t1019 VSS 0.028679f
C7099 VDPWR.t254 VSS 0.016792f
C7100 VDPWR.t562 VSS 0.006038f
C7101 VDPWR.n1109 VSS 0.037412f
C7102 VDPWR.n1110 VSS 0.017118f
C7103 VDPWR.n1111 VSS 0.002949f
C7104 VDPWR.n1112 VSS 0.012758f
C7105 VDPWR.n1113 VSS 0.002048f
C7106 VDPWR.n1114 VSS 0.001579f
C7107 VDPWR.n1115 VSS 0.00352f
C7108 VDPWR.n1116 VSS 0.116061f
C7109 VDPWR.n1117 VSS 0.003404f
C7110 VDPWR.n1118 VSS 0.00352f
C7111 VDPWR.n1119 VSS 0.002949f
C7112 VDPWR.n1120 VSS 0.001579f
C7113 VDPWR.n1121 VSS 0.002048f
C7114 VDPWR.n1122 VSS 0.002048f
C7115 VDPWR.n1123 VSS 0.003083f
C7116 VDPWR.n1124 VSS 0.002949f
C7117 VDPWR.n1125 VSS 0.012758f
C7118 VDPWR.n1126 VSS 0.015948f
C7119 VDPWR.t547 VSS 0.005499f
C7120 VDPWR.n1127 VSS 0.016304f
C7121 VDPWR.n1128 VSS 0.009681f
C7122 VDPWR.n1129 VSS 0.005888f
C7123 VDPWR.n1130 VSS 0.010659f
C7124 VDPWR.n1131 VSS 0.015934f
C7125 VDPWR.t1271 VSS 0.072626f
C7126 VDPWR.n1132 VSS 0.03993f
C7127 VDPWR.t449 VSS 0.004984f
C7128 VDPWR.n1133 VSS 0.005908f
C7129 VDPWR.t665 VSS 0.005483f
C7130 VDPWR.n1134 VSS 0.006928f
C7131 VDPWR.n1135 VSS 0.002048f
C7132 VDPWR.n1136 VSS 0.001973f
C7133 VDPWR.n1137 VSS 0.001579f
C7134 VDPWR.n1138 VSS 0.001579f
C7135 VDPWR.n1139 VSS 0.001973f
C7136 VDPWR.n1140 VSS 0.002048f
C7137 VDPWR.n1141 VSS 0.005888f
C7138 VDPWR.t1172 VSS 0.072626f
C7139 VDPWR.n1142 VSS 0.012342f
C7140 VDPWR.n1143 VSS 0.002944f
C7141 VDPWR.n1144 VSS 0.002112f
C7142 VDPWR.n1145 VSS 0.001973f
C7143 VDPWR.n1146 VSS 0.00288f
C7144 VDPWR.n1147 VSS 0.002048f
C7145 VDPWR.n1148 VSS 0.012758f
C7146 VDPWR.n1149 VSS 0.009777f
C7147 VDPWR.n1150 VSS 0.036592f
C7148 VDPWR.n1151 VSS 0.005756f
C7149 VDPWR.n1152 VSS 0.005888f
C7150 VDPWR.t644 VSS 0.005483f
C7151 VDPWR.n1153 VSS 0.006928f
C7152 VDPWR.t1184 VSS 0.072626f
C7153 VDPWR.n1154 VSS 0.036175f
C7154 VDPWR.t666 VSS 0.005483f
C7155 VDPWR.n1155 VSS 0.003531f
C7156 VDPWR.t659 VSS 0.005483f
C7157 VDPWR.n1156 VSS 0.006928f
C7158 VDPWR.n1157 VSS 0.005888f
C7159 VDPWR.t1174 VSS 0.072626f
C7160 VDPWR.n1158 VSS 0.036592f
C7161 VDPWR.n1159 VSS 0.00224f
C7162 VDPWR.n1160 VSS 0.001973f
C7163 VDPWR.n1161 VSS 0.00352f
C7164 VDPWR.n1162 VSS 0.116061f
C7165 VDPWR.n1163 VSS 0.00352f
C7166 VDPWR.n1164 VSS 0.001973f
C7167 VDPWR.n1165 VSS 0.002048f
C7168 VDPWR.t441 VSS 0.066226f
C7169 VDPWR.t616 VSS 0.072641f
C7170 VDPWR.t477 VSS 0.109622f
C7171 VDPWR.t577 VSS 0.063962f
C7172 VDPWR.t559 VSS 0.109622f
C7173 VDPWR.t545 VSS 0.098679f
C7174 VDPWR.n1166 VSS 0.072506f
C7175 VDPWR.t447 VSS 0.086792f
C7176 VDPWR.t749 VSS 0.109622f
C7177 VDPWR.t664 VSS 0.098679f
C7178 VDPWR.t643 VSS 0.109622f
C7179 VDPWR.t658 VSS 0.098679f
C7180 VDPWR.t513 VSS 0.052075f
C7181 VDPWR.t47 VSS 0.046226f
C7182 VDPWR.t932 VSS 0.033019f
C7183 VDPWR.t759 VSS 0.017358f
C7184 VDPWR.t605 VSS 0.006604f
C7185 VDPWR.t994 VSS 0.047358f
C7186 VDPWR.t992 VSS 0.038302f
C7187 VDPWR.t996 VSS 0.012264f
C7188 VDPWR.t934 VSS 0.021509f
C7189 VDPWR.t132 VSS 0.015849f
C7190 VDPWR.t1017 VSS 0.015849f
C7191 VDPWR.t135 VSS 0.017547f
C7192 VDPWR.t44 VSS 0.017924f
C7193 VDPWR.t65 VSS 0.017924f
C7194 VDPWR.t94 VSS 0.024906f
C7195 VDPWR.t1002 VSS 0.023208f
C7196 VDPWR.t1004 VSS 0.013019f
C7197 VDPWR.t134 VSS 0.017924f
C7198 VDPWR.t346 VSS 0.017924f
C7199 VDPWR.t133 VSS 0.015849f
C7200 VDPWR.t348 VSS 0.016038f
C7201 VDPWR.t918 VSS 0.023396f
C7202 VDPWR.t6 VSS 0.01283f
C7203 VDPWR.t136 VSS 0.013585f
C7204 VDPWR.t102 VSS 0.015849f
C7205 VDPWR.t1013 VSS 0.008868f
C7206 VDPWR.t739 VSS 0.072641f
C7207 VDPWR.n1167 VSS 0.060619f
C7208 VDPWR.n1168 VSS 0.009361f
C7209 VDPWR.n1169 VSS 0.002048f
C7210 VDPWR.n1170 VSS 0.001579f
C7211 VDPWR.n1171 VSS 0.001579f
C7212 VDPWR.n1172 VSS 0.001973f
C7213 VDPWR.n1173 VSS 0.002944f
C7214 VDPWR.n1174 VSS 0.002944f
C7215 VDPWR.n1175 VSS 0.002048f
C7216 VDPWR.n1176 VSS 0.012342f
C7217 VDPWR.t645 VSS 0.005483f
C7218 VDPWR.n1177 VSS 0.006928f
C7219 VDPWR.n1178 VSS 0.006017f
C7220 VDPWR.t740 VSS 0.004984f
C7221 VDPWR.n1179 VSS 0.006247f
C7222 VDPWR.n1180 VSS 0.005888f
C7223 VDPWR.t1275 VSS 0.020799f
C7224 VDPWR.n1181 VSS 0.021306f
C7225 VDPWR.t741 VSS 0.004984f
C7226 VDPWR.t103 VSS 0.007187f
C7227 VDPWR.n1182 VSS 0.012163f
C7228 VDPWR.n1183 VSS 0.003456f
C7229 VDPWR.t919 VSS 0.002754f
C7230 VDPWR.t349 VSS 0.006295f
C7231 VDPWR.n1184 VSS 0.005479f
C7232 VDPWR.n1185 VSS 0.004672f
C7233 VDPWR.n1186 VSS 0.001598f
C7234 VDPWR.n1187 VSS 0.002949f
C7235 VDPWR.n1188 VSS 0.003083f
C7236 VDPWR.n1189 VSS 0.001973f
C7237 VDPWR.n1190 VSS 0.00352f
C7238 VDPWR.n1191 VSS 0.140809f
C7239 VDPWR.n1192 VSS 0.281618f
C7240 VDPWR.n1193 VSS 0.116061f
C7241 VDPWR.n1194 VSS 0.003404f
C7242 VDPWR.n1195 VSS 0.003083f
C7243 VDPWR.n1196 VSS 0.00352f
C7244 VDPWR.n1197 VSS 0.001973f
C7245 VDPWR.n1198 VSS 0.002048f
C7246 VDPWR.t747 VSS 0.004984f
C7247 VDPWR.t1166 VSS 0.020982f
C7248 VDPWR.n1200 VSS 0.036453f
C7249 VDPWR.t748 VSS 0.004984f
C7250 VDPWR.n1201 VSS 0.020917f
C7251 VDPWR.t614 VSS 0.004984f
C7252 VDPWR.t1237 VSS 0.020982f
C7253 VDPWR.n1203 VSS 0.036453f
C7254 VDPWR.t615 VSS 0.004984f
C7255 VDPWR.n1204 VSS 0.020917f
C7256 VDPWR.n1205 VSS 0.018023f
C7257 VDPWR.t742 VSS 0.005024f
C7258 VDPWR.t1220 VSS 0.010664f
C7259 VDPWR.n1207 VSS 0.027341f
C7260 VDPWR.t743 VSS 0.005024f
C7261 VDPWR.n1208 VSS 0.014893f
C7262 VDPWR.n1209 VSS 0.001133f
C7263 VDPWR.n1210 VSS 0.005888f
C7264 VDPWR.t43 VSS 0.00632f
C7265 VDPWR.n1211 VSS 0.002085f
C7266 VDPWR.n1212 VSS 0.002405f
C7267 VDPWR.t455 VSS 0.005483f
C7268 VDPWR.n1213 VSS 0.002283f
C7269 VDPWR.n1214 VSS 0.002048f
C7270 VDPWR.n1215 VSS 0.001579f
C7271 VDPWR.n1216 VSS 0.001579f
C7272 VDPWR.n1217 VSS 0.002949f
C7273 VDPWR.n1218 VSS 0.007422f
C7274 VDPWR.n1219 VSS 0.005888f
C7275 VDPWR.t175 VSS 0.002754f
C7276 VDPWR.t826 VSS 0.001152f
C7277 VDPWR.t164 VSS 0.001152f
C7278 VDPWR.n1220 VSS 0.002373f
C7279 VDPWR.n1221 VSS 0.006065f
C7280 VDPWR.t454 VSS 0.0055f
C7281 VDPWR.t746 VSS 0.005055f
C7282 VDPWR.n1222 VSS 0.035589f
C7283 VDPWR.t602 VSS 0.052075f
C7284 VDPWR.t613 VSS 0.069811f
C7285 VDPWR.t46 VSS 0.014151f
C7286 VDPWR.t0 VSS 0.015849f
C7287 VDPWR.t940 VSS 0.015849f
C7288 VDPWR.t906 VSS 0.015849f
C7289 VDPWR.t936 VSS 0.031321f
C7290 VDPWR.t42 VSS 0.024151f
C7291 VDPWR.t2 VSS 0.029811f
C7292 VDPWR.t25 VSS 0.02717f
C7293 VDPWR.t857 VSS 0.015849f
C7294 VDPWR.t166 VSS 0.024717f
C7295 VDPWR.t26 VSS 0.028302f
C7296 VDPWR.t168 VSS 0.04434f
C7297 VDPWR.t165 VSS 0.037358f
C7298 VDPWR.t24 VSS 0.033962f
C7299 VDPWR.t174 VSS 0.033019f
C7300 VDPWR.t453 VSS 0.035472f
C7301 VDPWR.t163 VSS 0.03434f
C7302 VDPWR.t825 VSS 0.021698f
C7303 VDPWR.t744 VSS 0.052075f
C7304 VDPWR.n1223 VSS 0.037789f
C7305 VDPWR.n1224 VSS 0.006017f
C7306 VDPWR.n1225 VSS 0.002048f
C7307 VDPWR.n1226 VSS 0.001973f
C7308 VDPWR.n1227 VSS 0.00352f
C7309 VDPWR.n1228 VSS 0.116061f
C7310 VDPWR.n1229 VSS 0.00352f
C7311 VDPWR.n1230 VSS 0.002757f
C7312 VDPWR.n1231 VSS 0.001579f
C7313 VDPWR.n1232 VSS 0.001579f
C7314 VDPWR.n1233 VSS 0.001973f
C7315 VDPWR.n1234 VSS 0.002944f
C7316 VDPWR.n1235 VSS 0.012758f
C7317 VDPWR.n1236 VSS 0.005888f
C7318 VDPWR.t1177 VSS 0.072626f
C7319 VDPWR.t1223 VSS 0.072626f
C7320 VDPWR.n1237 VSS 0.036592f
C7321 VDPWR.n1238 VSS 0.005344f
C7322 VDPWR.t612 VSS 0.005501f
C7323 VDPWR.n1239 VSS 0.011251f
C7324 VDPWR.n1240 VSS 0.005888f
C7325 VDPWR.n1241 VSS 0.012758f
C7326 VDPWR.n1242 VSS 0.002048f
C7327 VDPWR.n1243 VSS 0.001973f
C7328 VDPWR.n1244 VSS 0.00352f
C7329 VDPWR.n1245 VSS 0.116061f
C7330 VDPWR.n1246 VSS 0.116061f
C7331 VDPWR.n1247 VSS 0.00352f
C7332 VDPWR.n1248 VSS 0.002949f
C7333 VDPWR.n1249 VSS 0.001579f
C7334 VDPWR.n1250 VSS 0.002048f
C7335 VDPWR.n1251 VSS 0.002112f
C7336 VDPWR.n1252 VSS 0.001579f
C7337 VDPWR.n1253 VSS 0.001973f
C7338 VDPWR.n1254 VSS 0.00288f
C7339 VDPWR.t1235 VSS 0.072626f
C7340 VDPWR.n1255 VSS 0.009361f
C7341 VDPWR.n1256 VSS 0.004416f
C7342 VDPWR.t726 VSS 0.005059f
C7343 VDPWR.n1257 VSS 0.01476f
C7344 VDPWR.n1258 VSS 0.015674f
C7345 VDPWR.t1189 VSS 0.021124f
C7346 VDPWR.n1259 VSS 0.020912f
C7347 VDPWR.t725 VSS 0.004984f
C7348 VDPWR.n1260 VSS 0.005999f
C7349 VDPWR.n1261 VSS 0.006f
C7350 VDPWR.t536 VSS 0.066226f
C7351 VDPWR.t519 VSS 0.072641f
C7352 VDPWR.t717 VSS 0.109622f
C7353 VDPWR.t580 VSS 0.063962f
C7354 VDPWR.t468 VSS 0.109622f
C7355 VDPWR.t550 VSS 0.098679f
C7356 VDPWR.t574 VSS 0.098679f
C7357 VDPWR.t650 VSS 0.109622f
C7358 VDPWR.t610 VSS 0.098679f
C7359 VDPWR.t752 VSS 0.109622f
C7360 VDPWR.t724 VSS 0.034717f
C7361 VDPWR.n1262 VSS 0.037412f
C7362 VDPWR.n1263 VSS 0.006017f
C7363 VDPWR.n1264 VSS 0.002048f
C7364 VDPWR.n1265 VSS 0.001973f
C7365 VDPWR.n1266 VSS 0.00352f
C7366 VDPWR.n1267 VSS 0.116061f
C7367 VDPWR.n1268 VSS 0.00352f
C7368 VDPWR.n1269 VSS 0.002949f
C7369 VDPWR.n1270 VSS 0.001579f
C7370 VDPWR.n1271 VSS 0.002048f
C7371 VDPWR.n1272 VSS 0.002944f
C7372 VDPWR.t1260 VSS 0.072626f
C7373 VDPWR.n1273 VSS 0.012758f
C7374 VDPWR.n1274 VSS 0.005344f
C7375 VDPWR.t1286 VSS 0.074001f
C7376 VDPWR.t582 VSS 0.005483f
C7377 VDPWR.n1275 VSS 0.006928f
C7378 VDPWR.n1276 VSS 0.005888f
C7379 VDPWR.n1277 VSS 0.008742f
C7380 VDPWR.n1278 VSS 0.005888f
C7381 VDPWR.t1246 VSS 0.072626f
C7382 VDPWR.n1279 VSS 0.040608f
C7383 VDPWR.n1280 VSS 0.00288f
C7384 VDPWR.n1281 VSS 0.001973f
C7385 VDPWR.n1282 VSS 0.00352f
C7386 VDPWR.n1283 VSS 0.155317f
C7387 VDPWR.n1284 VSS 0.167264f
C7388 VDPWR.n1285 VSS 0.003404f
C7389 VDPWR.n1286 VSS 0.00352f
C7390 VDPWR.n1287 VSS 0.001477f
C7391 VDPWR.n1288 VSS 0.001579f
C7392 VDPWR.n1289 VSS 0.002048f
C7393 VDPWR.n1290 VSS 0.003083f
C7394 VDPWR.t1088 VSS 0.001527f
C7395 VDPWR.t41 VSS 0.001527f
C7396 VDPWR.n1291 VSS 0.003322f
C7397 VDPWR.t686 VSS 0.004984f
C7398 VDPWR.n1292 VSS 0.011445f
C7399 VDPWR.n1293 VSS 0.005888f
C7400 VDPWR.n1294 VSS 0.015256f
C7401 VDPWR.n1295 VSS 0.005888f
C7402 VDPWR.t1171 VSS 0.036876f
C7403 VDPWR.t654 VSS 0.005483f
C7404 VDPWR.n1296 VSS 0.003947f
C7405 VDPWR.n1297 VSS 0.022156f
C7406 VDPWR.n1298 VSS 0.002048f
C7407 VDPWR.n1299 VSS 0.001973f
C7408 VDPWR.n1300 VSS 0.00352f
C7409 VDPWR.n1301 VSS 0.00352f
C7410 VDPWR.n1302 VSS 0.002757f
C7411 VDPWR.n1303 VSS 0.001579f
C7412 VDPWR.n1304 VSS 0.001579f
C7413 VDPWR.n1305 VSS 0.001973f
C7414 VDPWR.n1306 VSS 0.002944f
C7415 VDPWR.n1307 VSS 0.012758f
C7416 VDPWR.n1308 VSS 0.005888f
C7417 VDPWR.t1191 VSS 0.072626f
C7418 VDPWR.t1168 VSS 0.072626f
C7419 VDPWR.n1309 VSS 0.066804f
C7420 VDPWR.n1310 VSS 0.005888f
C7421 VDPWR.t466 VSS 0.005483f
C7422 VDPWR.t622 VSS 0.005483f
C7423 VDPWR.n1311 VSS 0.007477f
C7424 VDPWR.t567 VSS 0.005483f
C7425 VDPWR.t710 VSS 0.005483f
C7426 VDPWR.n1312 VSS 0.007477f
C7427 VDPWR.n1313 VSS 0.003904f
C7428 VDPWR.n1314 VSS 0.012758f
C7429 VDPWR.n1315 VSS 0.002112f
C7430 VDPWR.n1316 VSS 0.001973f
C7431 VDPWR.n1317 VSS 0.00352f
C7432 VDPWR.n1318 VSS 0.00352f
C7433 VDPWR.n1319 VSS 0.002949f
C7434 VDPWR.n1320 VSS 0.001579f
C7435 VDPWR.n1321 VSS 0.009361f
C7436 VDPWR.n1322 VSS 0.005888f
C7437 VDPWR.t566 VSS 0.005483f
C7438 VDPWR.t709 VSS 0.005483f
C7439 VDPWR.n1323 VSS 0.007477f
C7440 VDPWR.t487 VSS 0.005024f
C7441 VDPWR.t1244 VSS 0.010664f
C7442 VDPWR.n1325 VSS 0.027341f
C7443 VDPWR.t488 VSS 0.005024f
C7444 VDPWR.n1326 VSS 0.014893f
C7445 VDPWR.t675 VSS 0.005499f
C7446 VDPWR.n1327 VSS 0.016304f
C7447 VDPWR.t621 VSS 0.005483f
C7448 VDPWR.n1328 VSS 0.006928f
C7449 VDPWR.n1329 VSS 0.002048f
C7450 VDPWR.n1330 VSS 0.001973f
C7451 VDPWR.n1331 VSS 0.00352f
C7452 VDPWR.n1332 VSS 0.00352f
C7453 VDPWR.n1333 VSS 0.002949f
C7454 VDPWR.n1334 VSS 0.001579f
C7455 VDPWR.n1335 VSS 0.002048f
C7456 VDPWR.n1336 VSS 0.002944f
C7457 VDPWR.t1213 VSS 0.072626f
C7458 VDPWR.n1337 VSS 0.012758f
C7459 VDPWR.n1338 VSS 0.005344f
C7460 VDPWR.t1192 VSS 0.074001f
C7461 VDPWR.t524 VSS 0.005483f
C7462 VDPWR.n1339 VSS 0.006928f
C7463 VDPWR.n1340 VSS 0.005888f
C7464 VDPWR.n1341 VSS 0.008742f
C7465 VDPWR.n1342 VSS 0.005888f
C7466 VDPWR.t1272 VSS 0.072626f
C7467 VDPWR.n1343 VSS 0.040608f
C7468 VDPWR.n1344 VSS 0.00288f
C7469 VDPWR.n1345 VSS 0.001973f
C7470 VDPWR.n1346 VSS 0.00352f
C7471 VDPWR.n1347 VSS 0.001579f
C7472 VDPWR.n1348 VSS 0.002048f
C7473 VDPWR.t1239 VSS 0.036234f
C7474 VDPWR.n1349 VSS 0.027337f
C7475 VDPWR.t523 VSS 0.005483f
C7476 VDPWR.t505 VSS 0.004984f
C7477 VDPWR.n1350 VSS 0.011995f
C7478 VDPWR.t457 VSS 0.005024f
C7479 VDPWR.t1258 VSS 0.010664f
C7480 VDPWR.n1352 VSS 0.027341f
C7481 VDPWR.t458 VSS 0.005024f
C7482 VDPWR.n1353 VSS 0.014893f
C7483 VDPWR.t646 VSS 0.005024f
C7484 VDPWR.t1225 VSS 0.010664f
C7485 VDPWR.n1355 VSS 0.027341f
C7486 VDPWR.t647 VSS 0.005024f
C7487 VDPWR.n1356 VSS 0.014893f
C7488 VDPWR.n1357 VSS 0.01227f
C7489 VDPWR.t430 VSS 0.005024f
C7490 VDPWR.t1262 VSS 0.010664f
C7491 VDPWR.n1359 VSS 0.027341f
C7492 VDPWR.t431 VSS 0.005024f
C7493 VDPWR.n1360 VSS 0.014893f
C7494 VDPWR.n1361 VSS 0.003844f
C7495 VDPWR.n1362 VSS 0.004957f
C7496 VDPWR.t633 VSS 0.005024f
C7497 VDPWR.t1233 VSS 0.010664f
C7498 VDPWR.n1364 VSS 0.027341f
C7499 VDPWR.t634 VSS 0.005024f
C7500 VDPWR.n1365 VSS 0.014893f
C7501 VDPWR.n1366 VSS 0.013462f
C7502 VDPWR.n1367 VSS 0.00331f
C7503 VDPWR.n1368 VSS 0.003842f
C7504 VDPWR.n1369 VSS 0.004416f
C7505 VDPWR.n1370 VSS 0.002368f
C7506 VDPWR.n1371 VSS 0.001973f
C7507 VDPWR.n1372 VSS 0.003404f
C7508 VDPWR.n1373 VSS 0.003083f
C7509 VDPWR.n1374 VSS 0.002629f
C7510 VDPWR.n1375 VSS 0.00352f
C7511 VDPWR.n1376 VSS 0.015256f
C7512 VDPWR.n1377 VSS 0.025685f
C7513 VDPWR.n1378 VSS 0.015256f
C7514 VDPWR.n1379 VSS 0.015934f
C7515 VDPWR.n1380 VSS 0.002048f
C7516 VDPWR.n1381 VSS 0.002944f
C7517 VDPWR.n1382 VSS 0.001973f
C7518 VDPWR.n1383 VSS 0.001579f
C7519 VDPWR.n1384 VSS 0.00352f
C7520 VDPWR.n1385 VSS 0.003404f
C7521 VDPWR.n1386 VSS 0.003083f
C7522 VDPWR.n1387 VSS 0.002117f
C7523 VDPWR.n1388 VSS 0.003008f
C7524 VDPWR.n1389 VSS 0.015256f
C7525 VDPWR.n1390 VSS 0.020793f
C7526 VDPWR.t506 VSS 0.004984f
C7527 VDPWR.n1391 VSS 0.011445f
C7528 VDPWR.n1392 VSS 0.020115f
C7529 VDPWR.n1393 VSS 0.005888f
C7530 VDPWR.n1394 VSS 0.003488f
C7531 VDPWR.n1395 VSS 0.004416f
C7532 VDPWR.n1396 VSS 0.005612f
C7533 VDPWR.t620 VSS 0.005483f
C7534 VDPWR.n1397 VSS 0.006928f
C7535 VDPWR.n1398 VSS 0.012342f
C7536 VDPWR.n1399 VSS 0.012342f
C7537 VDPWR.n1400 VSS 0.005888f
C7538 VDPWR.n1401 VSS 0.003488f
C7539 VDPWR.n1402 VSS 0.003209f
C7540 VDPWR.n1403 VSS 0.034322f
C7541 VDPWR.n1404 VSS 0.002865f
C7542 VDPWR.t674 VSS 0.005483f
C7543 VDPWR.n1405 VSS 0.006928f
C7544 VDPWR.n1406 VSS 0.012342f
C7545 VDPWR.n1407 VSS 0.005888f
C7546 VDPWR.n1408 VSS 0.005888f
C7547 VDPWR.n1409 VSS 0.004544f
C7548 VDPWR.n1410 VSS 0.009777f
C7549 VDPWR.n1411 VSS 0.036592f
C7550 VDPWR.n1412 VSS 0.009361f
C7551 VDPWR.n1413 VSS 0.012342f
C7552 VDPWR.n1414 VSS 0.012758f
C7553 VDPWR.n1415 VSS 0.002048f
C7554 VDPWR.n1416 VSS 0.001579f
C7555 VDPWR.n1417 VSS 0.001973f
C7556 VDPWR.n1418 VSS 0.00224f
C7557 VDPWR.n1419 VSS 0.002752f
C7558 VDPWR.n1420 VSS 0.001973f
C7559 VDPWR.n1421 VSS 0.003083f
C7560 VDPWR.n1422 VSS 0.003404f
C7561 VDPWR.n1423 VSS 0.155317f
C7562 VDPWR.n1424 VSS 0.003404f
C7563 VDPWR.n1425 VSS 0.003083f
C7564 VDPWR.n1426 VSS 0.002949f
C7565 VDPWR.n1427 VSS 0.002528f
C7566 VDPWR.n1428 VSS 0.006017f
C7567 VDPWR.t456 VSS 0.066226f
C7568 VDPWR.t429 VSS 0.072641f
C7569 VDPWR.t504 VSS 0.109622f
C7570 VDPWR.t522 VSS 0.063962f
C7571 VDPWR.t619 VSS 0.109622f
C7572 VDPWR.t673 VSS 0.098679f
C7573 VDPWR.t450 VSS 0.052075f
C7574 VDPWR.t459 VSS 0.208301f
C7575 VDPWR.t40 VSS 0.028868f
C7576 VDPWR.t1087 VSS 0.022453f
C7577 VDPWR.t653 VSS 0.063962f
C7578 VDPWR.t684 VSS 0.092075f
C7579 VDPWR.n1429 VSS 0.040844f
C7580 VDPWR.t465 VSS 0.208301f
C7581 VDPWR.t565 VSS 0.208301f
C7582 VDPWR.t486 VSS 0.055283f
C7583 VDPWR.n1430 VSS 0.05194f
C7584 VDPWR.n1431 VSS 0.015948f
C7585 VDPWR.n1432 VSS 0.003168f
C7586 VDPWR.n1433 VSS 0.004953f
C7587 VDPWR.n1434 VSS 0.010348f
C7588 VDPWR.n1435 VSS 0.004425f
C7589 VDPWR.n1436 VSS 0.004416f
C7590 VDPWR.n1437 VSS 0.005888f
C7591 VDPWR.n1438 VSS 0.012342f
C7592 VDPWR.n1439 VSS 0.012758f
C7593 VDPWR.t1281 VSS 0.072626f
C7594 VDPWR.t1252 VSS 0.072626f
C7595 VDPWR.n1440 VSS 0.066804f
C7596 VDPWR.n1441 VSS 0.009777f
C7597 VDPWR.n1442 VSS 0.005888f
C7598 VDPWR.n1443 VSS 0.005888f
C7599 VDPWR.n1444 VSS 0.005568f
C7600 VDPWR.n1445 VSS 0.012758f
C7601 VDPWR.n1446 VSS 0.012758f
C7602 VDPWR.n1447 VSS 0.002048f
C7603 VDPWR.n1448 VSS 0.001579f
C7604 VDPWR.n1449 VSS 0.001973f
C7605 VDPWR.n1450 VSS 0.00288f
C7606 VDPWR.n1451 VSS 0.002048f
C7607 VDPWR.n1452 VSS 0.002944f
C7608 VDPWR.n1453 VSS 0.001973f
C7609 VDPWR.n1454 VSS 0.003083f
C7610 VDPWR.n1455 VSS 0.003404f
C7611 VDPWR.n1456 VSS 0.155317f
C7612 VDPWR.n1457 VSS 0.003404f
C7613 VDPWR.n1458 VSS 0.003083f
C7614 VDPWR.n1459 VSS 0.002949f
C7615 VDPWR.n1460 VSS 0.002048f
C7616 VDPWR.n1461 VSS 0.012758f
C7617 VDPWR.n1462 VSS 0.012758f
C7618 VDPWR.n1463 VSS 0.012342f
C7619 VDPWR.n1464 VSS 0.005888f
C7620 VDPWR.n1465 VSS 0.004818f
C7621 VDPWR.n1466 VSS 0.004712f
C7622 VDPWR.n1467 VSS 0.005344f
C7623 VDPWR.n1468 VSS 0.005888f
C7624 VDPWR.n1469 VSS 0.012342f
C7625 VDPWR.n1470 VSS 0.012758f
C7626 VDPWR.n1471 VSS 0.009777f
C7627 VDPWR.n1472 VSS 0.005888f
C7628 VDPWR.n1473 VSS 0.005888f
C7629 VDPWR.n1474 VSS 0.009361f
C7630 VDPWR.n1475 VSS 0.012758f
C7631 VDPWR.n1476 VSS 0.012758f
C7632 VDPWR.n1477 VSS 0.005888f
C7633 VDPWR.n1478 VSS 0.005888f
C7634 VDPWR.n1479 VSS 0.003648f
C7635 VDPWR.n1480 VSS 0.012758f
C7636 VDPWR.t467 VSS 0.005483f
C7637 VDPWR.n1481 VSS 0.00453f
C7638 VDPWR.t623 VSS 0.005483f
C7639 VDPWR.n1482 VSS 0.007477f
C7640 VDPWR.n1483 VSS 0.002944f
C7641 VDPWR.n1484 VSS 0.002048f
C7642 VDPWR.n1485 VSS 0.012342f
C7643 VDPWR.n1486 VSS 0.012758f
C7644 VDPWR.n1487 VSS 0.002048f
C7645 VDPWR.n1488 VSS 0.00224f
C7646 VDPWR.n1489 VSS 0.001973f
C7647 VDPWR.n1490 VSS 0.003083f
C7648 VDPWR.n1491 VSS 0.003404f
C7649 VDPWR.n1492 VSS 0.155317f
C7650 VDPWR.n1493 VSS 0.003404f
C7651 VDPWR.n1494 VSS 0.003083f
C7652 VDPWR.n1495 VSS 5.48e-19
C7653 VDPWR.n1496 VSS 0.003168f
C7654 VDPWR.n1497 VSS 0.00224f
C7655 VDPWR.n1498 VSS 0.001642f
C7656 VDPWR.n1499 VSS 0.003023f
C7657 VDPWR.n1500 VSS 0.002272f
C7658 VDPWR.n1501 VSS 0.004416f
C7659 VDPWR.n1502 VSS 0.008674f
C7660 VDPWR.t685 VSS 0.004984f
C7661 VDPWR.n1503 VSS 0.011445f
C7662 VDPWR.n1504 VSS 0.015143f
C7663 VDPWR.n1505 VSS 0.052403f
C7664 VDPWR.t1222 VSS 0.072626f
C7665 VDPWR.n1506 VSS 0.040608f
C7666 VDPWR.n1507 VSS 0.010509f
C7667 VDPWR.n1508 VSS 0.005888f
C7668 VDPWR.n1509 VSS 0.005888f
C7669 VDPWR.n1510 VSS 0.005888f
C7670 VDPWR.n1511 VSS 0.020793f
C7671 VDPWR.n1512 VSS 0.020793f
C7672 VDPWR.n1513 VSS 0.020115f
C7673 VDPWR.n1514 VSS 0.005888f
C7674 VDPWR.n1515 VSS 0.003488f
C7675 VDPWR.n1516 VSS 0.008952f
C7676 VDPWR.n1517 VSS 0.00176f
C7677 VDPWR.n1518 VSS 0.007073f
C7678 VDPWR.n1519 VSS 0.013601f
C7679 VDPWR.t655 VSS 0.005483f
C7680 VDPWR.n1520 VSS 0.00426f
C7681 VDPWR.t460 VSS 0.005483f
C7682 VDPWR.t608 VSS 0.005483f
C7683 VDPWR.n1521 VSS 0.007477f
C7684 VDPWR.n1522 VSS 9.32e-19
C7685 VDPWR.n1523 VSS 0.005888f
C7686 VDPWR.t1195 VSS 0.072626f
C7687 VDPWR.t1170 VSS 0.072626f
C7688 VDPWR.n1524 VSS 0.066804f
C7689 VDPWR.n1525 VSS 0.005888f
C7690 VDPWR.n1526 VSS 0.012758f
C7691 VDPWR.n1527 VSS 0.005888f
C7692 VDPWR.t461 VSS 0.005483f
C7693 VDPWR.t609 VSS 0.005483f
C7694 VDPWR.n1528 VSS 0.007477f
C7695 VDPWR.n1529 VSS 7.36e-19
C7696 VDPWR.n1530 VSS 0.001973f
C7697 VDPWR.n1531 VSS 0.155317f
C7698 VDPWR.n1532 VSS 0.00352f
C7699 VDPWR.n1533 VSS 0.001579f
C7700 VDPWR.n1534 VSS 0.0024f
C7701 VDPWR.n1535 VSS 0.002048f
C7702 VDPWR.n1536 VSS 0.002112f
C7703 VDPWR.n1537 VSS 0.00453f
C7704 VDPWR.t451 VSS 0.005024f
C7705 VDPWR.t1257 VSS 0.010664f
C7706 VDPWR.n1539 VSS 0.027341f
C7707 VDPWR.t452 VSS 0.005024f
C7708 VDPWR.n1540 VSS 0.014893f
C7709 VDPWR.t648 VSS 0.005024f
C7710 VDPWR.t1226 VSS 0.010664f
C7711 VDPWR.n1542 VSS 0.027341f
C7712 VDPWR.t649 VSS 0.005024f
C7713 VDPWR.n1543 VSS 0.014893f
C7714 VDPWR.n1544 VSS 0.001973f
C7715 VDPWR.n1545 VSS 0.003404f
C7716 VDPWR.n1546 VSS 0.003083f
C7717 VDPWR.n1547 VSS 0.002885f
C7718 VDPWR.n1548 VSS 0.001376f
C7719 VDPWR.n1549 VSS 0.012555f
C7720 VDPWR.n1550 VSS 0.002048f
C7721 VDPWR.n1551 VSS 0.002944f
C7722 VDPWR.n1552 VSS 0.001973f
C7723 VDPWR.n1553 VSS 0.001579f
C7724 VDPWR.n1554 VSS 0.00352f
C7725 VDPWR.n1555 VSS 0.003404f
C7726 VDPWR.n1556 VSS 0.003083f
C7727 VDPWR.n1557 VSS 0.002949f
C7728 VDPWR.n1558 VSS 0.005696f
C7729 VDPWR.n1559 VSS 0.012342f
C7730 VDPWR.n1560 VSS 0.012758f
C7731 VDPWR.n1561 VSS 0.012758f
C7732 VDPWR.n1562 VSS 0.005888f
C7733 VDPWR.n1563 VSS 0.005888f
C7734 VDPWR.n1564 VSS 0.005888f
C7735 VDPWR.n1565 VSS 0.012758f
C7736 VDPWR.n1566 VSS 0.012758f
C7737 VDPWR.n1567 VSS 0.009361f
C7738 VDPWR.n1568 VSS 0.005888f
C7739 VDPWR.n1569 VSS 0.005888f
C7740 VDPWR.n1570 VSS 0.009777f
C7741 VDPWR.n1571 VSS 0.012758f
C7742 VDPWR.n1572 VSS 0.012342f
C7743 VDPWR.n1573 VSS 0.005888f
C7744 VDPWR.n1574 VSS 0.004416f
C7745 VDPWR.n1575 VSS 0.004739f
C7746 VDPWR.n1576 VSS 0.002934f
C7747 VDPWR.n1577 VSS 0.001504f
C7748 VDPWR.n1578 VSS 0.002944f
C7749 VDPWR.n1579 VSS 0.001973f
C7750 VDPWR.n1580 VSS 0.00352f
C7751 VDPWR.n1581 VSS 0.001579f
C7752 VDPWR.n1582 VSS 0.001973f
C7753 VDPWR.n1583 VSS 0.002112f
C7754 VDPWR.n1584 VSS 0.002336f
C7755 VDPWR.n1585 VSS 0.001973f
C7756 VDPWR.n1586 VSS 0.003083f
C7757 VDPWR.n1587 VSS 0.003404f
C7758 VDPWR.n1588 VSS 0.155317f
C7759 VDPWR.n1589 VSS 0.116061f
C7760 VDPWR.n1590 VSS 0.281618f
C7761 VDPWR.n1591 VSS 0.281618f
C7762 VDPWR.n1592 VSS 0.281618f
C7763 VDPWR.n1593 VSS 0.532156f
C7764 VDPWR.n1594 VSS 0.194931f
C7765 VDPWR.n1595 VSS 0.003404f
C7766 VDPWR.n1596 VSS 0.194931f
C7767 VDPWR.n1597 VSS 0.00352f
C7768 VDPWR.n1598 VSS 0.002629f
C7769 VDPWR.n1599 VSS 0.001579f
C7770 VDPWR.n1600 VSS 0.002944f
C7771 VDPWR.n1601 VSS 0.015256f
C7772 VDPWR.t578 VSS 0.005483f
C7773 VDPWR.t478 VSS 0.004984f
C7774 VDPWR.n1602 VSS 0.011995f
C7775 VDPWR.n1603 VSS 0.003842f
C7776 VDPWR.t617 VSS 0.005024f
C7777 VDPWR.t1186 VSS 0.010664f
C7778 VDPWR.n1605 VSS 0.027341f
C7779 VDPWR.t618 VSS 0.005024f
C7780 VDPWR.n1606 VSS 0.014893f
C7781 VDPWR.n1607 VSS 0.00352f
C7782 VDPWR.n1608 VSS 0.004416f
C7783 VDPWR.n1609 VSS 0.004957f
C7784 VDPWR.t694 VSS 0.005024f
C7785 VDPWR.t1169 VSS 0.010664f
C7786 VDPWR.n1611 VSS 0.027341f
C7787 VDPWR.t695 VSS 0.005024f
C7788 VDPWR.n1612 VSS 0.014893f
C7789 VDPWR.t442 VSS 0.005024f
C7790 VDPWR.t1251 VSS 0.010664f
C7791 VDPWR.n1614 VSS 0.027341f
C7792 VDPWR.t443 VSS 0.005024f
C7793 VDPWR.n1615 VSS 0.014893f
C7794 VDPWR.n1616 VSS 0.003844f
C7795 VDPWR.t534 VSS 0.005024f
C7796 VDPWR.t1229 VSS 0.010664f
C7797 VDPWR.n1618 VSS 0.027341f
C7798 VDPWR.t535 VSS 0.005024f
C7799 VDPWR.n1619 VSS 0.014893f
C7800 VDPWR.n1620 VSS 0.01227f
C7801 VDPWR.n1621 VSS 0.013462f
C7802 VDPWR.n1622 VSS 0.00331f
C7803 VDPWR.t1241 VSS 0.036234f
C7804 VDPWR.n1623 VSS 0.027337f
C7805 VDPWR.n1624 VSS 0.025685f
C7806 VDPWR.t1210 VSS 0.072626f
C7807 VDPWR.n1625 VSS 0.040608f
C7808 VDPWR.n1626 VSS 0.005888f
C7809 VDPWR.t479 VSS 0.004984f
C7810 VDPWR.n1627 VSS 0.011445f
C7811 VDPWR.t560 VSS 0.005483f
C7812 VDPWR.n1628 VSS 0.006928f
C7813 VDPWR.n1629 VSS 0.005888f
C7814 VDPWR.t1208 VSS 0.074001f
C7815 VDPWR.n1630 VSS 0.034322f
C7816 VDPWR.n1631 VSS 0.005888f
C7817 VDPWR.t1224 VSS 0.072626f
C7818 VDPWR.n1632 VSS 0.009361f
C7819 VDPWR.n1633 VSS 0.036592f
C7820 VDPWR.n1634 VSS 0.009777f
C7821 VDPWR.n1635 VSS 0.004544f
C7822 VDPWR.n1636 VSS 0.005888f
C7823 VDPWR.n1637 VSS 0.012758f
C7824 VDPWR.n1638 VSS 0.012342f
C7825 VDPWR.t546 VSS 0.005483f
C7826 VDPWR.n1639 VSS 0.006928f
C7827 VDPWR.n1640 VSS 0.002865f
C7828 VDPWR.n1641 VSS 0.005344f
C7829 VDPWR.n1642 VSS 0.003488f
C7830 VDPWR.n1643 VSS 0.003209f
C7831 VDPWR.t579 VSS 0.005483f
C7832 VDPWR.n1644 VSS 0.006928f
C7833 VDPWR.n1645 VSS 0.012342f
C7834 VDPWR.n1646 VSS 0.012342f
C7835 VDPWR.n1647 VSS 0.005888f
C7836 VDPWR.n1648 VSS 0.004416f
C7837 VDPWR.n1649 VSS 0.005612f
C7838 VDPWR.n1650 VSS 0.008742f
C7839 VDPWR.n1651 VSS 0.003488f
C7840 VDPWR.n1652 VSS 0.005888f
C7841 VDPWR.n1653 VSS 0.020115f
C7842 VDPWR.n1654 VSS 0.020793f
C7843 VDPWR.n1655 VSS 0.015256f
C7844 VDPWR.n1656 VSS 0.003008f
C7845 VDPWR.n1657 VSS 0.002117f
C7846 VDPWR.n1658 VSS 0.001973f
C7847 VDPWR.n1659 VSS 0.00352f
C7848 VDPWR.n1660 VSS 0.001579f
C7849 VDPWR.n1661 VSS 0.003083f
C7850 VDPWR.n1662 VSS 0.001973f
C7851 VDPWR.n1663 VSS 0.00288f
C7852 VDPWR.n1664 VSS 0.002048f
C7853 VDPWR.n1665 VSS 0.015934f
C7854 VDPWR.n1666 VSS 0.015256f
C7855 VDPWR.n1667 VSS 0.002048f
C7856 VDPWR.n1668 VSS 0.002368f
C7857 VDPWR.n1669 VSS 0.001973f
C7858 VDPWR.n1670 VSS 0.003083f
C7859 VDPWR.n1671 VSS 0.003404f
C7860 VDPWR.n1672 VSS 0.140809f
C7861 VDPWR.n1673 VSS 0.281618f
C7862 VDPWR.n1674 VSS 0.532156f
C7863 VDPWR.n1675 VSS 0.194931f
C7864 VDPWR.n1676 VSS 0.00352f
C7865 VDPWR.n1677 VSS 0.002629f
C7866 VDPWR.n1678 VSS 0.001579f
C7867 VDPWR.n1679 VSS 0.001579f
C7868 VDPWR.n1680 VSS 0.001973f
C7869 VDPWR.n1681 VSS 0.002944f
C7870 VDPWR.t1199 VSS 0.036234f
C7871 VDPWR.n1682 VSS 0.027337f
C7872 VDPWR.t581 VSS 0.005483f
C7873 VDPWR.t718 VSS 0.004984f
C7874 VDPWR.n1683 VSS 0.011995f
C7875 VDPWR.t690 VSS 0.005024f
C7876 VDPWR.t1221 VSS 0.010664f
C7877 VDPWR.n1685 VSS 0.027341f
C7878 VDPWR.t691 VSS 0.005024f
C7879 VDPWR.n1686 VSS 0.014893f
C7880 VDPWR.t537 VSS 0.005024f
C7881 VDPWR.t1266 VSS 0.010664f
C7882 VDPWR.n1688 VSS 0.027341f
C7883 VDPWR.t538 VSS 0.005024f
C7884 VDPWR.n1689 VSS 0.014893f
C7885 VDPWR.n1690 VSS 0.01227f
C7886 VDPWR.t520 VSS 0.005024f
C7887 VDPWR.t1227 VSS 0.010664f
C7888 VDPWR.n1692 VSS 0.027341f
C7889 VDPWR.t521 VSS 0.005024f
C7890 VDPWR.n1693 VSS 0.014893f
C7891 VDPWR.n1694 VSS 0.003844f
C7892 VDPWR.n1695 VSS 0.004957f
C7893 VDPWR.t702 VSS 0.005024f
C7894 VDPWR.t1197 VSS 0.010664f
C7895 VDPWR.n1697 VSS 0.027341f
C7896 VDPWR.t703 VSS 0.005024f
C7897 VDPWR.n1698 VSS 0.014893f
C7898 VDPWR.n1699 VSS 0.013462f
C7899 VDPWR.n1700 VSS 0.00331f
C7900 VDPWR.n1701 VSS 0.003842f
C7901 VDPWR.n1702 VSS 0.004416f
C7902 VDPWR.n1703 VSS 0.00352f
C7903 VDPWR.n1704 VSS 0.015256f
C7904 VDPWR.n1705 VSS 0.025685f
C7905 VDPWR.n1706 VSS 0.002048f
C7906 VDPWR.n1707 VSS 0.015934f
C7907 VDPWR.n1708 VSS 0.015256f
C7908 VDPWR.n1709 VSS 0.002048f
C7909 VDPWR.n1710 VSS 0.002368f
C7910 VDPWR.n1711 VSS 0.001973f
C7911 VDPWR.n1712 VSS 0.003083f
C7912 VDPWR.n1713 VSS 0.003404f
C7913 VDPWR.n1714 VSS 0.140809f
C7914 VDPWR.n1715 VSS 0.003404f
C7915 VDPWR.n1716 VSS 0.003083f
C7916 VDPWR.n1717 VSS 0.002117f
C7917 VDPWR.n1718 VSS 0.003008f
C7918 VDPWR.n1719 VSS 0.015256f
C7919 VDPWR.n1720 VSS 0.020793f
C7920 VDPWR.t719 VSS 0.004984f
C7921 VDPWR.n1721 VSS 0.011445f
C7922 VDPWR.n1722 VSS 0.020115f
C7923 VDPWR.n1723 VSS 0.005888f
C7924 VDPWR.n1724 VSS 0.003488f
C7925 VDPWR.n1725 VSS 0.004416f
C7926 VDPWR.n1726 VSS 0.005612f
C7927 VDPWR.t469 VSS 0.005483f
C7928 VDPWR.n1727 VSS 0.006928f
C7929 VDPWR.n1728 VSS 0.012342f
C7930 VDPWR.n1729 VSS 0.012342f
C7931 VDPWR.n1730 VSS 0.005888f
C7932 VDPWR.n1731 VSS 0.003488f
C7933 VDPWR.n1732 VSS 0.003209f
C7934 VDPWR.n1733 VSS 0.034322f
C7935 VDPWR.n1734 VSS 0.002865f
C7936 VDPWR.t551 VSS 0.005483f
C7937 VDPWR.n1735 VSS 0.006928f
C7938 VDPWR.n1736 VSS 0.012342f
C7939 VDPWR.n1737 VSS 0.005888f
C7940 VDPWR.n1738 VSS 0.005888f
C7941 VDPWR.n1739 VSS 0.004544f
C7942 VDPWR.n1740 VSS 0.009777f
C7943 VDPWR.n1741 VSS 0.036592f
C7944 VDPWR.n1742 VSS 0.009361f
C7945 VDPWR.t470 VSS 0.005483f
C7946 VDPWR.n1743 VSS 0.006928f
C7947 VDPWR.n1744 VSS 0.012342f
C7948 VDPWR.n1745 VSS 0.012758f
C7949 VDPWR.n1746 VSS 0.002048f
C7950 VDPWR.n1747 VSS 0.001579f
C7951 VDPWR.n1748 VSS 0.001973f
C7952 VDPWR.n1749 VSS 0.00224f
C7953 VDPWR.n1750 VSS 0.002752f
C7954 VDPWR.n1751 VSS 0.001973f
C7955 VDPWR.n1752 VSS 0.003083f
C7956 VDPWR.n1753 VSS 0.003404f
C7957 VDPWR.n1754 VSS 0.140809f
C7958 VDPWR.n1755 VSS 0.003404f
C7959 VDPWR.n1756 VSS 0.003083f
C7960 VDPWR.n1757 VSS 0.002949f
C7961 VDPWR.n1758 VSS 0.002528f
C7962 VDPWR.n1759 VSS 0.003168f
C7963 VDPWR.n1760 VSS 0.017118f
C7964 VDPWR.t552 VSS 0.0055f
C7965 VDPWR.n1761 VSS 0.011274f
C7966 VDPWR.n1762 VSS 0.006252f
C7967 VDPWR.n1763 VSS 0.00224f
C7968 VDPWR.n1764 VSS 0.003146f
C7969 VDPWR.n1765 VSS 0.00425f
C7970 VDPWR.n1766 VSS 0.007049f
C7971 VDPWR.t753 VSS 0.0055f
C7972 VDPWR.n1767 VSS 0.011154f
C7973 VDPWR.n1768 VSS 0.004646f
C7974 VDPWR.t611 VSS 0.005483f
C7975 VDPWR.n1769 VSS 0.006928f
C7976 VDPWR.t1175 VSS 0.072626f
C7977 VDPWR.n1770 VSS 0.036592f
C7978 VDPWR.n1771 VSS 0.009361f
C7979 VDPWR.n1772 VSS 0.005888f
C7980 VDPWR.n1773 VSS 0.005888f
C7981 VDPWR.n1774 VSS 0.005568f
C7982 VDPWR.n1775 VSS 0.009777f
C7983 VDPWR.n1776 VSS 0.036592f
C7984 VDPWR.n1777 VSS 0.009361f
C7985 VDPWR.n1778 VSS 0.012758f
C7986 VDPWR.n1779 VSS 0.002048f
C7987 VDPWR.n1780 VSS 0.002944f
C7988 VDPWR.n1781 VSS 0.001973f
C7989 VDPWR.n1782 VSS 0.003083f
C7990 VDPWR.n1783 VSS 0.003404f
C7991 VDPWR.n1784 VSS 0.140809f
C7992 VDPWR.n1785 VSS 0.003404f
C7993 VDPWR.n1786 VSS 0.003083f
C7994 VDPWR.n1787 VSS 0.002949f
C7995 VDPWR.n1788 VSS 0.003904f
C7996 VDPWR.n1789 VSS 0.012758f
C7997 VDPWR.n1790 VSS 0.012342f
C7998 VDPWR.t754 VSS 0.005483f
C7999 VDPWR.n1791 VSS 0.006928f
C8000 VDPWR.n1792 VSS 0.004736f
C8001 VDPWR.n1793 VSS 0.003488f
C8002 VDPWR.n1794 VSS 0.00425f
C8003 VDPWR.n1795 VSS 0.004321f
C8004 VDPWR.t651 VSS 0.0055f
C8005 VDPWR.n1796 VSS 0.011154f
C8006 VDPWR.n1797 VSS 0.004646f
C8007 VDPWR.t575 VSS 0.005483f
C8008 VDPWR.n1798 VSS 0.006928f
C8009 VDPWR.n1799 VSS 0.009361f
C8010 VDPWR.n1800 VSS 0.005888f
C8011 VDPWR.n1801 VSS 0.005888f
C8012 VDPWR.n1802 VSS 0.009361f
C8013 VDPWR.n1803 VSS 0.009777f
C8014 VDPWR.n1804 VSS 0.036592f
C8015 VDPWR.n1805 VSS 0.009361f
C8016 VDPWR.n1806 VSS 0.005888f
C8017 VDPWR.n1807 VSS 0.005888f
C8018 VDPWR.n1808 VSS 0.003648f
C8019 VDPWR.n1809 VSS 0.012758f
C8020 VDPWR.t652 VSS 0.005483f
C8021 VDPWR.n1810 VSS 0.006928f
C8022 VDPWR.n1811 VSS 0.002944f
C8023 VDPWR.n1812 VSS 0.002048f
C8024 VDPWR.n1813 VSS 0.012342f
C8025 VDPWR.n1814 VSS 0.012758f
C8026 VDPWR.n1815 VSS 0.002048f
C8027 VDPWR.n1816 VSS 0.00224f
C8028 VDPWR.n1817 VSS 0.001973f
C8029 VDPWR.n1818 VSS 0.003083f
C8030 VDPWR.n1819 VSS 0.003404f
C8031 VDPWR.n1820 VSS 0.140809f
C8032 VDPWR.n1821 VSS 0.003404f
C8033 VDPWR.n1822 VSS 0.003083f
C8034 VDPWR.n1823 VSS 5.48e-19
C8035 VDPWR.n1824 VSS 0.003168f
C8036 VDPWR.n1825 VSS 0.015948f
C8037 VDPWR.t576 VSS 0.005504f
C8038 VDPWR.n1826 VSS 0.00626f
C8039 VDPWR.n1827 VSS 0.008018f
C8040 VDPWR.t1181 VSS 0.021195f
C8041 VDPWR.n1828 VSS 0.007844f
C8042 VDPWR.t745 VSS 0.004984f
C8043 VDPWR.n1829 VSS 0.003662f
C8044 VDPWR.n1830 VSS 0.002301f
C8045 VDPWR.n1831 VSS 0.002016f
C8046 VDPWR.n1832 VSS 0.006108f
C8047 VDPWR.n1833 VSS 0.012813f
C8048 VDPWR.n1834 VSS 0.016328f
C8049 VDPWR.t1219 VSS 0.072626f
C8050 VDPWR.n1835 VSS 0.033842f
C8051 VDPWR.n1836 VSS 0.004517f
C8052 VDPWR.n1837 VSS 0.002016f
C8053 VDPWR.n1838 VSS 0.005344f
C8054 VDPWR.n1839 VSS 0.003792f
C8055 VDPWR.n1840 VSS 0.007139f
C8056 VDPWR.n1841 VSS 0.007119f
C8057 VDPWR.n1842 VSS 0.003993f
C8058 VDPWR.n1843 VSS 0.005888f
C8059 VDPWR.n1844 VSS 0.005888f
C8060 VDPWR.n1845 VSS 0.004672f
C8061 VDPWR.n1846 VSS 0.007422f
C8062 VDPWR.t169 VSS 0.002785f
C8063 VDPWR.t27 VSS 0.00135f
C8064 VDPWR.n1847 VSS 0.00567f
C8065 VDPWR.n1848 VSS 0.006831f
C8066 VDPWR.n1849 VSS 0.005687f
C8067 VDPWR.n1850 VSS 0.007422f
C8068 VDPWR.n1851 VSS 0.002048f
C8069 VDPWR.n1852 VSS 0.001973f
C8070 VDPWR.n1853 VSS 0.002112f
C8071 VDPWR.n1854 VSS 0.00288f
C8072 VDPWR.n1855 VSS 0.001973f
C8073 VDPWR.n1856 VSS 0.003083f
C8074 VDPWR.n1857 VSS 0.003404f
C8075 VDPWR.n1858 VSS 0.00352f
C8076 VDPWR.n1859 VSS 0.00352f
C8077 VDPWR.n1860 VSS 0.003404f
C8078 VDPWR.n1861 VSS 0.003083f
C8079 VDPWR.n1862 VSS 0.001973f
C8080 VDPWR.n1863 VSS 0.002944f
C8081 VDPWR.n1864 VSS 0.001504f
C8082 VDPWR.n1865 VSS 0.003079f
C8083 VDPWR.n1866 VSS 0.001972f
C8084 VDPWR.n1867 VSS 0.0048f
C8085 VDPWR.n1868 VSS 0.005888f
C8086 VDPWR.n1869 VSS 0.005888f
C8087 VDPWR.n1870 VSS 0.001247f
C8088 VDPWR.n1871 VSS 0.00338f
C8089 VDPWR.t3 VSS 0.002834f
C8090 VDPWR.n1872 VSS 0.00693f
C8091 VDPWR.t937 VSS 0.0018f
C8092 VDPWR.t941 VSS 0.0018f
C8093 VDPWR.n1873 VSS 0.003905f
C8094 VDPWR.t907 VSS 0.0018f
C8095 VDPWR.t1 VSS 0.0018f
C8096 VDPWR.n1874 VSS 0.004032f
C8097 VDPWR.n1875 VSS 0.005167f
C8098 VDPWR.n1876 VSS 0.004501f
C8099 VDPWR.n1877 VSS 9.41e-19
C8100 VDPWR.n1878 VSS 0.005888f
C8101 VDPWR.n1879 VSS 0.005888f
C8102 VDPWR.n1880 VSS 0.003488f
C8103 VDPWR.n1881 VSS 0.002085f
C8104 VDPWR.n1882 VSS 0.001757f
C8105 VDPWR.n1883 VSS 0.00224f
C8106 VDPWR.n1884 VSS 0.007808f
C8107 VDPWR.n1885 VSS 7.36e-19
C8108 VDPWR.n1886 VSS 0.006896f
C8109 VDPWR.n1887 VSS 0.003083f
C8110 VDPWR.n1888 VSS 0.001579f
C8111 VDPWR.n1889 VSS 0.001973f
C8112 VDPWR.n1890 VSS 0.001472f
C8113 VDPWR.n1891 VSS 0.002944f
C8114 VDPWR.n1892 VSS 0.002048f
C8115 VDPWR.t603 VSS 0.005024f
C8116 VDPWR.t1242 VSS 0.010664f
C8117 VDPWR.n1894 VSS 0.027341f
C8118 VDPWR.t604 VSS 0.005024f
C8119 VDPWR.n1895 VSS 0.014893f
C8120 VDPWR.n1896 VSS 0.012262f
C8121 VDPWR.n1897 VSS 0.001376f
C8122 VDPWR.n1898 VSS 0.002885f
C8123 VDPWR.n1899 VSS 0.002112f
C8124 VDPWR.n1900 VSS 0.001973f
C8125 VDPWR.n1901 VSS 0.001579f
C8126 VDPWR.n1902 VSS 0.00352f
C8127 VDPWR.n1903 VSS 0.003404f
C8128 VDPWR.n1904 VSS 0.140809f
C8129 VDPWR.n1905 VSS 0.116061f
C8130 VDPWR.n1906 VSS 0.167264f
C8131 VDPWR.n1907 VSS 0.281618f
C8132 VDPWR.n1908 VSS 0.116061f
C8133 VDPWR.n1909 VSS 0.001579f
C8134 VDPWR.n1910 VSS 0.001973f
C8135 VDPWR.n1911 VSS 0.001472f
C8136 VDPWR.n1912 VSS 0.002048f
C8137 VDPWR.n1913 VSS 0.002944f
C8138 VDPWR.n1914 VSS 0.002048f
C8139 VDPWR.n1915 VSS 0.004863f
C8140 VDPWR.t45 VSS 0.00112f
C8141 VDPWR.t95 VSS -0.001177f
C8142 VDPWR.n1916 VSS 0.007456f
C8143 VDPWR.t1003 VSS 0.002785f
C8144 VDPWR.t66 VSS 0.00135f
C8145 VDPWR.n1917 VSS 0.00567f
C8146 VDPWR.n1918 VSS 0.004338f
C8147 VDPWR.n1919 VSS 0.00438f
C8148 VDPWR.n1920 VSS 0.001111f
C8149 VDPWR.t993 VSS 0.0018f
C8150 VDPWR.t995 VSS 0.0018f
C8151 VDPWR.n1921 VSS 0.004044f
C8152 VDPWR.n1922 VSS 0.017119f
C8153 VDPWR.t997 VSS 0.002834f
C8154 VDPWR.n1923 VSS 0.005888f
C8155 VDPWR.n1924 VSS 0.01283f
C8156 VDPWR.t1196 VSS 0.037391f
C8157 VDPWR.t606 VSS 0.004984f
C8158 VDPWR.n1925 VSS 0.06261f
C8159 VDPWR.n1926 VSS 0.016449f
C8160 VDPWR.t933 VSS 0.001867f
C8161 VDPWR.t48 VSS 0.002067f
C8162 VDPWR.n1927 VSS 0.003981f
C8163 VDPWR.t607 VSS 0.004984f
C8164 VDPWR.n1928 VSS 0.008777f
C8165 VDPWR.n1929 VSS 7.36e-19
C8166 VDPWR.n1930 VSS 0.001973f
C8167 VDPWR.n1931 VSS 0.00352f
C8168 VDPWR.n1932 VSS 0.001579f
C8169 VDPWR.n1933 VSS 0.001472f
C8170 VDPWR.n1934 VSS 0.002048f
C8171 VDPWR.n1935 VSS 0.002112f
C8172 VDPWR.n1936 VSS 0.005471f
C8173 VDPWR.t514 VSS 0.005024f
C8174 VDPWR.t1232 VSS 0.010664f
C8175 VDPWR.n1938 VSS 0.027341f
C8176 VDPWR.t515 VSS 0.005024f
C8177 VDPWR.n1939 VSS 0.014893f
C8178 VDPWR.t592 VSS 0.005024f
C8179 VDPWR.t1203 VSS 0.010664f
C8180 VDPWR.n1941 VSS 0.027341f
C8181 VDPWR.t593 VSS 0.005024f
C8182 VDPWR.n1942 VSS 0.014893f
C8183 VDPWR.n1943 VSS 0.001973f
C8184 VDPWR.n1944 VSS 0.003404f
C8185 VDPWR.n1945 VSS 0.003083f
C8186 VDPWR.n1946 VSS 0.002885f
C8187 VDPWR.n1947 VSS 0.001376f
C8188 VDPWR.n1948 VSS 0.012553f
C8189 VDPWR.n1949 VSS 0.002048f
C8190 VDPWR.n1950 VSS 0.002944f
C8191 VDPWR.n1951 VSS 0.001973f
C8192 VDPWR.n1952 VSS 0.001579f
C8193 VDPWR.n1953 VSS 0.00352f
C8194 VDPWR.n1954 VSS 0.003404f
C8195 VDPWR.n1955 VSS 0.003083f
C8196 VDPWR.n1956 VSS 0.001477f
C8197 VDPWR.n1957 VSS 0.004416f
C8198 VDPWR.n1958 VSS 0.014953f
C8199 VDPWR.n1959 VSS 0.007897f
C8200 VDPWR.n1960 VSS 0.009969f
C8201 VDPWR.n1961 VSS 0.012517f
C8202 VDPWR.n1962 VSS 0.005344f
C8203 VDPWR.n1963 VSS 0.002016f
C8204 VDPWR.n1964 VSS 0.006234f
C8205 VDPWR.n1965 VSS 0.00224f
C8206 VDPWR.n1966 VSS 0.006477f
C8207 VDPWR.t1018 VSS 7.56e-19
C8208 VDPWR.t935 VSS 7.56e-19
C8209 VDPWR.n1967 VSS 0.00175f
C8210 VDPWR.n1968 VSS 0.016544f
C8211 VDPWR.n1969 VSS 0.002085f
C8212 VDPWR.n1970 VSS 0.006766f
C8213 VDPWR.n1971 VSS 0.002949f
C8214 VDPWR.n1972 VSS 0.003083f
C8215 VDPWR.n1973 VSS 0.003404f
C8216 VDPWR.n1974 VSS 0.140809f
C8217 VDPWR.n1975 VSS 0.003404f
C8218 VDPWR.n1976 VSS 0.00352f
C8219 VDPWR.n1977 VSS 0.001579f
C8220 VDPWR.n1978 VSS 0.001973f
C8221 VDPWR.n1979 VSS 9.28e-19
C8222 VDPWR.n1980 VSS 0.001711f
C8223 VDPWR.t347 VSS 0.002467f
C8224 VDPWR.t1005 VSS 0.001867f
C8225 VDPWR.n1981 VSS 0.00469f
C8226 VDPWR.n1982 VSS 0.009342f
C8227 VDPWR.n1983 VSS 0.001643f
C8228 VDPWR.n1984 VSS 0.005888f
C8229 VDPWR.n1985 VSS 0.004416f
C8230 VDPWR.n1986 VSS 1.47e-19
C8231 VDPWR.n1987 VSS 0.004452f
C8232 VDPWR.n1988 VSS 0.001655f
C8233 VDPWR.t1014 VSS 0.001152f
C8234 VDPWR.t137 VSS 0.001152f
C8235 VDPWR.n1989 VSS 0.002399f
C8236 VDPWR.n1990 VSS 0.006697f
C8237 VDPWR.n1991 VSS 0.005344f
C8238 VDPWR.n1992 VSS 0.002016f
C8239 VDPWR.n1993 VSS 0.003488f
C8240 VDPWR.n1994 VSS 0.007364f
C8241 VDPWR.t660 VSS 0.005483f
C8242 VDPWR.n1995 VSS 0.011995f
C8243 VDPWR.n1996 VSS 0.020115f
C8244 VDPWR.n1997 VSS 0.015595f
C8245 VDPWR.n1998 VSS 0.005888f
C8246 VDPWR.n1999 VSS 0.004416f
C8247 VDPWR.n2000 VSS 0.008952f
C8248 VDPWR.n2001 VSS 0.016769f
C8249 VDPWR.n2002 VSS 0.003168f
C8250 VDPWR.n2003 VSS 5.48e-19
C8251 VDPWR.n2004 VSS 0.003083f
C8252 VDPWR.n2005 VSS 0.003404f
C8253 VDPWR.n2006 VSS 0.140809f
C8254 VDPWR.n2007 VSS 0.003404f
C8255 VDPWR.n2008 VSS 0.003083f
C8256 VDPWR.n2009 VSS 0.002757f
C8257 VDPWR.n2010 VSS 0.003648f
C8258 VDPWR.n2011 VSS 0.009777f
C8259 VDPWR.n2012 VSS 0.012758f
C8260 VDPWR.n2013 VSS 0.012342f
C8261 VDPWR.n2014 VSS 0.005888f
C8262 VDPWR.n2015 VSS 0.005344f
C8263 VDPWR.n2016 VSS 0.005756f
C8264 VDPWR.n2017 VSS 0.005803f
C8265 VDPWR.n2018 VSS 0.003488f
C8266 VDPWR.n2019 VSS 0.005888f
C8267 VDPWR.n2020 VSS 0.009777f
C8268 VDPWR.n2021 VSS 0.012758f
C8269 VDPWR.n2022 VSS 0.012342f
C8270 VDPWR.n2023 VSS 0.005888f
C8271 VDPWR.n2024 VSS 0.005344f
C8272 VDPWR.n2025 VSS 0.003488f
C8273 VDPWR.n2026 VSS 0.005803f
C8274 VDPWR.t751 VSS 0.005483f
C8275 VDPWR.n2027 VSS 0.006928f
C8276 VDPWR.n2028 VSS 0.012342f
C8277 VDPWR.n2029 VSS 0.009361f
C8278 VDPWR.n2030 VSS 0.003904f
C8279 VDPWR.n2031 VSS 0.002949f
C8280 VDPWR.n2032 VSS 0.003083f
C8281 VDPWR.n2033 VSS 0.003404f
C8282 VDPWR.n2034 VSS 0.00352f
C8283 VDPWR.n2035 VSS 0.00352f
C8284 VDPWR.n2036 VSS 0.003404f
C8285 VDPWR.n2037 VSS 0.003083f
C8286 VDPWR.n2038 VSS 0.002949f
C8287 VDPWR.n2039 VSS 0.004096f
C8288 VDPWR.n2040 VSS 0.005612f
C8289 VDPWR.n2041 VSS 0.008742f
C8290 VDPWR.n2042 VSS 0.003488f
C8291 VDPWR.n2043 VSS 0.005888f
C8292 VDPWR.n2044 VSS 0.005888f
C8293 VDPWR.n2045 VSS 0.020793f
C8294 VDPWR.n2046 VSS 0.020115f
C8295 VDPWR.t750 VSS 0.005483f
C8296 VDPWR.n2047 VSS 0.010606f
C8297 VDPWR.n2048 VSS 0.013537f
C8298 VDPWR.t448 VSS 0.004984f
C8299 VDPWR.n2049 VSS 0.029901f
C8300 VDPWR.t1249 VSS 0.017526f
C8301 VDPWR.n2050 VSS 0.03397f
C8302 VDPWR.n2051 VSS 0.007752f
C8303 VDPWR.n2052 VSS 0.001735f
C8304 VDPWR.n2053 VSS 0.009861f
C8305 VDPWR.n2054 VSS 0.005344f
C8306 VDPWR.n2055 VSS 0.004953f
C8307 VDPWR.n2056 VSS 0.003168f
C8308 VDPWR.n2057 VSS 0.002528f
C8309 VDPWR.n2058 VSS 0.006017f
C8310 VDPWR.t561 VSS 0.005483f
C8311 VDPWR.n2059 VSS 0.006928f
C8312 VDPWR.n2060 VSS 0.012342f
C8313 VDPWR.n2061 VSS 0.002048f
C8314 VDPWR.n2062 VSS 0.002944f
C8315 VDPWR.n2063 VSS 0.001973f
C8316 VDPWR.n2064 VSS 0.00352f
C8317 VDPWR.n2065 VSS 0.001579f
C8318 VDPWR.n2066 VSS 0.001973f
C8319 VDPWR.n2067 VSS 0.00224f
C8320 VDPWR.n2068 VSS 0.002752f
C8321 VDPWR.n2069 VSS 0.001973f
C8322 VDPWR.n2070 VSS 0.003083f
C8323 VDPWR.n2071 VSS 0.003404f
C8324 VDPWR.n2072 VSS 0.140809f
C8325 VDPWR.n2073 VSS 0.116061f
C8326 VDPWR.n2074 VSS 0.00352f
C8327 VDPWR.n2075 VSS 0.002949f
C8328 VDPWR.n2076 VSS 0.001579f
C8329 VDPWR.t1279 VSS 0.072626f
C8330 VDPWR.n2077 VSS 0.036592f
C8331 VDPWR.n2078 VSS 0.005888f
C8332 VDPWR.t1209 VSS 0.072626f
C8333 VDPWR.n2079 VSS 0.036175f
C8334 VDPWR.t494 VSS 0.005483f
C8335 VDPWR.n2080 VSS 0.006928f
C8336 VDPWR.n2081 VSS 0.004416f
C8337 VDPWR.t558 VSS 0.004984f
C8338 VDPWR.n2082 VSS 0.011445f
C8339 VDPWR.n2083 VSS 0.005888f
C8340 VDPWR.n2084 VSS 0.015256f
C8341 VDPWR.n2085 VSS 0.00288f
C8342 VDPWR.n2086 VSS 0.001973f
C8343 VDPWR.n2087 VSS 0.00352f
C8344 VDPWR.n2088 VSS 0.001579f
C8345 VDPWR.n2089 VSS 0.002368f
C8346 VDPWR.t1243 VSS 0.036876f
C8347 VDPWR.t557 VSS 0.004984f
C8348 VDPWR.n2090 VSS 0.011445f
C8349 VDPWR.t680 VSS 0.005101f
C8350 VDPWR.n2091 VSS 0.002138f
C8351 VDPWR.n2092 VSS 0.011656f
C8352 VDPWR.t1188 VSS 0.010699f
C8353 VDPWR.n2093 VSS 0.020574f
C8354 VDPWR.t679 VSS 0.005024f
C8355 VDPWR.n2094 VSS 0.007271f
C8356 VDPWR.n2095 VSS 0.007169f
C8357 VDPWR.t526 VSS 0.005024f
C8358 VDPWR.t1254 VSS 0.010664f
C8359 VDPWR.n2097 VSS 0.027341f
C8360 VDPWR.t527 VSS 0.005024f
C8361 VDPWR.n2098 VSS 0.014893f
C8362 VDPWR.t635 VSS 0.005024f
C8363 VDPWR.t1183 VSS 0.010664f
C8364 VDPWR.n2100 VSS 0.027341f
C8365 VDPWR.t636 VSS 0.005024f
C8366 VDPWR.n2101 VSS 0.014893f
C8367 VDPWR.n2102 VSS 0.01227f
C8368 VDPWR.n2103 VSS 0.003844f
C8369 VDPWR.n2104 VSS 0.003523f
C8370 VDPWR.n2105 VSS 0.002016f
C8371 VDPWR.n2106 VSS 0.002762f
C8372 VDPWR.t493 VSS 0.005503f
C8373 VDPWR.n2107 VSS 0.006102f
C8374 VDPWR.n2108 VSS 0.007518f
C8375 VDPWR.n2109 VSS 0.004416f
C8376 VDPWR.n2110 VSS 0.001973f
C8377 VDPWR.n2111 VSS 0.003404f
C8378 VDPWR.n2112 VSS 0.003083f
C8379 VDPWR.n2113 VSS 0.002629f
C8380 VDPWR.n2114 VSS 0.00352f
C8381 VDPWR.n2115 VSS 0.015143f
C8382 VDPWR.n2116 VSS 0.052403f
C8383 VDPWR.t1238 VSS 0.072626f
C8384 VDPWR.n2117 VSS 0.040608f
C8385 VDPWR.n2118 VSS 0.010509f
C8386 VDPWR.n2119 VSS 0.002048f
C8387 VDPWR.n2120 VSS 0.002048f
C8388 VDPWR.n2121 VSS 0.002944f
C8389 VDPWR.n2122 VSS 0.001973f
C8390 VDPWR.n2123 VSS 0.001579f
C8391 VDPWR.n2124 VSS 0.00352f
C8392 VDPWR.n2125 VSS 0.003404f
C8393 VDPWR.n2126 VSS 0.003083f
C8394 VDPWR.n2127 VSS 0.002117f
C8395 VDPWR.n2128 VSS 0.003008f
C8396 VDPWR.n2129 VSS 0.020793f
C8397 VDPWR.n2130 VSS 0.020793f
C8398 VDPWR.n2131 VSS 0.020115f
C8399 VDPWR.n2132 VSS 0.005888f
C8400 VDPWR.n2133 VSS 0.003488f
C8401 VDPWR.n2134 VSS 0.008742f
C8402 VDPWR.n2135 VSS 0.005612f
C8403 VDPWR.t641 VSS 0.005483f
C8404 VDPWR.n2136 VSS 0.006928f
C8405 VDPWR.n2137 VSS 0.011926f
C8406 VDPWR.n2138 VSS 0.005888f
C8407 VDPWR.n2139 VSS 0.003488f
C8408 VDPWR.n2140 VSS 0.005803f
C8409 VDPWR.t705 VSS 0.005483f
C8410 VDPWR.n2141 VSS 0.003947f
C8411 VDPWR.n2142 VSS 0.005756f
C8412 VDPWR.n2143 VSS 0.005344f
C8413 VDPWR.n2144 VSS 0.005888f
C8414 VDPWR.n2145 VSS 0.009361f
C8415 VDPWR.n2146 VSS 0.012758f
C8416 VDPWR.n2147 VSS 0.009777f
C8417 VDPWR.n2148 VSS 0.005888f
C8418 VDPWR.n2149 VSS 0.004544f
C8419 VDPWR.n2150 VSS 0.009361f
C8420 VDPWR.n2151 VSS 0.012758f
C8421 VDPWR.n2152 VSS 0.002048f
C8422 VDPWR.n2153 VSS 0.001973f
C8423 VDPWR.n2154 VSS 0.00224f
C8424 VDPWR.n2155 VSS 0.002752f
C8425 VDPWR.n2156 VSS 0.001973f
C8426 VDPWR.n2157 VSS 0.003083f
C8427 VDPWR.n2158 VSS 0.003404f
C8428 VDPWR.n2159 VSS 0.140809f
C8429 VDPWR.n2160 VSS 0.003404f
C8430 VDPWR.n2161 VSS 0.003083f
C8431 VDPWR.n2162 VSS 0.001973f
C8432 VDPWR.n2163 VSS 0.002944f
C8433 VDPWR.n2164 VSS 0.002048f
C8434 VDPWR.n2165 VSS 0.012342f
C8435 VDPWR.t642 VSS 0.005483f
C8436 VDPWR.n2166 VSS 0.006928f
C8437 VDPWR.n2167 VSS 0.006017f
C8438 VDPWR.n2168 VSS 0.002528f
C8439 VDPWR.n2169 VSS 0.003168f
C8440 VDPWR.n2170 VSS 0.00224f
C8441 VDPWR.n2171 VSS 0.006252f
C8442 VDPWR.t706 VSS 0.005503f
C8443 VDPWR.n2172 VSS 0.006241f
C8444 VDPWR.n2173 VSS 0.00232f
C8445 VDPWR.n2174 VSS 0.002016f
C8446 VDPWR.n2175 VSS 0.002944f
C8447 VDPWR.n2176 VSS 0.00168f
C8448 VDPWR.n2177 VSS 0.014269f
C8449 VDPWR.t1020 VSS 0.001867f
C8450 VDPWR.t259 VSS 0.001867f
C8451 VDPWR.n2178 VSS 0.004011f
C8452 VDPWR.t564 VSS 0.004984f
C8453 VDPWR.n2179 VSS 0.014116f
C8454 VDPWR.n2180 VSS 0.014701f
C8455 VDPWR.n2181 VSS 0.005344f
C8456 VDPWR.n2182 VSS 0.003488f
C8457 VDPWR.n2183 VSS 0.004416f
C8458 VDPWR.n2184 VSS 0.002878f
C8459 VDPWR.t433 VSS 0.005483f
C8460 VDPWR.n2185 VSS 0.003532f
C8461 VDPWR.n2186 VSS 0.008738f
C8462 VDPWR.n2187 VSS 0.004474f
C8463 VDPWR.n2188 VSS 0.006263f
C8464 VDPWR.n2189 VSS 0.005888f
C8465 VDPWR.n2190 VSS 0.005568f
C8466 VDPWR.n2191 VSS 0.003213f
C8467 VDPWR.n2192 VSS 0.033954f
C8468 VDPWR.n2193 VSS 0.003782f
C8469 VDPWR.n2194 VSS 0.008648f
C8470 VDPWR.t401 VSS 0.001867f
C8471 VDPWR.t423 VSS 0.001867f
C8472 VDPWR.n2195 VSS 0.003854f
C8473 VDPWR.n2196 VSS 0.008648f
C8474 VDPWR.n2197 VSS 0.002112f
C8475 VDPWR.n2198 VSS 0.005888f
C8476 VDPWR.t395 VSS 0.001867f
C8477 VDPWR.t399 VSS 0.0018f
C8478 VDPWR.n2199 VSS 0.003787f
C8479 VDPWR.n2200 VSS 0.00427f
C8480 VDPWR.t403 VSS 0.001867f
C8481 VDPWR.t413 VSS 0.001867f
C8482 VDPWR.n2201 VSS 0.003854f
C8483 VDPWR.n2202 VSS 0.008115f
C8484 VDPWR.t434 VSS 0.005483f
C8485 VDPWR.n2203 VSS 0.003762f
C8486 VDPWR.t407 VSS 0.001867f
C8487 VDPWR.t409 VSS 0.001867f
C8488 VDPWR.n2204 VSS 0.003854f
C8489 VDPWR.n2205 VSS 0.004861f
C8490 VDPWR.n2206 VSS 0.005888f
C8491 VDPWR.t737 VSS 0.005483f
C8492 VDPWR.n2207 VSS 0.00425f
C8493 VDPWR.t405 VSS 0.001867f
C8494 VDPWR.t415 VSS 0.001867f
C8495 VDPWR.n2208 VSS 0.003854f
C8496 VDPWR.t1173 VSS 0.072626f
C8497 VDPWR.n2209 VSS 0.033277f
C8498 VDPWR.t419 VSS 0.006558f
C8499 VDPWR.n2210 VSS 0.007607f
C8500 VDPWR.t728 VSS 0.004984f
C8501 VDPWR.n2211 VSS 0.006247f
C8502 VDPWR.n2212 VSS 0.008952f
C8503 VDPWR.n2213 VSS 0.002176f
C8504 VDPWR.n2214 VSS 0.00224f
C8505 VDPWR.n2215 VSS 0.007073f
C8506 VDPWR.n2216 VSS 0.004356f
C8507 VDPWR.n2217 VSS 0.004416f
C8508 VDPWR.n2218 VSS 0.005888f
C8509 VDPWR.n2219 VSS 0.005683f
C8510 VDPWR.n2220 VSS 0.004131f
C8511 VDPWR.n2221 VSS 0.008552f
C8512 VDPWR.n2222 VSS 0.006832f
C8513 VDPWR.n2223 VSS 0.005888f
C8514 VDPWR.n2224 VSS 0.005344f
C8515 VDPWR.n2225 VSS 0.002741f
C8516 VDPWR.n2226 VSS 0.002996f
C8517 VDPWR.n2227 VSS 0.003488f
C8518 VDPWR.n2228 VSS 0.005888f
C8519 VDPWR.n2229 VSS 0.005888f
C8520 VDPWR.n2230 VSS 0.006466f
C8521 VDPWR.n2231 VSS 0.008359f
C8522 VDPWR.n2232 VSS 0.004758f
C8523 VDPWR.n2233 VSS 0.005938f
C8524 VDPWR.n2234 VSS 0.003904f
C8525 VDPWR.n2235 VSS 0.001973f
C8526 VDPWR.n2236 VSS 0.00352f
C8527 VDPWR.n2237 VSS 0.001579f
C8528 VDPWR.n2238 VSS 0.001973f
C8529 VDPWR.n2239 VSS 0.003083f
C8530 VDPWR.n2240 VSS 0.002949f
C8531 VDPWR.n2241 VSS 0.002048f
C8532 VDPWR.n2242 VSS 0.005287f
C8533 VDPWR.n2243 VSS 0.00545f
C8534 VDPWR.n2244 VSS 0.002048f
C8535 VDPWR.n2245 VSS 0.002944f
C8536 VDPWR.n2246 VSS 0.001973f
C8537 VDPWR.n2247 VSS 0.003083f
C8538 VDPWR.n2248 VSS 0.003404f
C8539 VDPWR.n2249 VSS 0.140809f
C8540 VDPWR.n2250 VSS 0.116061f
C8541 VDPWR.n2251 VSS 0.281618f
C8542 VDPWR.n2252 VSS 0.281618f
C8543 VDPWR.n2253 VSS 0.281618f
C8544 VDPWR.n2254 VSS 0.167264f
C8545 VDPWR.n2255 VSS 0.116061f
C8546 VDPWR.n2256 VSS 0.140809f
C8547 VDPWR.n2257 VSS 0.003404f
C8548 VDPWR.n2258 VSS 0.00352f
C8549 VDPWR.n2259 VSS 0.00352f
C8550 VDPWR.n2260 VSS 0.001579f
C8551 VDPWR.n2261 VSS 0.001973f
C8552 VDPWR.n2262 VSS 0.001472f
C8553 VDPWR.n2263 VSS 7.36e-19
C8554 VDPWR.n2264 VSS 0.007329f
C8555 VDPWR.t591 VSS 0.005483f
C8556 VDPWR.n2265 VSS 0.011995f
C8557 VDPWR.n2266 VSS 0.020115f
C8558 VDPWR.n2267 VSS 0.015595f
C8559 VDPWR.n2268 VSS 0.005888f
C8560 VDPWR.n2269 VSS 0.004416f
C8561 VDPWR.n2270 VSS 0.008952f
C8562 VDPWR.n2271 VSS 0.004007f
C8563 VDPWR.n2272 VSS 0.004416f
C8564 VDPWR.n2273 VSS 0.005888f
C8565 VDPWR.n2274 VSS 0.006773f
C8566 VDPWR.n2275 VSS 0.004131f
C8567 VDPWR.n2276 VSS 0.008552f
C8568 VDPWR.n2277 VSS 0.005084f
C8569 VDPWR.n2278 VSS 0.005888f
C8570 VDPWR.n2279 VSS 0.005888f
C8571 VDPWR.n2280 VSS 0.005888f
C8572 VDPWR.n2281 VSS 0.006954f
C8573 VDPWR.n2282 VSS 0.008359f
C8574 VDPWR.n2283 VSS 0.004026f
C8575 VDPWR.t590 VSS 0.005483f
C8576 VDPWR.n2284 VSS 0.004291f
C8577 VDPWR.n2285 VSS 0.002441f
C8578 VDPWR.n2286 VSS 0.0048f
C8579 VDPWR.n2287 VSS 0.002405f
C8580 VDPWR.n2288 VSS 0.003083f
C8581 VDPWR.n2289 VSS 0.003404f
C8582 VDPWR.n2290 VSS 0.140809f
C8583 VDPWR.n2291 VSS 0.003404f
C8584 VDPWR.n2292 VSS 0.00352f
C8585 VDPWR.n2293 VSS 0.001579f
C8586 VDPWR.n2294 VSS 0.001973f
C8587 VDPWR.n2295 VSS 0.00288f
C8588 VDPWR.n2296 VSS 0.002048f
C8589 VDPWR.n2297 VSS 0.005287f
C8590 VDPWR.n2298 VSS 0.00545f
C8591 VDPWR.n2299 VSS 0.004672f
C8592 VDPWR.n2300 VSS 0.005888f
C8593 VDPWR.n2301 VSS 0.005888f
C8594 VDPWR.n2302 VSS 0.004962f
C8595 VDPWR.n2303 VSS 0.008648f
C8596 VDPWR.n2304 VSS 0.006263f
C8597 VDPWR.n2305 VSS 0.004474f
C8598 VDPWR.n2306 VSS 0.005888f
C8599 VDPWR.n2307 VSS 0.005888f
C8600 VDPWR.n2308 VSS 0.006418f
C8601 VDPWR.n2309 VSS 0.003953f
C8602 VDPWR.n2310 VSS 0.009049f
C8603 VDPWR.n2311 VSS 0.006938f
C8604 VDPWR.n2312 VSS 0.005344f
C8605 VDPWR.n2313 VSS 0.002016f
C8606 VDPWR.n2314 VSS 0.002016f
C8607 VDPWR.n2315 VSS 0.002963f
C8608 VDPWR.t738 VSS 0.005483f
C8609 VDPWR.n2316 VSS 0.00426f
C8610 VDPWR.n2317 VSS 0.016735f
C8611 VDPWR.n2318 VSS 0.00224f
C8612 VDPWR.n2319 VSS 5.48e-19
C8613 VDPWR.n2320 VSS 0.003083f
C8614 VDPWR.n2321 VSS 0.001973f
C8615 VDPWR.n2322 VSS 0.002944f
C8616 VDPWR.n2323 VSS 0.002048f
C8617 VDPWR.n2324 VSS 0.020115f
C8618 VDPWR.n2325 VSS 0.015595f
C8619 VDPWR.n2326 VSS 0.002048f
C8620 VDPWR.n2327 VSS 0.00224f
C8621 VDPWR.n2328 VSS 0.001973f
C8622 VDPWR.n2329 VSS 0.003083f
C8623 VDPWR.n2330 VSS 0.003404f
C8624 VDPWR.n2331 VSS 0.140809f
C8625 VDPWR.n2332 VSS 0.116061f
C8626 VDPWR.n2333 VSS 0.281618f
C8627 VDPWR.n2334 VSS 0.281618f
C8628 VDPWR.n2335 VSS 0.532156f
C8629 VDPWR.n2336 VSS 0.194931f
C8630 VDPWR.n2338 VSS 0.003432f
C8631 VDPWR.n2339 VSS 0.107527f
C8632 VDPWR.n2340 VSS 0.097681f
C8633 VDPWR.n2341 VSS 0.001579f
C8634 VDPWR.n2342 VSS 0.003054f
C8635 VDPWR.n2343 VSS 0.427843f
C8636 VDPWR.n2344 VSS 0.003054f
C8637 VDPWR.n2345 VSS 0.001973f
C8638 VDPWR.n2346 VSS 0.002949f
C8639 VDPWR.t802 VSS 0.001527f
C8640 VDPWR.t8 VSS 0.001527f
C8641 VDPWR.n2347 VSS 0.003322f
C8642 VDPWR.t1052 VSS 0.003924f
C8643 VDPWR.t374 VSS 0.002867f
C8644 VDPWR.n2348 VSS 0.010151f
C8645 VDPWR.n2349 VSS 0.005906f
C8646 VDPWR.n2350 VSS 0.005344f
C8647 VDPWR.t834 VSS 0.002741f
C8648 VDPWR.t1194 VSS 0.029301f
C8649 VDPWR.n2351 VSS 0.039775f
C8650 VDPWR.t353 VSS 0.0022f
C8651 VDPWR.t913 VSS 0.0022f
C8652 VDPWR.n2352 VSS 0.004485f
C8653 VDPWR.n2353 VSS 0.006511f
C8654 VDPWR.n2354 VSS 0.004416f
C8655 VDPWR.t296 VSS 0.001527f
C8656 VDPWR.t301 VSS 0.001527f
C8657 VDPWR.n2355 VSS 0.003394f
C8658 VDPWR.t21 VSS 0.002267f
C8659 VDPWR.t1050 VSS 0.002333f
C8660 VDPWR.n2356 VSS 0.005483f
C8661 VDPWR.t440 VSS 0.004984f
C8662 VDPWR.n2357 VSS 0.008777f
C8663 VDPWR.n2358 VSS 0.003008f
C8664 VDPWR.t1269 VSS 0.020799f
C8665 VDPWR.t389 VSS 0.00632f
C8666 VDPWR.n2359 VSS 0.005918f
C8667 VDPWR.n2360 VSS 0.001472f
C8668 VDPWR.n2361 VSS 0.002117f
C8669 VDPWR.n2362 VSS 0.001579f
C8670 VDPWR.n2363 VSS 0.001973f
C8671 VDPWR.n2364 VSS 0.001579f
C8672 VDPWR.n2365 VSS 0.002629f
C8673 VDPWR.t809 VSS 0.0018f
C8674 VDPWR.t806 VSS 0.0018f
C8675 VDPWR.n2366 VSS 0.003944f
C8676 VDPWR.n2367 VSS 0.00352f
C8677 VDPWR.t97 VSS 0.001527f
C8678 VDPWR.t808 VSS 0.001527f
C8679 VDPWR.n2368 VSS 0.003394f
C8680 VDPWR.n2369 VSS 0.001711f
C8681 VDPWR.t836 VSS 0.001527f
C8682 VDPWR.t141 VSS 0.001527f
C8683 VDPWR.n2370 VSS 0.003394f
C8684 VDPWR.t475 VSS 0.005024f
C8685 VDPWR.t1274 VSS 0.010664f
C8686 VDPWR.n2372 VSS 0.027341f
C8687 VDPWR.t476 VSS 0.005024f
C8688 VDPWR.n2373 VSS 0.014893f
C8689 VDPWR.t594 VSS 0.005024f
C8690 VDPWR.t1211 VSS 0.010664f
C8691 VDPWR.n2375 VSS 0.027341f
C8692 VDPWR.t595 VSS 0.005024f
C8693 VDPWR.n2376 VSS 0.014893f
C8694 VDPWR.n2377 VSS 0.012599f
C8695 VDPWR.n2378 VSS 0.003844f
C8696 VDPWR.n2379 VSS 0.002016f
C8697 VDPWR.n2380 VSS 0.001383f
C8698 VDPWR.n2381 VSS 0.009183f
C8699 VDPWR.n2382 VSS 0.0032f
C8700 VDPWR.n2383 VSS 0.002016f
C8701 VDPWR.n2384 VSS 0.004416f
C8702 VDPWR.n2385 VSS 0.001711f
C8703 VDPWR.n2386 VSS 0.012693f
C8704 VDPWR.n2387 VSS 8.61e-19
C8705 VDPWR.n2388 VSS 0.001792f
C8706 VDPWR.n2389 VSS 0.002368f
C8707 VDPWR.n2390 VSS 0.001973f
C8708 VDPWR.n2391 VSS 0.003054f
C8709 VDPWR.n2392 VSS 0.24535f
C8710 VDPWR.n2393 VSS 0.003054f
C8711 VDPWR.n2394 VSS 0.001973f
C8712 VDPWR.n2395 VSS 0.00288f
C8713 VDPWR.n2396 VSS 0.002048f
C8714 VDPWR.n2397 VSS 0.002847f
C8715 VDPWR.t439 VSS 0.004984f
C8716 VDPWR.n2398 VSS 0.004913f
C8717 VDPWR.n2399 VSS 0.018812f
C8718 VDPWR.n2400 VSS 0.011593f
C8719 VDPWR.n2401 VSS 0.014953f
C8720 VDPWR.n2402 VSS 0.004416f
C8721 VDPWR.n2403 VSS 0.002016f
C8722 VDPWR.n2404 VSS 0.005635f
C8723 VDPWR.n2405 VSS 0.008623f
C8724 VDPWR.n2406 VSS 0.008617f
C8725 VDPWR.n2407 VSS 0.005888f
C8726 VDPWR.n2408 VSS 0.004416f
C8727 VDPWR.n2409 VSS 0.00224f
C8728 VDPWR.n2410 VSS 0.001408f
C8729 VDPWR.t638 VSS 0.004984f
C8730 VDPWR.n2411 VSS 0.008777f
C8731 VDPWR.n2412 VSS 0.005906f
C8732 VDPWR.n2413 VSS 0.004416f
C8733 VDPWR.n2414 VSS 0.004416f
C8734 VDPWR.n2415 VSS 0.002016f
C8735 VDPWR.n2416 VSS 0.008233f
C8736 VDPWR.n2417 VSS 0.011294f
C8737 VDPWR.n2418 VSS 0.014953f
C8738 VDPWR.t1041 VSS 0.001036f
C8739 VDPWR.t357 VSS 0.001036f
C8740 VDPWR.n2419 VSS 0.002169f
C8741 VDPWR.t639 VSS 0.004984f
C8742 VDPWR.n2420 VSS 0.007433f
C8743 VDPWR.n2421 VSS 0.013464f
C8744 VDPWR.n2422 VSS 0.009073f
C8745 VDPWR.n2423 VSS 0.004544f
C8746 VDPWR.n2424 VSS 0.002949f
C8747 VDPWR.n2425 VSS 0.001888f
C8748 VDPWR.n2426 VSS 0.001973f
C8749 VDPWR.n2427 VSS 9.28e-19
C8750 VDPWR.n2428 VSS 0.001472f
C8751 VDPWR.n2429 VSS 7.36e-19
C8752 VDPWR.n2430 VSS 0.001782f
C8753 VDPWR.n2431 VSS 0.007807f
C8754 VDPWR.t474 VSS 0.052075f
C8755 VDPWR.t835 VSS 0.017547f
C8756 VDPWR.t140 VSS 0.01717f
C8757 VDPWR.t387 VSS 0.023208f
C8758 VDPWR.t96 VSS 0.031698f
C8759 VDPWR.t805 VSS 0.016604f
C8760 VDPWR.t807 VSS 0.013019f
C8761 VDPWR.t388 VSS 0.038302f
C8762 VDPWR.t167 VSS 0.037358f
C8763 VDPWR.t438 VSS 0.031132f
C8764 VDPWR.t20 VSS 0.01717f
C8765 VDPWR.t295 VSS 0.007358f
C8766 VDPWR.t1049 VSS 0.016604f
C8767 VDPWR.t300 VSS 0.017736f
C8768 VDPWR.t352 VSS 0.020755f
C8769 VDPWR.t912 VSS 0.026604f
C8770 VDPWR.t837 VSS 0.052453f
C8771 VDPWR.t637 VSS 0.005849f
C8772 VDPWR.t833 VSS 0.019245f
C8773 VDPWR.t1040 VSS 0.038491f
C8774 VDPWR.t356 VSS 0.027358f
C8775 VDPWR.t1051 VSS 0.017358f
C8776 VDPWR.t801 VSS 0.022453f
C8777 VDPWR.t7 VSS 0.043019f
C8778 VDPWR.t51 VSS 0.019057f
C8779 VDPWR.t870 VSS 0.016604f
C8780 VDPWR.t124 VSS 0.01566f
C8781 VDPWR.t126 VSS 0.017358f
C8782 VDPWR.t846 VSS 0.029245f
C8783 VDPWR.t733 VSS 0.031509f
C8784 VDPWR.t63 VSS 0.045849f
C8785 VDPWR.t159 VSS 0.022453f
C8786 VDPWR.t510 VSS 0.017358f
C8787 VDPWR.t670 VSS 0.103962f
C8788 VDPWR.t922 VSS 0.045849f
C8789 VDPWR.t223 VSS 0.017358f
C8790 VDPWR.t229 VSS 0.005849f
C8791 VDPWR.t297 VSS 0.025094f
C8792 VDPWR.t799 VSS 0.035849f
C8793 VDPWR.t227 VSS 0.021509f
C8794 VDPWR.t480 VSS 0.018868f
C8795 VDPWR.t324 VSS 0.02283f
C8796 VDPWR.n2432 VSS 0.053108f
C8797 VDPWR.n2433 VSS 0.022154f
C8798 VDPWR.t1255 VSS 0.029301f
C8799 VDPWR.t325 VSS 0.002741f
C8800 VDPWR.n2434 VSS 0.011294f
C8801 VDPWR.n2435 VSS 0.005888f
C8802 VDPWR.t228 VSS 0.001036f
C8803 VDPWR.t800 VSS 0.001036f
C8804 VDPWR.n2436 VSS 0.002169f
C8805 VDPWR.t482 VSS 0.004984f
C8806 VDPWR.n2437 VSS 0.008777f
C8807 VDPWR.t298 VSS 0.003924f
C8808 VDPWR.t230 VSS 0.002867f
C8809 VDPWR.n2438 VSS 0.010226f
C8810 VDPWR.n2439 VSS 0.002016f
C8811 VDPWR.n2440 VSS 0.003872f
C8812 VDPWR.t224 VSS 0.001527f
C8813 VDPWR.t923 VSS 0.001527f
C8814 VDPWR.n2441 VSS 0.003394f
C8815 VDPWR.n2442 VSS 0.002505f
C8816 VDPWR.n2443 VSS 0.001088f
C8817 VDPWR.n2444 VSS 0.001973f
C8818 VDPWR.n2445 VSS 0.001579f
C8819 VDPWR.n2446 VSS 0.003054f
C8820 VDPWR.n2447 VSS 0.001472f
C8821 VDPWR.n2448 VSS 0.002048f
C8822 VDPWR.n2449 VSS 0.002949f
C8823 VDPWR.t671 VSS 0.004984f
C8824 VDPWR.t511 VSS 0.005483f
C8825 VDPWR.n2450 VSS 0.011995f
C8826 VDPWR.n2451 VSS 0.003842f
C8827 VDPWR.n2452 VSS 0.003295f
C8828 VDPWR.t1182 VSS 0.029107f
C8829 VDPWR.n2453 VSS 0.015278f
C8830 VDPWR.n2454 VSS 0.015934f
C8831 VDPWR.n2455 VSS 0.003488f
C8832 VDPWR.t1264 VSS 0.072626f
C8833 VDPWR.n2456 VSS 0.040608f
C8834 VDPWR.n2457 VSS 0.004416f
C8835 VDPWR.t160 VSS 0.001527f
C8836 VDPWR.t64 VSS 0.001527f
C8837 VDPWR.n2458 VSS 0.003322f
C8838 VDPWR.t512 VSS 0.005501f
C8839 VDPWR.n2459 VSS 0.011323f
C8840 VDPWR.n2460 VSS 0.00425f
C8841 VDPWR.t127 VSS 0.001513f
C8842 VDPWR.t847 VSS 5.64e-19
C8843 VDPWR.n2461 VSS 0.006953f
C8844 VDPWR.t125 VSS 0.001527f
C8845 VDPWR.t52 VSS 0.001527f
C8846 VDPWR.n2462 VSS 0.003322f
C8847 VDPWR.n2463 VSS 0.008065f
C8848 VDPWR.n2464 VSS 9.32e-19
C8849 VDPWR.n2465 VSS 0.001973f
C8850 VDPWR.n2466 VSS 0.001472f
C8851 VDPWR.n2467 VSS 0.0024f
C8852 VDPWR.n2468 VSS 7.36e-19
C8853 VDPWR.n2469 VSS 0.001235f
C8854 VDPWR.n2470 VSS 0.015495f
C8855 VDPWR.t735 VSS 0.005058f
C8856 VDPWR.n2471 VSS 0.005913f
C8857 VDPWR.n2472 VSS 0.023007f
C8858 VDPWR.t1280 VSS 0.021124f
C8859 VDPWR.n2473 VSS 0.020912f
C8860 VDPWR.t734 VSS 0.004984f
C8861 VDPWR.n2474 VSS 0.005999f
C8862 VDPWR.n2475 VSS 0.00595f
C8863 VDPWR.n2476 VSS 0.003146f
C8864 VDPWR.n2477 VSS 0.00224f
C8865 VDPWR.n2478 VSS 0.006252f
C8866 VDPWR.n2479 VSS 0.007422f
C8867 VDPWR.n2480 VSS 0.013157f
C8868 VDPWR.n2481 VSS 0.005888f
C8869 VDPWR.n2482 VSS 0.004416f
C8870 VDPWR.n2483 VSS 0.004047f
C8871 VDPWR.n2484 VSS 0.008952f
C8872 VDPWR.t672 VSS 0.004984f
C8873 VDPWR.n2485 VSS 0.011445f
C8874 VDPWR.n2486 VSS 0.014578f
C8875 VDPWR.n2487 VSS 0.005888f
C8876 VDPWR.n2488 VSS 0.005888f
C8877 VDPWR.n2489 VSS 0.003904f
C8878 VDPWR.n2490 VSS 0.02068f
C8879 VDPWR.n2491 VSS 0.020136f
C8880 VDPWR.n2492 VSS 0.009831f
C8881 VDPWR.n2493 VSS 0.002048f
C8882 VDPWR.n2494 VSS 0.001973f
C8883 VDPWR.n2495 VSS 0.002112f
C8884 VDPWR.n2496 VSS 0.00288f
C8885 VDPWR.n2497 VSS 0.001973f
C8886 VDPWR.n2498 VSS 0.001579f
C8887 VDPWR.n2499 VSS 0.116061f
C8888 VDPWR.n2500 VSS 0.097057f
C8889 VDPWR.n2501 VSS 0.139727f
C8890 VDPWR.n2502 VSS 0.293684f
C8891 VDPWR.n2503 VSS 0.061977f
C8892 VDPWR.n2504 VSS 0.532156f
C8893 VDPWR.n2505 VSS 0.281618f
C8894 VDPWR.n2506 VSS 0.063151f
C8895 VDPWR.n2507 VSS 0.140809f
C8896 VDPWR.n2508 VSS 0.078917f
C8897 VDPWR.n2509 VSS 0.003054f
C8898 VDPWR.n2510 VSS 0.001477f
C8899 VDPWR.n2511 VSS 0.002944f
C8900 VDPWR.n2512 VSS 0.001711f
C8901 VDPWR.n2513 VSS 0.008968f
C8902 VDPWR.n2514 VSS 0.009333f
C8903 VDPWR.n2515 VSS 0.005043f
C8904 VDPWR.n2516 VSS 0.003488f
C8905 VDPWR.n2517 VSS 0.005888f
C8906 VDPWR.n2518 VSS 0.013609f
C8907 VDPWR.n2519 VSS 0.013968f
C8908 VDPWR.n2520 VSS 0.009073f
C8909 VDPWR.n2521 VSS 0.014953f
C8910 VDPWR.n2522 VSS 0.005344f
C8911 VDPWR.n2523 VSS 0.002016f
C8912 VDPWR.n2524 VSS 0.03255f
C8913 VDPWR.t481 VSS 0.004984f
C8914 VDPWR.n2525 VSS 0.008777f
C8915 VDPWR.n2526 VSS 0.005471f
C8916 VDPWR.n2527 VSS 0.00224f
C8917 VDPWR.n2528 VSS 0.00224f
C8918 VDPWR.n2529 VSS 0.003456f
C8919 VDPWR.n2530 VSS 0.001757f
C8920 VDPWR.n2531 VSS 0.007623f
C8921 VDPWR.n2532 VSS 0.002048f
C8922 VDPWR.n2533 VSS 0.0024f
C8923 VDPWR.n2534 VSS 0.001973f
C8924 VDPWR.n2535 VSS 0.001579f
C8925 VDPWR.n2536 VSS 0.081339f
C8926 VDPWR.n2537 VSS 0.107527f
C8927 VDPWR.n2538 VSS 0.116061f
C8928 VDPWR.n2539 VSS 0.532156f
C8929 VDPWR.n2540 VSS 0.194931f
C8930 VDPWR.n2541 VSS 0.00352f
C8931 VDPWR.n2542 VSS 0.001973f
C8932 VDPWR.n2543 VSS 0.00288f
C8933 VDPWR.n2544 VSS 0.005888f
C8934 VDPWR.t832 VSS 0.0018f
C8935 VDPWR.t321 VSS 0.0018f
C8936 VDPWR.n2545 VSS 0.004032f
C8937 VDPWR.t1144 VSS 0.0018f
C8938 VDPWR.t330 VSS 0.0018f
C8939 VDPWR.n2546 VSS 0.004032f
C8940 VDPWR.n2547 VSS 0.009337f
C8941 VDPWR.n2548 VSS 0.002048f
C8942 VDPWR.n2549 VSS 0.003054f
C8943 VDPWR.t707 VSS 0.005024f
C8944 VDPWR.t1179 VSS 0.010664f
C8945 VDPWR.n2551 VSS 0.027341f
C8946 VDPWR.t708 VSS 0.005024f
C8947 VDPWR.n2552 VSS 0.014893f
C8948 VDPWR.t490 VSS 0.005024f
C8949 VDPWR.t1278 VSS 0.010664f
C8950 VDPWR.n2554 VSS 0.027341f
C8951 VDPWR.t491 VSS 0.005024f
C8952 VDPWR.n2555 VSS 0.014893f
C8953 VDPWR.n2556 VSS 0.01227f
C8954 VDPWR.t720 VSS 0.004984f
C8955 VDPWR.t1176 VSS 0.020982f
C8956 VDPWR.n2558 VSS 0.036453f
C8957 VDPWR.t721 VSS 0.004984f
C8958 VDPWR.n2559 VSS 0.020917f
C8959 VDPWR.n2560 VSS 0.003844f
C8960 VDPWR.n2561 VSS 0.006902f
C8961 VDPWR.t499 VSS 0.004984f
C8962 VDPWR.t1276 VSS 0.020982f
C8963 VDPWR.n2563 VSS 0.036453f
C8964 VDPWR.t500 VSS 0.004984f
C8965 VDPWR.n2564 VSS 0.020917f
C8966 VDPWR.n2565 VSS 0.018023f
C8967 VDPWR.n2566 VSS 0.001133f
C8968 VDPWR.n2567 VSS 0.001757f
C8969 VDPWR.n2568 VSS 0.002048f
C8970 VDPWR.n2569 VSS 0.002629f
C8971 VDPWR.n2570 VSS 0.002368f
C8972 VDPWR.n2571 VSS 0.001973f
C8973 VDPWR.n2572 VSS 0.00352f
C8974 VDPWR.n2573 VSS 0.001579f
C8975 VDPWR.n2574 VSS 0.001579f
C8976 VDPWR.n2575 VSS 0.001973f
C8977 VDPWR.n2576 VSS 0.002944f
C8978 VDPWR.n2577 VSS 0.002048f
C8979 VDPWR.n2578 VSS 0.00187f
C8980 VDPWR.t830 VSS 0.002834f
C8981 VDPWR.t1145 VSS 0.002834f
C8982 VDPWR.n2579 VSS 0.002085f
C8983 VDPWR.n2580 VSS 0.005888f
C8984 VDPWR.t818 VSS 0.00135f
C8985 VDPWR.t794 VSS 0.002785f
C8986 VDPWR.n2581 VSS 0.00567f
C8987 VDPWR.t199 VSS 0.00135f
C8988 VDPWR.t201 VSS 0.002785f
C8989 VDPWR.n2582 VSS 0.00567f
C8990 VDPWR.n2583 VSS 0.002085f
C8991 VDPWR.n2584 VSS 0.005888f
C8992 VDPWR.t12 VSS 0.002776f
C8993 VDPWR.t264 VSS 0.002776f
C8994 VDPWR.t770 VSS 0.001152f
C8995 VDPWR.t787 VSS 0.001152f
C8996 VDPWR.n2585 VSS 0.002399f
C8997 VDPWR.t148 VSS 0.001152f
C8998 VDPWR.t784 VSS 0.001152f
C8999 VDPWR.n2586 VSS 0.002399f
C9000 VDPWR.n2587 VSS 0.011445f
C9001 VDPWR.n2588 VSS 0.001888f
C9002 VDPWR.n2589 VSS 0.001973f
C9003 VDPWR.n2590 VSS 0.001579f
C9004 VDPWR.n2591 VSS 0.001579f
C9005 VDPWR.n2592 VSS 0.001973f
C9006 VDPWR.n2593 VSS 0.002048f
C9007 VDPWR.n2594 VSS 0.00136f
C9008 VDPWR.t496 VSS 0.005024f
C9009 VDPWR.t1267 VSS 0.010664f
C9010 VDPWR.n2596 VSS 0.027341f
C9011 VDPWR.t497 VSS 0.005024f
C9012 VDPWR.n2597 VSS 0.014893f
C9013 VDPWR.n2598 VSS 9.28e-19
C9014 VDPWR.n2599 VSS 0.001973f
C9015 VDPWR.n2600 VSS 0.001472f
C9016 VDPWR.n2601 VSS 0.002944f
C9017 VDPWR.n2602 VSS 0.002048f
C9018 VDPWR.t319 VSS 0.0018f
C9019 VDPWR.t769 VSS 0.0018f
C9020 VDPWR.n2603 VSS 0.004047f
C9021 VDPWR.n2604 VSS 0.00224f
C9022 VDPWR.t317 VSS 0.00281f
C9023 VDPWR.n2605 VSS 0.001133f
C9024 VDPWR.n2606 VSS 0.005888f
C9025 VDPWR.t384 VSS 0.0018f
C9026 VDPWR.t1140 VSS 0.0018f
C9027 VDPWR.n2607 VSS 0.004032f
C9028 VDPWR.n2608 VSS 0.00519f
C9029 VDPWR.t382 VSS 0.00281f
C9030 VDPWR.t284 VSS 0.00135f
C9031 VDPWR.t376 VSS 0.002785f
C9032 VDPWR.n2609 VSS 0.00567f
C9033 VDPWR.n2610 VSS 0.002085f
C9034 VDPWR.n2611 VSS 0.005888f
C9035 VDPWR.t139 VSS 0.00135f
C9036 VDPWR.t1001 VSS 0.002785f
C9037 VDPWR.n2612 VSS 0.00567f
C9038 VDPWR.n2613 VSS 0.001349f
C9039 VDPWR.n2614 VSS 0.002048f
C9040 VDPWR.n2615 VSS 0.001973f
C9041 VDPWR.n2616 VSS 0.001579f
C9042 VDPWR.n2617 VSS 0.001579f
C9043 VDPWR.n2618 VSS 0.001973f
C9044 VDPWR.t82 VSS 0.001152f
C9045 VDPWR.t786 VSS 0.001152f
C9046 VDPWR.n2619 VSS 0.002399f
C9047 VDPWR.n2620 VSS 0.006924f
C9048 VDPWR.t35 VSS 0.002765f
C9049 VDPWR.n2621 VSS 0.001723f
C9050 VDPWR.n2622 VSS 0.007854f
C9051 VDPWR.t359 VSS 0.002333f
C9052 VDPWR.t193 VSS 0.002267f
C9053 VDPWR.n2623 VSS 0.005406f
C9054 VDPWR.n2624 VSS 0.004863f
C9055 VDPWR.t351 VSS 7.56e-19
C9056 VDPWR.t101 VSS 7.56e-19
C9057 VDPWR.n2625 VSS 0.00175f
C9058 VDPWR.t355 VSS 0.001513f
C9059 VDPWR.t1133 VSS 5.64e-19
C9060 VDPWR.n2626 VSS 0.006904f
C9061 VDPWR.n2627 VSS 0.009598f
C9062 VDPWR.t484 VSS 0.004984f
C9063 VDPWR.n2628 VSS 0.004577f
C9064 VDPWR.n2629 VSS 0.005906f
C9065 VDPWR.n2630 VSS 0.002176f
C9066 VDPWR.n2631 VSS 0.001984f
C9067 VDPWR.n2632 VSS 0.001612f
C9068 VDPWR.n2633 VSS 0.023712f
C9069 VDPWR.t1026 VSS 0.0022f
C9070 VDPWR.t99 VSS 0.0022f
C9071 VDPWR.n2634 VSS 0.004485f
C9072 VDPWR.n2635 VSS 0.006669f
C9073 VDPWR.t756 VSS 0.00112f
C9074 VDPWR.t33 VSS -0.001177f
C9075 VDPWR.n2636 VSS 0.007481f
C9076 VDPWR.n2637 VSS 0.005999f
C9077 VDPWR.n2638 VSS 0.005888f
C9078 VDPWR.n2639 VSS 0.004416f
C9079 VDPWR.n2640 VSS 0.002944f
C9080 VDPWR.n2641 VSS 0.001723f
C9081 VDPWR.t798 VSS 0.00112f
C9082 VDPWR.t791 VSS -0.001177f
C9083 VDPWR.n2642 VSS 0.007481f
C9084 VDPWR.n2643 VSS 0.006135f
C9085 VDPWR.n2644 VSS 0.003488f
C9086 VDPWR.n2645 VSS 0.005888f
C9087 VDPWR.n2646 VSS 0.005344f
C9088 VDPWR.t1030 VSS 7.56e-19
C9089 VDPWR.t222 VSS 7.56e-19
C9090 VDPWR.n2647 VSS 0.00175f
C9091 VDPWR.t144 VSS 0.001152f
C9092 VDPWR.t323 VSS 0.001152f
C9093 VDPWR.n2648 VSS 0.002399f
C9094 VDPWR.n2649 VSS 0.007139f
C9095 VDPWR.n2650 VSS 0.002944f
C9096 VDPWR.n2651 VSS 0.002048f
C9097 VDPWR.n2652 VSS 0.001973f
C9098 VDPWR.n2653 VSS 0.00288f
C9099 VDPWR.n2654 VSS 0.002112f
C9100 VDPWR.n2655 VSS 6.08e-19
C9101 VDPWR.n2656 VSS 0.00136f
C9102 VDPWR.n2657 VSS 0.020179f
C9103 VDPWR.n2658 VSS 0.001504f
C9104 VDPWR.n2659 VSS 0.001477f
C9105 VDPWR.n2660 VSS 0.003083f
C9106 VDPWR.n2661 VSS 0.003404f
C9107 VDPWR.n2662 VSS 0.00352f
C9108 VDPWR.n2663 VSS 0.00352f
C9109 VDPWR.n2664 VSS 0.003404f
C9110 VDPWR.n2665 VSS 0.003083f
C9111 VDPWR.n2666 VSS 0.002949f
C9112 VDPWR.n2667 VSS 0.005568f
C9113 VDPWR.t1161 VSS 0.002776f
C9114 VDPWR.n2668 VSS 0.005585f
C9115 VDPWR.n2669 VSS 0.00419f
C9116 VDPWR.n2670 VSS 0.00153f
C9117 VDPWR.n2671 VSS 0.002085f
C9118 VDPWR.n2672 VSS 0.005888f
C9119 VDPWR.n2673 VSS 0.005888f
C9120 VDPWR.n2674 VSS 0.005888f
C9121 VDPWR.n2675 VSS 0.001598f
C9122 VDPWR.n2676 VSS 0.004168f
C9123 VDPWR.n2677 VSS 0.004846f
C9124 VDPWR.n2678 VSS 0.001281f
C9125 VDPWR.n2679 VSS 0.001995f
C9126 VDPWR.n2680 VSS 0.005888f
C9127 VDPWR.n2681 VSS 0.005888f
C9128 VDPWR.n2682 VSS 0.004416f
C9129 VDPWR.n2683 VSS 0.001847f
C9130 VDPWR.n2684 VSS 0.005401f
C9131 VDPWR.t489 VSS 0.074905f
C9132 VDPWR.t498 VSS 0.09f
C9133 VDPWR.t831 VSS 0.040943f
C9134 VDPWR.t320 VSS 0.055472f
C9135 VDPWR.t829 VSS 0.061132f
C9136 VDPWR.t152 VSS 0.037358f
C9137 VDPWR.t150 VSS 0.033774f
C9138 VDPWR.t198 VSS 0.04283f
C9139 VDPWR.t200 VSS 0.04434f
C9140 VDPWR.t149 VSS 0.037358f
C9141 VDPWR.t151 VSS 0.033962f
C9142 VDPWR.t11 VSS 0.051509f
C9143 VDPWR.t147 VSS 0.051321f
C9144 VDPWR.t783 VSS 0.024906f
C9145 VDPWR.t318 VSS 0.031509f
C9146 VDPWR.t495 VSS 0.015849f
C9147 VDPWR.t768 VSS 0.020566f
C9148 VDPWR.t914 VSS 0.029245f
C9149 VDPWR.t483 VSS 0.015849f
C9150 VDPWR.t354 VSS 0.026038f
C9151 VDPWR.t1132 VSS 0.034717f
C9152 VDPWR.t192 VSS 0.01717f
C9153 VDPWR.t100 VSS 0.013774f
C9154 VDPWR.t358 VSS 0.015849f
C9155 VDPWR.t350 VSS 0.017736f
C9156 VDPWR.t98 VSS 0.017547f
C9157 VDPWR.t755 VSS 0.018113f
C9158 VDPWR.t1025 VSS 0.017924f
C9159 VDPWR.t32 VSS 0.018113f
C9160 VDPWR.t220 VSS 0.035472f
C9161 VDPWR.t790 VSS 0.036415f
C9162 VDPWR.t785 VSS 0.009623f
C9163 VDPWR.t797 VSS 0.015849f
C9164 VDPWR.t81 VSS 0.017547f
C9165 VDPWR.t221 VSS 0.018113f
C9166 VDPWR.t1029 VSS 0.021698f
C9167 VDPWR.t34 VSS 0.017358f
C9168 VDPWR.t816 VSS 0.009057f
C9169 VDPWR.t322 VSS 0.017924f
C9170 VDPWR.t80 VSS 0.035283f
C9171 VDPWR.t1000 VSS 0.035472f
C9172 VDPWR.t1160 VSS 0.024906f
C9173 VDPWR.t138 VSS 0.016038f
C9174 VDPWR.t766 VSS 0.017924f
C9175 VDPWR.t83 VSS 0.017924f
C9176 VDPWR.t143 VSS 0.015849f
C9177 VDPWR.t817 VSS 0.019434f
C9178 VDPWR.t375 VSS 0.021509f
C9179 VDPWR.t381 VSS 0.024906f
C9180 VDPWR.t283 VSS 0.032075f
C9181 VDPWR.t142 VSS 0.025472f
C9182 VDPWR.t1139 VSS 0.015849f
C9183 VDPWR.t767 VSS 0.015849f
C9184 VDPWR.t383 VSS 0.021509f
C9185 VDPWR.t316 VSS 0.028302f
C9186 VDPWR.n2685 VSS 0.031563f
C9187 VDPWR.n2686 VSS 0.010857f
C9188 VDPWR.n2687 VSS 0.014434f
C9189 VDPWR.n2688 VSS 0.002528f
C9190 VDPWR.n2689 VSS 0.002949f
C9191 VDPWR.n2690 VSS 0.003083f
C9192 VDPWR.n2691 VSS 0.003404f
C9193 VDPWR.n2692 VSS 0.00352f
C9194 VDPWR.n2693 VSS 0.00352f
C9195 VDPWR.n2694 VSS 0.003404f
C9196 VDPWR.n2695 VSS 0.003083f
C9197 VDPWR.n2696 VSS 0.002949f
C9198 VDPWR.n2697 VSS 0.004544f
C9199 VDPWR.n2698 VSS 0.005888f
C9200 VDPWR.n2699 VSS 0.001349f
C9201 VDPWR.n2700 VSS 0.009459f
C9202 VDPWR.n2701 VSS 0.00187f
C9203 VDPWR.n2702 VSS 0.005888f
C9204 VDPWR.n2703 VSS 0.005888f
C9205 VDPWR.n2704 VSS 0.005888f
C9206 VDPWR.n2705 VSS 0.002085f
C9207 VDPWR.n2706 VSS 0.001598f
C9208 VDPWR.n2707 VSS 0.007769f
C9209 VDPWR.n2708 VSS 0.00153f
C9210 VDPWR.n2709 VSS 0.005888f
C9211 VDPWR.n2710 VSS 0.005888f
C9212 VDPWR.n2711 VSS 0.005888f
C9213 VDPWR.n2712 VSS 0.002085f
C9214 VDPWR.n2713 VSS 0.001496f
C9215 VDPWR.n2714 VSS 0.011469f
C9216 VDPWR.n2715 VSS 0.003008f
C9217 VDPWR.n2716 VSS 0.002117f
C9218 VDPWR.n2717 VSS 0.003054f
C9219 VDPWR.n2718 VSS 0.003432f
C9220 VDPWR.n2719 VSS 0.128008f
C9221 VDPWR.n2720 VSS 0.00352f
C9222 VDPWR.n2721 VSS 0.007212f
C9223 VDPWR.n2722 VSS 0.001579f
C9224 VDPWR.n2723 VSS 0.001579f
C9225 VDPWR.n2724 VSS 0.001973f
C9226 VDPWR.n2725 VSS 0.002944f
C9227 VDPWR.n2726 VSS 0.016028f
C9228 VDPWR.t1204 VSS 0.037597f
C9229 VDPWR.n2727 VSS 0.067773f
C9230 VDPWR.t572 VSS 0.004984f
C9231 VDPWR.n2728 VSS 0.016028f
C9232 VDPWR.t625 VSS 0.005024f
C9233 VDPWR.t1218 VSS 0.010664f
C9234 VDPWR.n2730 VSS 0.027341f
C9235 VDPWR.t626 VSS 0.005024f
C9236 VDPWR.n2731 VSS 0.014893f
C9237 VDPWR.t722 VSS 0.005024f
C9238 VDPWR.t1277 VSS 0.010664f
C9239 VDPWR.n2733 VSS 0.027341f
C9240 VDPWR.t723 VSS 0.005024f
C9241 VDPWR.n2734 VSS 0.014893f
C9242 VDPWR.n2735 VSS 0.012599f
C9243 VDPWR.n2736 VSS 0.003844f
C9244 VDPWR.n2737 VSS 0.00224f
C9245 VDPWR.n2738 VSS 0.001428f
C9246 VDPWR.n2739 VSS 0.017613f
C9247 VDPWR.t588 VSS 0.004984f
C9248 VDPWR.n2740 VSS 0.030163f
C9249 VDPWR.t1231 VSS 0.028799f
C9250 VDPWR.n2741 VSS 0.019432f
C9251 VDPWR.n2742 VSS 0.00833f
C9252 VDPWR.t587 VSS 0.004984f
C9253 VDPWR.n2743 VSS 0.003892f
C9254 VDPWR.n2744 VSS 0.004088f
C9255 VDPWR.n2745 VSS 0.002272f
C9256 VDPWR.n2746 VSS 0.005f
C9257 VDPWR.n2747 VSS 9.28e-19
C9258 VDPWR.n2748 VSS 0.00176f
C9259 VDPWR.n2749 VSS 0.021585f
C9260 VDPWR.n2750 VSS 0.002048f
C9261 VDPWR.n2751 VSS 0.002368f
C9262 VDPWR.n2752 VSS 0.001973f
C9263 VDPWR.n2753 VSS 0.003083f
C9264 VDPWR.n2754 VSS 0.003404f
C9265 VDPWR.n2755 VSS 0.128862f
C9266 VDPWR.n2756 VSS 0.003404f
C9267 VDPWR.n2757 VSS 0.003083f
C9268 VDPWR.n2758 VSS 0.001477f
C9269 VDPWR.n2759 VSS 6.08e-19
C9270 VDPWR.n2760 VSS 0.013021f
C9271 VDPWR.n2761 VSS 0.021375f
C9272 VDPWR.t573 VSS 0.004984f
C9273 VDPWR.n2762 VSS 0.008777f
C9274 VDPWR.n2763 VSS 0.005754f
C9275 VDPWR.n2764 VSS 0.003488f
C9276 VDPWR.n2765 VSS 0.004416f
C9277 VDPWR.n2766 VSS 0.005888f
C9278 VDPWR.n2767 VSS 0.00245f
C9279 VDPWR.n2768 VSS 0.003286f
C9280 VDPWR.t268 VSS 0.004259f
C9281 VDPWR.n2769 VSS 0.00392f
C9282 VDPWR.t969 VSS 0.001036f
C9283 VDPWR.n2770 VSS 0.002948f
C9284 VDPWR.n2771 VSS 0.005781f
C9285 VDPWR.t1113 VSS 0.001867f
C9286 VDPWR.t1115 VSS 0.001867f
C9287 VDPWR.n2772 VSS 0.003889f
C9288 VDPWR.n2773 VSS 0.006022f
C9289 VDPWR.n2774 VSS 0.001365f
C9290 VDPWR.n2775 VSS 0.005888f
C9291 VDPWR.t867 VSS 0.001148f
C9292 VDPWR.t386 VSS 7.56e-19
C9293 VDPWR.n2776 VSS 0.001983f
C9294 VDPWR.n2777 VSS 0.004651f
C9295 VDPWR.n2778 VSS 0.005888f
C9296 VDPWR.n2779 VSS 0.003488f
C9297 VDPWR.n2780 VSS 0.001306f
C9298 VDPWR.t1127 VSS 0.001867f
C9299 VDPWR.t1117 VSS 0.001867f
C9300 VDPWR.n2781 VSS 0.003889f
C9301 VDPWR.n2782 VSS 0.007282f
C9302 VDPWR.t263 VSS 0.002867f
C9303 VDPWR.t361 VSS 0.003924f
C9304 VDPWR.n2783 VSS 0.010151f
C9305 VDPWR.n2784 VSS 0.007557f
C9306 VDPWR.n2785 VSS 0.001096f
C9307 VDPWR.n2786 VSS 0.005888f
C9308 VDPWR.n2787 VSS 0.004544f
C9309 VDPWR.n2788 VSS 0.001353f
C9310 VDPWR.n2789 VSS 0.001703f
C9311 VDPWR.n2790 VSS 0.005793f
C9312 VDPWR.n2791 VSS 0.006683f
C9313 VDPWR.t1101 VSS 0.001867f
C9314 VDPWR.t1111 VSS 0.001867f
C9315 VDPWR.n2792 VSS 0.003854f
C9316 VDPWR.t162 VSS 0.002741f
C9317 VDPWR.n2793 VSS 0.004148f
C9318 VDPWR.n2794 VSS 0.005921f
C9319 VDPWR.n2795 VSS 0.001563f
C9320 VDPWR.n2796 VSS 0.001259f
C9321 VDPWR.n2797 VSS 0.002048f
C9322 VDPWR.n2798 VSS 0.001579f
C9323 VDPWR.n2799 VSS 0.001973f
C9324 VDPWR.n2800 VSS 0.00224f
C9325 VDPWR.n2801 VSS 0.002752f
C9326 VDPWR.n2802 VSS 0.001973f
C9327 VDPWR.n2803 VSS 0.003083f
C9328 VDPWR.n2804 VSS 0.003404f
C9329 VDPWR.n2805 VSS 0.128862f
C9330 VDPWR.n2806 VSS 0.003404f
C9331 VDPWR.n2807 VSS 0.003083f
C9332 VDPWR.n2808 VSS 0.002949f
C9333 VDPWR.n2809 VSS 0.002528f
C9334 VDPWR.n2810 VSS 0.00224f
C9335 VDPWR.t624 VSS 0.051698f
C9336 VDPWR.t586 VSS 0.074717f
C9337 VDPWR.t571 VSS 0.046604f
C9338 VDPWR.t900 VSS 0.022453f
C9339 VDPWR.t954 VSS 0.028868f
C9340 VDPWR.t267 VSS 0.026604f
C9341 VDPWR.t1118 VSS 0.019623f
C9342 VDPWR.t1112 VSS 0.030189f
C9343 VDPWR.t968 VSS 0.016226f
C9344 VDPWR.t1114 VSS 0.016604f
C9345 VDPWR.t866 VSS 0.016226f
C9346 VDPWR.t1130 VSS 0.018113f
C9347 VDPWR.t1122 VSS 0.016604f
C9348 VDPWR.t385 VSS 0.012641f
C9349 VDPWR.t1126 VSS 0.019811f
C9350 VDPWR.t1116 VSS 0.019623f
C9351 VDPWR.t262 VSS 0.016226f
C9352 VDPWR.t1120 VSS 0.028868f
C9353 VDPWR.t1124 VSS 0.01849f
C9354 VDPWR.t360 VSS 0.016226f
C9355 VDPWR.t1128 VSS 0.016226f
C9356 VDPWR.t1042 VSS 0.016226f
C9357 VDPWR.t1102 VSS 0.019623f
C9358 VDPWR.t225 VSS 0.016226f
C9359 VDPWR.t1100 VSS 0.018868f
C9360 VDPWR.t161 VSS 0.016226f
C9361 VDPWR.t1110 VSS 0.012264f
C9362 VDPWR.t1104 VSS 0.014151f
C9363 VDPWR.t444 VSS 0.052075f
C9364 VDPWR.t462 VSS 0.098679f
C9365 VDPWR.t687 VSS 0.057736f
C9366 VDPWR.t1044 VSS 0.02566f
C9367 VDPWR.t872 VSS 0.039811f
C9368 VDPWR.t390 VSS 0.024906f
C9369 VDPWR.t153 VSS 0.039811f
C9370 VDPWR.t977 VSS 0.027547f
C9371 VDPWR.t804 VSS 0.033962f
C9372 VDPWR.t155 VSS 0.037358f
C9373 VDPWR.t1053 VSS 0.04434f
C9374 VDPWR.t920 VSS 0.033774f
C9375 VDPWR.t714 VSS 0.017924f
C9376 VDPWR.t156 VSS 0.024906f
C9377 VDPWR.t803 VSS 0.037358f
C9378 VDPWR.t812 VSS 0.061132f
C9379 VDPWR.t157 VSS 0.055472f
C9380 VDPWR.t810 VSS 0.023396f
C9381 VDPWR.n2811 VSS 0.038158f
C9382 VDPWR.t1141 VSS 0.029245f
C9383 VDPWR.t501 VSS 0.01849f
C9384 VDPWR.t22 VSS 0.018113f
C9385 VDPWR.t194 VSS 0.039057f
C9386 VDPWR.t14 VSS 0.036981f
C9387 VDPWR.t795 VSS 0.037358f
C9388 VDPWR.t377 VSS 0.013585f
C9389 VDPWR.t1143 VSS 0.015849f
C9390 VDPWR.t53 VSS 0.018113f
C9391 VDPWR.t308 VSS 0.039623f
C9392 VDPWR.t379 VSS 0.042641f
C9393 VDPWR.t362 VSS 0.021509f
C9394 VDPWR.t828 VSS 0.021321f
C9395 VDPWR.t1006 VSS 0.013019f
C9396 VDPWR.t986 VSS 0.020755f
C9397 VDPWR.t190 VSS 0.026792f
C9398 VDPWR.t364 VSS 0.022453f
C9399 VDPWR.t299 VSS 0.016038f
C9400 VDPWR.t231 VSS 0.017736f
C9401 VDPWR.t92 VSS 0.019434f
C9402 VDPWR.t983 VSS 0.022075f
C9403 VDPWR.t827 VSS 0.028868f
C9404 VDPWR.t1047 VSS 0.016038f
C9405 VDPWR.t1134 VSS 0.020755f
C9406 VDPWR.t1148 VSS 0.033962f
C9407 VDPWR.t366 VSS 0.019811f
C9408 VDPWR.t984 VSS 0.00566f
C9409 VDPWR.t1158 VSS 0.017547f
C9410 VDPWR.t773 VSS 0.025472f
C9411 VDPWR.t775 VSS 0.01717f
C9412 VDPWR.t331 VSS 0.016226f
C9413 VDPWR.t781 VSS 0.016604f
C9414 VDPWR.t16 VSS 0.00717f
C9415 VDPWR.t777 VSS 0.01717f
C9416 VDPWR.t1108 VSS 0.02434f
C9417 VDPWR.t1106 VSS 0.03f
C9418 VDPWR.n2812 VSS 0.019299f
C9419 VDPWR.n2813 VSS 0.011327f
C9420 VDPWR.n2814 VSS 0.00598f
C9421 VDPWR.t1109 VSS 0.001867f
C9422 VDPWR.t778 VSS 0.001867f
C9423 VDPWR.n2815 VSS 0.004076f
C9424 VDPWR.n2816 VSS 0.006757f
C9425 VDPWR.n2817 VSS 0.001703f
C9426 VDPWR.n2818 VSS 0.004416f
C9427 VDPWR.n2819 VSS 0.003744f
C9428 VDPWR.n2820 VSS 0.002016f
C9429 VDPWR.n2821 VSS 0.001213f
C9430 VDPWR.t17 VSS 0.001527f
C9431 VDPWR.t332 VSS 0.001527f
C9432 VDPWR.n2822 VSS 0.003394f
C9433 VDPWR.t782 VSS 0.001867f
C9434 VDPWR.t776 VSS 0.001867f
C9435 VDPWR.n2823 VSS 0.004071f
C9436 VDPWR.n2824 VSS 0.014462f
C9437 VDPWR.n2825 VSS 0.005344f
C9438 VDPWR.n2826 VSS 0.004416f
C9439 VDPWR.n2827 VSS 0.002016f
C9440 VDPWR.t774 VSS 0.006972f
C9441 VDPWR.n2828 VSS 0.008825f
C9442 VDPWR.t1159 VSS 0.001152f
C9443 VDPWR.t985 VSS 0.001152f
C9444 VDPWR.n2829 VSS 0.002399f
C9445 VDPWR.n2830 VSS 0.006436f
C9446 VDPWR.n2831 VSS 0.002048f
C9447 VDPWR.n2832 VSS 0.005312f
C9448 VDPWR.n2833 VSS 0.005568f
C9449 VDPWR.n2834 VSS 0.005721f
C9450 VDPWR.t1048 VSS 0.002195f
C9451 VDPWR.t93 VSS 0.002658f
C9452 VDPWR.n2835 VSS 0.006308f
C9453 VDPWR.n2836 VSS 0.003819f
C9454 VDPWR.n2837 VSS 0.001702f
C9455 VDPWR.n2838 VSS 0.002048f
C9456 VDPWR.n2839 VSS 0.002048f
C9457 VDPWR.n2840 VSS 0.002944f
C9458 VDPWR.n2841 VSS 0.001973f
C9459 VDPWR.n2842 VSS 0.003083f
C9460 VDPWR.n2843 VSS 0.003404f
C9461 VDPWR.n2844 VSS 0.128862f
C9462 VDPWR.n2845 VSS 0.003404f
C9463 VDPWR.n2846 VSS 0.003083f
C9464 VDPWR.n2847 VSS 0.001973f
C9465 VDPWR.n2848 VSS 0.002112f
C9466 VDPWR.n2849 VSS 0.002048f
C9467 VDPWR.n2850 VSS 0.002024f
C9468 VDPWR.t232 VSS 0.002785f
C9469 VDPWR.t191 VSS 0.00135f
C9470 VDPWR.n2851 VSS 0.00567f
C9471 VDPWR.t365 VSS 0.002864f
C9472 VDPWR.n2852 VSS 0.008079f
C9473 VDPWR.n2853 VSS 0.004349f
C9474 VDPWR.n2854 VSS 0.001598f
C9475 VDPWR.n2855 VSS 0.003904f
C9476 VDPWR.n2856 VSS 0.004416f
C9477 VDPWR.n2857 VSS 0.002016f
C9478 VDPWR.n2858 VSS 0.00187f
C9479 VDPWR.t363 VSS 0.001372f
C9480 VDPWR.t1007 VSS 0.002267f
C9481 VDPWR.n2859 VSS 0.006283f
C9482 VDPWR.n2860 VSS 0.007702f
C9483 VDPWR.n2861 VSS 7.82e-19
C9484 VDPWR.n2862 VSS 0.005888f
C9485 VDPWR.n2863 VSS 0.005888f
C9486 VDPWR.n2864 VSS 0.005888f
C9487 VDPWR.t309 VSS 0.007351f
C9488 VDPWR.n2865 VSS 0.006963f
C9489 VDPWR.n2866 VSS 0.005167f
C9490 VDPWR.n2867 VSS 0.001133f
C9491 VDPWR.n2868 VSS 0.001179f
C9492 VDPWR.n2869 VSS 0.004416f
C9493 VDPWR.n2870 VSS 0.002944f
C9494 VDPWR.n2871 VSS 0.001089f
C9495 VDPWR.t15 VSS 0.004259f
C9496 VDPWR.t195 VSS 0.001036f
C9497 VDPWR.n2872 VSS 0.002948f
C9498 VDPWR.n2873 VSS 0.00392f
C9499 VDPWR.n2874 VSS 0.002688f
C9500 VDPWR.n2875 VSS 0.003005f
C9501 VDPWR.n2876 VSS 0.00224f
C9502 VDPWR.n2877 VSS 0.00224f
C9503 VDPWR.n2878 VSS 0.001973f
C9504 VDPWR.n2879 VSS 0.003404f
C9505 VDPWR.n2880 VSS 0.003083f
C9506 VDPWR.n2881 VSS 0.002757f
C9507 VDPWR.n2882 VSS 0.002176f
C9508 VDPWR.n2883 VSS 0.003702f
C9509 VDPWR.t502 VSS 0.004984f
C9510 VDPWR.n2884 VSS 0.004913f
C9511 VDPWR.n2885 VSS 0.018812f
C9512 VDPWR.n2886 VSS 0.011593f
C9513 VDPWR.t23 VSS 0.001148f
C9514 VDPWR.t1142 VSS 7.56e-19
C9515 VDPWR.n2887 VSS 0.00196f
C9516 VDPWR.n2888 VSS 0.005471f
C9517 VDPWR.t503 VSS 0.004984f
C9518 VDPWR.n2889 VSS 0.008609f
C9519 VDPWR.n2890 VSS 0.011129f
C9520 VDPWR.n2891 VSS 0.007897f
C9521 VDPWR.n2892 VSS 0.002048f
C9522 VDPWR.n2893 VSS 0.002944f
C9523 VDPWR.n2894 VSS 0.001973f
C9524 VDPWR.n2895 VSS 0.001579f
C9525 VDPWR.n2896 VSS 0.00352f
C9526 VDPWR.n2897 VSS 0.003404f
C9527 VDPWR.n2898 VSS 0.003083f
C9528 VDPWR.n2899 VSS 5.48e-19
C9529 VDPWR.n2900 VSS 0.00224f
C9530 VDPWR.n2901 VSS 0.002272f
C9531 VDPWR.n2902 VSS 0.001642f
C9532 VDPWR.t715 VSS 0.005483f
C9533 VDPWR.n2903 VSS 8.72e-19
C9534 VDPWR.n2904 VSS 0.003023f
C9535 VDPWR.n2905 VSS 0.004416f
C9536 VDPWR.n2906 VSS 0.005888f
C9537 VDPWR.n2907 VSS 0.007099f
C9538 VDPWR.n2908 VSS 0.004558f
C9539 VDPWR.n2909 VSS 0.008069f
C9540 VDPWR.n2910 VSS 0.00484f
C9541 VDPWR.n2911 VSS 0.005888f
C9542 VDPWR.n2912 VSS 0.005888f
C9543 VDPWR.n2913 VSS 0.005445f
C9544 VDPWR.n2914 VSS 0.007422f
C9545 VDPWR.t921 VSS 0.00135f
C9546 VDPWR.t1054 VSS 0.002785f
C9547 VDPWR.n2915 VSS 0.00567f
C9548 VDPWR.n2916 VSS 0.007073f
C9549 VDPWR.n2917 VSS 0.005445f
C9550 VDPWR.n2918 VSS 0.005888f
C9551 VDPWR.n2919 VSS 0.005888f
C9552 VDPWR.n2920 VSS 0.004672f
C9553 VDPWR.n2921 VSS 0.007422f
C9554 VDPWR.n2922 VSS 0.007422f
C9555 VDPWR.n2923 VSS 0.00718f
C9556 VDPWR.n2924 VSS 0.002048f
C9557 VDPWR.n2925 VSS 0.001579f
C9558 VDPWR.n2926 VSS 0.001973f
C9559 VDPWR.n2927 VSS 0.002112f
C9560 VDPWR.n2928 VSS 0.00288f
C9561 VDPWR.n2929 VSS 0.001973f
C9562 VDPWR.n2930 VSS 0.003083f
C9563 VDPWR.n2931 VSS 0.003404f
C9564 VDPWR.n2932 VSS 0.128862f
C9565 VDPWR.n2933 VSS 0.003404f
C9566 VDPWR.n2934 VSS 0.003083f
C9567 VDPWR.n2935 VSS 0.002405f
C9568 VDPWR.n2936 VSS 0.001504f
C9569 VDPWR.n2937 VSS 9.22e-19
C9570 VDPWR.n2938 VSS 0.005576f
C9571 VDPWR.n2939 VSS 0.002784f
C9572 VDPWR.t688 VSS 0.005483f
C9573 VDPWR.n2940 VSS 0.00426f
C9574 VDPWR.n2941 VSS 0.00355f
C9575 VDPWR.n2942 VSS 0.005888f
C9576 VDPWR.n2943 VSS 0.003488f
C9577 VDPWR.n2944 VSS 0.007341f
C9578 VDPWR.t873 VSS 0.007047f
C9579 VDPWR.t1187 VSS 0.072626f
C9580 VDPWR.n2945 VSS 0.033681f
C9581 VDPWR.n2946 VSS 0.011895f
C9582 VDPWR.n2947 VSS 0.003953f
C9583 VDPWR.n2948 VSS 0.004416f
C9584 VDPWR.n2949 VSS 0.005888f
C9585 VDPWR.n2950 VSS 0.003456f
C9586 VDPWR.n2951 VSS 0.007073f
C9587 VDPWR.t463 VSS 0.004984f
C9588 VDPWR.n2952 VSS 0.011445f
C9589 VDPWR.n2953 VSS 0.008952f
C9590 VDPWR.n2954 VSS 0.004416f
C9591 VDPWR.n2955 VSS 0.005888f
C9592 VDPWR.n2956 VSS 0.005888f
C9593 VDPWR.n2957 VSS 0.020793f
C9594 VDPWR.n2958 VSS 0.020793f
C9595 VDPWR.t464 VSS 0.004984f
C9596 VDPWR.t689 VSS 0.005483f
C9597 VDPWR.n2959 VSS 0.011995f
C9598 VDPWR.n2960 VSS 0.020115f
C9599 VDPWR.n2961 VSS 0.005696f
C9600 VDPWR.n2962 VSS 7.36e-19
C9601 VDPWR.n2963 VSS 0.002949f
C9602 VDPWR.n2964 VSS 0.003083f
C9603 VDPWR.n2965 VSS 0.001579f
C9604 VDPWR.n2966 VSS 0.001973f
C9605 VDPWR.n2967 VSS 0.001472f
C9606 VDPWR.n2968 VSS 0.002944f
C9607 VDPWR.n2969 VSS 0.002048f
C9608 VDPWR.t445 VSS 0.005024f
C9609 VDPWR.t1253 VSS 0.010664f
C9610 VDPWR.n2971 VSS 0.027341f
C9611 VDPWR.t446 VSS 0.005024f
C9612 VDPWR.n2972 VSS 0.014893f
C9613 VDPWR.n2973 VSS 0.012551f
C9614 VDPWR.n2974 VSS 0.001376f
C9615 VDPWR.n2975 VSS 0.002885f
C9616 VDPWR.n2976 VSS 0.002112f
C9617 VDPWR.n2977 VSS 0.001973f
C9618 VDPWR.n2978 VSS 0.001579f
C9619 VDPWR.n2979 VSS 0.00352f
C9620 VDPWR.n2980 VSS 0.003404f
C9621 VDPWR.n2981 VSS 0.128862f
C9622 VDPWR.n2982 VSS 0.128008f
C9623 VDPWR.n2983 VSS 0.001579f
C9624 VDPWR.n2984 VSS 0.001579f
C9625 VDPWR.n2985 VSS 0.001973f
C9626 VDPWR.n2986 VSS 0.002112f
C9627 VDPWR.t877 VSS 0.007047f
C9628 VDPWR.t555 VSS 0.004984f
C9629 VDPWR.n2987 VSS 0.018696f
C9630 VDPWR.n2988 VSS 0.005471f
C9631 VDPWR.t427 VSS 0.005024f
C9632 VDPWR.t1285 VSS 0.010664f
C9633 VDPWR.n2990 VSS 0.027341f
C9634 VDPWR.t428 VSS 0.005024f
C9635 VDPWR.n2991 VSS 0.014893f
C9636 VDPWR.n2992 VSS 0.001472f
C9637 VDPWR.n2993 VSS 0.002048f
C9638 VDPWR.n2994 VSS 0.001973f
C9639 VDPWR.n2995 VSS 0.002944f
C9640 VDPWR.n2996 VSS 0.002048f
C9641 VDPWR.t548 VSS 0.005024f
C9642 VDPWR.t1256 VSS 0.010664f
C9643 VDPWR.n2998 VSS 0.027341f
C9644 VDPWR.t549 VSS 0.005024f
C9645 VDPWR.n2999 VSS 0.014893f
C9646 VDPWR.n3000 VSS 0.012553f
C9647 VDPWR.n3001 VSS 0.001376f
C9648 VDPWR.n3002 VSS 0.002885f
C9649 VDPWR.n3003 VSS 0.003083f
C9650 VDPWR.n3004 VSS 0.003404f
C9651 VDPWR.n3005 VSS 0.00352f
C9652 VDPWR.n3006 VSS 0.00352f
C9653 VDPWR.n3007 VSS 0.003404f
C9654 VDPWR.n3008 VSS 0.003083f
C9655 VDPWR.n3009 VSS 0.002949f
C9656 VDPWR.n3010 VSS 0.00512f
C9657 VDPWR.n3011 VSS 0.002048f
C9658 VDPWR.n3012 VSS 0.015457f
C9659 VDPWR.n3013 VSS 0.015289f
C9660 VDPWR.n3014 VSS 0.01206f
C9661 VDPWR.n3015 VSS 0.032215f
C9662 VDPWR.n3016 VSS 0.005888f
C9663 VDPWR.n3017 VSS 0.004416f
C9664 VDPWR.n3018 VSS 0.005376f
C9665 VDPWR.n3019 VSS 0.005676f
C9666 VDPWR.n3020 VSS 0.003488f
C9667 VDPWR.n3021 VSS 0.005888f
C9668 VDPWR.n3022 VSS 0.005888f
C9669 VDPWR.n3023 VSS 0.001349f
C9670 VDPWR.n3024 VSS 0.006073f
C9671 VDPWR.n3025 VSS 0.001383f
C9672 VDPWR.n3026 VSS 0.004406f
C9673 VDPWR.n3027 VSS 0.00153f
C9674 VDPWR.n3028 VSS 0.0048f
C9675 VDPWR.n3029 VSS 0.002949f
C9676 VDPWR.n3030 VSS 0.003083f
C9677 VDPWR.n3031 VSS 0.003404f
C9678 VDPWR.n3032 VSS 0.00352f
C9679 VDPWR.n3033 VSS 0.003404f
C9680 VDPWR.n3034 VSS 0.00352f
C9681 VDPWR.n3035 VSS 0.001579f
C9682 VDPWR.n3036 VSS 0.001973f
C9683 VDPWR.n3037 VSS 0.00288f
C9684 VDPWR.n3038 VSS 0.002048f
C9685 VDPWR.n3039 VSS 9.41e-19
C9686 VDPWR.n3040 VSS 0.007134f
C9687 VDPWR.n3041 VSS 0.00187f
C9688 VDPWR.n3042 VSS 0.005888f
C9689 VDPWR.n3043 VSS 0.005888f
C9690 VDPWR.n3044 VSS 5.44e-19
C9691 VDPWR.n3045 VSS 0.007134f
C9692 VDPWR.n3046 VSS 0.00187f
C9693 VDPWR.n3047 VSS 0.004416f
C9694 VDPWR.n3048 VSS 0.005888f
C9695 VDPWR.n3049 VSS 0.004416f
C9696 VDPWR.n3050 VSS 0.001247f
C9697 VDPWR.n3051 VSS 0.00364f
C9698 VDPWR.n3052 VSS 0.013305f
C9699 VDPWR.n3053 VSS 0.012101f
C9700 VDPWR.n3054 VSS 0.002016f
C9701 VDPWR.n3055 VSS 5.48e-19
C9702 VDPWR.n3056 VSS 0.003083f
C9703 VDPWR.n3057 VSS 0.001973f
C9704 VDPWR.n3058 VSS 0.002944f
C9705 VDPWR.n3059 VSS 0.002048f
C9706 VDPWR.n3060 VSS 0.012181f
C9707 VDPWR.n3061 VSS 0.011593f
C9708 VDPWR.n3062 VSS 0.002048f
C9709 VDPWR.n3063 VSS 0.00224f
C9710 VDPWR.n3064 VSS 0.001973f
C9711 VDPWR.n3065 VSS 0.003083f
C9712 VDPWR.n3066 VSS 0.003404f
C9713 VDPWR.n3067 VSS 0.128008f
C9714 VDPWR.n3068 VSS 0.116061f
C9715 VDPWR.n3069 VSS 0.281618f
C9716 VDPWR.n3070 VSS 0.167264f
C9717 VDPWR.n3071 VSS 0.281618f
C9718 VDPWR.n3072 VSS 0.116061f
C9719 VDPWR.n3073 VSS 0.107527f
C9720 VDPWR.n3074 VSS 0.078829f
C9721 VDPWR.n3075 VSS 0.003054f
C9722 VDPWR.n3076 VSS 0.002949f
C9723 VDPWR.n3077 VSS 0.004128f
C9724 VDPWR.n3078 VSS 0.002016f
C9725 VDPWR.n3079 VSS 0.001941f
C9726 VDPWR.n3080 VSS 0.005906f
C9727 VDPWR.n3081 VSS 0.003488f
C9728 VDPWR.n3082 VSS 0.004416f
C9729 VDPWR.n3083 VSS 0.011677f
C9730 VDPWR.n3084 VSS 0.015457f
C9731 VDPWR.n3085 VSS 0.011257f
C9732 VDPWR.n3086 VSS 0.005888f
C9733 VDPWR.n3087 VSS 0.005888f
C9734 VDPWR.n3088 VSS 0.005344f
C9735 VDPWR.n3089 VSS 0.011425f
C9736 VDPWR.n3090 VSS 0.046459f
C9737 VDPWR.n3091 VSS 0.009153f
C9738 VDPWR.n3092 VSS 0.010501f
C9739 VDPWR.n3093 VSS 0.002016f
C9740 VDPWR.n3094 VSS 0.002272f
C9741 VDPWR.n3095 VSS 0.005471f
C9742 VDPWR.n3096 VSS 0.01243f
C9743 VDPWR.n3097 VSS 0.001156f
C9744 VDPWR.n3098 VSS 0.002048f
C9745 VDPWR.n3099 VSS 0.002944f
C9746 VDPWR.n3100 VSS 0.001973f
C9747 VDPWR.n3101 VSS 0.001579f
C9748 VDPWR.n3102 VSS 0.078408f
C9749 VDPWR.n3103 VSS 0.272304f
C9750 VDPWR.n3104 VSS 0.13926f
C9751 VDPWR.n3105 VSS 0.13926f
C9752 VDPWR.n3106 VSS 0.209943f
C9753 VDPWR.n3107 VSS 0.292729f
C9754 VDPWR.n3108 VSS 0.060111f
C9755 VDPWR.n3109 VSS 0.281618f
C9756 VDPWR.n3110 VSS 0.167264f
C9757 VDPWR.n3111 VSS 0.060111f
C9758 VDPWR.n3112 VSS 0.096641f
C9759 VDPWR.n3113 VSS 0.107527f
C9760 VDPWR.n3114 VSS 0.02543f
C9761 VDPWR.n3115 VSS 0.067982f
C9762 VDPWR.n3116 VSS 1.57447f
C9763 VDPWR.n3117 VSS 3.32341f
C9764 VDPWR.n3118 VSS 0.390779f
C9765 VDPWR.n3119 VSS 0.035269f
C9766 VDPWR.n3120 VSS 0.114487f
C9767 VDPWR.n3121 VSS 0.055474f
C9768 VDPWR.n3122 VSS 0.055474f
C9769 VDPWR.n3123 VSS 0.055293f
C9770 VDPWR.n3124 VSS 0.076656f
C9771 VDPWR.n3125 VSS 0.247132f
C9772 VDPWR.t1094 VSS 0.356671f
C9773 VDPWR.n3126 VSS 0.344366f
C9774 VDPWR.t1095 VSS 0.356671f
C9775 VDPWR.n3127 VSS 0.247132f
C9776 VDPWR.n3128 VSS 2.38e-19
C9777 VDPWR.n3129 VSS 0.006274f
C9778 VDPWR.n3130 VSS 0.060635f
C9779 VDPWR.n3131 VSS 0.018181f
C9780 VDPWR.n3132 VSS 0.030678f
C9781 VDPWR.n3133 VSS 0.156059f
C9782 VDPWR.n3134 VSS 0.169072f
C9783 VDPWR.n3135 VSS 0.035235f
C9784 VDPWR.n3136 VSS 0.114487f
C9785 VDPWR.n3137 VSS 0.00445f
C9786 VDPWR.n3138 VSS 0.055474f
C9787 VDPWR.n3139 VSS 0.055474f
C9788 VDPWR.n3140 VSS 0.055293f
C9789 VDPWR.n3141 VSS 0.076656f
C9790 VDPWR.n3142 VSS 0.247132f
C9791 VDPWR.t49 VSS 0.356671f
C9792 VDPWR.n3143 VSS 0.344366f
C9793 VDPWR.t50 VSS 0.356671f
C9794 VDPWR.n3144 VSS 0.247132f
C9795 VDPWR.n3145 VSS 0.002025f
C9796 VDPWR.n3146 VSS 0.060694f
C9797 VDPWR.n3147 VSS 0.018181f
C9798 VDPWR.n3148 VSS 0.029169f
C9799 VDPWR.n3149 VSS 0.160902f
C9800 VDPWR.n3150 VSS 0.183546f
C9801 VDPWR.n3151 VSS 0.035121f
C9802 VDPWR.n3152 VSS 0.114487f
C9803 VDPWR.n3153 VSS 0.004458f
C9804 VDPWR.n3154 VSS 0.055474f
C9805 VDPWR.n3155 VSS 0.055474f
C9806 VDPWR.n3156 VSS 0.055293f
C9807 VDPWR.n3157 VSS 0.076656f
C9808 VDPWR.n3158 VSS 0.247132f
C9809 VDPWR.t239 VSS 0.356671f
C9810 VDPWR.n3159 VSS 0.344366f
C9811 VDPWR.t1093 VSS 0.356671f
C9812 VDPWR.n3160 VSS 0.247132f
C9813 VDPWR.n3161 VSS 0.002138f
C9814 VDPWR.n3162 VSS 0.060694f
C9815 VDPWR.n3163 VSS 0.018181f
C9816 VDPWR.n3164 VSS 0.029169f
C9817 VDPWR.n3165 VSS 0.162708f
C9818 VDPWR.n3166 VSS 0.166655f
C9819 VDPWR.n3167 VSS 0.006257f
C9820 VDPWR.n3168 VSS 0.060659f
C9821 VDPWR.n3169 VSS 0.018181f
C9822 VDPWR.n3170 VSS 0.029432f
C9823 VDPWR.n3171 VSS 0.060236f
C9824 VDPWR.n3172 VSS 0.674934f
C9825 VDPWR.t945 VSS 0.0028f
C9826 VDPWR.t1212 VSS 0.00165f
C9827 VDPWR.t948 VSS 0.0028f
C9828 VDPWR.t1206 VSS 0.00165f
C9829 VDPWR.n3173 VSS 0.004698f
C9830 VDPWR.n3174 VSS 0.006946f
C9831 VDPWR.n3175 VSS 0.006899f
C9832 VDPWR.n3176 VSS 0.030149f
C9833 VDPWR.n3177 VSS 0.092595f
C9834 VDPWR.n3178 VSS 0.037419f
C9835 ringtest_0.x4.net2.t7 VSS 0.015381f
C9836 ringtest_0.x4.net2.t8 VSS 0.026101f
C9837 ringtest_0.x4.net2.n0 VSS 0.037026f
C9838 ringtest_0.x4.net2.t4 VSS 0.015381f
C9839 ringtest_0.x4.net2.t3 VSS 0.026101f
C9840 ringtest_0.x4.net2.n1 VSS 0.033335f
C9841 ringtest_0.x4.net2.n2 VSS 0.017289f
C9842 ringtest_0.x4.net2.n3 VSS 0.0837f
C9843 ringtest_0.x4.net2.t5 VSS 0.026101f
C9844 ringtest_0.x4.net2.t2 VSS 0.016278f
C9845 ringtest_0.x4.net2.n4 VSS 0.052479f
C9846 ringtest_0.x4.net2.n5 VSS 0.259642f
C9847 ringtest_0.x4.net2.t9 VSS 0.013842f
C9848 ringtest_0.x4.net2.t11 VSS 0.011454f
C9849 ringtest_0.x4.net2.n6 VSS 0.060494f
C9850 ringtest_0.x4.net2.n7 VSS 0.03533f
C9851 ringtest_0.x4.net2.n8 VSS 0.650991f
C9852 ringtest_0.x4.net2.t6 VSS 0.017756f
C9853 ringtest_0.x4.net2.t10 VSS 0.028277f
C9854 ringtest_0.x4.net2.n9 VSS 0.038818f
C9855 ringtest_0.x4.net2.n10 VSS 0.03575f
C9856 ringtest_0.x4.net2.n11 VSS 0.11929f
C9857 ringtest_0.x4.net2.n12 VSS 0.278364f
C9858 ringtest_0.x4.net2.n13 VSS 0.037886f
C9859 ringtest_0.x4.net2.t1 VSS 0.08709f
C9860 ringtest_0.x4.net2.n14 VSS 0.10636f
C9861 ringtest_0.x4.net2.t0 VSS 0.032833f
.ends

