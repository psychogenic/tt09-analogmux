magic
tech sky130A
magscale 1 2
timestamp 1729136797
<< locali >>
rect 14472 -1376 14810 -1352
rect 7090 -1378 14810 -1376
rect 6608 -1380 14810 -1378
rect 6608 -1470 15696 -1380
rect 6608 -2024 6668 -1470
rect 7016 -1590 15696 -1470
rect 7016 -2024 7124 -1590
rect 6608 -2112 7124 -2024
rect 14472 -1936 15696 -1590
rect 14472 -2180 15706 -1936
rect 14622 -2196 15706 -2180
rect 15446 -2662 15706 -2196
rect 7932 -2922 15706 -2662
<< viali >>
rect 6668 -2024 7016 -1470
<< metal1 >>
rect 6648 -1470 7042 -1434
rect 6648 -1678 6668 -1470
rect 6638 -1964 6668 -1678
rect 6648 -2024 6668 -1964
rect 7016 -1678 7042 -1470
rect 7016 -1964 7606 -1678
rect 7016 -2024 7042 -1964
rect 6648 -2064 7042 -2024
rect 6696 -2290 6886 -2064
rect 6646 -2490 6886 -2290
rect 8098 -2386 8298 -1680
rect 9052 -2296 9252 -1664
rect 6696 -2545 6886 -2490
rect 6696 -3020 6886 -2735
rect 7011 -2586 7694 -2386
rect 7894 -2586 8298 -2386
rect 8784 -2496 9252 -2296
rect 10034 -2474 10234 -1672
rect 6703 -3039 6881 -3020
rect 7011 -4363 7211 -2586
rect 8784 -2992 8984 -2496
rect 9722 -2674 10234 -2474
rect 9722 -2956 9922 -2674
rect 11014 -2876 11214 -1664
rect 8067 -3192 8984 -2992
rect 9111 -3156 9922 -2956
rect 10141 -3076 11214 -2876
rect 12040 -2698 12240 -1672
rect 13102 -2876 13302 -1664
rect 8067 -4365 8267 -3192
rect 9111 -4369 9311 -3156
rect 10141 -4355 10341 -3076
rect 12040 -3348 12240 -2898
rect 11325 -3548 12240 -3348
rect 12381 -3076 13302 -2876
rect 11325 -4361 11525 -3548
rect 12381 -4363 12581 -3076
rect 14100 -3196 14300 -1664
rect 14998 -2005 16520 -2004
rect 14998 -2300 16709 -2005
rect 14998 -2588 15294 -2300
rect 16495 -2347 16709 -2300
rect 16489 -2561 16495 -2347
rect 16709 -2561 16715 -2347
rect 15046 -3020 15246 -2588
rect 13425 -3396 14300 -3196
rect 14455 -3220 15246 -3020
rect 13425 -4367 13625 -3396
rect 14455 -4353 14655 -3220
rect 4090 -5262 4290 -5126
rect 4090 -5326 4215 -5262
rect 4281 -5326 4290 -5262
rect 4215 -5334 4281 -5328
rect 4091 -5366 4525 -5364
rect 4086 -5430 4525 -5366
rect 4086 -5566 4286 -5430
rect 4086 -5643 4316 -5600
rect 4086 -5649 4379 -5643
rect 4086 -5715 4313 -5649
rect 4086 -5721 4379 -5715
rect 4086 -5752 4316 -5721
rect 4086 -5800 4286 -5752
rect 4870 -6138 4876 -5826
rect 5084 -6138 5242 -5826
rect 16074 -8846 16084 -8530
rect 16504 -8626 16514 -8530
rect 16504 -8846 18479 -8626
rect 16431 -8857 18479 -8846
rect 16200 -8863 16431 -8857
rect 15100 -9522 15106 -9322
rect 15306 -9522 15312 -9322
rect 15650 -9340 15660 -9048
rect 16062 -9092 16072 -9048
rect 16062 -9328 17446 -9092
rect 16062 -9340 16072 -9328
rect 12159 -10150 12359 -10144
rect 12159 -10716 12359 -10350
rect 15118 -10404 15294 -9522
rect 16198 -10358 16208 -10238
rect 16360 -10358 16370 -10238
rect 17230 -10402 17426 -9328
rect 18277 -10398 18449 -8857
rect 12159 -12316 12359 -11170
rect 12528 -12091 12728 -12038
rect 12528 -12176 12922 -12091
rect 12528 -12238 12728 -12176
rect 12972 -12270 13047 -12048
rect 13090 -12091 13156 -11979
rect 13090 -12163 13156 -12157
rect 12158 -12478 12359 -12316
rect 12922 -12470 13122 -12270
rect 12158 -12516 12358 -12478
rect 15096 -15340 15296 -14990
rect 16174 -15340 16374 -14942
rect 17244 -15340 17444 -14978
rect 18302 -15340 18502 -14980
rect 15096 -15358 18502 -15340
rect 15092 -15540 18502 -15358
rect 15092 -15558 15292 -15540
<< via1 >>
rect 6696 -2735 6886 -2545
rect 7694 -2586 7894 -2386
rect 12040 -2898 12240 -2698
rect 16495 -2561 16709 -2347
rect 4215 -5328 4281 -5262
rect 4313 -5715 4379 -5649
rect 4876 -6138 5084 -5826
rect 16084 -8846 16504 -8530
rect 16200 -8857 16431 -8846
rect 15106 -9522 15306 -9322
rect 15660 -9340 16062 -9048
rect 12159 -10350 12359 -10150
rect 16208 -10358 16360 -10238
rect 13090 -12157 13156 -12091
<< metal2 >>
rect 16495 -2347 16709 -2341
rect 7694 -2374 8038 -2362
rect 16069 -2372 16290 -2369
rect 7694 -2386 7992 -2374
rect 6690 -2735 6696 -2545
rect 6886 -2735 6892 -2545
rect 7894 -2586 7992 -2386
rect 7694 -2605 7992 -2586
rect 8223 -2605 8232 -2374
rect 16064 -2378 16295 -2372
rect 16064 -2599 16069 -2378
rect 16290 -2552 16295 -2378
rect 16290 -2599 16296 -2552
rect 16495 -2567 16709 -2561
rect 7694 -2606 8038 -2605
rect 16064 -2608 16296 -2599
rect 12026 -2680 12476 -2678
rect 15649 -2680 15875 -2676
rect 12026 -2698 12424 -2680
rect 6696 -2861 6886 -2735
rect 6694 -3039 6703 -2861
rect 6881 -3039 6890 -2861
rect 12026 -2898 12040 -2698
rect 12240 -2898 12424 -2698
rect 12026 -2916 12424 -2898
rect 12660 -2916 12669 -2680
rect 15644 -2685 15880 -2680
rect 15644 -2911 15649 -2685
rect 15875 -2911 15880 -2685
rect 6696 -3051 6886 -3039
rect 4209 -5328 4215 -5262
rect 4281 -5328 4397 -5262
rect 4313 -5649 4379 -5464
rect 4307 -5715 4313 -5649
rect 4379 -5715 4385 -5649
rect 4876 -5826 5084 -5820
rect 4856 -6138 4865 -5826
rect 5096 -6138 5105 -5826
rect 4876 -6144 5084 -6138
rect 15644 -9038 15880 -2911
rect 16064 -2968 16294 -2608
rect 16064 -8520 16295 -2968
rect 16498 -3062 16705 -2567
rect 16494 -3259 16503 -3062
rect 16700 -3259 16709 -3062
rect 16498 -3263 16705 -3259
rect 16064 -8530 16504 -8520
rect 16064 -8846 16084 -8530
rect 16064 -8857 16200 -8846
rect 16431 -8856 16504 -8846
rect 16431 -8857 16437 -8856
rect 15644 -9048 16062 -9038
rect 15106 -9215 15306 -9210
rect 15102 -9322 15111 -9215
rect 15301 -9322 15310 -9215
rect 15102 -9405 15106 -9322
rect 15306 -9405 15310 -9322
rect 15644 -9328 15660 -9048
rect 15660 -9350 16062 -9340
rect 15106 -9528 15306 -9522
rect 12150 -9838 12159 -9638
rect 12359 -9838 12368 -9638
rect 12159 -10150 12359 -9838
rect 12153 -10350 12159 -10150
rect 12359 -10350 12365 -10150
rect 16208 -10238 16360 -10228
rect 16208 -10368 16360 -10358
rect 6311 -12039 6320 -12009
rect 6308 -12173 6320 -12039
rect 6311 -12175 6320 -12173
rect 6486 -12039 6495 -12009
rect 6486 -12058 13857 -12039
rect 6486 -12091 14256 -12058
rect 6486 -12157 13090 -12091
rect 13156 -12154 14256 -12091
rect 13156 -12157 13857 -12154
rect 6486 -12173 13857 -12157
rect 6486 -12175 6495 -12173
<< via2 >>
rect 7992 -2605 8223 -2374
rect 16069 -2599 16290 -2378
rect 6703 -3039 6881 -2861
rect 12424 -2916 12660 -2680
rect 15649 -2911 15875 -2685
rect 4865 -6138 4876 -5826
rect 4876 -6138 5084 -5826
rect 5084 -6138 5096 -5826
rect 16503 -3259 16700 -3062
rect 15111 -9322 15301 -9215
rect 15111 -9405 15301 -9322
rect 12159 -9838 12359 -9638
rect 16208 -10358 16360 -10238
rect 6320 -12175 6486 -12009
<< metal3 >>
rect 7987 -2373 8228 -2369
rect 7987 -2374 16295 -2373
rect 7987 -2605 7992 -2374
rect 8223 -2378 16295 -2374
rect 8223 -2599 16069 -2378
rect 16290 -2599 16295 -2378
rect 8223 -2604 16295 -2599
rect 8223 -2605 8228 -2604
rect 7987 -2610 8228 -2605
rect 12419 -2680 12665 -2675
rect 6698 -2861 6886 -2856
rect 6698 -3039 6703 -2861
rect 6881 -3039 6886 -2861
rect 12419 -2916 12424 -2680
rect 12660 -2685 15880 -2680
rect 12660 -2911 15649 -2685
rect 15875 -2911 15880 -2685
rect 12660 -2916 15880 -2911
rect 12419 -2921 12665 -2916
rect 6698 -3094 6886 -3039
rect 16498 -3062 16705 -3057
rect 6693 -3280 6699 -3094
rect 6885 -3280 6891 -3094
rect 16498 -3259 16503 -3062
rect 16700 -3259 16705 -3062
rect 6698 -3281 6886 -3280
rect 16498 -3632 16705 -3259
rect 16344 -3833 16705 -3632
rect 11982 -4125 16077 -3937
rect 15890 -4735 16077 -4125
rect 4860 -5826 5101 -5821
rect 4860 -6138 4865 -5826
rect 5096 -5866 5101 -5826
rect 5096 -5873 5815 -5866
rect 5177 -6097 5815 -5873
rect 6046 -6097 6491 -5866
rect 5096 -6108 5177 -6102
rect 5096 -6138 5101 -6108
rect 4860 -6143 5101 -6138
rect 6315 -12009 6491 -8562
rect 12159 -9215 15306 -9096
rect 12159 -9296 15111 -9215
rect 12159 -9633 12359 -9296
rect 15106 -9405 15111 -9296
rect 15301 -9405 15306 -9215
rect 15106 -9410 15306 -9405
rect 12154 -9638 12364 -9633
rect 12154 -9838 12159 -9638
rect 12359 -9838 12364 -9638
rect 12154 -9843 12364 -9838
rect 15890 -10111 16076 -4735
rect 16344 -9066 16541 -3833
rect 16208 -9240 16541 -9066
rect 15899 -10155 16069 -10111
rect 16208 -10233 16360 -9240
rect 16198 -10238 16370 -10233
rect 16198 -10358 16208 -10238
rect 16360 -10358 16370 -10238
rect 16198 -10363 16370 -10358
rect 6315 -12175 6320 -12009
rect 6486 -12175 6491 -12009
rect 6315 -12180 6491 -12175
<< via3 >>
rect 6699 -3280 6885 -3094
rect 4948 -6102 5096 -5873
rect 5096 -6102 5177 -5873
rect 5815 -6097 6046 -5866
<< metal4 >>
rect 6442 -3094 6886 -3093
rect 6442 -3280 6699 -3094
rect 6885 -3280 6886 -3094
rect 6442 -3281 6886 -3280
rect 5815 -5865 6046 -5741
rect 5814 -5866 6047 -5865
rect 5814 -5872 5815 -5866
rect 4947 -5873 5815 -5872
rect 4947 -6102 4948 -5873
rect 5177 -6097 5815 -5873
rect 6046 -6097 6047 -5866
rect 5177 -6098 6047 -6097
rect 5177 -6102 6046 -6098
rect 4947 -6103 6046 -6102
use mux8onehot  x1
timestamp 1729136797
transform 1 0 -683 0 1 -10513
box 4991 -1147 16155 7524
use mux4onehot_b  x2
timestamp 1729136797
transform 1 0 7994 0 1 -7186
box 4658 -8054 11287 -2405
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR1 std
timestamp 1728357323
transform 0 -1 14757 1 0 -2427
box -307 -757 307 757
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR2
timestamp 1728357323
transform 0 -1 13799 1 0 -1815
box -307 -757 307 757
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR3
timestamp 1728357323
transform 0 -1 12721 1 0 -2425
box -307 -757 307 757
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR4
timestamp 1728357323
transform 0 -1 11731 1 0 -1803
box -307 -757 307 757
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR5
timestamp 1728357323
transform 0 -1 10653 1 0 -2425
box -307 -757 307 757
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR6
timestamp 1728357323
transform 0 -1 9733 1 0 -1803
box -307 -757 307 757
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR7
timestamp 1728357323
transform 0 -1 8671 1 0 -2425
box -307 -757 307 757
use sky130_fd_pr__res_high_po_1p41_DV8LAQ  XR8
timestamp 1728357323
transform 0 -1 7811 1 0 -1827
box -307 -757 307 757
<< labels >>
flabel metal1 12922 -12470 13122 -12270 0 FreeSans 256 0 0 0 SELECT0
port 2 nsew
flabel metal1 12528 -12238 12728 -12038 0 FreeSans 256 0 0 0 SELECT1
port 3 nsew
flabel metal1 4090 -5326 4290 -5126 0 FreeSans 256 0 0 0 RSEL0
port 5 nsew
flabel metal1 4086 -5566 4286 -5366 0 FreeSans 256 0 0 0 RSEL1
port 6 nsew
flabel metal1 4086 -5800 4286 -5600 0 FreeSans 256 0 0 0 RSEL2
port 7 nsew
flabel metal1 15092 -15558 15292 -15358 0 FreeSans 256 0 0 0 OUT
port 8 nsew
flabel metal1 12158 -12516 12358 -12316 0 FreeSans 256 0 0 0 LADDEROUT
port 9 nsew
flabel metal1 6646 -2490 6846 -2290 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 4966 -6072 5166 -5872 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 16224 -2300 16520 -2004 0 FreeSans 1600 0 0 0 VRES
port 4 nsew
flabel metal1 14028 -3366 14210 -3226 0 FreeSans 240 0 0 0 R1R2
flabel metal1 12396 -3118 12578 -2978 0 FreeSans 240 0 0 0 R2R3
flabel metal1 11992 -3518 12174 -3378 0 FreeSans 240 0 0 0 R3R4
flabel metal1 10156 -3084 10338 -2944 0 FreeSans 240 0 0 0 R4R5
flabel metal1 9172 -3122 9354 -2982 0 FreeSans 240 0 0 0 R5R6
flabel metal1 8718 -3170 8900 -3030 0 FreeSans 240 0 0 0 R6R7
flabel metal1 7098 -2546 7280 -2406 0 FreeSans 240 0 0 0 R7R8
<< end >>
