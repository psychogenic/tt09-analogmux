* NGSPICE file created from passgatex4_parax.ext - technology: sky130A

.subckt passgatex4_parax VCC GN1 A1 GN2 GP3 GN3 GN4 A4 Z2 Z4 A3 GP2 Z1 Z3 VSS A2 GP4
+ GP1
X0 A1.t3 GP1.t0 Z1.t3 VCC.t2 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1 Z2.t3 GN2.t0 A2.t2 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X2 A3.t1 GP3.t0 Z3.t0 VCC.t3 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X3 Z4 GN4.t0 A4.t3 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X4 A2.t0 GP2.t0 Z2.t0 VCC.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X5 Z3.t3 GN3.t0 A3.t3 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X6 Z2.t2 GN2.t1 A2.t3 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X7 A1.t2 GP1.t1 Z1.t2 VCC.t2 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X8 Z3.t2 GN3.t1 A3.t2 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X9 Z1.t0 GN1.t0 A1.t0 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X10 A2.t1 GP2.t1 Z2.t1 VCC.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X11 A4.t1 GP4.t0 Z4 VCC.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X12 Z1.t1 GN1.t1 A1.t1 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X13 A4.t0 GP4.t1 Z4 VCC.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X14 Z4 GN4.t1 A4.t2 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X15 A3.t0 GP3.t1 Z3.t1 VCC.t3 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
R0 GP1.n0 GP1.t1 450.938
R1 GP1.n0 GP1.t0 445.666
R2 GP1.n1 GP1.n0 2.90754
R3 GP1 GP1.n1 0.214408
R4 GP1.n1 GP1 0.16816
R5 Z1.n1 Z1.t3 23.6581
R6 Z1.n3 Z1.t2 23.3739
R7 Z1.n1 Z1.t0 10.7528
R8 Z1.n0 Z1.t1 10.6417
R9 Z1.n2 Z1.n1 1.30064
R10 Z1 Z1.n4 0.983856
R11 Z1.n3 Z1.n2 0.726502
R12 Z1.n2 Z1.n0 0.512491
R13 Z1.n4 Z1.n0 0.359663
R14 Z1.n4 Z1.n3 0.216071
R15 A1.n1 A1.t2 26.3998
R16 A1.n1 A1.t3 23.5483
R17 A1.n0 A1.t1 12.7127
R18 A1.n0 A1.t0 10.8578
R19 A1.n2 A1.n1 3.12177
R20 A1.n2 A1.n0 1.81453
R21 A1.n3 A1.n2 1.1255
R22 A1.n3 A1 0.21549
R23 A1 A1.n3 0.0655
R24 VCC.n45 VCC.n39 8629.41
R25 VCC.n42 VCC.n41 8629.41
R26 VCC.n32 VCC.n26 8629.41
R27 VCC.n29 VCC.n28 8629.41
R28 VCC.n19 VCC.n13 8629.41
R29 VCC.n16 VCC.n15 8629.41
R30 VCC.n7 VCC.n1 8629.41
R31 VCC.n4 VCC.n3 8629.41
R32 VCC.n46 VCC.n40 920.471
R33 VCC.n33 VCC.n27 920.471
R34 VCC.n20 VCC.n14 920.471
R35 VCC.n8 VCC.n2 920.471
R36 VCC.n47 VCC.n46 917.46
R37 VCC.n34 VCC.n33 917.46
R38 VCC.n21 VCC.n20 917.46
R39 VCC.n9 VCC.n8 917.46
R40 VCC.n40 VCC.n38 480.764
R41 VCC.n27 VCC.n25 480.764
R42 VCC.n14 VCC.n12 480.764
R43 VCC.n2 VCC.n0 480.764
R44 VCC.n48 VCC.n38 379.2
R45 VCC.n35 VCC.n25 379.2
R46 VCC.n22 VCC.n12 379.2
R47 VCC.n10 VCC.n0 379.2
R48 VCC.n47 VCC.n39 64.4072
R49 VCC.n34 VCC.n26 64.4072
R50 VCC.n21 VCC.n13 64.4072
R51 VCC.n9 VCC.n1 64.4072
R52 VCC.n41 VCC.n40 61.6672
R53 VCC.n28 VCC.n27 61.6672
R54 VCC.n15 VCC.n14 61.6672
R55 VCC.n3 VCC.n2 61.6672
R56 VCC.n43 VCC.n39 60.9564
R57 VCC.n44 VCC.n41 60.9564
R58 VCC.n30 VCC.n26 60.9564
R59 VCC.n31 VCC.n28 60.9564
R60 VCC.n17 VCC.n13 60.9564
R61 VCC.n18 VCC.n15 60.9564
R62 VCC.n5 VCC.n1 60.9564
R63 VCC.n6 VCC.n3 60.9564
R64 VCC.n45 VCC.n44 38.5759
R65 VCC.n43 VCC.n42 38.5759
R66 VCC.n32 VCC.n31 38.5759
R67 VCC.n30 VCC.n29 38.5759
R68 VCC.n19 VCC.n18 38.5759
R69 VCC.n17 VCC.n16 38.5759
R70 VCC.n7 VCC.n6 38.5759
R71 VCC.n5 VCC.n4 38.5759
R72 VCC.n48 VCC.n47 32.5881
R73 VCC.n35 VCC.n34 32.5881
R74 VCC.n22 VCC.n21 32.5881
R75 VCC.n10 VCC.n9 32.5881
R76 VCC.n49 VCC.n48 11.3235
R77 VCC.n36 VCC.n35 11.3235
R78 VCC.n23 VCC.n22 11.3235
R79 VCC.n11 VCC.n10 11.3235
R80 VCC.n46 VCC.n45 2.84665
R81 VCC.n42 VCC.n38 2.84665
R82 VCC.n33 VCC.n32 2.84665
R83 VCC.n29 VCC.n25 2.84665
R84 VCC.n20 VCC.n19 2.84665
R85 VCC.n16 VCC.n12 2.84665
R86 VCC.n8 VCC.n7 2.84665
R87 VCC.n4 VCC.n0 2.84665
R88 VCC.n49 VCC.n37 2.44889
R89 VCC.n24 VCC.n11 2.42357
R90 VCC.n37 VCC.n24 1.31329
R91 VCC.n37 VCC.n36 1.143
R92 VCC.n24 VCC.n23 1.143
R93 VCC.n44 VCC.t2 0.27666
R94 VCC.t2 VCC.n43 0.27666
R95 VCC.n31 VCC.t1 0.27666
R96 VCC.t1 VCC.n30 0.27666
R97 VCC.n18 VCC.t3 0.27666
R98 VCC.t3 VCC.n17 0.27666
R99 VCC.n6 VCC.t0 0.27666
R100 VCC.t0 VCC.n5 0.27666
R101 VCC.n36 VCC 0.06425
R102 VCC.n23 VCC 0.06425
R103 VCC.n11 VCC 0.06425
R104 VCC VCC.n49 0.06425
R105 GN2.n0 GN2.t1 377.486
R106 GN2.n0 GN2.t0 374.202
R107 GN2 GN2.n0 18.2232
R108 A2.n1 A2.t1 26.3998
R109 A2.n1 A2.t0 23.5483
R110 A2.n0 A2.t3 12.7127
R111 A2.n0 A2.t2 10.8578
R112 A2.n2 A2.n1 3.12177
R113 A2.n2 A2.n0 1.81453
R114 A2.n3 A2.n2 1.1255
R115 A2.n3 A2 0.219402
R116 A2 A2.n3 0.0655
R117 Z2.n1 Z2.t0 23.6581
R118 Z2.n3 Z2.t1 23.3739
R119 Z2.n1 Z2.t3 10.7528
R120 Z2.n0 Z2.t2 10.6417
R121 Z2.n2 Z2.n1 1.30064
R122 Z2.n5 Z2.n4 0.936641
R123 Z2.n3 Z2.n2 0.726502
R124 Z2.n2 Z2.n0 0.512491
R125 Z2.n4 Z2.n0 0.359663
R126 Z2.n4 Z2.n3 0.216071
R127 Z2.n5 Z2 0.0776605
R128 Z2 Z2.n5 0.0561931
R129 VSS.n44 VSS.n6 11744.7
R130 VSS.n48 VSS.n6 11744.7
R131 VSS.n44 VSS.n7 11744.7
R132 VSS.n48 VSS.n7 11744.7
R133 VSS.n37 VSS.n11 11744.7
R134 VSS.n41 VSS.n11 11744.7
R135 VSS.n37 VSS.n12 11744.7
R136 VSS.n41 VSS.n12 11744.7
R137 VSS.n34 VSS.n16 11744.7
R138 VSS.n30 VSS.n17 11744.7
R139 VSS.n34 VSS.n17 11744.7
R140 VSS.n54 VSS.n4 11744.7
R141 VSS.n51 VSS.n5 11744.7
R142 VSS.n51 VSS.n4 11744.7
R143 VSS.n43 VSS.n42 5804.7
R144 VSS.n52 VSS.n49 5804.7
R145 VSS.n36 VSS.n35 5792.48
R146 VSS.n39 VSS.n38 767.294
R147 VSS.n50 VSS.n3 767.294
R148 VSS.n46 VSS.n45 763.106
R149 VSS.n32 VSS.n31 763.106
R150 VSS.n45 VSS.n10 732.236
R151 VSS.n38 VSS.n15 732.236
R152 VSS.n31 VSS.n28 732.236
R153 VSS.n50 VSS.n1 732.236
R154 VSS.n40 VSS.n39 325.502
R155 VSS.n55 VSS.n3 325.502
R156 VSS.n47 VSS.n46 304.204
R157 VSS.n33 VSS.n32 304.204
R158 VSS.n47 VSS.n8 242.448
R159 VSS.n40 VSS.n13 242.448
R160 VSS.n33 VSS.n18 242.448
R161 VSS.n56 VSS.n55 242.448
R162 VSS.n32 VSS.n17 195
R163 VSS.n17 VSS.t1 195
R164 VSS.n27 VSS.n16 195
R165 VSS.n39 VSS.n12 195
R166 VSS.n12 VSS.t3 195
R167 VSS.n14 VSS.n11 195
R168 VSS.n11 VSS.t3 195
R169 VSS.n46 VSS.n7 195
R170 VSS.n7 VSS.t2 195
R171 VSS.n9 VSS.n6 195
R172 VSS.n6 VSS.t2 195
R173 VSS.n4 VSS.n2 195
R174 VSS.t0 VSS.n4 195
R175 VSS.n5 VSS.n3 195
R176 VSS.n29 VSS.n16 189.179
R177 VSS.n53 VSS.n5 189.179
R178 VSS.n30 VSS.n29 161.525
R179 VSS.n54 VSS.n53 161.525
R180 VSS.n35 VSS.t1 155.459
R181 VSS.n36 VSS.t3 155.459
R182 VSS.n42 VSS.t3 155.459
R183 VSS.n43 VSS.t2 155.459
R184 VSS.n49 VSS.t2 155.459
R185 VSS.t0 VSS.n52 155.459
R186 VSS.n10 VSS.n9 30.8711
R187 VSS.n15 VSS.n14 30.8711
R188 VSS.n28 VSS.n27 30.8711
R189 VSS.n2 VSS.n1 30.8711
R190 VSS.n34 VSS.n33 11.0382
R191 VSS.n35 VSS.n34 11.0382
R192 VSS.n31 VSS.n30 11.0382
R193 VSS.n41 VSS.n40 11.0382
R194 VSS.n42 VSS.n41 11.0382
R195 VSS.n38 VSS.n37 11.0382
R196 VSS.n37 VSS.n36 11.0382
R197 VSS.n48 VSS.n47 11.0382
R198 VSS.n49 VSS.n48 11.0382
R199 VSS.n45 VSS.n44 11.0382
R200 VSS.n44 VSS.n43 11.0382
R201 VSS.n51 VSS.n50 11.0382
R202 VSS.n52 VSS.n51 11.0382
R203 VSS.n55 VSS.n54 11.0382
R204 VSS.n9 VSS.n8 10.9181
R205 VSS.n14 VSS.n13 10.9181
R206 VSS.n27 VSS.n18 10.9181
R207 VSS.n56 VSS.n2 10.9181
R208 VSS.n19 VSS.n10 10.4476
R209 VSS.n22 VSS.n15 10.4476
R210 VSS.n28 VSS.n26 10.4476
R211 VSS.n57 VSS.n1 10.4476
R212 VSS.n25 VSS.n24 8.74451
R213 VSS.n58 VSS.n0 8.52409
R214 VSS.n21 VSS.n20 8.00143
R215 VSS.n24 VSS.n23 7.99855
R216 VSS.n20 VSS.n19 7.16724
R217 VSS.n23 VSS.n22 7.16724
R218 VSS.n26 VSS.n25 7.16724
R219 VSS.n58 VSS.n57 7.16724
R220 VSS.n19 VSS.n8 4.73093
R221 VSS.n22 VSS.n13 4.73093
R222 VSS.n26 VSS.n18 4.73093
R223 VSS.n57 VSS.n56 4.73093
R224 VSS.n0 VSS 4.20526
R225 VSS.n29 VSS.t1 2.68284
R226 VSS.n53 VSS.t0 2.68284
R227 VSS.n24 VSS.n21 0.738855
R228 VSS.n21 VSS.n0 0.0960161
R229 VSS.n20 VSS 0.064875
R230 VSS.n23 VSS 0.064875
R231 VSS VSS.n58 0.064875
R232 VSS.n25 VSS 0.063625
R233 GP3.n0 GP3.t0 450.938
R234 GP3.n0 GP3.t1 445.666
R235 GP3.n1 GP3.n0 2.92815
R236 GP3 GP3.n1 0.201889
R237 GP3.n1 GP3 0.172091
R238 Z3.n1 Z3.t1 23.6581
R239 Z3.n3 Z3.t0 23.3739
R240 Z3.n1 Z3.t3 10.7528
R241 Z3.n0 Z3.t2 10.6417
R242 Z3.n2 Z3.n1 1.30064
R243 Z3.n5 Z3.n4 0.924585
R244 Z3.n3 Z3.n2 0.726502
R245 Z3.n2 Z3.n0 0.512491
R246 Z3.n4 Z3.n0 0.359663
R247 Z3.n4 Z3.n3 0.216071
R248 Z3.n5 Z3 0.0656042
R249 Z3 Z3.n5 0.0376287
R250 A3.n1 A3.t1 26.3998
R251 A3.n1 A3.t0 23.5483
R252 A3.n0 A3.t2 12.7127
R253 A3.n0 A3.t3 10.8578
R254 A3.n2 A3.n1 3.12177
R255 A3.n2 A3.n0 1.81453
R256 A3.n3 A3.n2 1.1255
R257 A3.n3 A3 0.210543
R258 A3 A3.n3 0.0655
R259 GN4.n0 GN4.t1 377.486
R260 GN4.n0 GN4.t0 374.202
R261 GN4 GN4.n0 14.8467
R262 A4.n1 A4.t1 26.3998
R263 A4.n1 A4.t0 23.5483
R264 A4.n0 A4.t2 12.7127
R265 A4.n0 A4.t3 10.8578
R266 A4.n2 A4.n1 3.12177
R267 A4.n2 A4.n0 1.81453
R268 A4.n3 A4.n2 1.1255
R269 A4.n3 A4 0.212013
R270 A4 A4.n3 0.0655
R271 GP2.n0 GP2.t1 450.938
R272 GP2.n0 GP2.t0 445.666
R273 GP2.n1 GP2.n0 2.94361
R274 GP2 GP2.n1 0.194849
R275 GP2.n1 GP2 0.165901
R276 GN3.n0 GN3.t1 377.486
R277 GN3.n0 GN3.t0 374.202
R278 GN3 GN3.n0 18.2186
R279 GN1.n0 GN1.t1 377.486
R280 GN1.n0 GN1.t0 374.202
R281 GN1 GN1.n0 18.2364
R282 GP4.n0 GP4.t0 450.938
R283 GP4.n0 GP4.t1 445.666
R284 GP4.n1 GP4.n0 2.95993
R285 GP4.n2 GP4 0.231981
R286 GP4.n2 GP4.n1 0.137486
R287 GP4.n1 GP4 0.133242
R288 GP4 GP4.n2 0.0861164
C0 GP2 Z3 0.063817f
C1 GN4 Z4 0.443708f
C2 GN3 Z4 1.95e-20
C3 GN3 GN2 0.049403f
C4 GP3 VCC 1.3339f
C5 GN3 GP1 8.02e-21
C6 A1 Z1 4.51652f
C7 GN4 A2 1.12e-20
C8 GN3 A2 0.137623f
C9 A3 GN4 0.164499f
C10 A3 GN3 3.78496f
C11 A4 GP2 2.06e-19
C12 Z4 GP3 0.071646f
C13 Z4 VCC 2.71929f
C14 GN2 GP3 4.86e-19
C15 GN2 VCC 0.111197f
C16 Z2 GN3 0.00126f
C17 GN1 Z1 0.427952f
C18 GP1 VCC 1.33304f
C19 A2 GP3 0.001381f
C20 A2 VCC 1.60611f
C21 A3 GP3 3.95861f
C22 A3 VCC 1.61166f
C23 GP2 Z1 3.73e-21
C24 GN1 A1 3.78938f
C25 GN4 Z3 0.00128f
C26 GN3 Z3 0.427085f
C27 GN2 GP1 0.963716f
C28 Z2 GP3 1.03e-20
C29 Z2 VCC 2.76335f
C30 GN2 A2 3.77855f
C31 A3 Z4 0.005563f
C32 GP1 A2 0.122954f
C33 GP2 A1 0.001388f
C34 A3 GN2 0.006579f
C35 A3 GP1 2.46e-21
C36 A3 A2 1.81997f
C37 Z3 GP3 0.278332f
C38 Z3 VCC 2.77127f
C39 GN4 A4 3.82631f
C40 Z2 GN2 0.427019f
C41 GN3 A4 0.007063f
C42 Z2 GP1 0.065749f
C43 GP4 GN4 0.328236f
C44 GN3 GP4 2.62e-19
C45 Z2 A2 4.51569f
C46 A3 Z2 1.49e-20
C47 Z4 Z3 0.002229f
C48 GN2 Z3 2.12e-20
C49 GP1 Z3 1.86e-21
C50 A4 GP3 0.160779f
C51 A4 VCC 1.51968f
C52 Z3 A2 0.004565f
C53 GP4 GP3 0.006538f
C54 GP4 VCC 1.17956f
C55 A3 Z3 4.51555f
C56 GN3 A1 1.74e-20
C57 A4 Z4 4.51497f
C58 Z2 Z3 7.65e-19
C59 GP4 Z4 0.278468f
C60 Z1 VCC 2.57564f
C61 A4 A2 2.39e-19
C62 A3 A4 2.08862f
C63 A3 GP4 0.001458f
C64 A1 VCC 1.56879f
C65 GN2 Z1 6.82e-19
C66 GP1 Z1 0.278468f
C67 GN4 GP2 4.67e-21
C68 GN3 GP2 0.973561f
C69 GN2 A1 0.131325f
C70 GN1 VCC 0.086074f
C71 GP1 A1 3.95876f
C72 A2 A1 1.81909f
C73 GP2 GP3 0.00647f
C74 GP4 Z3 1.58e-20
C75 GP2 VCC 1.33274f
C76 GN2 GN1 0.005648f
C77 GP1 GN1 0.338174f
C78 Z2 A1 0.004942f
C79 GN1 A2 1.17e-19
C80 Z4 GP2 6e-21
C81 GN2 GP2 0.344354f
C82 GP2 GP1 0.006857f
C83 GP4 A4 3.96061f
C84 GP2 A2 3.95592f
C85 GN3 GN4 0.049952f
C86 Z3 A1 4.74e-21
C87 A3 GP2 0.144934f
C88 Z2 GN1 4.77e-21
C89 Z2 GP2 0.278333f
C90 GN4 GP3 1.06141f
C91 GN3 GP3 0.342495f
C92 GN4 VCC 0.11928f
C93 GN3 VCC 0.118245f
C94 GP4 VSS 1.683101f
C95 Z4 VSS 2.21497f
C96 A4 VSS 3.720489f
C97 GN4 VSS 3.102249f
C98 GP3 VSS 1.288311f
C99 Z3 VSS 2.488353f
C100 A3 VSS 3.173578f
C101 GN3 VSS 3.09235f
C102 GP2 VSS 1.293998f
C103 Z2 VSS 2.454255f
C104 A2 VSS 3.299938f
C105 GN2 VSS 3.155516f
C106 GP1 VSS 1.41263f
C107 Z1 VSS 2.811708f
C108 A1 VSS 4.255557f
C109 GN1 VSS 3.876651f
C110 VCC VSS 40.664856f
C111 GP4.t1 VSS 0.49038f
C112 GP4.t0 VSS 0.504054f
C113 GP4.n0 VSS 1.79195f
C114 GP4.n1 VSS 0.821938f
C115 GP4.n2 VSS 0.149514f
C116 GN1.t1 VSS 0.384049f
C117 GN1.t0 VSS 0.374783f
C118 GN1.n0 VSS 2.50763f
C119 GN3.t1 VSS 0.381287f
C120 GN3.t0 VSS 0.372088f
C121 GN3.n0 VSS 2.50166f
C122 GP2.t0 VSS 0.493574f
C123 GP2.t1 VSS 0.507337f
C124 GP2.n0 VSS 1.79995f
C125 GP2.n1 VSS 0.827626f
C126 A4.t2 VSS 0.893325f
C127 A4.t3 VSS 0.512841f
C128 A4.n0 VSS 4.96695f
C129 A4.t1 VSS 0.924602f
C130 A4.t0 VSS 0.65407f
C131 A4.n1 VSS 5.0783f
C132 A4.n2 VSS 0.803255f
C133 A4.n3 VSS 0.268546f
C134 GN4.t1 VSS 0.371267f
C135 GN4.t0 VSS 0.362309f
C136 GN4.n0 VSS 2.53592f
C137 A3.t2 VSS 0.893857f
C138 A3.t3 VSS 0.513146f
C139 A3.n0 VSS 4.9699f
C140 A3.t1 VSS 0.925152f
C141 A3.t0 VSS 0.654459f
C142 A3.n1 VSS 5.08132f
C143 A3.n2 VSS 0.803733f
C144 A3.n3 VSS 0.264783f
C145 Z3.t2 VSS 0.357224f
C146 Z3.n0 VSS 0.533399f
C147 Z3.t3 VSS 0.364394f
C148 Z3.t1 VSS 0.483559f
C149 Z3.n1 VSS 2.44018f
C150 Z3.n2 VSS 0.825656f
C151 Z3.t0 VSS 0.470601f
C152 Z3.n3 VSS 0.585287f
C153 Z3.n4 VSS 0.719041f
C154 Z3.n5 VSS 0.327501f
C155 GP3.t1 VSS 0.492441f
C156 GP3.t0 VSS 0.506172f
C157 GP3.n0 VSS 1.79256f
C158 GP3.n1 VSS 0.851069f
C159 Z2.t2 VSS 0.358514f
C160 Z2.n0 VSS 0.535326f
C161 Z2.t3 VSS 0.365711f
C162 Z2.t0 VSS 0.485306f
C163 Z2.n1 VSS 2.449f
C164 Z2.n2 VSS 0.828639f
C165 Z2.t1 VSS 0.472301f
C166 Z2.n3 VSS 0.587401f
C167 Z2.n4 VSS 0.723878f
C168 Z2.n5 VSS 0.319918f
C169 A2.t3 VSS 0.763965f
C170 A2.t2 VSS 0.438578f
C171 A2.n0 VSS 4.2477f
C172 A2.t1 VSS 0.790712f
C173 A2.t0 VSS 0.559356f
C174 A2.n1 VSS 4.34292f
C175 A2.n2 VSS 0.686937f
C176 A2.n3 VSS 0.222065f
C177 GN2.t1 VSS 0.38601f
C178 GN2.t0 VSS 0.376697f
C179 GN2.n0 VSS 2.5115f
C180 VCC.n0 VSS 0.146622f
C181 VCC.n1 VSS 0.072002f
C182 VCC.n2 VSS 0.098158f
C183 VCC.n3 VSS 0.071893f
C184 VCC.n4 VSS 0.596403f
C185 VCC.t0 VSS 0.793007f
C186 VCC.n7 VSS 0.596403f
C187 VCC.n8 VSS 0.070957f
C188 VCC.n9 VSS 0.046534f
C189 VCC.n10 VSS 0.09375f
C190 VCC.n11 VSS 0.078237f
C191 VCC.n12 VSS 0.146622f
C192 VCC.n13 VSS 0.072002f
C193 VCC.n14 VSS 0.098158f
C194 VCC.n15 VSS 0.071893f
C195 VCC.n16 VSS 0.596403f
C196 VCC.t3 VSS 0.793007f
C197 VCC.n19 VSS 0.596403f
C198 VCC.n20 VSS 0.070957f
C199 VCC.n21 VSS 0.046534f
C200 VCC.n22 VSS 0.09375f
C201 VCC.n23 VSS 0.045778f
C202 VCC.n24 VSS 0.127428f
C203 VCC.n25 VSS 0.146622f
C204 VCC.n26 VSS 0.072002f
C205 VCC.n27 VSS 0.098158f
C206 VCC.n28 VSS 0.071893f
C207 VCC.n29 VSS 0.596403f
C208 VCC.t1 VSS 0.793007f
C209 VCC.n32 VSS 0.596403f
C210 VCC.n33 VSS 0.070957f
C211 VCC.n34 VSS 0.046534f
C212 VCC.n35 VSS 0.09375f
C213 VCC.n36 VSS 0.045778f
C214 VCC.n37 VSS 0.127169f
C215 VCC.n38 VSS 0.146622f
C216 VCC.n39 VSS 0.072002f
C217 VCC.n40 VSS 0.098158f
C218 VCC.n41 VSS 0.071893f
C219 VCC.n42 VSS 0.596403f
C220 VCC.t2 VSS 0.793007f
C221 VCC.n45 VSS 0.596403f
C222 VCC.n46 VSS 0.070957f
C223 VCC.n47 VSS 0.046534f
C224 VCC.n48 VSS 0.09375f
C225 VCC.n49 VSS 0.078735f
C226 A1.t1 VSS 0.764072f
C227 A1.t0 VSS 0.438639f
C228 A1.n0 VSS 4.24829f
C229 A1.t2 VSS 0.790823f
C230 A1.t3 VSS 0.559434f
C231 A1.n1 VSS 4.34353f
C232 A1.n2 VSS 0.687033f
C233 A1.n3 VSS 0.214444f
C234 Z1.t1 VSS 0.348645f
C235 Z1.n0 VSS 0.52059f
C236 Z1.t0 VSS 0.355644f
C237 Z1.t3 VSS 0.471947f
C238 Z1.n1 VSS 2.38159f
C239 Z1.n2 VSS 0.805829f
C240 Z1.t2 VSS 0.4593f
C241 Z1.n3 VSS 0.571232f
C242 Z1.n4 VSS 0.72588f
C243 GP1.t0 VSS 0.491835f
C244 GP1.t1 VSS 0.50555f
C245 GP1.n0 VSS 1.78594f
C246 GP1.n1 VSS 0.835837f
.ends

