magic
tech sky130A
magscale 1 2
timestamp 1728249049
<< viali >>
rect 1409 5185 1443 5219
rect 3617 5185 3651 5219
rect 1685 5117 1719 5151
rect 3341 5117 3375 5151
rect 1685 4709 1719 4743
rect 1869 4641 1903 4675
rect 1961 4573 1995 4607
rect 1409 4505 1443 4539
rect 2145 4437 2179 4471
rect 2329 4165 2363 4199
rect 1593 4097 1627 4131
rect 3065 4097 3099 4131
rect 2789 4029 2823 4063
rect 2697 3961 2731 3995
rect 1409 3893 1443 3927
rect 2881 3893 2915 3927
rect 2145 3621 2179 3655
rect 1593 3553 1627 3587
rect 1501 3485 1535 3519
rect 1685 3485 1719 3519
rect 2053 3485 2087 3519
rect 2329 3485 2363 3519
rect 1869 3349 1903 3383
rect 1593 3077 1627 3111
rect 1409 3009 1443 3043
rect 1869 3009 1903 3043
rect 2605 3009 2639 3043
rect 2881 3009 2915 3043
rect 3617 3009 3651 3043
rect 3801 3009 3835 3043
rect 4077 3009 4111 3043
rect 2329 2941 2363 2975
rect 3433 2941 3467 2975
rect 3893 2873 3927 2907
rect 1777 2805 1811 2839
rect 1961 2805 1995 2839
rect 2421 2805 2455 2839
rect 2973 2805 3007 2839
rect 3341 2805 3375 2839
rect 1593 2601 1627 2635
rect 2513 2533 2547 2567
rect 3341 2533 3375 2567
rect 3801 2533 3835 2567
rect 3525 2465 3559 2499
rect 1777 2397 1811 2431
rect 2053 2397 2087 2431
rect 2329 2397 2363 2431
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 3157 2397 3191 2431
rect 3433 2397 3467 2431
rect 3617 2397 3651 2431
rect 3985 2397 4019 2431
rect 2237 2261 2271 2295
rect 2789 2261 2823 2295
rect 3065 2261 3099 2295
<< metal1 >>
rect 1104 5466 4416 5488
rect 1104 5414 1810 5466
rect 1862 5414 1874 5466
rect 1926 5414 1938 5466
rect 1990 5414 2002 5466
rect 2054 5414 2066 5466
rect 2118 5414 3130 5466
rect 3182 5414 3194 5466
rect 3246 5414 3258 5466
rect 3310 5414 3322 5466
rect 3374 5414 3386 5466
rect 3438 5414 4416 5466
rect 1104 5392 4416 5414
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 4062 5216 4068 5228
rect 3651 5188 4068 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 1670 5108 1676 5160
rect 1728 5108 1734 5160
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 3108 5120 3341 5148
rect 3108 5108 3114 5120
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 1104 4922 4416 4944
rect 1104 4870 1150 4922
rect 1202 4870 1214 4922
rect 1266 4870 1278 4922
rect 1330 4870 1342 4922
rect 1394 4870 1406 4922
rect 1458 4870 2470 4922
rect 2522 4870 2534 4922
rect 2586 4870 2598 4922
rect 2650 4870 2662 4922
rect 2714 4870 2726 4922
rect 2778 4870 3790 4922
rect 3842 4870 3854 4922
rect 3906 4870 3918 4922
rect 3970 4870 3982 4922
rect 4034 4870 4046 4922
rect 4098 4870 4416 4922
rect 1104 4848 4416 4870
rect 1670 4700 1676 4752
rect 1728 4700 1734 4752
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 1903 4644 1992 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 1964 4613 1992 4644
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 1397 4539 1455 4545
rect 1397 4505 1409 4539
rect 1443 4536 1455 4539
rect 3050 4536 3056 4548
rect 1443 4508 3056 4536
rect 1443 4505 1455 4508
rect 1397 4499 1455 4505
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 2130 4428 2136 4480
rect 2188 4428 2194 4480
rect 1104 4378 4416 4400
rect 1104 4326 1810 4378
rect 1862 4326 1874 4378
rect 1926 4326 1938 4378
rect 1990 4326 2002 4378
rect 2054 4326 2066 4378
rect 2118 4326 3130 4378
rect 3182 4326 3194 4378
rect 3246 4326 3258 4378
rect 3310 4326 3322 4378
rect 3374 4326 3386 4378
rect 3438 4326 4416 4378
rect 1104 4304 4416 4326
rect 1670 4156 1676 4208
rect 1728 4196 1734 4208
rect 2317 4199 2375 4205
rect 2317 4196 2329 4199
rect 1728 4168 2329 4196
rect 1728 4156 1734 4168
rect 2317 4165 2329 4168
rect 2363 4165 2375 4199
rect 2317 4159 2375 4165
rect 1578 4088 1584 4140
rect 1636 4088 1642 4140
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 3068 4060 3096 4091
rect 2823 4032 3096 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 2685 3995 2743 4001
rect 2685 3961 2697 3995
rect 2731 3992 2743 3995
rect 3050 3992 3056 4004
rect 2731 3964 3056 3992
rect 2731 3961 2743 3964
rect 2685 3955 2743 3961
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 1026 3884 1032 3936
rect 1084 3924 1090 3936
rect 1397 3927 1455 3933
rect 1397 3924 1409 3927
rect 1084 3896 1409 3924
rect 1084 3884 1090 3896
rect 1397 3893 1409 3896
rect 1443 3893 1455 3927
rect 1397 3887 1455 3893
rect 2869 3927 2927 3933
rect 2869 3893 2881 3927
rect 2915 3924 2927 3927
rect 2958 3924 2964 3936
rect 2915 3896 2964 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 1104 3834 4416 3856
rect 1104 3782 1150 3834
rect 1202 3782 1214 3834
rect 1266 3782 1278 3834
rect 1330 3782 1342 3834
rect 1394 3782 1406 3834
rect 1458 3782 2470 3834
rect 2522 3782 2534 3834
rect 2586 3782 2598 3834
rect 2650 3782 2662 3834
rect 2714 3782 2726 3834
rect 2778 3782 3790 3834
rect 3842 3782 3854 3834
rect 3906 3782 3918 3834
rect 3970 3782 3982 3834
rect 4034 3782 4046 3834
rect 4098 3782 4416 3834
rect 1104 3760 4416 3782
rect 784 3610 790 3662
rect 842 3652 848 3662
rect 2133 3655 2191 3661
rect 2133 3652 2145 3655
rect 842 3624 2145 3652
rect 842 3622 1059 3624
rect 842 3610 848 3622
rect 2133 3621 2145 3624
rect 2179 3621 2191 3655
rect 2133 3615 2191 3621
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1627 3556 2360 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 1489 3519 1547 3525
rect 1489 3516 1501 3519
rect 1452 3488 1501 3516
rect 1452 3476 1458 3488
rect 1489 3485 1501 3488
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 1670 3476 1676 3528
rect 1728 3476 1734 3528
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2130 3516 2136 3528
rect 2087 3488 2136 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2332 3525 2360 3556
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 1688 3448 1716 3476
rect 1504 3420 1716 3448
rect 1504 3392 1532 3420
rect 1486 3340 1492 3392
rect 1544 3340 1550 3392
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1728 3352 1869 3380
rect 1728 3340 1734 3352
rect 1857 3349 1869 3352
rect 1903 3349 1915 3383
rect 1857 3343 1915 3349
rect 1104 3290 4416 3312
rect 1104 3238 1810 3290
rect 1862 3238 1874 3290
rect 1926 3238 1938 3290
rect 1990 3238 2002 3290
rect 2054 3238 2066 3290
rect 2118 3238 3130 3290
rect 3182 3238 3194 3290
rect 3246 3238 3258 3290
rect 3310 3238 3322 3290
rect 3374 3238 3386 3290
rect 3438 3238 4416 3290
rect 1104 3216 4416 3238
rect 1486 3068 1492 3120
rect 1544 3108 1550 3120
rect 1581 3111 1639 3117
rect 1581 3108 1593 3111
rect 1544 3080 1593 3108
rect 1544 3068 1550 3080
rect 1581 3077 1593 3080
rect 1627 3077 1639 3111
rect 1581 3071 1639 3077
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 1360 3012 1409 3040
rect 1360 3000 1366 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1596 3040 1624 3071
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2004 3080 2912 3108
rect 2004 3068 2010 3080
rect 2884 3049 2912 3080
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1596 3012 1869 3040
rect 1397 3003 1455 3009
rect 1857 3009 1869 3012
rect 1903 3040 1915 3043
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 1903 3012 2268 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 1412 2972 1440 3003
rect 1946 2972 1952 2984
rect 1412 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 2240 2904 2268 3012
rect 2332 3012 2605 3040
rect 2332 2981 2360 3012
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3050 3040 3056 3052
rect 2915 3012 3056 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3050 3000 3056 3012
rect 3108 3040 3114 3052
rect 3510 3040 3516 3052
rect 3108 3012 3516 3040
rect 3108 3000 3114 3012
rect 3510 3000 3516 3012
rect 3568 3040 3574 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3568 3012 3617 3040
rect 3568 3000 3574 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 3835 3012 4077 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4065 3009 4077 3012
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2941 2375 2975
rect 3418 2972 3424 2984
rect 2317 2935 2375 2941
rect 2792 2944 3424 2972
rect 2240 2876 2544 2904
rect 1762 2796 1768 2848
rect 1820 2796 1826 2848
rect 1946 2796 1952 2848
rect 2004 2796 2010 2848
rect 2038 2796 2044 2848
rect 2096 2836 2102 2848
rect 2409 2839 2467 2845
rect 2409 2836 2421 2839
rect 2096 2808 2421 2836
rect 2096 2796 2102 2808
rect 2409 2805 2421 2808
rect 2455 2805 2467 2839
rect 2516 2836 2544 2876
rect 2792 2836 2820 2944
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 3881 2907 3939 2913
rect 3881 2904 3893 2907
rect 2924 2876 3893 2904
rect 2924 2864 2930 2876
rect 3881 2873 3893 2876
rect 3927 2873 3939 2907
rect 3881 2867 3939 2873
rect 2961 2839 3019 2845
rect 2961 2836 2973 2839
rect 2516 2808 2973 2836
rect 2409 2799 2467 2805
rect 2961 2805 2973 2808
rect 3007 2805 3019 2839
rect 2961 2799 3019 2805
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 3602 2836 3608 2848
rect 3375 2808 3608 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 3602 2796 3608 2808
rect 3660 2796 3666 2848
rect 1104 2746 4416 2768
rect 1104 2694 1150 2746
rect 1202 2694 1214 2746
rect 1266 2694 1278 2746
rect 1330 2694 1342 2746
rect 1394 2694 1406 2746
rect 1458 2694 2470 2746
rect 2522 2694 2534 2746
rect 2586 2694 2598 2746
rect 2650 2694 2662 2746
rect 2714 2694 2726 2746
rect 2778 2694 3790 2746
rect 3842 2694 3854 2746
rect 3906 2694 3918 2746
rect 3970 2694 3982 2746
rect 4034 2694 4046 2746
rect 4098 2694 4416 2746
rect 1104 2672 4416 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3660 2604 4016 2632
rect 3660 2592 3666 2604
rect 2501 2567 2559 2573
rect 2501 2533 2513 2567
rect 2547 2564 2559 2567
rect 3050 2564 3056 2576
rect 2547 2536 3056 2564
rect 2547 2533 2559 2536
rect 2501 2527 2559 2533
rect 3050 2524 3056 2536
rect 3108 2524 3114 2576
rect 3329 2567 3387 2573
rect 3329 2533 3341 2567
rect 3375 2564 3387 2567
rect 3694 2564 3700 2576
rect 3375 2536 3700 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 3789 2567 3847 2573
rect 3789 2533 3801 2567
rect 3835 2533 3847 2567
rect 3789 2527 3847 2533
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 2884 2468 3525 2496
rect 1762 2388 1768 2440
rect 1820 2388 1826 2440
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2774 2428 2780 2440
rect 2639 2400 2780 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2332 2360 2360 2391
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 2884 2437 2912 2468
rect 3513 2465 3525 2468
rect 3559 2465 3571 2499
rect 3513 2459 3571 2465
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 2958 2360 2964 2372
rect 2332 2332 2964 2360
rect 2958 2320 2964 2332
rect 3016 2320 3022 2372
rect 3160 2360 3188 2391
rect 3418 2388 3424 2440
rect 3476 2388 3482 2440
rect 3602 2388 3608 2440
rect 3660 2388 3666 2440
rect 3804 2428 3832 2527
rect 3988 2437 4016 2604
rect 3712 2400 3832 2428
rect 3973 2431 4031 2437
rect 3712 2360 3740 2400
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 3160 2332 3740 2360
rect 2225 2295 2283 2301
rect 2225 2261 2237 2295
rect 2271 2292 2283 2295
rect 2406 2292 2412 2304
rect 2271 2264 2412 2292
rect 2271 2261 2283 2264
rect 2225 2255 2283 2261
rect 2406 2252 2412 2264
rect 2464 2252 2470 2304
rect 2774 2252 2780 2304
rect 2832 2252 2838 2304
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 4636 2292 4642 2304
rect 3099 2264 4642 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 4636 2252 4642 2264
rect 4694 2252 4700 2304
rect 1104 2202 4416 2224
rect 1104 2150 1810 2202
rect 1862 2150 1874 2202
rect 1926 2150 1938 2202
rect 1990 2150 2002 2202
rect 2054 2150 2066 2202
rect 2118 2150 3130 2202
rect 3182 2150 3194 2202
rect 3246 2150 3258 2202
rect 3310 2150 3322 2202
rect 3374 2150 3386 2202
rect 3438 2150 4416 2202
rect 1104 2128 4416 2150
rect 2774 2048 2780 2100
rect 2832 2088 2838 2100
rect 4338 2088 4344 2100
rect 2832 2060 4344 2088
rect 2832 2048 2838 2060
rect 4338 2048 4344 2060
rect 4396 2048 4402 2100
<< via1 >>
rect 1810 5414 1862 5466
rect 1874 5414 1926 5466
rect 1938 5414 1990 5466
rect 2002 5414 2054 5466
rect 2066 5414 2118 5466
rect 3130 5414 3182 5466
rect 3194 5414 3246 5466
rect 3258 5414 3310 5466
rect 3322 5414 3374 5466
rect 3386 5414 3438 5466
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 4068 5176 4120 5228
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 3056 5108 3108 5160
rect 1150 4870 1202 4922
rect 1214 4870 1266 4922
rect 1278 4870 1330 4922
rect 1342 4870 1394 4922
rect 1406 4870 1458 4922
rect 2470 4870 2522 4922
rect 2534 4870 2586 4922
rect 2598 4870 2650 4922
rect 2662 4870 2714 4922
rect 2726 4870 2778 4922
rect 3790 4870 3842 4922
rect 3854 4870 3906 4922
rect 3918 4870 3970 4922
rect 3982 4870 4034 4922
rect 4046 4870 4098 4922
rect 1676 4743 1728 4752
rect 1676 4709 1685 4743
rect 1685 4709 1719 4743
rect 1719 4709 1728 4743
rect 1676 4700 1728 4709
rect 3056 4496 3108 4548
rect 2136 4471 2188 4480
rect 2136 4437 2145 4471
rect 2145 4437 2179 4471
rect 2179 4437 2188 4471
rect 2136 4428 2188 4437
rect 1810 4326 1862 4378
rect 1874 4326 1926 4378
rect 1938 4326 1990 4378
rect 2002 4326 2054 4378
rect 2066 4326 2118 4378
rect 3130 4326 3182 4378
rect 3194 4326 3246 4378
rect 3258 4326 3310 4378
rect 3322 4326 3374 4378
rect 3386 4326 3438 4378
rect 1676 4156 1728 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 3056 3952 3108 4004
rect 1032 3884 1084 3936
rect 2964 3884 3016 3936
rect 1150 3782 1202 3834
rect 1214 3782 1266 3834
rect 1278 3782 1330 3834
rect 1342 3782 1394 3834
rect 1406 3782 1458 3834
rect 2470 3782 2522 3834
rect 2534 3782 2586 3834
rect 2598 3782 2650 3834
rect 2662 3782 2714 3834
rect 2726 3782 2778 3834
rect 3790 3782 3842 3834
rect 3854 3782 3906 3834
rect 3918 3782 3970 3834
rect 3982 3782 4034 3834
rect 4046 3782 4098 3834
rect 790 3610 842 3662
rect 1400 3476 1452 3528
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 2136 3476 2188 3528
rect 1492 3340 1544 3392
rect 1676 3340 1728 3392
rect 1810 3238 1862 3290
rect 1874 3238 1926 3290
rect 1938 3238 1990 3290
rect 2002 3238 2054 3290
rect 2066 3238 2118 3290
rect 3130 3238 3182 3290
rect 3194 3238 3246 3290
rect 3258 3238 3310 3290
rect 3322 3238 3374 3290
rect 3386 3238 3438 3290
rect 1492 3068 1544 3120
rect 1308 3000 1360 3052
rect 1952 3068 2004 3120
rect 1952 2932 2004 2984
rect 3056 3000 3108 3052
rect 3516 3000 3568 3052
rect 3424 2975 3476 2984
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 1952 2839 2004 2848
rect 1952 2805 1961 2839
rect 1961 2805 1995 2839
rect 1995 2805 2004 2839
rect 1952 2796 2004 2805
rect 2044 2796 2096 2848
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 2872 2864 2924 2916
rect 3608 2796 3660 2848
rect 1150 2694 1202 2746
rect 1214 2694 1266 2746
rect 1278 2694 1330 2746
rect 1342 2694 1394 2746
rect 1406 2694 1458 2746
rect 2470 2694 2522 2746
rect 2534 2694 2586 2746
rect 2598 2694 2650 2746
rect 2662 2694 2714 2746
rect 2726 2694 2778 2746
rect 3790 2694 3842 2746
rect 3854 2694 3906 2746
rect 3918 2694 3970 2746
rect 3982 2694 4034 2746
rect 4046 2694 4098 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 3608 2592 3660 2644
rect 3056 2524 3108 2576
rect 3700 2524 3752 2576
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2780 2388 2832 2440
rect 2964 2320 3016 2372
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3424 2388 3476 2397
rect 3608 2431 3660 2440
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 2412 2252 2464 2304
rect 2780 2295 2832 2304
rect 2780 2261 2789 2295
rect 2789 2261 2823 2295
rect 2823 2261 2832 2295
rect 2780 2252 2832 2261
rect 4642 2252 4694 2304
rect 1810 2150 1862 2202
rect 1874 2150 1926 2202
rect 1938 2150 1990 2202
rect 2002 2150 2054 2202
rect 2066 2150 2118 2202
rect 3130 2150 3182 2202
rect 3194 2150 3246 2202
rect 3258 2150 3310 2202
rect 3322 2150 3374 2202
rect 3386 2150 3438 2202
rect 2780 2048 2832 2100
rect 4344 2048 4396 2100
<< metal2 >>
rect 1306 5699 1362 6262
rect 1776 5709 1832 6262
rect 1320 5522 1348 5699
rect 1790 5604 1818 5709
rect 1790 5576 4108 5604
rect 1320 5494 1440 5522
rect 1412 5234 1440 5494
rect 1810 5468 2118 5477
rect 1810 5466 1816 5468
rect 1872 5466 1896 5468
rect 1952 5466 1976 5468
rect 2032 5466 2056 5468
rect 2112 5466 2118 5468
rect 1872 5414 1874 5466
rect 2054 5414 2056 5466
rect 1810 5412 1816 5414
rect 1872 5412 1896 5414
rect 1952 5412 1976 5414
rect 2032 5412 2056 5414
rect 2112 5412 2118 5414
rect 1810 5403 2118 5412
rect 3130 5468 3438 5477
rect 3130 5466 3136 5468
rect 3192 5466 3216 5468
rect 3272 5466 3296 5468
rect 3352 5466 3376 5468
rect 3432 5466 3438 5468
rect 3192 5414 3194 5466
rect 3374 5414 3376 5466
rect 3130 5412 3136 5414
rect 3192 5412 3216 5414
rect 3272 5412 3296 5414
rect 3352 5412 3376 5414
rect 3432 5412 3438 5414
rect 3130 5403 3438 5412
rect 4080 5234 4108 5576
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 1150 4924 1458 4933
rect 1150 4922 1156 4924
rect 1212 4922 1236 4924
rect 1292 4922 1316 4924
rect 1372 4922 1396 4924
rect 1452 4922 1458 4924
rect 1212 4870 1214 4922
rect 1394 4870 1396 4922
rect 1150 4868 1156 4870
rect 1212 4868 1236 4870
rect 1292 4868 1316 4870
rect 1372 4868 1396 4870
rect 1452 4868 1458 4870
rect 1150 4859 1458 4868
rect 1688 4758 1716 5102
rect 2470 4924 2778 4933
rect 2470 4922 2476 4924
rect 2532 4922 2556 4924
rect 2612 4922 2636 4924
rect 2692 4922 2716 4924
rect 2772 4922 2778 4924
rect 2532 4870 2534 4922
rect 2714 4870 2716 4922
rect 2470 4868 2476 4870
rect 2532 4868 2556 4870
rect 2612 4868 2636 4870
rect 2692 4868 2716 4870
rect 2772 4868 2778 4870
rect 2470 4859 2778 4868
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1688 4214 1716 4694
rect 3068 4554 3096 5102
rect 3790 4924 4098 4933
rect 3790 4922 3796 4924
rect 3852 4922 3876 4924
rect 3932 4922 3956 4924
rect 4012 4922 4036 4924
rect 4092 4922 4098 4924
rect 3852 4870 3854 4922
rect 4034 4870 4036 4922
rect 3790 4868 3796 4870
rect 3852 4868 3876 4870
rect 3932 4868 3956 4870
rect 4012 4868 4036 4870
rect 4092 4868 4098 4870
rect 3790 4859 4098 4868
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 1810 4380 2118 4389
rect 1810 4378 1816 4380
rect 1872 4378 1896 4380
rect 1952 4378 1976 4380
rect 2032 4378 2056 4380
rect 2112 4378 2118 4380
rect 1872 4326 1874 4378
rect 2054 4326 2056 4378
rect 1810 4324 1816 4326
rect 1872 4324 1896 4326
rect 1952 4324 1976 4326
rect 2032 4324 2056 4326
rect 2112 4324 2118 4326
rect 1810 4315 2118 4324
rect 1676 4208 1728 4214
rect 1676 4150 1728 4156
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1032 3936 1084 3942
rect 1032 3878 1084 3884
rect 790 3662 842 3668
rect 790 3604 842 3610
rect 802 2028 830 3604
rect 802 1930 832 2028
rect 1044 1934 1072 3878
rect 1150 3836 1458 3845
rect 1150 3834 1156 3836
rect 1212 3834 1236 3836
rect 1292 3834 1316 3836
rect 1372 3834 1396 3836
rect 1452 3834 1458 3836
rect 1212 3782 1214 3834
rect 1394 3782 1396 3834
rect 1150 3780 1156 3782
rect 1212 3780 1236 3782
rect 1292 3780 1316 3782
rect 1372 3780 1396 3782
rect 1452 3780 1458 3782
rect 1150 3771 1458 3780
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1412 3210 1440 3470
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1320 3182 1440 3210
rect 1320 3058 1348 3182
rect 1504 3126 1532 3334
rect 1492 3120 1544 3126
rect 1492 3062 1544 3068
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1150 2748 1458 2757
rect 1150 2746 1156 2748
rect 1212 2746 1236 2748
rect 1292 2746 1316 2748
rect 1372 2746 1396 2748
rect 1452 2746 1458 2748
rect 1212 2694 1214 2746
rect 1394 2694 1396 2746
rect 1150 2692 1156 2694
rect 1212 2692 1236 2694
rect 1292 2692 1316 2694
rect 1372 2692 1396 2694
rect 1452 2692 1458 2694
rect 1150 2683 1458 2692
rect 1596 2650 1624 4082
rect 1688 3534 1716 4150
rect 2148 3534 2176 4422
rect 3068 4010 3096 4490
rect 3130 4380 3438 4389
rect 3130 4378 3136 4380
rect 3192 4378 3216 4380
rect 3272 4378 3296 4380
rect 3352 4378 3376 4380
rect 3432 4378 3438 4380
rect 3192 4326 3194 4378
rect 3374 4326 3376 4378
rect 3130 4324 3136 4326
rect 3192 4324 3216 4326
rect 3272 4324 3296 4326
rect 3352 4324 3376 4326
rect 3432 4324 3438 4326
rect 3130 4315 3438 4324
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2470 3836 2778 3845
rect 2470 3834 2476 3836
rect 2532 3834 2556 3836
rect 2612 3834 2636 3836
rect 2692 3834 2716 3836
rect 2772 3834 2778 3836
rect 2532 3782 2534 3834
rect 2714 3782 2716 3834
rect 2470 3780 2476 3782
rect 2532 3780 2556 3782
rect 2612 3780 2636 3782
rect 2692 3780 2716 3782
rect 2772 3780 2778 3782
rect 2470 3771 2778 3780
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1688 2060 1716 3334
rect 1810 3292 2118 3301
rect 1810 3290 1816 3292
rect 1872 3290 1896 3292
rect 1952 3290 1976 3292
rect 2032 3290 2056 3292
rect 2112 3290 2118 3292
rect 1872 3238 1874 3290
rect 2054 3238 2056 3290
rect 1810 3236 1816 3238
rect 1872 3236 1896 3238
rect 1952 3236 1976 3238
rect 2032 3236 2056 3238
rect 2112 3236 2118 3238
rect 1810 3227 2118 3236
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1964 2990 1992 3062
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 1964 2854 1992 2926
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1780 2446 1808 2790
rect 2056 2446 2084 2790
rect 2470 2748 2778 2757
rect 2470 2746 2476 2748
rect 2532 2746 2556 2748
rect 2612 2746 2636 2748
rect 2692 2746 2716 2748
rect 2772 2746 2778 2748
rect 2532 2694 2534 2746
rect 2714 2694 2716 2746
rect 2470 2692 2476 2694
rect 2532 2692 2556 2694
rect 2612 2692 2636 2694
rect 2692 2692 2716 2694
rect 2772 2692 2778 2694
rect 2470 2683 2778 2692
rect 2884 2530 2912 2858
rect 2792 2502 2912 2530
rect 2792 2446 2820 2502
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2976 2378 3004 3878
rect 3068 3058 3096 3946
rect 3790 3836 4098 3845
rect 3790 3834 3796 3836
rect 3852 3834 3876 3836
rect 3932 3834 3956 3836
rect 4012 3834 4036 3836
rect 4092 3834 4098 3836
rect 3852 3782 3854 3834
rect 4034 3782 4036 3834
rect 3790 3780 3796 3782
rect 3852 3780 3876 3782
rect 3932 3780 3956 3782
rect 4012 3780 4036 3782
rect 4092 3780 4098 3782
rect 3790 3771 4098 3780
rect 3130 3292 3438 3301
rect 3130 3290 3136 3292
rect 3192 3290 3216 3292
rect 3272 3290 3296 3292
rect 3352 3290 3376 3292
rect 3432 3290 3438 3292
rect 3192 3238 3194 3290
rect 3374 3238 3376 3290
rect 3130 3236 3136 3238
rect 3192 3236 3216 3238
rect 3272 3236 3296 3238
rect 3352 3236 3376 3238
rect 3432 3236 3438 3238
rect 3130 3227 3438 3236
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 1810 2204 2118 2213
rect 1810 2202 1816 2204
rect 1872 2202 1896 2204
rect 1952 2202 1976 2204
rect 2032 2202 2056 2204
rect 2112 2202 2118 2204
rect 1872 2150 1874 2202
rect 2054 2150 2056 2202
rect 1810 2148 1816 2150
rect 1872 2148 1896 2150
rect 1952 2148 1976 2150
rect 2032 2148 2056 2150
rect 2112 2148 2118 2150
rect 1810 2139 2118 2148
rect 1688 2032 1810 2060
rect 790 1432 846 1930
rect 1044 1906 1180 1934
rect 1782 1932 1810 2032
rect 2424 2030 2452 2246
rect 2792 2106 2820 2246
rect 2780 2100 2832 2106
rect 2780 2042 2832 2048
rect 3068 2030 3096 2518
rect 3436 2446 3464 2926
rect 3528 2530 3556 2994
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3620 2650 3648 2790
rect 3790 2748 4098 2757
rect 3790 2746 3796 2748
rect 3852 2746 3876 2748
rect 3932 2746 3956 2748
rect 4012 2746 4036 2748
rect 4092 2746 4098 2748
rect 3852 2694 3854 2746
rect 4034 2694 4036 2746
rect 3790 2692 3796 2694
rect 3852 2692 3876 2694
rect 3932 2692 3956 2694
rect 4012 2692 4036 2694
rect 4092 2692 4098 2694
rect 3790 2683 4098 2692
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3700 2576 3752 2582
rect 3528 2502 3648 2530
rect 3700 2518 3752 2524
rect 3620 2446 3648 2502
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3130 2204 3438 2213
rect 3130 2202 3136 2204
rect 3192 2202 3216 2204
rect 3272 2202 3296 2204
rect 3352 2202 3376 2204
rect 3432 2202 3438 2204
rect 3192 2150 3194 2202
rect 3374 2150 3376 2202
rect 3130 2148 3136 2150
rect 3192 2148 3216 2150
rect 3272 2148 3296 2150
rect 3352 2148 3376 2150
rect 3432 2148 3438 2150
rect 3130 2139 3438 2148
rect 3712 2030 3740 2518
rect 4642 2304 4694 2310
rect 4642 2246 4694 2252
rect 4344 2102 4396 2106
rect 4344 2100 4400 2102
rect 4396 2048 4400 2100
rect 2424 1932 2454 2030
rect 3068 1932 3098 2030
rect 3712 1932 3742 2030
rect 1124 1434 1180 1906
rect 1768 1434 1824 1932
rect 2412 1434 2468 1932
rect 3056 1434 3112 1932
rect 3700 1434 3756 1932
rect 4344 1434 4400 2048
rect 4654 2030 4682 2246
rect 4654 1932 4684 2030
rect 4642 1434 4698 1932
<< via2 >>
rect 1816 5466 1872 5468
rect 1896 5466 1952 5468
rect 1976 5466 2032 5468
rect 2056 5466 2112 5468
rect 1816 5414 1862 5466
rect 1862 5414 1872 5466
rect 1896 5414 1926 5466
rect 1926 5414 1938 5466
rect 1938 5414 1952 5466
rect 1976 5414 1990 5466
rect 1990 5414 2002 5466
rect 2002 5414 2032 5466
rect 2056 5414 2066 5466
rect 2066 5414 2112 5466
rect 1816 5412 1872 5414
rect 1896 5412 1952 5414
rect 1976 5412 2032 5414
rect 2056 5412 2112 5414
rect 3136 5466 3192 5468
rect 3216 5466 3272 5468
rect 3296 5466 3352 5468
rect 3376 5466 3432 5468
rect 3136 5414 3182 5466
rect 3182 5414 3192 5466
rect 3216 5414 3246 5466
rect 3246 5414 3258 5466
rect 3258 5414 3272 5466
rect 3296 5414 3310 5466
rect 3310 5414 3322 5466
rect 3322 5414 3352 5466
rect 3376 5414 3386 5466
rect 3386 5414 3432 5466
rect 3136 5412 3192 5414
rect 3216 5412 3272 5414
rect 3296 5412 3352 5414
rect 3376 5412 3432 5414
rect 1156 4922 1212 4924
rect 1236 4922 1292 4924
rect 1316 4922 1372 4924
rect 1396 4922 1452 4924
rect 1156 4870 1202 4922
rect 1202 4870 1212 4922
rect 1236 4870 1266 4922
rect 1266 4870 1278 4922
rect 1278 4870 1292 4922
rect 1316 4870 1330 4922
rect 1330 4870 1342 4922
rect 1342 4870 1372 4922
rect 1396 4870 1406 4922
rect 1406 4870 1452 4922
rect 1156 4868 1212 4870
rect 1236 4868 1292 4870
rect 1316 4868 1372 4870
rect 1396 4868 1452 4870
rect 2476 4922 2532 4924
rect 2556 4922 2612 4924
rect 2636 4922 2692 4924
rect 2716 4922 2772 4924
rect 2476 4870 2522 4922
rect 2522 4870 2532 4922
rect 2556 4870 2586 4922
rect 2586 4870 2598 4922
rect 2598 4870 2612 4922
rect 2636 4870 2650 4922
rect 2650 4870 2662 4922
rect 2662 4870 2692 4922
rect 2716 4870 2726 4922
rect 2726 4870 2772 4922
rect 2476 4868 2532 4870
rect 2556 4868 2612 4870
rect 2636 4868 2692 4870
rect 2716 4868 2772 4870
rect 3796 4922 3852 4924
rect 3876 4922 3932 4924
rect 3956 4922 4012 4924
rect 4036 4922 4092 4924
rect 3796 4870 3842 4922
rect 3842 4870 3852 4922
rect 3876 4870 3906 4922
rect 3906 4870 3918 4922
rect 3918 4870 3932 4922
rect 3956 4870 3970 4922
rect 3970 4870 3982 4922
rect 3982 4870 4012 4922
rect 4036 4870 4046 4922
rect 4046 4870 4092 4922
rect 3796 4868 3852 4870
rect 3876 4868 3932 4870
rect 3956 4868 4012 4870
rect 4036 4868 4092 4870
rect 1816 4378 1872 4380
rect 1896 4378 1952 4380
rect 1976 4378 2032 4380
rect 2056 4378 2112 4380
rect 1816 4326 1862 4378
rect 1862 4326 1872 4378
rect 1896 4326 1926 4378
rect 1926 4326 1938 4378
rect 1938 4326 1952 4378
rect 1976 4326 1990 4378
rect 1990 4326 2002 4378
rect 2002 4326 2032 4378
rect 2056 4326 2066 4378
rect 2066 4326 2112 4378
rect 1816 4324 1872 4326
rect 1896 4324 1952 4326
rect 1976 4324 2032 4326
rect 2056 4324 2112 4326
rect 1156 3834 1212 3836
rect 1236 3834 1292 3836
rect 1316 3834 1372 3836
rect 1396 3834 1452 3836
rect 1156 3782 1202 3834
rect 1202 3782 1212 3834
rect 1236 3782 1266 3834
rect 1266 3782 1278 3834
rect 1278 3782 1292 3834
rect 1316 3782 1330 3834
rect 1330 3782 1342 3834
rect 1342 3782 1372 3834
rect 1396 3782 1406 3834
rect 1406 3782 1452 3834
rect 1156 3780 1212 3782
rect 1236 3780 1292 3782
rect 1316 3780 1372 3782
rect 1396 3780 1452 3782
rect 1156 2746 1212 2748
rect 1236 2746 1292 2748
rect 1316 2746 1372 2748
rect 1396 2746 1452 2748
rect 1156 2694 1202 2746
rect 1202 2694 1212 2746
rect 1236 2694 1266 2746
rect 1266 2694 1278 2746
rect 1278 2694 1292 2746
rect 1316 2694 1330 2746
rect 1330 2694 1342 2746
rect 1342 2694 1372 2746
rect 1396 2694 1406 2746
rect 1406 2694 1452 2746
rect 1156 2692 1212 2694
rect 1236 2692 1292 2694
rect 1316 2692 1372 2694
rect 1396 2692 1452 2694
rect 3136 4378 3192 4380
rect 3216 4378 3272 4380
rect 3296 4378 3352 4380
rect 3376 4378 3432 4380
rect 3136 4326 3182 4378
rect 3182 4326 3192 4378
rect 3216 4326 3246 4378
rect 3246 4326 3258 4378
rect 3258 4326 3272 4378
rect 3296 4326 3310 4378
rect 3310 4326 3322 4378
rect 3322 4326 3352 4378
rect 3376 4326 3386 4378
rect 3386 4326 3432 4378
rect 3136 4324 3192 4326
rect 3216 4324 3272 4326
rect 3296 4324 3352 4326
rect 3376 4324 3432 4326
rect 2476 3834 2532 3836
rect 2556 3834 2612 3836
rect 2636 3834 2692 3836
rect 2716 3834 2772 3836
rect 2476 3782 2522 3834
rect 2522 3782 2532 3834
rect 2556 3782 2586 3834
rect 2586 3782 2598 3834
rect 2598 3782 2612 3834
rect 2636 3782 2650 3834
rect 2650 3782 2662 3834
rect 2662 3782 2692 3834
rect 2716 3782 2726 3834
rect 2726 3782 2772 3834
rect 2476 3780 2532 3782
rect 2556 3780 2612 3782
rect 2636 3780 2692 3782
rect 2716 3780 2772 3782
rect 1816 3290 1872 3292
rect 1896 3290 1952 3292
rect 1976 3290 2032 3292
rect 2056 3290 2112 3292
rect 1816 3238 1862 3290
rect 1862 3238 1872 3290
rect 1896 3238 1926 3290
rect 1926 3238 1938 3290
rect 1938 3238 1952 3290
rect 1976 3238 1990 3290
rect 1990 3238 2002 3290
rect 2002 3238 2032 3290
rect 2056 3238 2066 3290
rect 2066 3238 2112 3290
rect 1816 3236 1872 3238
rect 1896 3236 1952 3238
rect 1976 3236 2032 3238
rect 2056 3236 2112 3238
rect 2476 2746 2532 2748
rect 2556 2746 2612 2748
rect 2636 2746 2692 2748
rect 2716 2746 2772 2748
rect 2476 2694 2522 2746
rect 2522 2694 2532 2746
rect 2556 2694 2586 2746
rect 2586 2694 2598 2746
rect 2598 2694 2612 2746
rect 2636 2694 2650 2746
rect 2650 2694 2662 2746
rect 2662 2694 2692 2746
rect 2716 2694 2726 2746
rect 2726 2694 2772 2746
rect 2476 2692 2532 2694
rect 2556 2692 2612 2694
rect 2636 2692 2692 2694
rect 2716 2692 2772 2694
rect 3796 3834 3852 3836
rect 3876 3834 3932 3836
rect 3956 3834 4012 3836
rect 4036 3834 4092 3836
rect 3796 3782 3842 3834
rect 3842 3782 3852 3834
rect 3876 3782 3906 3834
rect 3906 3782 3918 3834
rect 3918 3782 3932 3834
rect 3956 3782 3970 3834
rect 3970 3782 3982 3834
rect 3982 3782 4012 3834
rect 4036 3782 4046 3834
rect 4046 3782 4092 3834
rect 3796 3780 3852 3782
rect 3876 3780 3932 3782
rect 3956 3780 4012 3782
rect 4036 3780 4092 3782
rect 3136 3290 3192 3292
rect 3216 3290 3272 3292
rect 3296 3290 3352 3292
rect 3376 3290 3432 3292
rect 3136 3238 3182 3290
rect 3182 3238 3192 3290
rect 3216 3238 3246 3290
rect 3246 3238 3258 3290
rect 3258 3238 3272 3290
rect 3296 3238 3310 3290
rect 3310 3238 3322 3290
rect 3322 3238 3352 3290
rect 3376 3238 3386 3290
rect 3386 3238 3432 3290
rect 3136 3236 3192 3238
rect 3216 3236 3272 3238
rect 3296 3236 3352 3238
rect 3376 3236 3432 3238
rect 1816 2202 1872 2204
rect 1896 2202 1952 2204
rect 1976 2202 2032 2204
rect 2056 2202 2112 2204
rect 1816 2150 1862 2202
rect 1862 2150 1872 2202
rect 1896 2150 1926 2202
rect 1926 2150 1938 2202
rect 1938 2150 1952 2202
rect 1976 2150 1990 2202
rect 1990 2150 2002 2202
rect 2002 2150 2032 2202
rect 2056 2150 2066 2202
rect 2066 2150 2112 2202
rect 1816 2148 1872 2150
rect 1896 2148 1952 2150
rect 1976 2148 2032 2150
rect 2056 2148 2112 2150
rect 3796 2746 3852 2748
rect 3876 2746 3932 2748
rect 3956 2746 4012 2748
rect 4036 2746 4092 2748
rect 3796 2694 3842 2746
rect 3842 2694 3852 2746
rect 3876 2694 3906 2746
rect 3906 2694 3918 2746
rect 3918 2694 3932 2746
rect 3956 2694 3970 2746
rect 3970 2694 3982 2746
rect 3982 2694 4012 2746
rect 4036 2694 4046 2746
rect 4046 2694 4092 2746
rect 3796 2692 3852 2694
rect 3876 2692 3932 2694
rect 3956 2692 4012 2694
rect 4036 2692 4092 2694
rect 3136 2202 3192 2204
rect 3216 2202 3272 2204
rect 3296 2202 3352 2204
rect 3376 2202 3432 2204
rect 3136 2150 3182 2202
rect 3182 2150 3192 2202
rect 3216 2150 3246 2202
rect 3246 2150 3258 2202
rect 3258 2150 3272 2202
rect 3296 2150 3310 2202
rect 3310 2150 3322 2202
rect 3322 2150 3352 2202
rect 3376 2150 3386 2202
rect 3386 2150 3432 2202
rect 3136 2148 3192 2150
rect 3216 2148 3272 2150
rect 3296 2148 3352 2150
rect 3376 2148 3432 2150
<< metal3 >>
rect 1806 5472 2122 5473
rect 1806 5408 1812 5472
rect 1876 5408 1892 5472
rect 1956 5408 1972 5472
rect 2036 5408 2052 5472
rect 2116 5408 2122 5472
rect 1806 5407 2122 5408
rect 3126 5472 3442 5473
rect 3126 5408 3132 5472
rect 3196 5408 3212 5472
rect 3276 5408 3292 5472
rect 3356 5408 3372 5472
rect 3436 5408 3442 5472
rect 3126 5407 3442 5408
rect 1146 4928 1462 4929
rect 1146 4864 1152 4928
rect 1216 4864 1232 4928
rect 1296 4864 1312 4928
rect 1376 4864 1392 4928
rect 1456 4864 1462 4928
rect 1146 4863 1462 4864
rect 2466 4928 2782 4929
rect 2466 4864 2472 4928
rect 2536 4864 2552 4928
rect 2616 4864 2632 4928
rect 2696 4864 2712 4928
rect 2776 4864 2782 4928
rect 2466 4863 2782 4864
rect 3786 4928 4102 4929
rect 3786 4864 3792 4928
rect 3856 4864 3872 4928
rect 3936 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4102 4928
rect 3786 4863 4102 4864
rect 1806 4384 2122 4385
rect 1806 4320 1812 4384
rect 1876 4320 1892 4384
rect 1956 4320 1972 4384
rect 2036 4320 2052 4384
rect 2116 4320 2122 4384
rect 1806 4319 2122 4320
rect 3126 4384 3442 4385
rect 3126 4320 3132 4384
rect 3196 4320 3212 4384
rect 3276 4320 3292 4384
rect 3356 4320 3372 4384
rect 3436 4320 3442 4384
rect 3126 4319 3442 4320
rect 1146 3840 1462 3841
rect 1146 3776 1152 3840
rect 1216 3776 1232 3840
rect 1296 3776 1312 3840
rect 1376 3776 1392 3840
rect 1456 3776 1462 3840
rect 1146 3775 1462 3776
rect 2466 3840 2782 3841
rect 2466 3776 2472 3840
rect 2536 3776 2552 3840
rect 2616 3776 2632 3840
rect 2696 3776 2712 3840
rect 2776 3776 2782 3840
rect 2466 3775 2782 3776
rect 3786 3840 4102 3841
rect 3786 3776 3792 3840
rect 3856 3776 3872 3840
rect 3936 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4102 3840
rect 3786 3775 4102 3776
rect 1806 3296 2122 3297
rect 1806 3232 1812 3296
rect 1876 3232 1892 3296
rect 1956 3232 1972 3296
rect 2036 3232 2052 3296
rect 2116 3232 2122 3296
rect 1806 3231 2122 3232
rect 3126 3296 3442 3297
rect 3126 3232 3132 3296
rect 3196 3232 3212 3296
rect 3276 3232 3292 3296
rect 3356 3232 3372 3296
rect 3436 3232 3442 3296
rect 3126 3231 3442 3232
rect 1146 2752 1462 2753
rect 1146 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1462 2752
rect 1146 2687 1462 2688
rect 2466 2752 2782 2753
rect 2466 2688 2472 2752
rect 2536 2688 2552 2752
rect 2616 2688 2632 2752
rect 2696 2688 2712 2752
rect 2776 2688 2782 2752
rect 2466 2687 2782 2688
rect 3786 2752 4102 2753
rect 3786 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4102 2752
rect 3786 2687 4102 2688
rect 1806 2208 2122 2209
rect 1806 2144 1812 2208
rect 1876 2144 1892 2208
rect 1956 2144 1972 2208
rect 2036 2144 2052 2208
rect 2116 2144 2122 2208
rect 1806 2143 2122 2144
rect 3126 2208 3442 2209
rect 3126 2144 3132 2208
rect 3196 2144 3212 2208
rect 3276 2144 3292 2208
rect 3356 2144 3372 2208
rect 3436 2144 3442 2208
rect 3126 2143 3442 2144
<< via3 >>
rect 1812 5468 1876 5472
rect 1812 5412 1816 5468
rect 1816 5412 1872 5468
rect 1872 5412 1876 5468
rect 1812 5408 1876 5412
rect 1892 5468 1956 5472
rect 1892 5412 1896 5468
rect 1896 5412 1952 5468
rect 1952 5412 1956 5468
rect 1892 5408 1956 5412
rect 1972 5468 2036 5472
rect 1972 5412 1976 5468
rect 1976 5412 2032 5468
rect 2032 5412 2036 5468
rect 1972 5408 2036 5412
rect 2052 5468 2116 5472
rect 2052 5412 2056 5468
rect 2056 5412 2112 5468
rect 2112 5412 2116 5468
rect 2052 5408 2116 5412
rect 3132 5468 3196 5472
rect 3132 5412 3136 5468
rect 3136 5412 3192 5468
rect 3192 5412 3196 5468
rect 3132 5408 3196 5412
rect 3212 5468 3276 5472
rect 3212 5412 3216 5468
rect 3216 5412 3272 5468
rect 3272 5412 3276 5468
rect 3212 5408 3276 5412
rect 3292 5468 3356 5472
rect 3292 5412 3296 5468
rect 3296 5412 3352 5468
rect 3352 5412 3356 5468
rect 3292 5408 3356 5412
rect 3372 5468 3436 5472
rect 3372 5412 3376 5468
rect 3376 5412 3432 5468
rect 3432 5412 3436 5468
rect 3372 5408 3436 5412
rect 1152 4924 1216 4928
rect 1152 4868 1156 4924
rect 1156 4868 1212 4924
rect 1212 4868 1216 4924
rect 1152 4864 1216 4868
rect 1232 4924 1296 4928
rect 1232 4868 1236 4924
rect 1236 4868 1292 4924
rect 1292 4868 1296 4924
rect 1232 4864 1296 4868
rect 1312 4924 1376 4928
rect 1312 4868 1316 4924
rect 1316 4868 1372 4924
rect 1372 4868 1376 4924
rect 1312 4864 1376 4868
rect 1392 4924 1456 4928
rect 1392 4868 1396 4924
rect 1396 4868 1452 4924
rect 1452 4868 1456 4924
rect 1392 4864 1456 4868
rect 2472 4924 2536 4928
rect 2472 4868 2476 4924
rect 2476 4868 2532 4924
rect 2532 4868 2536 4924
rect 2472 4864 2536 4868
rect 2552 4924 2616 4928
rect 2552 4868 2556 4924
rect 2556 4868 2612 4924
rect 2612 4868 2616 4924
rect 2552 4864 2616 4868
rect 2632 4924 2696 4928
rect 2632 4868 2636 4924
rect 2636 4868 2692 4924
rect 2692 4868 2696 4924
rect 2632 4864 2696 4868
rect 2712 4924 2776 4928
rect 2712 4868 2716 4924
rect 2716 4868 2772 4924
rect 2772 4868 2776 4924
rect 2712 4864 2776 4868
rect 3792 4924 3856 4928
rect 3792 4868 3796 4924
rect 3796 4868 3852 4924
rect 3852 4868 3856 4924
rect 3792 4864 3856 4868
rect 3872 4924 3936 4928
rect 3872 4868 3876 4924
rect 3876 4868 3932 4924
rect 3932 4868 3936 4924
rect 3872 4864 3936 4868
rect 3952 4924 4016 4928
rect 3952 4868 3956 4924
rect 3956 4868 4012 4924
rect 4012 4868 4016 4924
rect 3952 4864 4016 4868
rect 4032 4924 4096 4928
rect 4032 4868 4036 4924
rect 4036 4868 4092 4924
rect 4092 4868 4096 4924
rect 4032 4864 4096 4868
rect 1812 4380 1876 4384
rect 1812 4324 1816 4380
rect 1816 4324 1872 4380
rect 1872 4324 1876 4380
rect 1812 4320 1876 4324
rect 1892 4380 1956 4384
rect 1892 4324 1896 4380
rect 1896 4324 1952 4380
rect 1952 4324 1956 4380
rect 1892 4320 1956 4324
rect 1972 4380 2036 4384
rect 1972 4324 1976 4380
rect 1976 4324 2032 4380
rect 2032 4324 2036 4380
rect 1972 4320 2036 4324
rect 2052 4380 2116 4384
rect 2052 4324 2056 4380
rect 2056 4324 2112 4380
rect 2112 4324 2116 4380
rect 2052 4320 2116 4324
rect 3132 4380 3196 4384
rect 3132 4324 3136 4380
rect 3136 4324 3192 4380
rect 3192 4324 3196 4380
rect 3132 4320 3196 4324
rect 3212 4380 3276 4384
rect 3212 4324 3216 4380
rect 3216 4324 3272 4380
rect 3272 4324 3276 4380
rect 3212 4320 3276 4324
rect 3292 4380 3356 4384
rect 3292 4324 3296 4380
rect 3296 4324 3352 4380
rect 3352 4324 3356 4380
rect 3292 4320 3356 4324
rect 3372 4380 3436 4384
rect 3372 4324 3376 4380
rect 3376 4324 3432 4380
rect 3432 4324 3436 4380
rect 3372 4320 3436 4324
rect 1152 3836 1216 3840
rect 1152 3780 1156 3836
rect 1156 3780 1212 3836
rect 1212 3780 1216 3836
rect 1152 3776 1216 3780
rect 1232 3836 1296 3840
rect 1232 3780 1236 3836
rect 1236 3780 1292 3836
rect 1292 3780 1296 3836
rect 1232 3776 1296 3780
rect 1312 3836 1376 3840
rect 1312 3780 1316 3836
rect 1316 3780 1372 3836
rect 1372 3780 1376 3836
rect 1312 3776 1376 3780
rect 1392 3836 1456 3840
rect 1392 3780 1396 3836
rect 1396 3780 1452 3836
rect 1452 3780 1456 3836
rect 1392 3776 1456 3780
rect 2472 3836 2536 3840
rect 2472 3780 2476 3836
rect 2476 3780 2532 3836
rect 2532 3780 2536 3836
rect 2472 3776 2536 3780
rect 2552 3836 2616 3840
rect 2552 3780 2556 3836
rect 2556 3780 2612 3836
rect 2612 3780 2616 3836
rect 2552 3776 2616 3780
rect 2632 3836 2696 3840
rect 2632 3780 2636 3836
rect 2636 3780 2692 3836
rect 2692 3780 2696 3836
rect 2632 3776 2696 3780
rect 2712 3836 2776 3840
rect 2712 3780 2716 3836
rect 2716 3780 2772 3836
rect 2772 3780 2776 3836
rect 2712 3776 2776 3780
rect 3792 3836 3856 3840
rect 3792 3780 3796 3836
rect 3796 3780 3852 3836
rect 3852 3780 3856 3836
rect 3792 3776 3856 3780
rect 3872 3836 3936 3840
rect 3872 3780 3876 3836
rect 3876 3780 3932 3836
rect 3932 3780 3936 3836
rect 3872 3776 3936 3780
rect 3952 3836 4016 3840
rect 3952 3780 3956 3836
rect 3956 3780 4012 3836
rect 4012 3780 4016 3836
rect 3952 3776 4016 3780
rect 4032 3836 4096 3840
rect 4032 3780 4036 3836
rect 4036 3780 4092 3836
rect 4092 3780 4096 3836
rect 4032 3776 4096 3780
rect 1812 3292 1876 3296
rect 1812 3236 1816 3292
rect 1816 3236 1872 3292
rect 1872 3236 1876 3292
rect 1812 3232 1876 3236
rect 1892 3292 1956 3296
rect 1892 3236 1896 3292
rect 1896 3236 1952 3292
rect 1952 3236 1956 3292
rect 1892 3232 1956 3236
rect 1972 3292 2036 3296
rect 1972 3236 1976 3292
rect 1976 3236 2032 3292
rect 2032 3236 2036 3292
rect 1972 3232 2036 3236
rect 2052 3292 2116 3296
rect 2052 3236 2056 3292
rect 2056 3236 2112 3292
rect 2112 3236 2116 3292
rect 2052 3232 2116 3236
rect 3132 3292 3196 3296
rect 3132 3236 3136 3292
rect 3136 3236 3192 3292
rect 3192 3236 3196 3292
rect 3132 3232 3196 3236
rect 3212 3292 3276 3296
rect 3212 3236 3216 3292
rect 3216 3236 3272 3292
rect 3272 3236 3276 3292
rect 3212 3232 3276 3236
rect 3292 3292 3356 3296
rect 3292 3236 3296 3292
rect 3296 3236 3352 3292
rect 3352 3236 3356 3292
rect 3292 3232 3356 3236
rect 3372 3292 3436 3296
rect 3372 3236 3376 3292
rect 3376 3236 3432 3292
rect 3432 3236 3436 3292
rect 3372 3232 3436 3236
rect 1152 2748 1216 2752
rect 1152 2692 1156 2748
rect 1156 2692 1212 2748
rect 1212 2692 1216 2748
rect 1152 2688 1216 2692
rect 1232 2748 1296 2752
rect 1232 2692 1236 2748
rect 1236 2692 1292 2748
rect 1292 2692 1296 2748
rect 1232 2688 1296 2692
rect 1312 2748 1376 2752
rect 1312 2692 1316 2748
rect 1316 2692 1372 2748
rect 1372 2692 1376 2748
rect 1312 2688 1376 2692
rect 1392 2748 1456 2752
rect 1392 2692 1396 2748
rect 1396 2692 1452 2748
rect 1452 2692 1456 2748
rect 1392 2688 1456 2692
rect 2472 2748 2536 2752
rect 2472 2692 2476 2748
rect 2476 2692 2532 2748
rect 2532 2692 2536 2748
rect 2472 2688 2536 2692
rect 2552 2748 2616 2752
rect 2552 2692 2556 2748
rect 2556 2692 2612 2748
rect 2612 2692 2616 2748
rect 2552 2688 2616 2692
rect 2632 2748 2696 2752
rect 2632 2692 2636 2748
rect 2636 2692 2692 2748
rect 2692 2692 2696 2748
rect 2632 2688 2696 2692
rect 2712 2748 2776 2752
rect 2712 2692 2716 2748
rect 2716 2692 2772 2748
rect 2772 2692 2776 2748
rect 2712 2688 2776 2692
rect 3792 2748 3856 2752
rect 3792 2692 3796 2748
rect 3796 2692 3852 2748
rect 3852 2692 3856 2748
rect 3792 2688 3856 2692
rect 3872 2748 3936 2752
rect 3872 2692 3876 2748
rect 3876 2692 3932 2748
rect 3932 2692 3936 2748
rect 3872 2688 3936 2692
rect 3952 2748 4016 2752
rect 3952 2692 3956 2748
rect 3956 2692 4012 2748
rect 4012 2692 4016 2748
rect 3952 2688 4016 2692
rect 4032 2748 4096 2752
rect 4032 2692 4036 2748
rect 4036 2692 4092 2748
rect 4092 2692 4096 2748
rect 4032 2688 4096 2692
rect 1812 2204 1876 2208
rect 1812 2148 1816 2204
rect 1816 2148 1872 2204
rect 1872 2148 1876 2204
rect 1812 2144 1876 2148
rect 1892 2204 1956 2208
rect 1892 2148 1896 2204
rect 1896 2148 1952 2204
rect 1952 2148 1956 2204
rect 1892 2144 1956 2148
rect 1972 2204 2036 2208
rect 1972 2148 1976 2204
rect 1976 2148 2032 2204
rect 2032 2148 2036 2204
rect 1972 2144 2036 2148
rect 2052 2204 2116 2208
rect 2052 2148 2056 2204
rect 2056 2148 2112 2204
rect 2112 2148 2116 2204
rect 2052 2144 2116 2148
rect 3132 2204 3196 2208
rect 3132 2148 3136 2204
rect 3136 2148 3192 2204
rect 3192 2148 3196 2204
rect 3132 2144 3196 2148
rect 3212 2204 3276 2208
rect 3212 2148 3216 2204
rect 3216 2148 3272 2204
rect 3272 2148 3276 2204
rect 3212 2144 3276 2148
rect 3292 2204 3356 2208
rect 3292 2148 3296 2204
rect 3296 2148 3352 2204
rect 3352 2148 3356 2204
rect 3292 2144 3356 2148
rect 3372 2204 3436 2208
rect 3372 2148 3376 2204
rect 3376 2148 3432 2204
rect 3432 2148 3436 2204
rect 3372 2144 3436 2148
<< metal4 >>
rect 1144 5134 1464 5488
rect 1144 4928 1186 5134
rect 1422 4928 1464 5134
rect 1144 4864 1152 4928
rect 1216 4864 1232 4898
rect 1296 4864 1312 4898
rect 1376 4864 1392 4898
rect 1456 4864 1464 4928
rect 1144 3840 1464 4864
rect 1144 3776 1152 3840
rect 1216 3814 1232 3840
rect 1296 3814 1312 3840
rect 1376 3814 1392 3840
rect 1456 3776 1464 3840
rect 1144 3578 1186 3776
rect 1422 3578 1464 3776
rect 1144 2752 1464 3578
rect 1144 2688 1152 2752
rect 1216 2688 1232 2752
rect 1296 2688 1312 2752
rect 1376 2688 1392 2752
rect 1456 2688 1464 2752
rect 1144 2494 1464 2688
rect 1144 2258 1186 2494
rect 1422 2258 1464 2494
rect 1144 2128 1464 2258
rect 1804 5472 2124 5488
rect 1804 5408 1812 5472
rect 1876 5408 1892 5472
rect 1956 5408 1972 5472
rect 2036 5408 2052 5472
rect 2116 5408 2124 5472
rect 1804 4474 2124 5408
rect 1804 4384 1846 4474
rect 2082 4384 2124 4474
rect 1804 4320 1812 4384
rect 2116 4320 2124 4384
rect 1804 4238 1846 4320
rect 2082 4238 2124 4320
rect 1804 3296 2124 4238
rect 1804 3232 1812 3296
rect 1876 3232 1892 3296
rect 1956 3232 1972 3296
rect 2036 3232 2052 3296
rect 2116 3232 2124 3296
rect 1804 3154 2124 3232
rect 1804 2918 1846 3154
rect 2082 2918 2124 3154
rect 1804 2208 2124 2918
rect 1804 2144 1812 2208
rect 1876 2144 1892 2208
rect 1956 2144 1972 2208
rect 2036 2144 2052 2208
rect 2116 2144 2124 2208
rect 1804 2128 2124 2144
rect 2464 5134 2784 5488
rect 2464 4928 2506 5134
rect 2742 4928 2784 5134
rect 2464 4864 2472 4928
rect 2536 4864 2552 4898
rect 2616 4864 2632 4898
rect 2696 4864 2712 4898
rect 2776 4864 2784 4928
rect 2464 3840 2784 4864
rect 2464 3776 2472 3840
rect 2536 3814 2552 3840
rect 2616 3814 2632 3840
rect 2696 3814 2712 3840
rect 2776 3776 2784 3840
rect 2464 3578 2506 3776
rect 2742 3578 2784 3776
rect 2464 2752 2784 3578
rect 2464 2688 2472 2752
rect 2536 2688 2552 2752
rect 2616 2688 2632 2752
rect 2696 2688 2712 2752
rect 2776 2688 2784 2752
rect 2464 2494 2784 2688
rect 2464 2258 2506 2494
rect 2742 2258 2784 2494
rect 2464 2128 2784 2258
rect 3124 5472 3444 5488
rect 3124 5408 3132 5472
rect 3196 5408 3212 5472
rect 3276 5408 3292 5472
rect 3356 5408 3372 5472
rect 3436 5408 3444 5472
rect 3124 4474 3444 5408
rect 3124 4384 3166 4474
rect 3402 4384 3444 4474
rect 3124 4320 3132 4384
rect 3436 4320 3444 4384
rect 3124 4238 3166 4320
rect 3402 4238 3444 4320
rect 3124 3296 3444 4238
rect 3124 3232 3132 3296
rect 3196 3232 3212 3296
rect 3276 3232 3292 3296
rect 3356 3232 3372 3296
rect 3436 3232 3444 3296
rect 3124 3154 3444 3232
rect 3124 2918 3166 3154
rect 3402 2918 3444 3154
rect 3124 2208 3444 2918
rect 3124 2144 3132 2208
rect 3196 2144 3212 2208
rect 3276 2144 3292 2208
rect 3356 2144 3372 2208
rect 3436 2144 3444 2208
rect 3124 2128 3444 2144
rect 3784 5134 4104 5488
rect 3784 4928 3826 5134
rect 4062 4928 4104 5134
rect 3784 4864 3792 4928
rect 3856 4864 3872 4898
rect 3936 4864 3952 4898
rect 4016 4864 4032 4898
rect 4096 4864 4104 4928
rect 3784 3840 4104 4864
rect 3784 3776 3792 3840
rect 3856 3814 3872 3840
rect 3936 3814 3952 3840
rect 4016 3814 4032 3840
rect 4096 3776 4104 3840
rect 3784 3578 3826 3776
rect 4062 3578 4104 3776
rect 3784 2752 4104 3578
rect 3784 2688 3792 2752
rect 3856 2688 3872 2752
rect 3936 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4104 2752
rect 3784 2494 4104 2688
rect 3784 2258 3826 2494
rect 4062 2258 4104 2494
rect 3784 2128 4104 2258
<< via4 >>
rect 1186 4928 1422 5134
rect 1186 4898 1216 4928
rect 1216 4898 1232 4928
rect 1232 4898 1296 4928
rect 1296 4898 1312 4928
rect 1312 4898 1376 4928
rect 1376 4898 1392 4928
rect 1392 4898 1422 4928
rect 1186 3776 1216 3814
rect 1216 3776 1232 3814
rect 1232 3776 1296 3814
rect 1296 3776 1312 3814
rect 1312 3776 1376 3814
rect 1376 3776 1392 3814
rect 1392 3776 1422 3814
rect 1186 3578 1422 3776
rect 1186 2258 1422 2494
rect 1846 4384 2082 4474
rect 1846 4320 1876 4384
rect 1876 4320 1892 4384
rect 1892 4320 1956 4384
rect 1956 4320 1972 4384
rect 1972 4320 2036 4384
rect 2036 4320 2052 4384
rect 2052 4320 2082 4384
rect 1846 4238 2082 4320
rect 1846 2918 2082 3154
rect 2506 4928 2742 5134
rect 2506 4898 2536 4928
rect 2536 4898 2552 4928
rect 2552 4898 2616 4928
rect 2616 4898 2632 4928
rect 2632 4898 2696 4928
rect 2696 4898 2712 4928
rect 2712 4898 2742 4928
rect 2506 3776 2536 3814
rect 2536 3776 2552 3814
rect 2552 3776 2616 3814
rect 2616 3776 2632 3814
rect 2632 3776 2696 3814
rect 2696 3776 2712 3814
rect 2712 3776 2742 3814
rect 2506 3578 2742 3776
rect 2506 2258 2742 2494
rect 3166 4384 3402 4474
rect 3166 4320 3196 4384
rect 3196 4320 3212 4384
rect 3212 4320 3276 4384
rect 3276 4320 3292 4384
rect 3292 4320 3356 4384
rect 3356 4320 3372 4384
rect 3372 4320 3402 4384
rect 3166 4238 3402 4320
rect 3166 2918 3402 3154
rect 3826 4928 4062 5134
rect 3826 4898 3856 4928
rect 3856 4898 3872 4928
rect 3872 4898 3936 4928
rect 3936 4898 3952 4928
rect 3952 4898 4016 4928
rect 4016 4898 4032 4928
rect 4032 4898 4062 4928
rect 3826 3776 3856 3814
rect 3856 3776 3872 3814
rect 3872 3776 3936 3814
rect 3936 3776 3952 3814
rect 3952 3776 4016 3814
rect 4016 3776 4032 3814
rect 4032 3776 4062 3814
rect 3826 3578 4062 3776
rect 3826 2258 4062 2494
<< metal5 >>
rect 1056 5134 4464 5176
rect 1056 4898 1186 5134
rect 1422 4898 2506 5134
rect 2742 4898 3826 5134
rect 4062 4898 4464 5134
rect 1056 4856 4464 4898
rect 1056 4474 4464 4516
rect 1056 4238 1846 4474
rect 2082 4238 3166 4474
rect 3402 4238 4464 4474
rect 1056 4196 4464 4238
rect 1056 3814 4464 3856
rect 1056 3578 1186 3814
rect 1422 3578 2506 3814
rect 2742 3578 3826 3814
rect 4062 3578 4464 3814
rect 1056 3536 4464 3578
rect 1056 3154 4464 3196
rect 1056 2918 1846 3154
rect 2082 2918 3166 3154
rect 3402 2918 4464 3154
rect 1056 2876 4464 2918
rect 1056 2494 4464 2536
rect 1056 2258 1186 2494
rect 1422 2258 2506 2494
rect 2742 2258 3826 2494
rect 4062 2258 4464 2494
rect 1056 2216 4464 2258
use sky130_fd_sc_hd__or2b_1  _06_ std
timestamp 1728241097
transform 1 0 2852 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _07_ std
timestamp 1728241097
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _08_
timestamp 1728241097
transform 1 0 1840 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1728241097
transform 1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _10_ std
timestamp 1728241097
transform -1 0 3680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _11_ std
timestamp 1728241097
transform 1 0 1380 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1728241097
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _13_ std
timestamp 1728241097
transform 1 0 2300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1728241097
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _15_
timestamp 1728241097
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1728241097
transform -1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _17_ std
timestamp 1728241097
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _18_ std
timestamp 1728241097
transform 1 0 3404 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1728241097
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 std
timestamp 1728241097
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_8
timestamp 1728241097
transform 1 0 1840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_32 std
timestamp 1728241097
transform 1 0 4048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_17
timestamp 1728241097
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1728241097
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_7
timestamp 1728241097
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_14 std
timestamp 1728241097
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1728241097
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29 std
timestamp 1728241097
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_6 std
timestamp 1728241097
transform 1 0 1656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_12
timestamp 1728241097
transform 1 0 2208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_22 std
timestamp 1728241097
transform 1 0 3128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_30 std
timestamp 1728241097
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_12
timestamp 1728241097
transform 1 0 2208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_24
timestamp 1728241097
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1728241097
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_13
timestamp 1728241097
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_17
timestamp 1728241097
transform 1 0 2668 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_29
timestamp 1728241097
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 std
timestamp 1728241097
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1728241097
transform -1 0 3680 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  output3 std
timestamp 1728241097
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output4
timestamp 1728241097
transform -1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1728241097
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output6
timestamp 1728241097
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1728241097
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1728241097
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1728241097
transform 1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output10
timestamp 1728241097
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_6
timestamp 1728241097
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1728241097
transform -1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_7
timestamp 1728241097
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1728241097
transform -1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_8
timestamp 1728241097
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1728241097
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_9
timestamp 1728241097
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1728241097
transform -1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_10
timestamp 1728241097
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1728241097
transform -1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_11
timestamp 1728241097
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1728241097
transform -1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_12 std
timestamp 1728241097
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_13
timestamp 1728241097
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_14
timestamp 1728241097
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_15
timestamp 1728241097
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
<< labels >>
rlabel metal1 s 2760 5440 2760 5440 4 VGND
rlabel metal2 s 2760 4896 2760 4896 4 VPWR
rlabel metal1 s 4002 2516 4002 2516 4 _00_
rlabel metal1 s 2484 3026 2484 3026 4 _01_
rlabel metal2 s 1794 2618 1794 2618 4 _02_
rlabel metal1 s 3082 4080 3082 4080 4 _03_
rlabel metal1 s 1978 4624 1978 4624 4 _04_
rlabel metal1 s 3956 3026 3956 3026 4 _05_
rlabel metal2 s 3082 1656 3082 1656 4 gno2
rlabel metal2 s 2438 1520 2438 1520 4 gpo1
rlabel metal2 s 3726 1656 3726 1656 4 gpo2
rlabel metal2 s 1702 4930 1702 4930 4 net1
rlabel metal1 s 2898 2448 2898 2448 4 net10
rlabel metal1 s 2898 3978 2898 3978 4 net2
rlabel metal1 s 2346 3536 2346 3536 4 net3
rlabel metal1 s 2116 3502 2116 3502 4 net4
rlabel metal1 s 2346 2380 2346 2380 4 net5
rlabel metal1 s 2714 2414 2714 2414 4 net6
rlabel metal2 s 1610 3366 1610 3366 4 net7
rlabel metal2 s 2070 2618 2070 2618 4 net8
rlabel metal1 s 3174 2380 3174 2380 4 net9
rlabel metal2 s 1426 5355 1426 5355 4 select[0]
rlabel metal1 s 3864 5202 3864 5202 4 select[1]
flabel metal5 s 1056 4196 4464 4516 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 2876 4464 3196 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 3124 2128 3444 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1804 2128 2124 5488 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4856 4464 5176 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3536 4464 3856 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 2216 4464 2536 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 3784 2128 4104 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2464 2128 2784 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1144 2128 1464 5488 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 1776 5709 1832 6200 0 FreeSans 280 90 0 0 select[1]
port 12 nsew
flabel metal2 s 1306 5699 1362 6200 0 FreeSans 280 90 0 0 select[0]
port 11 nsew
flabel metal2 s 1768 1450 1824 1932 0 FreeSans 280 90 0 0 gno1
port 4 nsew
flabel metal2 s 3056 1450 3112 1932 0 FreeSans 280 90 0 0 gno2
port 5 nsew
flabel metal2 s 4344 1450 4400 1932 0 FreeSans 280 90 0 0 gno3
port 6 nsew
flabel metal2 s 1124 1450 1180 1932 0 FreeSans 280 90 0 0 gpo0
port 7 nsew
flabel metal2 s 2412 1450 2468 1932 0 FreeSans 280 90 0 0 gpo1
port 8 nsew
flabel metal2 s 3700 1450 3756 1932 0 FreeSans 280 90 0 0 gpo2
port 9 nsew
rlabel metal2 s 816 2198 816 2198 4 gno0
flabel metal2 s 790 1450 846 1930 0 FreeSans 280 90 0 0 gno0
port 3 nsew
rlabel metal2 s 4668 1520 4668 1520 4 gpo3
flabel metal2 s 4642 1450 4698 1932 0 FreeSans 280 90 0 0 gpo3
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 5551 7695
string GDS_END 119538
string GDS_FILE /tmp/passgatesCtrl.gds
string GDS_START 63214
<< end >>
