* NGSPICE file created from mux8onehot_parax.ext - technology: sky130A

.subckt mux8onehot_parax select1 select2 A1 A3 A2 A4 Z A8 select0 A7 A6 VPWR A5 VGND
X0 a_5645_5909# a_5645_6085# a_5671_6037# VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X1 VGND.t6 select1.t0 a_5645_6085# VGND.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X2 x5.A select2.t0 Z.t5 VPWR.t31 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X3 x3.Z3 x1.gno0.t2 A5.t3 VGND.t15 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X4 VGND.t50 a_5645_6461# x1.gno2 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X5 x1.gpo3.t3 x1.gno3.t2 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X6 x1.nSEL2 select2.t1 VPWR.t30 VPWR.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X7 VGND.t38 a_5645_5909# x1.gno1 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X8 VPWR.t59 select0.t0 x1.nSEL0 VPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X9 x5.A select2.t2 Z.t4 VPWR.t28 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X10 A1.t1 x1.gpo0.t4 x5.A VPWR.t60 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X11 x5.A x1.gno1 A2.t2 VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X12 VPWR.t74 VGND.t76 VPWR.t73 VPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X13 x3.Z3 x1.nSEL2 Z.t3 VPWR.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X14 x1.nSEL0 select0.t1 VPWR.t53 VPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X15 x5.A x1.gno3.t3 A4.t1 VGND.t22 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X16 VGND.t67 VPWR.t79 VGND.t66 VGND.t65 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X17 a_5671_6037# select0.t2 VGND.t36 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X18 A7.t3 x1.gpo2 x3.Z3 VPWR.t77 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X19 x3.Z3 x1.nSEL2 Z.t2 VPWR.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X20 Z.t1 x1.nSEL2 x5.A VGND.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X21 A3.t3 x1.gpo2 x5.A VPWR.t78 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X22 VGND.t75 select1.t1 x1.nSEL1 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X23 x1.gpo3.t1 x1.gno3.t4 VPWR.t33 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X24 Z.t7 select2.t3 x3.Z3 VGND.t70 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X25 VGND.t3 a_5645_7149# x1.gno3.t1 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X26 VPWR.t57 a_5645_6637# a_5645_6461# VPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X27 x3.Z3 x1.gno1 A6.t3 VGND.t44 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X28 a_5645_7149# select1.t2 a_5699_7287# VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X29 x3.Z3 x1.gno0.t3 A5.t2 VGND.t15 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X30 a_5645_6637# select0.t3 VPWR.t21 VPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X31 VGND.t24 x1.gno0.t4 x1.gpo0.t3 VGND.t23 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X32 a_5699_7287# select0.t4 VGND.t62 VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X33 VGND.t9 VPWR.t80 VGND.t8 VGND.t7 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X34 x5.A x1.gno2 A3.t1 VGND.t30 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X35 A8.t3 x1.gpo3.t4 x3.Z3 VPWR.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X36 A1.t0 x1.gpo0.t5 x5.A VPWR.t60 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X37 a_5645_6461# a_5645_6637# a_5671_6589# VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X38 x5.A x1.gno3.t5 A4.t0 VGND.t22 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X39 VGND.t32 x1.gno2 x1.gpo2 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X40 x1.gpo0.t2 x1.gno0.t5 VGND.t34 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X41 VGND.t64 select0.t5 a_5645_6637# VGND.t63 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X42 Z.t0 x1.nSEL2 x5.A VGND.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X43 VPWR.t19 select1.t3 x1.nSEL1 VPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X44 VPWR.t17 select1.t4 a_5645_7149# VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X45 A5.t1 x1.gpo0.t6 x3.Z3 VPWR.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X46 VPWR.t71 VGND.t77 VPWR.t70 VPWR.t69 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X47 Z.t6 select2.t4 x3.Z3 VGND.t57 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X48 VPWR.t41 a_5645_5493# x1.gno0.t0 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X49 a_5645_7149# select0.t6 VPWR.t62 VPWR.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X50 VPWR.t76 x1.gno0.t6 x1.gpo0.t1 VPWR.t75 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X51 x3.Z3 x1.gno2 A7.t1 VGND.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X52 x3.Z3 x1.gno1 A6.t2 VGND.t44 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X53 A4.t3 x1.gpo3.t5 x5.A VPWR.t22 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X54 VGND.t19 select2.t5 x1.nSEL2 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X55 a_5645_5493# x1.nSEL0 a_5699_5631# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X56 x1.nSEL1 select1.t5 VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X57 x5.A x1.gno0.t7 A1.t3 VGND.t4 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X58 VPWR.t25 x1.gno2 x1.gpo2 VPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X59 x1.gpo0.t0 x1.gno0.t8 VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X60 a_5645_5909# select0.t7 VPWR.t43 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X61 x5.A x1.gno2 A3.t0 VGND.t30 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X62 A2.t3 x1.gpo1.t4 x5.A VPWR.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X63 x5.A x1.gno0.t9 A1.t2 VGND.t4 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X64 A3.t2 x1.gpo2 x5.A VPWR.t78 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X65 VPWR.t68 VGND.t78 VPWR.t67 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X66 a_5699_5631# x1.nSEL1 VGND.t52 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X67 VGND.t73 VPWR.t81 VGND.t72 VGND.t71 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X68 x3.Z3 x1.gno3.t6 A8.t1 VGND.t14 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X69 VPWR.t45 a_5645_6461# x1.gno2 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X70 VGND.t43 x1.gno1 x1.gpo1.t3 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X71 A6.t1 x1.gpo1.t5 x3.Z3 VPWR.t6 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X72 A5.t0 x1.gpo0.t7 x3.Z3 VPWR.t4 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X73 VPWR.t51 x1.nSEL0 a_5645_5493# VPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X74 x1.gpo1.t2 x1.gno1 VGND.t41 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X75 VGND.t69 x1.gno3.t7 x1.gpo3.t2 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X76 VPWR.t35 a_5645_5909# x1.gno1 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X77 x1.gpo2 x1.gno2 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X78 A7.t2 x1.gpo2 x3.Z3 VPWR.t77 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X79 x1.nSEL1 select1.t6 VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X80 VPWR.t27 select2.t6 x1.nSEL2 VPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X81 a_5671_6589# select1.t7 VGND.t21 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X82 x3.Z3 x1.gno2 A7.t0 VGND.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X83 A8.t2 x1.gpo3.t6 x3.Z3 VPWR.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X84 A4.t2 x1.gpo3.t7 x5.A VPWR.t22 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X85 a_5645_5493# x1.nSEL1 VPWR.t47 VPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X86 VGND.t46 a_5645_5493# x1.gno0.t1 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X87 VGND.t55 VPWR.t82 VGND.t54 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X88 x5.A x1.gno1 A2.t1 VGND.t39 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X89 VPWR.t39 x1.gno1 x1.gpo1.t1 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X90 A2.t0 x1.gpo1.t6 x5.A VPWR.t5 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X91 VPWR.t3 a_5645_7149# x1.gno3.t0 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X92 x1.nSEL2 select2.t7 VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X93 VGND.t48 select0.t8 x1.nSEL0 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X94 x1.gpo1.t0 x1.gno1 VPWR.t37 VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X95 VPWR.t49 x1.gno3.t8 x1.gpo3.t0 VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X96 x3.Z3 x1.gno3.t9 A8.t0 VGND.t14 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X97 VPWR.t55 a_5645_6085# a_5645_5909# VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X98 x1.gpo2 x1.gno2 VPWR.t24 VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X99 VPWR.t65 VGND.t79 VPWR.t64 VPWR.t63 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X100 a_5645_6085# select1.t8 VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X101 x1.nSEL0 select0.t9 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X102 a_5645_6461# select1.t9 VPWR.t11 VPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X103 A6.t0 x1.gpo1.t7 x3.Z3 VPWR.t6 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
R0 VGND.n237 VGND.n236 587674
R1 VGND.n171 VGND.n170 153375
R2 VGND.n193 VGND.n178 117542
R3 VGND.n249 VGND.n172 71206.2
R4 VGND.n249 VGND.n248 64736.2
R5 VGND.n238 VGND.n9 16580.8
R6 VGND.n242 VGND.n173 11744.7
R7 VGND.n247 VGND.n173 11744.7
R8 VGND.n242 VGND.n174 11744.7
R9 VGND.n247 VGND.n174 11744.7
R10 VGND.n253 VGND.n28 11744.7
R11 VGND.n253 VGND.n29 11744.7
R12 VGND.n257 VGND.n29 11744.7
R13 VGND.n257 VGND.n28 11744.7
R14 VGND.n264 VGND.n22 11744.7
R15 VGND.n260 VGND.n22 11744.7
R16 VGND.n264 VGND.n23 11744.7
R17 VGND.n260 VGND.n23 11744.7
R18 VGND.n271 VGND.n16 11744.7
R19 VGND.n267 VGND.n16 11744.7
R20 VGND.n271 VGND.n17 11744.7
R21 VGND.n267 VGND.n17 11744.7
R22 VGND.n278 VGND.n10 11744.7
R23 VGND.n274 VGND.n10 11744.7
R24 VGND.n278 VGND.n11 11744.7
R25 VGND.n274 VGND.n11 11744.7
R26 VGND.n190 VGND.n179 11744.7
R27 VGND.n185 VGND.n179 11744.7
R28 VGND.n190 VGND.n181 11744.7
R29 VGND.n185 VGND.n181 11744.7
R30 VGND.n205 VGND.n204 11744.7
R31 VGND.n201 VGND.n200 11744.7
R32 VGND.n204 VGND.n201 11744.7
R33 VGND.n234 VGND.n194 11744.7
R34 VGND.n230 VGND.n195 11744.7
R35 VGND.n234 VGND.n195 11744.7
R36 VGND.n218 VGND.n217 11744.7
R37 VGND.n214 VGND.n213 11744.7
R38 VGND.n217 VGND.n214 11744.7
R39 VGND.n281 VGND.n4 11744.7
R40 VGND.n281 VGND.n5 11744.7
R41 VGND.n7 VGND.n4 11744.7
R42 VGND.n237 VGND.n178 10428.2
R43 VGND.n238 VGND.n191 7573.12
R44 VGND.n191 VGND.t0 7065.1
R45 VGND.t1 VGND.n172 7065.1
R46 VGND.n180 VGND.t0 6710.74
R47 VGND.n180 VGND.t1 6710.74
R48 VGND.n241 VGND.n239 6647.5
R49 VGND.n273 VGND.n272 6049.9
R50 VGND.n241 VGND.t70 6006.85
R51 VGND.n248 VGND.t57 6006.85
R52 VGND.n259 VGND.n258 6004.3
R53 VGND.n280 VGND.n279 5972.7
R54 VGND.n266 VGND.n265 5963.12
R55 VGND.t70 VGND.n240 5705.56
R56 VGND.n240 VGND.t57 5705.56
R57 VGND.n239 VGND.n178 4796.58
R58 VGND.n238 VGND.n237 3666.67
R59 VGND.n192 VGND.n9 3385.09
R60 VGND.n15 VGND.n9 3361.58
R61 VGND.n27 VGND.n21 3305.56
R62 VGND.n235 VGND.n193 3279.94
R63 VGND.n21 VGND.n15 3275.35
R64 VGND.n62 VGND.n27 2366.85
R65 VGND.n250 VGND.n249 2235.82
R66 VGND.n236 VGND.n235 1652.78
R67 VGND.n236 VGND.n192 1652.78
R68 VGND.t2 VGND.n169 1550.96
R69 VGND VGND.t63 1289.66
R70 VGND.n137 VGND.n136 1198.25
R71 VGND.n159 VGND.n40 1198.25
R72 VGND.n169 VGND.n168 1194.5
R73 VGND.n140 VGND.n139 1171.32
R74 VGND.n251 VGND.n250 1006.48
R75 VGND.n169 VGND 918.774
R76 VGND.t45 VGND 918.774
R77 VGND.t61 VGND.t2 910.346
R78 VGND.t20 VGND.t49 826.054
R79 VGND.t35 VGND.t37 826.054
R80 VGND.t5 VGND.t74 792.337
R81 VGND.n256 VGND.n255 767.294
R82 VGND.n270 VGND.n269 767.294
R83 VGND.n232 VGND.n231 767.294
R84 VGND.n6 VGND.n3 767.294
R85 VGND.n263 VGND.n262 763.106
R86 VGND.n277 VGND.n276 763.106
R87 VGND.n202 VGND.n198 763.106
R88 VGND.n215 VGND.n211 763.106
R89 VGND.n243 VGND.n177 763.09
R90 VGND.n189 VGND.n182 763.09
R91 VGND.n177 VGND.n175 732.236
R92 VGND.n256 VGND.n30 732.236
R93 VGND.n270 VGND.n18 732.236
R94 VGND.n263 VGND.n24 732.236
R95 VGND.n277 VGND.n12 732.236
R96 VGND.n184 VGND.n182 732.236
R97 VGND.n207 VGND.n198 732.236
R98 VGND.n231 VGND.n228 732.236
R99 VGND.n220 VGND.n211 732.236
R100 VGND.n6 VGND.n1 732.236
R101 VGND.n250 VGND.n171 709.912
R102 VGND.t18 VGND.t25 708.047
R103 VGND.t74 VGND.t16 708.047
R104 VGND.t47 VGND.t10 708.047
R105 VGND.t58 VGND.t51 708.047
R106 VGND.n139 VGND.t65 606.351
R107 VGND.t56 VGND 564.751
R108 VGND.t25 VGND 564.751
R109 VGND.t10 VGND 564.751
R110 VGND VGND.t58 564.751
R111 VGND.n171 VGND 564.751
R112 VGND.n170 VGND.t56 522.606
R113 VGND.t51 VGND.t71 522.606
R114 VGND.t59 VGND 480.461
R115 VGND VGND.t53 408.628
R116 VGND.t71 VGND.t45 387.74
R117 VGND.n138 VGND 384.901
R118 VGND.t42 VGND.n137 374.356
R119 VGND.n40 VGND.t60 337.166
R120 VGND.n252 VGND.n251 332.642
R121 VGND.t68 VGND 329.539
R122 VGND.t31 VGND 329.539
R123 VGND.t23 VGND 329.539
R124 VGND.n255 VGND.n254 325.502
R125 VGND.n269 VGND.n268 325.502
R126 VGND.n233 VGND.n232 325.502
R127 VGND.n282 VGND.n3 325.502
R128 VGND.n40 VGND.t20 320.307
R129 VGND.n244 VGND.n243 304.553
R130 VGND.n189 VGND.n188 304.553
R131 VGND.n262 VGND.n261 304.204
R132 VGND.n276 VGND.n275 304.204
R133 VGND.n203 VGND.n202 304.204
R134 VGND.n216 VGND.n215 304.204
R135 VGND.t60 VGND 295.019
R136 VGND.n245 VGND.n244 266.349
R137 VGND.n188 VGND.n187 266.349
R138 VGND VGND.t5 261.303
R139 VGND.t7 VGND 244.445
R140 VGND.n254 VGND.n32 242.448
R141 VGND.n268 VGND.n20 242.448
R142 VGND.n261 VGND.n26 242.448
R143 VGND.n275 VGND.n14 242.448
R144 VGND.n203 VGND.n197 242.448
R145 VGND.n233 VGND.n196 242.448
R146 VGND.n216 VGND.n210 242.448
R147 VGND.n283 VGND.n282 242.448
R148 VGND.n152 VGND.t6 240.575
R149 VGND.n164 VGND.t64 237.327
R150 VGND.t12 VGND.t68 221.451
R151 VGND.t28 VGND.t31 221.451
R152 VGND.t40 VGND.t42 221.451
R153 VGND.t33 VGND.t23 221.451
R154 VGND.n106 VGND.t79 218.308
R155 VGND.n82 VGND.t78 218.308
R156 VGND.n50 VGND.t77 218.308
R157 VGND.n36 VGND.t76 218.308
R158 VGND.n103 VGND.t66 214.456
R159 VGND.n105 VGND.t67 214.456
R160 VGND.n80 VGND.t54 214.456
R161 VGND.n67 VGND.t55 214.456
R162 VGND.n45 VGND.t72 214.456
R163 VGND.n49 VGND.t73 214.456
R164 VGND.n34 VGND.t8 214.456
R165 VGND.n37 VGND.t9 214.456
R166 VGND.n74 VGND.n70 204.457
R167 VGND.n146 VGND.n44 200.231
R168 VGND.n39 VGND.n38 200.231
R169 VGND.n52 VGND.n47 200.105
R170 VGND.n137 VGND 197.724
R171 VGND.n139 VGND 197.724
R172 VGND.n276 VGND.n11 195
R173 VGND.n11 VGND.t22 195
R174 VGND.n13 VGND.n10 195
R175 VGND.n10 VGND.t22 195
R176 VGND.n269 VGND.n17 195
R177 VGND.n17 VGND.t30 195
R178 VGND.n19 VGND.n16 195
R179 VGND.n16 VGND.t30 195
R180 VGND.n262 VGND.n23 195
R181 VGND.n23 VGND.t39 195
R182 VGND.n25 VGND.n22 195
R183 VGND.n22 VGND.t39 195
R184 VGND.n31 VGND.n28 195
R185 VGND.n138 VGND.n28 195
R186 VGND.n255 VGND.n29 195
R187 VGND.n29 VGND.t4 195
R188 VGND.n186 VGND.n185 195
R189 VGND.n185 VGND.n172 195
R190 VGND.n190 VGND.n189 195
R191 VGND.n191 VGND.n190 195
R192 VGND.n247 VGND.n246 195
R193 VGND.n248 VGND.n247 195
R194 VGND.n243 VGND.n242 195
R195 VGND.n242 VGND.n241 195
R196 VGND.n202 VGND.n201 195
R197 VGND.n201 VGND.t14 195
R198 VGND.n206 VGND.n205 195
R199 VGND.n232 VGND.n195 195
R200 VGND.n195 VGND.t27 195
R201 VGND.n227 VGND.n194 195
R202 VGND.n215 VGND.n214 195
R203 VGND.n214 VGND.t44 195
R204 VGND.n219 VGND.n218 195
R205 VGND.n4 VGND.n2 195
R206 VGND.t15 VGND.n4 195
R207 VGND.n5 VGND.n3 195
R208 VGND.n8 VGND.n5 188.989
R209 VGND.n218 VGND.n212 188.988
R210 VGND.n229 VGND.n194 188.986
R211 VGND.n205 VGND.n199 188.984
R212 VGND.n170 VGND.t61 185.441
R213 VGND.n258 VGND.t4 183.936
R214 VGND VGND.t35 177.012
R215 VGND VGND.t28 176.633
R216 VGND VGND.t40 176.633
R217 VGND VGND.t33 176.633
R218 VGND.n251 VGND 176.633
R219 VGND.n200 VGND.n199 173.373
R220 VGND.n230 VGND.n229 173.304
R221 VGND.n213 VGND.n212 173.167
R222 VGND.n8 VGND.n7 173.097
R223 VGND.n115 VGND.t69 162.471
R224 VGND.n120 VGND.t32 162.471
R225 VGND.n64 VGND.t43 162.471
R226 VGND.n130 VGND.t24 162.471
R227 VGND.n41 VGND.t75 162.471
R228 VGND.n146 VGND.t48 160.046
R229 VGND.n39 VGND.t19 160.046
R230 VGND.n119 VGND.t13 160.017
R231 VGND.n63 VGND.t29 160.017
R232 VGND.n131 VGND.t41 160.017
R233 VGND.n126 VGND.t34 160.017
R234 VGND.n57 VGND.t11 160.017
R235 VGND.n147 VGND.t17 160.017
R236 VGND.n152 VGND.t26 158.534
R237 VGND.n279 VGND.t22 155.954
R238 VGND.n272 VGND.t30 155.954
R239 VGND.n265 VGND.t39 155.831
R240 VGND.n252 VGND.t4 139.648
R241 VGND.n204 VGND.n193 118.54
R242 VGND.n235 VGND.n234 111.895
R243 VGND.n217 VGND.n192 111.808
R244 VGND.n273 VGND.n15 99.881
R245 VGND.n266 VGND.n21 93.748
R246 VGND.n259 VGND.n27 93.6734
R247 VGND.n62 VGND.t12 89.635
R248 VGND.n9 VGND.t15 89.4314
R249 VGND VGND.n62 86.9987
R250 VGND.t16 VGND.t59 84.2917
R251 VGND.n239 VGND.n238 79.0175
R252 VGND.n47 VGND.t52 72.8576
R253 VGND.n70 VGND.t62 72.8576
R254 VGND.n280 VGND.n9 72.6343
R255 VGND.n235 VGND.t27 66.9242
R256 VGND.t44 VGND.n192 66.8669
R257 VGND.n21 VGND.t30 62.2068
R258 VGND.n27 VGND.t39 62.1573
R259 VGND.t14 VGND.n193 60.352
R260 VGND.n44 VGND.t36 58.5719
R261 VGND.n38 VGND.t21 58.5719
R262 VGND.n15 VGND.t22 56.0738
R263 VGND.n246 VGND.n245 54.2123
R264 VGND.n187 VGND.n186 54.2123
R265 VGND.t49 VGND.t18 50.5752
R266 VGND.t37 VGND.t47 50.5752
R267 VGND.n76 VGND 43.9579
R268 VGND.n253 VGND.n252 42.2329
R269 VGND.n76 VGND.n75 34.6358
R270 VGND.n73 VGND.n33 34.6358
R271 VGND.n246 VGND.n175 30.8711
R272 VGND.n31 VGND.n30 30.8711
R273 VGND.n19 VGND.n18 30.8711
R274 VGND.n25 VGND.n24 30.8711
R275 VGND.n13 VGND.n12 30.8711
R276 VGND.n186 VGND.n184 30.8711
R277 VGND.n207 VGND.n206 30.8711
R278 VGND.n228 VGND.n227 30.8711
R279 VGND.n220 VGND.n219 30.8711
R280 VGND.n2 VGND.n1 30.8711
R281 VGND.n140 VGND.n61 26.9246
R282 VGND.n168 VGND.n33 25.6926
R283 VGND.n44 VGND.t38 25.4291
R284 VGND.n38 VGND.t50 25.4291
R285 VGND.n115 VGND.n66 25.224
R286 VGND.n119 VGND.n66 25.224
R287 VGND.n121 VGND.n120 25.224
R288 VGND.n121 VGND.n63 25.224
R289 VGND.n132 VGND.n64 25.224
R290 VGND.n132 VGND.n131 25.224
R291 VGND.n130 VGND.n129 25.224
R292 VGND.n129 VGND.n126 25.224
R293 VGND.n57 VGND.n43 25.224
R294 VGND.n148 VGND.n41 25.224
R295 VGND.n148 VGND.n147 25.224
R296 VGND.n153 VGND.n152 24.0946
R297 VGND.t65 VGND.n138 23.7273
R298 VGND.n47 VGND.t46 22.3257
R299 VGND.n70 VGND.t3 22.3257
R300 VGND.n146 VGND.n43 21.4593
R301 VGND.n153 VGND.n39 21.4593
R302 VGND.n120 VGND.n119 20.3299
R303 VGND.n131 VGND.n130 20.3299
R304 VGND.n115 VGND.n114 19.2926
R305 VGND.n57 VGND.n56 17.7867
R306 VGND.n136 VGND.n64 17.3181
R307 VGND.t63 VGND.t7 16.8587
R308 VGND.n136 VGND.n63 15.8123
R309 VGND.n126 VGND.n61 15.8123
R310 VGND.n281 VGND.n280 15.1478
R311 VGND.n102 VGND.n61 14.775
R312 VGND.n160 VGND.n159 14.775
R313 VGND.n152 VGND.n41 13.5534
R314 VGND.n79 VGND.n78 11.2844
R315 VGND.n275 VGND.n274 11.0382
R316 VGND.n274 VGND.n273 11.0382
R317 VGND.n278 VGND.n277 11.0382
R318 VGND.n279 VGND.n278 11.0382
R319 VGND.n268 VGND.n267 11.0382
R320 VGND.n267 VGND.n266 11.0382
R321 VGND.n271 VGND.n270 11.0382
R322 VGND.n272 VGND.n271 11.0382
R323 VGND.n261 VGND.n260 11.0382
R324 VGND.n260 VGND.n259 11.0382
R325 VGND.n264 VGND.n263 11.0382
R326 VGND.n265 VGND.n264 11.0382
R327 VGND.n254 VGND.n253 11.0382
R328 VGND.n257 VGND.n256 11.0382
R329 VGND.n258 VGND.n257 11.0382
R330 VGND.n188 VGND.n181 11.0382
R331 VGND.n181 VGND.n180 11.0382
R332 VGND.n182 VGND.n179 11.0382
R333 VGND.n180 VGND.n179 11.0382
R334 VGND.n244 VGND.n174 11.0382
R335 VGND.n240 VGND.n174 11.0382
R336 VGND.n177 VGND.n173 11.0382
R337 VGND.n240 VGND.n173 11.0382
R338 VGND.n204 VGND.n203 11.0382
R339 VGND.n200 VGND.n198 11.0382
R340 VGND.n234 VGND.n233 11.0382
R341 VGND.n231 VGND.n230 11.0382
R342 VGND.n217 VGND.n216 11.0382
R343 VGND.n213 VGND.n211 11.0382
R344 VGND.n7 VGND.n6 11.0382
R345 VGND.n282 VGND.n281 11.0382
R346 VGND.n32 VGND.n31 10.9181
R347 VGND.n20 VGND.n19 10.9181
R348 VGND.n26 VGND.n25 10.9181
R349 VGND.n14 VGND.n13 10.9181
R350 VGND.n206 VGND.n197 10.9181
R351 VGND.n227 VGND.n196 10.9181
R352 VGND.n219 VGND.n210 10.9181
R353 VGND.n283 VGND.n2 10.9181
R354 VGND.n176 VGND.n175 10.4476
R355 VGND.n85 VGND.n30 10.4476
R356 VGND.n89 VGND.n18 10.4476
R357 VGND.n87 VGND.n24 10.4476
R358 VGND.n91 VGND.n12 10.4476
R359 VGND.n184 VGND.n183 10.4476
R360 VGND.n208 VGND.n207 10.4476
R361 VGND.n228 VGND.n226 10.4476
R362 VGND.n221 VGND.n220 10.4476
R363 VGND.n284 VGND.n1 10.4476
R364 VGND.n147 VGND.n146 10.1652
R365 VGND.n105 VGND.n100 9.70901
R366 VGND.n80 VGND.n79 9.70901
R367 VGND.n49 VGND.n48 9.70901
R368 VGND.n74 VGND.n73 9.41227
R369 VGND.n141 VGND.n140 9.3005
R370 VGND.n127 VGND.n126 9.3005
R371 VGND.n131 VGND.n124 9.3005
R372 VGND.n136 VGND.n135 9.3005
R373 VGND.n123 VGND.n63 9.3005
R374 VGND.n119 VGND.n118 9.3005
R375 VGND.n114 VGND.n113 9.3005
R376 VGND.n84 VGND.n83 9.3005
R377 VGND.n81 VGND.n68 9.3005
R378 VGND.n116 VGND.n115 9.3005
R379 VGND.n117 VGND.n66 9.3005
R380 VGND.n120 VGND.n65 9.3005
R381 VGND.n122 VGND.n121 9.3005
R382 VGND.n134 VGND.n64 9.3005
R383 VGND.n133 VGND.n132 9.3005
R384 VGND.n130 VGND.n125 9.3005
R385 VGND.n129 VGND.n128 9.3005
R386 VGND.n108 VGND.n107 9.3005
R387 VGND.n104 VGND.n99 9.3005
R388 VGND.n102 VGND.n101 9.3005
R389 VGND.n61 VGND.n59 9.3005
R390 VGND.n168 VGND.n167 9.3005
R391 VGND.n166 VGND.n165 9.3005
R392 VGND.n157 VGND.n39 9.3005
R393 VGND.n152 VGND.n151 9.3005
R394 VGND.n146 VGND.n145 9.3005
R395 VGND.n51 VGND.n46 9.3005
R396 VGND.n54 VGND.n53 9.3005
R397 VGND.n56 VGND.n55 9.3005
R398 VGND.n58 VGND.n57 9.3005
R399 VGND.n144 VGND.n43 9.3005
R400 VGND.n147 VGND.n42 9.3005
R401 VGND.n149 VGND.n148 9.3005
R402 VGND.n150 VGND.n41 9.3005
R403 VGND.n154 VGND.n153 9.3005
R404 VGND.n161 VGND.n160 9.3005
R405 VGND.n163 VGND.n162 9.3005
R406 VGND.n71 VGND.n33 9.3005
R407 VGND.n73 VGND.n72 9.3005
R408 VGND.n75 VGND.n69 9.3005
R409 VGND.n77 VGND.n76 9.3005
R410 VGND.n159 VGND.n158 9.3005
R411 VGND.n93 VGND.n92 8.45078
R412 VGND.n224 VGND.n209 8.45078
R413 VGND.n95 VGND.n86 8.30267
R414 VGND.n285 VGND.n0 8.30267
R415 VGND.n94 VGND.n88 7.97888
R416 VGND.n223 VGND.n222 7.97888
R417 VGND.n93 VGND.n90 7.97601
R418 VGND.n225 VGND.n224 7.97601
R419 VGND.n176 VGND 7.23036
R420 VGND.n183 VGND 7.23036
R421 VGND.n86 VGND.n85 7.16724
R422 VGND.n90 VGND.n89 7.16724
R423 VGND.n88 VGND.n87 7.16724
R424 VGND.n92 VGND.n91 7.16724
R425 VGND.n209 VGND.n208 7.16724
R426 VGND.n226 VGND.n225 7.16724
R427 VGND.n222 VGND.n221 7.16724
R428 VGND.n285 VGND.n284 7.16724
R429 VGND.n159 VGND.n39 7.15344
R430 VGND.n143 VGND.n142 6.50373
R431 VGND.n75 VGND.n74 6.4005
R432 VGND.n107 VGND.n104 6.26433
R433 VGND.n83 VGND.n81 6.26433
R434 VGND.n104 VGND.n103 5.85582
R435 VGND.n81 VGND.n80 5.85582
R436 VGND.n53 VGND.n45 5.85582
R437 VGND.n165 VGND.n34 5.85582
R438 VGND.n164 VGND.n163 5.85582
R439 VGND.n142 VGND.n59 4.788
R440 VGND.n85 VGND.n32 4.73093
R441 VGND.n89 VGND.n20 4.73093
R442 VGND.n87 VGND.n26 4.73093
R443 VGND.n91 VGND.n14 4.73093
R444 VGND.n208 VGND.n197 4.73093
R445 VGND.n226 VGND.n196 4.73093
R446 VGND.n221 VGND.n210 4.73093
R447 VGND.n284 VGND.n283 4.73093
R448 VGND.n142 VGND.n141 4.50726
R449 VGND.n97 VGND 4.01425
R450 VGND.n96 VGND 4.01425
R451 VGND.n245 VGND.n176 3.78485
R452 VGND.n187 VGND.n183 3.78485
R453 VGND.n52 VGND.n51 3.40476
R454 VGND.n107 VGND.n106 3.13241
R455 VGND.n83 VGND.n82 3.13241
R456 VGND.n51 VGND.n50 3.13241
R457 VGND.n163 VGND.n36 3.13241
R458 VGND.n155 VGND.n35 2.88636
R459 VGND.t14 VGND.n199 2.87953
R460 VGND.n229 VGND.t27 2.87839
R461 VGND.t44 VGND.n212 2.87611
R462 VGND.t15 VGND.n8 2.87497
R463 VGND.n53 VGND.n52 2.86007
R464 VGND.n106 VGND.n105 2.7239
R465 VGND.n82 VGND.n67 2.7239
R466 VGND.n50 VGND.n49 2.7239
R467 VGND.n37 VGND.n36 2.7239
R468 VGND.n112 VGND.n111 1.753
R469 VGND.n110 VGND.n109 1.753
R470 VGND VGND.n98 1.48125
R471 VGND.n156 VGND.n155 1.21169
R472 VGND.n98 VGND.n97 1.11894
R473 VGND.n111 VGND 0.95037
R474 VGND.n111 VGND.n110 0.761313
R475 VGND.n155 VGND 0.531208
R476 VGND.n94 VGND.n93 0.467019
R477 VGND.n224 VGND.n223 0.467019
R478 VGND.n103 VGND.n102 0.409011
R479 VGND.n114 VGND.n67 0.409011
R480 VGND.n56 VGND.n45 0.409011
R481 VGND.n168 VGND.n34 0.409011
R482 VGND.n165 VGND.n164 0.409011
R483 VGND.n160 VGND.n37 0.409011
R484 VGND.n97 VGND.n0 0.198729
R485 VGND.n96 VGND.n95 0.194976
R486 VGND.n141 VGND.n60 0.1255
R487 VGND.n79 VGND.n68 0.120292
R488 VGND.n84 VGND.n68 0.120292
R489 VGND.n117 VGND.n116 0.120292
R490 VGND.n118 VGND.n117 0.120292
R491 VGND.n122 VGND.n65 0.120292
R492 VGND.n123 VGND.n122 0.120292
R493 VGND.n134 VGND.n133 0.120292
R494 VGND.n133 VGND.n124 0.120292
R495 VGND.n128 VGND.n125 0.120292
R496 VGND.n128 VGND.n127 0.120292
R497 VGND.n101 VGND.n99 0.120292
R498 VGND.n108 VGND.n100 0.120292
R499 VGND.n77 VGND.n69 0.120292
R500 VGND.n72 VGND.n69 0.120292
R501 VGND.n72 VGND.n71 0.120292
R502 VGND.n162 VGND.n161 0.120292
R503 VGND.n150 VGND.n149 0.120292
R504 VGND.n149 VGND.n42 0.120292
R505 VGND.n145 VGND.n144 0.120292
R506 VGND.n55 VGND.n54 0.120292
R507 VGND.n54 VGND.n46 0.120292
R508 VGND.n48 VGND.n46 0.120292
R509 VGND.n162 VGND 0.0981562
R510 VGND.n78 VGND 0.09425
R511 VGND.n110 VGND 0.0881354
R512 VGND.n95 VGND.n94 0.0766574
R513 VGND.n223 VGND.n0 0.0766574
R514 VGND.n109 VGND.n108 0.0721146
R515 VGND.n156 VGND.n154 0.0708125
R516 VGND.n86 VGND 0.064875
R517 VGND.n90 VGND 0.064875
R518 VGND.n88 VGND 0.064875
R519 VGND.n225 VGND 0.064875
R520 VGND.n222 VGND 0.064875
R521 VGND VGND.n285 0.064875
R522 VGND.n92 VGND 0.063625
R523 VGND.n209 VGND 0.063625
R524 VGND.n112 VGND.n84 0.0616979
R525 VGND.n116 VGND 0.0603958
R526 VGND VGND.n65 0.0603958
R527 VGND.n135 VGND 0.0603958
R528 VGND VGND.n134 0.0603958
R529 VGND.n125 VGND 0.0603958
R530 VGND VGND.n59 0.0603958
R531 VGND.n101 VGND 0.0603958
R532 VGND.n71 VGND 0.0603958
R533 VGND VGND.n166 0.0603958
R534 VGND.n158 VGND 0.0603958
R535 VGND VGND.n157 0.0603958
R536 VGND.n154 VGND 0.0603958
R537 VGND.n151 VGND 0.0603958
R538 VGND VGND.n150 0.0603958
R539 VGND.n145 VGND 0.0603958
R540 VGND.n144 VGND 0.0603958
R541 VGND.n55 VGND 0.0603958
R542 VGND.n113 VGND.n112 0.0590938
R543 VGND VGND.n143 0.0590938
R544 VGND.n157 VGND.n156 0.0499792
R545 VGND.n109 VGND.n99 0.0486771
R546 VGND VGND.n35 0.0460729
R547 VGND.n98 VGND.n96 0.040297
R548 VGND.n167 VGND 0.0343542
R549 VGND.n135 VGND 0.0330521
R550 VGND.n158 VGND 0.0330521
R551 VGND VGND.n60 0.03175
R552 VGND.n113 VGND 0.0226354
R553 VGND.n118 VGND 0.0226354
R554 VGND VGND.n123 0.0226354
R555 VGND VGND.n124 0.0226354
R556 VGND.n127 VGND 0.0226354
R557 VGND.n100 VGND 0.0226354
R558 VGND.n166 VGND 0.0226354
R559 VGND.n161 VGND 0.0226354
R560 VGND.n151 VGND 0.0226354
R561 VGND VGND.n42 0.0226354
R562 VGND.n58 VGND 0.0226354
R563 VGND.n48 VGND 0.0226354
R564 VGND.n167 VGND.n35 0.0148229
R565 VGND.n78 VGND.n77 0.00440625
R566 VGND.n60 VGND.n59 0.00180208
R567 VGND.n143 VGND.n58 0.00180208
R568 select1.n10 select1.t8 327.99
R569 select1.n3 select1.t7 293.969
R570 select1.n6 select1.t4 256.07
R571 select1.n1 select1.t6 212.081
R572 select1.n0 select1.t3 212.081
R573 select1.n10 select1.t0 199.457
R574 select1.n2 select1.n1 182.929
R575 select1 select1.n3 154.065
R576 select1.n11 select1.n10 152
R577 select1.n7 select1.n6 152
R578 select1.n6 select1.t2 150.03
R579 select1.n1 select1.t5 139.78
R580 select1.n0 select1.t1 139.78
R581 select1.n3 select1.t9 138.338
R582 select1.n1 select1.n0 61.346
R583 select1.n5 select1 22.1096
R584 select1.n14 select1.n13 14.6836
R585 select1.n13 select1.n12 14.6704
R586 select1.n12 select1 13.8672
R587 select1.n4 select1 13.8328
R588 select1.n11 select1 12.1605
R589 select1.n14 select1.n2 10.6811
R590 select1.n7 select1.n5 10.4374
R591 select1.n9 select1.n8 8.15359
R592 select1.n2 select1 6.1445
R593 select1.n4 select1 5.16179
R594 select1.n9 select1.n4 4.65206
R595 select1.n8 select1 3.93896
R596 select1 select1.n11 2.34717
R597 select1.n5 select1 2.16665
R598 select1.n8 select1.n7 1.57588
R599 select1.n13 select1.n9 0.79438
R600 select1.n12 select1 0.6405
R601 select1 select1.n14 0.248606
R602 select2.n5 select2.t0 450.938
R603 select2.n5 select2.t2 445.666
R604 select2.n0 select2.t3 377.486
R605 select2.n0 select2.t4 374.202
R606 select2.n2 select2.t1 212.081
R607 select2.n1 select2.t6 212.081
R608 select2.n3 select2.n2 183.441
R609 select2.n2 select2.t7 139.78
R610 select2.n1 select2.t5 139.78
R611 select2.n2 select2.n1 61.346
R612 select2.n8 select2.n7 12.4093
R613 select2 select2.n3 11.4331
R614 select2.n7 select2.n6 9.10647
R615 select2.n7 select2.n4 8.98648
R616 select2.n3 select2 5.6325
R617 select2.n4 select2 5.02323
R618 select2.n6 select2.n5 3.1748
R619 select2.n8 select2.n0 2.10165
R620 select2.n9 select2 1.09425
R621 select2.n4 select2 0.941788
R622 select2.n6 select2 0.063625
R623 select2.n9 select2.n8 0.062375
R624 select2 select2.n9 0.003
R625 Z.n1 Z.t4 23.6581
R626 Z.n7 Z.t3 23.6581
R627 Z.n0 Z.t5 23.3739
R628 Z.n6 Z.t2 23.3739
R629 Z.n1 Z.t1 10.7528
R630 Z.n7 Z.t6 10.7528
R631 Z.n3 Z.t0 10.6417
R632 Z.n9 Z.t7 10.6417
R633 Z.n2 Z.n1 1.30064
R634 Z.n8 Z.n7 1.30064
R635 Z.n11 Z.n10 1.04212
R636 Z Z.n5 0.919875
R637 Z.n5 Z.n4 0.859481
R638 Z.n11 Z 0.754624
R639 Z.n2 Z.n0 0.726502
R640 Z.n8 Z.n6 0.726502
R641 Z.n3 Z.n2 0.512491
R642 Z.n9 Z.n8 0.512491
R643 Z.n4 Z.n3 0.359663
R644 Z.n10 Z.n9 0.359663
R645 Z.n4 Z.n0 0.216071
R646 Z.n10 Z.n6 0.216071
R647 Z Z.n11 0.0100278
R648 Z.n5 Z 0.001125
R649 VPWR.n190 VPWR.n188 8629.41
R650 VPWR.n193 VPWR.n187 8629.41
R651 VPWR.n206 VPWR.n205 8629.41
R652 VPWR.n208 VPWR.n203 8629.41
R653 VPWR.n226 VPWR.n220 8629.41
R654 VPWR.n229 VPWR.n219 8629.41
R655 VPWR.n242 VPWR.n241 8629.41
R656 VPWR.n244 VPWR.n238 8629.41
R657 VPWR.n259 VPWR.n252 8629.41
R658 VPWR.n256 VPWR.n253 8629.41
R659 VPWR.n53 VPWR.n52 8629.41
R660 VPWR.n55 VPWR.n50 8629.41
R661 VPWR.n36 VPWR.n35 8629.41
R662 VPWR.n38 VPWR.n33 8629.41
R663 VPWR.n19 VPWR.n17 8629.41
R664 VPWR.n22 VPWR.n16 8629.41
R665 VPWR.n8 VPWR.n2 8629.41
R666 VPWR.n8 VPWR.n3 8629.41
R667 VPWR.n6 VPWR.n2 8629.41
R668 VPWR.n6 VPWR.n3 8629.41
R669 VPWR.n276 VPWR.n270 8629.41
R670 VPWR.n276 VPWR.n271 8629.41
R671 VPWR.n274 VPWR.n270 8629.41
R672 VPWR.n274 VPWR.n271 8629.41
R673 VPWR.n8 VPWR.t0 2459.29
R674 VPWR.t1 VPWR.n6 2459.29
R675 VPWR.n276 VPWR.t31 2459.29
R676 VPWR.t28 VPWR.n274 2459.29
R677 VPWR.t0 VPWR.n7 2298.92
R678 VPWR.n7 VPWR.t1 2298.92
R679 VPWR.t31 VPWR.n275 2298.92
R680 VPWR.n275 VPWR.t28 2298.92
R681 VPWR.n189 VPWR.n186 920.471
R682 VPWR.n209 VPWR.n202 920.471
R683 VPWR.n225 VPWR.n221 920.471
R684 VPWR.n245 VPWR.n237 920.471
R685 VPWR.n255 VPWR.n254 920.471
R686 VPWR.n56 VPWR.n49 920.471
R687 VPWR.n39 VPWR.n32 920.471
R688 VPWR.n18 VPWR.n15 920.471
R689 VPWR.n5 VPWR.n4 920.471
R690 VPWR.n273 VPWR.n272 920.471
R691 VPWR.n195 VPWR.n186 914.447
R692 VPWR.n210 VPWR.n209 914.447
R693 VPWR.n221 VPWR.n217 914.447
R694 VPWR.n246 VPWR.n245 914.447
R695 VPWR.n254 VPWR.n251 914.447
R696 VPWR.n58 VPWR.n56 914.447
R697 VPWR.n41 VPWR.n39 914.447
R698 VPWR.n24 VPWR.n15 914.447
R699 VPWR.n4 VPWR.n0 914.447
R700 VPWR.n272 VPWR.n268 914.447
R701 VPWR.t70 VPWR.n124 804.731
R702 VPWR.n126 VPWR.t70 751.692
R703 VPWR.n98 VPWR.t17 671.408
R704 VPWR.n87 VPWR.t51 671.408
R705 VPWR VPWR.t69 630.375
R706 VPWR.n157 VPWR.n156 602.456
R707 VPWR.n179 VPWR.n67 602.456
R708 VPWR.n71 VPWR.n70 585
R709 VPWR.n73 VPWR.n72 585
R710 VPWR.n5 VPWR.n1 480.764
R711 VPWR.n273 VPWR.n269 480.764
R712 VPWR.n189 VPWR.n184 480.764
R713 VPWR.n202 VPWR.n200 480.764
R714 VPWR.n225 VPWR.n224 480.764
R715 VPWR.n239 VPWR.n237 480.764
R716 VPWR.n255 VPWR.n250 480.764
R717 VPWR.n49 VPWR.n47 480.764
R718 VPWR.n32 VPWR.n30 480.764
R719 VPWR.n18 VPWR.n14 480.764
R720 VPWR VPWR.t72 458.724
R721 VPWR.t69 VPWR 458.724
R722 VPWR.n119 VPWR.t26 420.25
R723 VPWR.n115 VPWR.t73 388.656
R724 VPWR.n150 VPWR.t74 388.656
R725 VPWR.n128 VPWR.t71 388.656
R726 VPWR.n101 VPWR.t67 388.656
R727 VPWR.n110 VPWR.t68 388.656
R728 VPWR.n75 VPWR.t64 388.656
R729 VPWR.n80 VPWR.t65 388.656
R730 VPWR.n197 VPWR.n184 379.2
R731 VPWR.n212 VPWR.n200 379.2
R732 VPWR.n224 VPWR.n223 379.2
R733 VPWR.n239 VPWR.n236 379.2
R734 VPWR.n263 VPWR.n250 379.2
R735 VPWR.n60 VPWR.n47 379.2
R736 VPWR.n43 VPWR.n30 379.2
R737 VPWR.n26 VPWR.n14 379.2
R738 VPWR.n10 VPWR.n1 379.2
R739 VPWR.n278 VPWR.n269 379.2
R740 VPWR VPWR.t18 369.938
R741 VPWR VPWR.t58 369.938
R742 VPWR.n104 VPWR.n97 322.329
R743 VPWR.n82 VPWR.n78 322.329
R744 VPWR.n161 VPWR.n159 259.697
R745 VPWR.n137 VPWR.t59 255.905
R746 VPWR.n142 VPWR.t19 255.905
R747 VPWR.n118 VPWR.t27 255.905
R748 VPWR.n158 VPWR.t25 255.905
R749 VPWR.n108 VPWR.t49 254.475
R750 VPWR.n133 VPWR.t53 252.95
R751 VPWR.n138 VPWR.t15 252.95
R752 VPWR.n143 VPWR.t30 252.95
R753 VPWR.n178 VPWR.t37 252.95
R754 VPWR.n157 VPWR.t33 251.516
R755 VPWR.n68 VPWR.t76 250.724
R756 VPWR.n66 VPWR.t39 250.724
R757 VPWR.t26 VPWR.t29 248.599
R758 VPWR.t18 VPWR.t14 248.599
R759 VPWR.t58 VPWR.t52 248.599
R760 VPWR.n173 VPWR.t9 248.219
R761 VPWR.n160 VPWR.t24 248.219
R762 VPWR.n119 VPWR 221.964
R763 VPWR.n126 VPWR.t81 215.827
R764 VPWR.n108 VPWR.n107 213.119
R765 VPWR.n148 VPWR.n119 213.119
R766 VPWR.n116 VPWR.t80 210.964
R767 VPWR.n102 VPWR.t82 210.964
R768 VPWR.n77 VPWR.t79 210.964
R769 VPWR.n168 VPWR.n167 209.368
R770 VPWR.t29 VPWR 198.287
R771 VPWR.t14 VPWR 198.287
R772 VPWR.t52 VPWR 198.287
R773 VPWR.n170 VPWR.n169 183.673
R774 VPWR VPWR.t2 182.952
R775 VPWR VPWR.n168 182.952
R776 VPWR.t40 VPWR 182.952
R777 VPWR.n72 VPWR.n71 159.476
R778 VPWR.n159 VPWR.t11 157.014
R779 VPWR.t75 VPWR.t42 154.417
R780 VPWR.t56 VPWR.t10 147.703
R781 VPWR.t61 VPWR.t16 140.989
R782 VPWR.t10 VPWR.t23 140.989
R783 VPWR.t36 VPWR.t38 140.989
R784 VPWR.t8 VPWR.t75 140.989
R785 VPWR.t50 VPWR.t46 140.989
R786 VPWR.n159 VPWR.t45 137.079
R787 VPWR.n107 VPWR 125.883
R788 VPWR.n169 VPWR 125.883
R789 VPWR.n97 VPWR.t62 116.341
R790 VPWR.n78 VPWR.t47 116.341
R791 VPWR.t16 VPWR 112.457
R792 VPWR.t23 VPWR 112.457
R793 VPWR VPWR.t50 112.457
R794 VPWR VPWR.t34 109.1
R795 VPWR.n11 VPWR.n0 105.788
R796 VPWR.n279 VPWR.n268 105.788
R797 VPWR.t66 VPWR.t61 104.064
R798 VPWR.t46 VPWR.t63 104.064
R799 VPWR.t20 VPWR 102.385
R800 VPWR.t48 VPWR 99.0288
R801 VPWR.n156 VPWR.t57 96.1553
R802 VPWR.n67 VPWR.t55 96.1553
R803 VPWR VPWR.t54 92.315
R804 VPWR.n71 VPWR.t43 86.7743
R805 VPWR.n107 VPWR.t48 83.9228
R806 VPWR.n168 VPWR.t44 80.5659
R807 VPWR.t2 VPWR.t66 77.209
R808 VPWR.t63 VPWR.t40 77.209
R809 VPWR.n72 VPWR.t35 66.8398
R810 VPWR.n196 VPWR.n195 66.6358
R811 VPWR.n211 VPWR.n210 66.6358
R812 VPWR.n218 VPWR.n217 66.6358
R813 VPWR.n247 VPWR.n246 66.6358
R814 VPWR.n262 VPWR.n251 66.6358
R815 VPWR.n59 VPWR.n58 66.6358
R816 VPWR.n42 VPWR.n41 66.6358
R817 VPWR.n25 VPWR.n24 66.6358
R818 VPWR.n10 VPWR.n9 63.3551
R819 VPWR.n278 VPWR.n277 63.3551
R820 VPWR.n156 VPWR.t21 63.3219
R821 VPWR.n67 VPWR.t13 63.3219
R822 VPWR VPWR.t56 62.103
R823 VPWR.n190 VPWR.n189 61.6672
R824 VPWR.n194 VPWR.n193 61.6672
R825 VPWR.n206 VPWR.n202 61.6672
R826 VPWR.n203 VPWR.n201 61.6672
R827 VPWR.n226 VPWR.n225 61.6672
R828 VPWR.n230 VPWR.n229 61.6672
R829 VPWR.n242 VPWR.n237 61.6672
R830 VPWR.n238 VPWR.n234 61.6672
R831 VPWR.n260 VPWR.n259 61.6672
R832 VPWR.n256 VPWR.n255 61.6672
R833 VPWR.n53 VPWR.n49 61.6672
R834 VPWR.n50 VPWR.n48 61.6672
R835 VPWR.n36 VPWR.n32 61.6672
R836 VPWR.n33 VPWR.n31 61.6672
R837 VPWR.n19 VPWR.n18 61.6672
R838 VPWR.n23 VPWR.n22 61.6672
R839 VPWR.n6 VPWR.n5 61.6672
R840 VPWR.n9 VPWR.n8 61.6672
R841 VPWR.n274 VPWR.n273 61.6672
R842 VPWR.n277 VPWR.n276 61.6672
R843 VPWR.n191 VPWR.n190 60.9564
R844 VPWR.n193 VPWR.n192 60.9564
R845 VPWR.n207 VPWR.n206 60.9564
R846 VPWR.n204 VPWR.n203 60.9564
R847 VPWR.n227 VPWR.n226 60.9564
R848 VPWR.n229 VPWR.n228 60.9564
R849 VPWR.n243 VPWR.n242 60.9564
R850 VPWR.n240 VPWR.n238 60.9564
R851 VPWR.n259 VPWR.n258 60.9564
R852 VPWR.n257 VPWR.n256 60.9564
R853 VPWR.n54 VPWR.n53 60.9564
R854 VPWR.n51 VPWR.n50 60.9564
R855 VPWR.n37 VPWR.n36 60.9564
R856 VPWR.n34 VPWR.n33 60.9564
R857 VPWR.n20 VPWR.n19 60.9564
R858 VPWR.n22 VPWR.n21 60.9564
R859 VPWR.n211 VPWR.n201 60.6123
R860 VPWR.n230 VPWR.n218 60.6123
R861 VPWR.n59 VPWR.n48 60.6123
R862 VPWR.n42 VPWR.n31 60.6123
R863 VPWR.n196 VPWR.n185 59.4829
R864 VPWR.n262 VPWR.n261 59.4829
R865 VPWR.n248 VPWR.n247 58.7299
R866 VPWR.n25 VPWR.n13 58.7299
R867 VPWR.t42 VPWR 55.3892
R868 VPWR.t12 VPWR 52.0323
R869 VPWR VPWR.t44 45.3185
R870 VPWR VPWR.t32 41.9616
R871 VPWR.n191 VPWR.n187 38.5759
R872 VPWR.n192 VPWR.n188 38.5759
R873 VPWR.n208 VPWR.n207 38.5759
R874 VPWR.n205 VPWR.n204 38.5759
R875 VPWR.n227 VPWR.n219 38.5759
R876 VPWR.n228 VPWR.n220 38.5759
R877 VPWR.n244 VPWR.n243 38.5759
R878 VPWR.n241 VPWR.n240 38.5759
R879 VPWR.n257 VPWR.n252 38.5759
R880 VPWR.n258 VPWR.n253 38.5759
R881 VPWR.n55 VPWR.n54 38.5759
R882 VPWR.n52 VPWR.n51 38.5759
R883 VPWR.n38 VPWR.n37 38.5759
R884 VPWR.n35 VPWR.n34 38.5759
R885 VPWR.n20 VPWR.n16 38.5759
R886 VPWR.n21 VPWR.n17 38.5759
R887 VPWR.n167 VPWR.n89 34.6358
R888 VPWR.n167 VPWR.n90 34.6358
R889 VPWR.n172 VPWR.n171 34.6358
R890 VPWR.n169 VPWR 28.5341
R891 VPWR.n97 VPWR.t3 28.4453
R892 VPWR.n78 VPWR.t41 28.4453
R893 VPWR.n174 VPWR.n173 28.3534
R894 VPWR.n171 VPWR.n170 25.6953
R895 VPWR.n137 VPWR.n122 25.224
R896 VPWR.n133 VPWR.n122 25.224
R897 VPWR.n142 VPWR.n121 25.224
R898 VPWR.n138 VPWR.n121 25.224
R899 VPWR.n144 VPWR.n118 25.224
R900 VPWR.n144 VPWR.n143 25.224
R901 VPWR.n162 VPWR.n158 25.224
R902 VPWR.n108 VPWR.n92 23.7181
R903 VPWR VPWR.n98 23.252
R904 VPWR.n157 VPWR.n92 21.4593
R905 VPWR.n138 VPWR.n137 20.3299
R906 VPWR.n143 VPWR.n142 20.3299
R907 VPWR.t54 VPWR.t36 20.1418
R908 VPWR.n179 VPWR.n66 19.9534
R909 VPWR.n178 VPWR.n177 19.8181
R910 VPWR.n148 VPWR.n118 17.3181
R911 VPWR.n161 VPWR.n160 17.3181
R912 VPWR.n158 VPWR.n157 16.5652
R913 VPWR.n162 VPWR.n161 16.5652
R914 VPWR.n133 VPWR.n132 15.8123
R915 VPWR.n149 VPWR.n148 14.2735
R916 VPWR.n109 VPWR.n108 14.2735
R917 VPWR.n171 VPWR.n87 13.9299
R918 VPWR.n179 VPWR.n178 13.5534
R919 VPWR.n114 VPWR.n113 11.4366
R920 VPWR.n198 VPWR.n197 11.3235
R921 VPWR.n213 VPWR.n212 11.3235
R922 VPWR.n223 VPWR.n222 11.3235
R923 VPWR.n236 VPWR.n235 11.3235
R924 VPWR.n264 VPWR.n263 11.3235
R925 VPWR.n61 VPWR.n60 11.3235
R926 VPWR.n44 VPWR.n43 11.3235
R927 VPWR.n27 VPWR.n26 11.3235
R928 VPWR.n170 VPWR.n88 11.2937
R929 VPWR.n154 VPWR.n153 11.2737
R930 VPWR.t32 VPWR.t20 10.0712
R931 VPWR.n128 VPWR.n125 9.60526
R932 VPWR.n115 VPWR.n114 9.60526
R933 VPWR.n80 VPWR.n79 9.60526
R934 VPWR.n117 VPWR.n93 9.3005
R935 VPWR.n152 VPWR.n151 9.3005
R936 VPWR.n149 VPWR.n94 9.3005
R937 VPWR.n148 VPWR.n147 9.3005
R938 VPWR.n143 VPWR.n120 9.3005
R939 VPWR.n139 VPWR.n138 9.3005
R940 VPWR.n134 VPWR.n133 9.3005
R941 VPWR.n130 VPWR.n129 9.3005
R942 VPWR.n135 VPWR.n122 9.3005
R943 VPWR.n137 VPWR.n136 9.3005
R944 VPWR.n140 VPWR.n121 9.3005
R945 VPWR.n142 VPWR.n141 9.3005
R946 VPWR.n145 VPWR.n144 9.3005
R947 VPWR.n146 VPWR.n118 9.3005
R948 VPWR.n175 VPWR.n174 9.3005
R949 VPWR.n180 VPWR.n179 9.3005
R950 VPWR.n164 VPWR.n89 9.3005
R951 VPWR.n157 VPWR.n155 9.3005
R952 VPWR.n108 VPWR.n106 9.3005
R953 VPWR.n100 VPWR.n99 9.3005
R954 VPWR.n103 VPWR.n95 9.3005
R955 VPWR.n112 VPWR.n111 9.3005
R956 VPWR.n109 VPWR.n96 9.3005
R957 VPWR.n105 VPWR.n92 9.3005
R958 VPWR.n158 VPWR.n91 9.3005
R959 VPWR.n163 VPWR.n162 9.3005
R960 VPWR.n167 VPWR.n166 9.3005
R961 VPWR.n165 VPWR.n90 9.3005
R962 VPWR.n178 VPWR.n65 9.3005
R963 VPWR.n177 VPWR.n176 9.3005
R964 VPWR.n172 VPWR.n69 9.3005
R965 VPWR.n171 VPWR.n74 9.3005
R966 VPWR.n86 VPWR.n85 9.3005
R967 VPWR.n84 VPWR.n83 9.3005
R968 VPWR.n81 VPWR.n76 9.3005
R969 VPWR.n28 VPWR.n13 8.23557
R970 VPWR.n12 VPWR.n11 7.54844
R971 VPWR.n280 VPWR.n279 7.54407
R972 VPWR.n185 VPWR.n183 6.88686
R973 VPWR.n73 VPWR.n70 6.8005
R974 VPWR.n132 VPWR.n124 6.48583
R975 VPWR.n195 VPWR.n194 6.02403
R976 VPWR.n246 VPWR.n234 6.02403
R977 VPWR.n260 VPWR.n251 6.02403
R978 VPWR.n24 VPWR.n23 6.02403
R979 VPWR.n9 VPWR.n0 6.02403
R980 VPWR.n277 VPWR.n268 6.02403
R981 VPWR.n127 VPWR.n126 5.8885
R982 VPWR.n11 VPWR.n10 5.18145
R983 VPWR.n279 VPWR.n278 5.18145
R984 VPWR.n201 VPWR.n64 4.89462
R985 VPWR.n231 VPWR.n217 4.89462
R986 VPWR.n57 VPWR.n48 4.89462
R987 VPWR.n41 VPWR.n40 4.89462
R988 VPWR.n151 VPWR.n117 4.67352
R989 VPWR.n132 VPWR.n131 4.62124
R990 VPWR.n129 VPWR.n128 4.36875
R991 VPWR.n151 VPWR.n150 4.36875
R992 VPWR.n111 VPWR.n110 4.36875
R993 VPWR.n81 VPWR.n80 4.36875
R994 VPWR.t38 VPWR.t12 3.35739
R995 VPWR.t34 VPWR.t8 3.35739
R996 VPWR.n183 VPWR 3.29986
R997 VPWR.n215 VPWR.n64 3.25464
R998 VPWR.n249 VPWR.n248 3.24308
R999 VPWR.n57 VPWR.n46 3.23917
R1000 VPWR.n232 VPWR.n231 3.23136
R1001 VPWR.n40 VPWR.n29 3.23136
R1002 VPWR.n261 VPWR.n63 3.22655
R1003 VPWR.n129 VPWR.n127 3.2005
R1004 VPWR.n187 VPWR.n186 2.84665
R1005 VPWR.n188 VPWR.n184 2.84665
R1006 VPWR.n209 VPWR.n208 2.84665
R1007 VPWR.n205 VPWR.n200 2.84665
R1008 VPWR.n221 VPWR.n219 2.84665
R1009 VPWR.n224 VPWR.n220 2.84665
R1010 VPWR.n245 VPWR.n244 2.84665
R1011 VPWR.n241 VPWR.n239 2.84665
R1012 VPWR.n254 VPWR.n252 2.84665
R1013 VPWR.n253 VPWR.n250 2.84665
R1014 VPWR.n56 VPWR.n55 2.84665
R1015 VPWR.n52 VPWR.n47 2.84665
R1016 VPWR.n39 VPWR.n38 2.84665
R1017 VPWR.n35 VPWR.n30 2.84665
R1018 VPWR.n16 VPWR.n15 2.84665
R1019 VPWR.n17 VPWR.n14 2.84665
R1020 VPWR.n3 VPWR.n1 2.84665
R1021 VPWR.n7 VPWR.n3 2.84665
R1022 VPWR.n4 VPWR.n2 2.84665
R1023 VPWR.n7 VPWR.n2 2.84665
R1024 VPWR.n271 VPWR.n269 2.84665
R1025 VPWR.n275 VPWR.n271 2.84665
R1026 VPWR.n272 VPWR.n270 2.84665
R1027 VPWR.n275 VPWR.n270 2.84665
R1028 VPWR.n127 VPWR.n124 2.8165
R1029 VPWR.n104 VPWR.n103 2.54018
R1030 VPWR.n83 VPWR.n82 2.54018
R1031 VPWR.n117 VPWR.n116 2.33701
R1032 VPWR.n103 VPWR.n102 2.33701
R1033 VPWR.n83 VPWR.n77 2.33701
R1034 VPWR.n197 VPWR.n196 2.28169
R1035 VPWR.n212 VPWR.n211 2.28169
R1036 VPWR.n223 VPWR.n218 2.28169
R1037 VPWR.n247 VPWR.n236 2.28169
R1038 VPWR.n263 VPWR.n262 2.28169
R1039 VPWR.n60 VPWR.n59 2.28169
R1040 VPWR.n43 VPWR.n42 2.28169
R1041 VPWR.n26 VPWR.n25 2.28169
R1042 VPWR.n233 VPWR.n232 2.13544
R1043 VPWR.n111 VPWR.n104 2.13383
R1044 VPWR.n82 VPWR.n81 2.13383
R1045 VPWR.n267 VPWR.n12 2.06883
R1046 VPWR.n116 VPWR.n115 2.03225
R1047 VPWR.n102 VPWR.n101 2.03225
R1048 VPWR.n77 VPWR.n75 2.03225
R1049 VPWR.n249 VPWR.n233 1.95379
R1050 VPWR.n248 VPWR.n234 1.88285
R1051 VPWR.n23 VPWR.n13 1.88285
R1052 VPWR.n182 VPWR.n181 1.753
R1053 VPWR VPWR.n182 1.64258
R1054 VPWR.n90 VPWR.n66 1.50638
R1055 VPWR.n174 VPWR.n73 1.4005
R1056 VPWR.n100 VPWR.n98 1.37193
R1057 VPWR.n87 VPWR.n86 1.37193
R1058 VPWR.n280 VPWR.n267 1.33758
R1059 VPWR.n214 VPWR.n213 1.143
R1060 VPWR.n222 VPWR.n216 1.143
R1061 VPWR.n62 VPWR.n61 1.143
R1062 VPWR.n45 VPWR.n44 1.143
R1063 VPWR.n199 VPWR.n198 1.13925
R1064 VPWR.n265 VPWR.n264 1.13925
R1065 VPWR.n235 VPWR.n233 1.13675
R1066 VPWR.n28 VPWR.n27 1.13675
R1067 VPWR.n194 VPWR.n185 1.12991
R1068 VPWR.n210 VPWR.n64 1.12991
R1069 VPWR.n231 VPWR.n230 1.12991
R1070 VPWR.n261 VPWR.n260 1.12991
R1071 VPWR.n58 VPWR.n57 1.12991
R1072 VPWR.n40 VPWR.n31 1.12991
R1073 VPWR.n123 VPWR 1.06099
R1074 VPWR.n46 VPWR.n45 0.862816
R1075 VPWR.n214 VPWR.n199 0.854667
R1076 VPWR.n29 VPWR.n28 0.770881
R1077 VPWR.n160 VPWR.n89 0.753441
R1078 VPWR.n173 VPWR.n172 0.753441
R1079 VPWR.n63 VPWR.n62 0.747859
R1080 VPWR.n267 VPWR.n266 0.704667
R1081 VPWR.n70 VPWR.n68 0.6005
R1082 VPWR.n216 VPWR.n215 0.588641
R1083 VPWR.n265 VPWR.n249 0.518882
R1084 VPWR.n182 VPWR 0.460219
R1085 VPWR.n177 VPWR.n68 0.4005
R1086 VPWR.n45 VPWR.n29 0.392323
R1087 VPWR.n62 VPWR.n46 0.360318
R1088 VPWR.n150 VPWR.n149 0.305262
R1089 VPWR.n101 VPWR.n100 0.305262
R1090 VPWR.n110 VPWR.n109 0.305262
R1091 VPWR.n86 VPWR.n75 0.305262
R1092 VPWR.t60 VPWR.n191 0.27666
R1093 VPWR.n192 VPWR.t60 0.27666
R1094 VPWR.n207 VPWR.t5 0.27666
R1095 VPWR.n204 VPWR.t5 0.27666
R1096 VPWR.t78 VPWR.n227 0.27666
R1097 VPWR.n228 VPWR.t78 0.27666
R1098 VPWR.n243 VPWR.t22 0.27666
R1099 VPWR.n240 VPWR.t22 0.27666
R1100 VPWR.t4 VPWR.n257 0.27666
R1101 VPWR.n258 VPWR.t4 0.27666
R1102 VPWR.n54 VPWR.t6 0.27666
R1103 VPWR.n51 VPWR.t6 0.27666
R1104 VPWR.n37 VPWR.t77 0.27666
R1105 VPWR.n34 VPWR.t77 0.27666
R1106 VPWR.t7 VPWR.n20 0.27666
R1107 VPWR.n21 VPWR.t7 0.27666
R1108 VPWR.n215 VPWR.n214 0.268128
R1109 VPWR.n232 VPWR.n216 0.223986
R1110 VPWR.n199 VPWR.n183 0.202423
R1111 VPWR.n131 VPWR.n130 0.180304
R1112 VPWR.n131 VPWR 0.120408
R1113 VPWR.n114 VPWR.n93 0.120292
R1114 VPWR.n152 VPWR.n94 0.120292
R1115 VPWR.n146 VPWR.n145 0.120292
R1116 VPWR.n145 VPWR.n120 0.120292
R1117 VPWR.n141 VPWR.n140 0.120292
R1118 VPWR.n140 VPWR.n139 0.120292
R1119 VPWR.n136 VPWR.n135 0.120292
R1120 VPWR.n135 VPWR.n134 0.120292
R1121 VPWR.n130 VPWR.n125 0.120292
R1122 VPWR.n99 VPWR.n95 0.120292
R1123 VPWR.n112 VPWR.n96 0.120292
R1124 VPWR.n163 VPWR.n91 0.120292
R1125 VPWR.n164 VPWR.n163 0.120292
R1126 VPWR.n180 VPWR.n65 0.120292
R1127 VPWR.n176 VPWR.n175 0.120292
R1128 VPWR.n175 VPWR.n69 0.120292
R1129 VPWR.n85 VPWR.n84 0.120292
R1130 VPWR.n84 VPWR.n76 0.120292
R1131 VPWR.n79 VPWR.n76 0.120292
R1132 VPWR.n153 VPWR.n93 0.11899
R1133 VPWR.n266 VPWR.n63 0.1125
R1134 VPWR.n99 VPWR 0.0981562
R1135 VPWR.n154 VPWR 0.0955521
R1136 VPWR.n113 VPWR.n95 0.0916458
R1137 VPWR.n198 VPWR 0.06425
R1138 VPWR.n213 VPWR 0.06425
R1139 VPWR.n222 VPWR 0.06425
R1140 VPWR.n235 VPWR 0.06425
R1141 VPWR.n264 VPWR 0.06425
R1142 VPWR.n61 VPWR 0.06425
R1143 VPWR.n44 VPWR 0.06425
R1144 VPWR.n27 VPWR 0.06425
R1145 VPWR VPWR.n280 0.06425
R1146 VPWR.n147 VPWR 0.0603958
R1147 VPWR VPWR.n146 0.0603958
R1148 VPWR.n141 VPWR 0.0603958
R1149 VPWR.n136 VPWR 0.0603958
R1150 VPWR.n106 VPWR 0.0603958
R1151 VPWR VPWR.n105 0.0603958
R1152 VPWR VPWR.n91 0.0603958
R1153 VPWR.n166 VPWR 0.0603958
R1154 VPWR VPWR.n165 0.0603958
R1155 VPWR.n176 VPWR 0.0603958
R1156 VPWR.n85 VPWR 0.0603958
R1157 VPWR.n12 VPWR 0.059875
R1158 VPWR.n88 VPWR 0.0590938
R1159 VPWR.n266 VPWR.n265 0.054
R1160 VPWR.n181 VPWR 0.0525833
R1161 VPWR.n181 VPWR.n180 0.0460729
R1162 VPWR.n106 VPWR 0.0382604
R1163 VPWR VPWR.n123 0.0369583
R1164 VPWR.n147 VPWR 0.03175
R1165 VPWR.n166 VPWR 0.03175
R1166 VPWR.n113 VPWR.n112 0.0291458
R1167 VPWR VPWR.n94 0.0226354
R1168 VPWR VPWR.n120 0.0226354
R1169 VPWR.n139 VPWR 0.0226354
R1170 VPWR.n134 VPWR 0.0226354
R1171 VPWR.n125 VPWR 0.0226354
R1172 VPWR VPWR.n96 0.0226354
R1173 VPWR.n105 VPWR 0.0226354
R1174 VPWR.n155 VPWR 0.0226354
R1175 VPWR VPWR.n164 0.0226354
R1176 VPWR.n165 VPWR 0.0226354
R1177 VPWR VPWR.n65 0.0226354
R1178 VPWR VPWR.n69 0.0226354
R1179 VPWR VPWR.n74 0.0226354
R1180 VPWR.n79 VPWR 0.0226354
R1181 VPWR.n155 VPWR.n154 0.00310417
R1182 VPWR.n153 VPWR.n152 0.00180208
R1183 VPWR.n123 VPWR 0.00180208
R1184 VPWR.n88 VPWR.n74 0.00180208
R1185 x1.gno0.n2 x1.gno0.t9 377.486
R1186 x1.gno0.n3 x1.gno0.t2 377.486
R1187 x1.gno0.n2 x1.gno0.t7 374.202
R1188 x1.gno0.n3 x1.gno0.t3 374.202
R1189 x1.gno0.n10 x1.gno0.t0 339.418
R1190 x1.gno0.n1 x1.gno0.t1 274.06
R1191 x1.gno0.n7 x1.gno0.t8 212.081
R1192 x1.gno0.n6 x1.gno0.t6 212.081
R1193 x1.gno0.n8 x1.gno0.n7 182.673
R1194 x1.gno0.n7 x1.gno0.t5 139.78
R1195 x1.gno0.n6 x1.gno0.t4 139.78
R1196 x1.gno0.n7 x1.gno0.n6 61.346
R1197 x1.gno0.n5 x1.gno0.n8 15.8606
R1198 x1.gno0 x1.gno0.n9 13.8044
R1199 x1.gno0.n0 x1.gno0.n4 13.4101
R1200 x1.gno0.n0 x1.gno0 11.5859
R1201 x1.gno0.n4 x1.gno0 11.5859
R1202 x1.gno0 x1.gno0.n1 11.0989
R1203 x1.gno0.n9 x1.gno0.n5 6.94768
R1204 x1.gno0 x1.gno0.n0 6.73859
R1205 x1.gno0.n11 x1.gno0 6.6565
R1206 x1.gno0.n8 x1.gno0 6.4005
R1207 x1.gno0.n1 x1.gno0 6.1445
R1208 x1.gno0.n0 x1.gno0 5.13959
R1209 x1.gno0.n4 x1.gno0 4.55738
R1210 x1.gno0.n11 x1.gno0.n10 4.0914
R1211 x1.gno0 x1.gno0.n11 3.61789
R1212 x1.gno0.n9 x1.gno0 3.26325
R1213 x1.gno0.n1 x1.gno0 2.86947
R1214 x1.gno0 x1.gno0.n2 2.04102
R1215 x1.gno0 x1.gno0.n3 2.04102
R1216 x1.gno0.n10 x1.gno0 1.74382
R1217 x1.gno0.n5 x1.gno0 1.47326
R1218 A5.n1 A5.t0 26.3998
R1219 A5.n1 A5.t1 23.5483
R1220 A5.n0 A5.t3 12.7127
R1221 A5.n0 A5.t2 10.8578
R1222 A5.n2 A5.n1 3.12177
R1223 A5.n2 A5.n0 1.81453
R1224 A5.n3 A5.n2 1.1255
R1225 A5.n3 A5 0.21549
R1226 A5 A5.n3 0.0655
R1227 x1.gno3.n3 x1.gno3.t3 377.486
R1228 x1.gno3.n1 x1.gno3.t6 377.486
R1229 x1.gno3.n3 x1.gno3.t5 374.202
R1230 x1.gno3.n1 x1.gno3.t9 374.202
R1231 x1.gno3.n9 x1.gno3.t0 339.418
R1232 x1.gno3.n0 x1.gno3.t1 274.06
R1233 x1.gno3.n6 x1.gno3.t4 212.081
R1234 x1.gno3.n5 x1.gno3.t8 212.081
R1235 x1.gno3.n7 x1.gno3.n6 184.977
R1236 x1.gno3.n6 x1.gno3.t2 139.78
R1237 x1.gno3.n5 x1.gno3.t7 139.78
R1238 x1.gno3.n6 x1.gno3.n5 61.346
R1239 x1.gno3.n8 x1.gno3 18.2601
R1240 x1.gno3 x1.gno3.n7 13.8193
R1241 x1.gno3 x1.gno3.n4 11.7568
R1242 x1.gno3.n4 x1.gno3.n2 11.6628
R1243 x1.gno3 x1.gno3.n0 11.2645
R1244 x1.gno3 x1.gno3.n8 8.9605
R1245 x1.gno3.n8 x1.gno3 8.4485
R1246 x1.gno3.n2 x1.gno3 8.16743
R1247 x1.gno3.n10 x1.gno3 6.6565
R1248 x1.gno3.n0 x1.gno3 6.1445
R1249 x1.gno3.n4 x1.gno3 5.8185
R1250 x1.gno3.n2 x1.gno3 4.58237
R1251 x1.gno3.n7 x1.gno3 4.0965
R1252 x1.gno3.n10 x1.gno3.n9 4.0914
R1253 x1.gno3 x1.gno3.n10 3.61789
R1254 x1.gno3.n0 x1.gno3 2.86947
R1255 x1.gno3 x1.gno3.n3 2.04102
R1256 x1.gno3 x1.gno3.n1 2.04102
R1257 x1.gno3.n9 x1.gno3 1.74382
R1258 x1.gpo3.n3 x1.gpo3.t7 450.938
R1259 x1.gpo3.n2 x1.gpo3.t4 450.938
R1260 x1.gpo3.n3 x1.gpo3.t5 445.666
R1261 x1.gpo3.n2 x1.gpo3.t6 445.666
R1262 x1.gpo3 x1.gpo3.n7 203.923
R1263 x1.gpo3.n1 x1.gpo3.n0 101.49
R1264 x1.gpo3.n7 x1.gpo3.t0 26.5955
R1265 x1.gpo3.n7 x1.gpo3.t1 26.5955
R1266 x1.gpo3.n0 x1.gpo3.t2 24.9236
R1267 x1.gpo3.n0 x1.gpo3.t3 24.9236
R1268 x1.gpo3.n4 x1.gpo3 11.0619
R1269 x1.gpo3.n6 x1.gpo3 10.7525
R1270 x1.gpo3 x1.gpo3.n4 9.34192
R1271 x1.gpo3.n5 x1.gpo3 7.73829
R1272 x1.gpo3.n6 x1.gpo3 6.6565
R1273 x1.gpo3.n4 x1.gpo3 5.84951
R1274 x1.gpo3 x1.gpo3.n6 5.04292
R1275 x1.gpo3 x1.gpo3.n3 2.95993
R1276 x1.gpo3 x1.gpo3.n2 2.95993
R1277 x1.gpo3.n1 x1.gpo3 1.93989
R1278 x1.gpo3 x1.gpo3.n5 1.5365
R1279 x1.gpo3.n5 x1.gpo3.n1 1.0245
R1280 select0.n5 select0.t3 327.99
R1281 select0.n9 select0.t2 293.969
R1282 select0.n3 select0.t6 261.887
R1283 select0.n1 select0.t1 212.081
R1284 select0.n0 select0.t0 212.081
R1285 select0.n5 select0.t5 199.457
R1286 select0.n2 select0.n1 183.185
R1287 select0.n3 select0.t4 155.847
R1288 select0 select0.n9 154.065
R1289 select0.n6 select0.n5 152
R1290 select0.n4 select0.n3 152
R1291 select0.n1 select0.t9 139.78
R1292 select0.n0 select0.t8 139.78
R1293 select0.n9 select0.t7 138.338
R1294 select0.n1 select0.n0 61.346
R1295 select0.n10 select0 13.4199
R1296 select0.n8 select0.n4 11.9062
R1297 select0.n11 select0.n8 11.7395
R1298 select0.n12 select0.n11 11.5949
R1299 select0.n12 select0.n2 9.68118
R1300 select0.n7 select0 9.17383
R1301 select0.n2 select0 5.8885
R1302 select0.n10 select0 5.57469
R1303 select0.n8 select0.n7 4.6505
R1304 select0.n11 select0.n10 4.6505
R1305 select0.n7 select0.n6 2.98717
R1306 select0.n6 select0 2.34717
R1307 select0.n4 select0 2.07109
R1308 select0 select0.n12 0.559212
R1309 x1.gpo0.n4 x1.gpo0.t5 450.938
R1310 x1.gpo0.n3 x1.gpo0.t7 450.938
R1311 x1.gpo0.n4 x1.gpo0.t4 445.666
R1312 x1.gpo0.n3 x1.gpo0.t6 445.666
R1313 x1.gpo0.n7 x1.gpo0.n6 195.832
R1314 x1.gpo0.n1 x1.gpo0.n0 101.49
R1315 x1.gpo0.n6 x1.gpo0.t1 26.5955
R1316 x1.gpo0.n6 x1.gpo0.t0 26.5955
R1317 x1.gpo0.n0 x1.gpo0.t3 24.9236
R1318 x1.gpo0.n0 x1.gpo0.t2 24.9236
R1319 x1.gpo0.n5 x1.gpo0 13.3282
R1320 x1.gpo0.n7 x1.gpo0 11.8923
R1321 x1.gpo0.n2 x1.gpo0 10.7525
R1322 x1.gpo0 x1.gpo0.n7 8.09215
R1323 x1.gpo0.n2 x1.gpo0 6.6565
R1324 x1.gpo0 x1.gpo0.n5 5.46644
R1325 x1.gpo0.n5 x1.gpo0 5.31412
R1326 x1.gpo0 x1.gpo0.n2 5.04292
R1327 x1.gpo0 x1.gpo0.n4 3.18415
R1328 x1.gpo0 x1.gpo0.n3 2.90754
R1329 x1.gpo0 x1.gpo0.n1 2.5605
R1330 x1.gpo0.n1 x1.gpo0 1.93989
R1331 A1.n1 A1.t0 26.3998
R1332 A1.n1 A1.t1 23.5483
R1333 A1.n0 A1.t2 12.7127
R1334 A1.n0 A1.t3 10.8578
R1335 A1.n2 A1.n1 3.12177
R1336 A1.n2 A1.n0 1.81453
R1337 A1.n3 A1.n2 1.1255
R1338 A1.n3 A1 0.21549
R1339 A1 A1.n3 0.0655
R1340 A2.n1 A2.t0 26.3998
R1341 A2.n1 A2.t3 23.5483
R1342 A2.n0 A2.t1 12.7127
R1343 A2.n0 A2.t2 10.8578
R1344 A2.n2 A2.n1 3.12177
R1345 A2.n2 A2.n0 1.81453
R1346 A2.n3 A2.n2 1.1255
R1347 A2.n3 A2 0.219402
R1348 A2 A2.n3 0.0655
R1349 A4.n1 A4.t2 26.3998
R1350 A4.n1 A4.t3 23.5483
R1351 A4.n0 A4.t1 12.7127
R1352 A4.n0 A4.t0 10.8578
R1353 A4.n2 A4.n1 3.12177
R1354 A4.n2 A4.n0 1.81453
R1355 A4.n3 A4.n2 1.1255
R1356 A4 A4.n3 0.203263
R1357 A4.n3 A4 0.0655
R1358 A7.n1 A7.t2 26.3998
R1359 A7.n1 A7.t3 23.5483
R1360 A7.n0 A7.t1 12.7127
R1361 A7.n0 A7.t0 10.8578
R1362 A7.n2 A7.n1 3.12177
R1363 A7.n2 A7.n0 1.81453
R1364 A7.n3 A7.n2 1.1255
R1365 A7.n3 A7 0.210543
R1366 A7 A7.n3 0.0655
R1367 A3.n1 A3.t3 26.3998
R1368 A3.n1 A3.t2 23.5483
R1369 A3.n0 A3.t1 12.7127
R1370 A3.n0 A3.t0 10.8578
R1371 A3.n2 A3.n1 3.12177
R1372 A3.n2 A3.n0 1.81453
R1373 A3.n3 A3.n2 1.1255
R1374 A3.n3 A3 0.210543
R1375 A3 A3.n3 0.0655
R1376 A6.n1 A6.t0 26.3998
R1377 A6.n1 A6.t1 23.5483
R1378 A6.n0 A6.t3 12.7127
R1379 A6.n0 A6.t2 10.8578
R1380 A6.n2 A6.n1 3.12177
R1381 A6.n2 A6.n0 1.81453
R1382 A6.n3 A6.n2 1.1255
R1383 A6.n3 A6 0.219402
R1384 A6 A6.n3 0.0655
R1385 A8.n1 A8.t3 26.3998
R1386 A8.n1 A8.t2 23.5483
R1387 A8.n0 A8.t1 12.7127
R1388 A8.n0 A8.t0 10.8578
R1389 A8.n2 A8.n1 3.12177
R1390 A8.n2 A8.n0 1.81453
R1391 A8.n3 A8.n2 1.1255
R1392 A8 A8.n3 0.203263
R1393 A8.n3 A8 0.0655
R1394 x1.gpo1.n4 x1.gpo1.t6 450.938
R1395 x1.gpo1.n3 x1.gpo1.t7 450.938
R1396 x1.gpo1.n4 x1.gpo1.t4 445.666
R1397 x1.gpo1.n3 x1.gpo1.t5 445.666
R1398 x1.gpo1.n7 x1.gpo1.n6 195.958
R1399 x1.gpo1.n1 x1.gpo1.n0 101.49
R1400 x1.gpo1.n6 x1.gpo1.t1 26.5955
R1401 x1.gpo1.n6 x1.gpo1.t0 26.5955
R1402 x1.gpo1.n0 x1.gpo1.t3 24.9236
R1403 x1.gpo1.n0 x1.gpo1.t2 24.9236
R1404 x1.gpo1.n5 x1.gpo1 14.964
R1405 x1.gpo1.n7 x1.gpo1 11.8408
R1406 x1.gpo1.n2 x1.gpo1 10.7525
R1407 x1.gpo1 x1.gpo1.n5 8.86265
R1408 x1.gpo1 x1.gpo1.n7 7.96524
R1409 x1.gpo1.n2 x1.gpo1 6.6565
R1410 x1.gpo1.n5 x1.gpo1 5.75481
R1411 x1.gpo1 x1.gpo1.n2 5.04292
R1412 x1.gpo1 x1.gpo1.n4 2.94361
R1413 x1.gpo1 x1.gpo1.n3 2.94361
R1414 x1.gpo1 x1.gpo1.n1 2.5605
R1415 x1.gpo1.n1 x1.gpo1 1.93989
C0 x1.gno1 x1.gno2 0.179257f
C1 x1.gno2 x1.gpo2 5.02054f
C2 x1.gno1 x1.gpo2 0.060968f
C3 A8 A7 2.08862f
C4 A8 A6 2.39e-19
C5 A6 A7 1.81997f
C6 A6 A4 7.47e-20
C7 A5 A6 1.81909f
C8 select2 Z 0.799881f
C9 A5 A4 1.27332f
C10 A3 A4 2.08862f
C11 VPWR Z 5.306779f
C12 A2 A4 2.39e-19
C13 A8 VPWR 1.54289f
C14 A3 A2 1.81997f
C15 select2 A4 6.76e-20
C16 A5 select2 2.94e-19
C17 VPWR A7 1.61205f
C18 x3.Z3 Z 5.48465f
C19 select2 A3 2.39e-19
C20 A6 VPWR 1.60651f
C21 x5.A Z 4.51604f
C22 A2 A1 1.81909f
C23 A8 x3.Z3 4.51511f
C24 A5 VPWR 1.60179f
C25 A4 VPWR 1.56602f
C26 select2 A1 0.054741f
C27 A3 VPWR 1.61205f
C28 select0 A1 2.25e-21
C29 x3.Z3 A7 4.5214f
C30 A6 x3.Z3 4.52053f
C31 select2 select0 0.446748f
C32 A2 VPWR 1.60691f
C33 x1.gpo0 Z 2.38e-19
C34 A5 x3.Z3 4.52088f
C35 A4 x3.Z3 0.003925f
C36 select1 A1 4.98e-22
C37 x5.A A5 4.07e-21
C38 VPWR A1 1.6325f
C39 x5.A A4 4.5151f
C40 select1 select2 0.289185f
C41 select1 select0 1.85585f
C42 A3 x3.Z3 1.64e-20
C43 select2 VPWR 3.46438f
C44 x5.A A3 4.5214f
C45 x1.gno0 Z 4.27e-20
C46 select0 VPWR 1.13942f
C47 x5.A A2 4.52052f
C48 x1.gpo0 A7 2.46e-21
C49 A6 x1.gpo0 0.12311f
C50 select1 VPWR 2.65613f
C51 x5.A A1 4.52065f
C52 x1.gpo1 Z 2.41e-19
C53 m2_5776_5494# select0 0.130999f
C54 m2_5776_5494# select2 4.4e-19
C55 A8 x1.gpo1 2.07e-19
C56 x1.gpo0 A4 0.002819f
C57 A5 x1.gpo0 4.0165f
C58 select2 x3.Z3 5.00334f
C59 x5.A select2 5.67997f
C60 x1.nSEL2 Z 0.833318f
C61 x1.gno0 A6 3.66e-20
C62 a_5699_5631# select0 9.55e-19
C63 A3 x1.gpo0 0.001407f
C64 m2_5776_5494# select1 0.183786f
C65 x1.gno0 A4 0.218459f
C66 x1.gno0 A5 3.85224f
C67 x1.gpo1 A7 0.145249f
C68 m2_5776_5494# VPWR 0.139797f
C69 A2 x1.gpo0 0.124367f
C70 x3.Z3 VPWR 14.4075f
C71 select2 x1.nSEL0 0.131256f
C72 a_5645_5493# select2 4.33e-19
C73 x5.A VPWR 14.1327f
C74 A6 x1.gpo1 4.01113f
C75 x1.nSEL0 select0 0.325123f
C76 a_5645_5493# select0 0.048888f
C77 x1.gno0 A3 0.131584f
C78 A5 x1.gpo1 0.001763f
C79 x1.gpo0 A1 3.9665f
C80 a_5699_5631# VPWR 9.09e-19
C81 x1.gpo1 A4 4.15e-19
C82 x1.gno0 A2 0.135398f
C83 select2 x1.gpo0 5.94e-19
C84 select0 x1.gpo0 8.18e-19
C85 x1.gpo3 Z 1.68e-19
C86 select1 x1.nSEL0 0.137595f
C87 a_5645_5493# select1 0.02803f
C88 A3 x1.gpo1 0.1453f
C89 a_5645_5493# VPWR 0.21052f
C90 x1.nSEL0 VPWR 0.386805f
C91 A8 x1.gpo3 4.00906f
C92 x5.A x3.Z3 2.05508f
C93 x1.gno0 A1 4.31208f
C94 x1.gno0 select2 0.054258f
C95 A2 x1.gpo1 3.95776f
C96 x1.gno0 select0 0.020289f
C97 select1 x1.gpo0 8.43e-19
C98 x1.nSEL2 A3 7.03e-21
C99 x1.gno3 Z 9.07e-20
C100 x1.gpo0 VPWR 3.28453f
C101 a_5645_5909# select2 8.66e-20
C102 a_5645_5909# select0 0.246189f
C103 x1.gpo3 A7 0.00162f
C104 m2_5776_5494# a_5645_5493# 0.01297f
C105 x1.gpo1 A1 0.002755f
C106 A8 x1.gno3 3.84592f
C107 m2_5776_5494# x1.nSEL0 3.43e-19
C108 x1.nSEL2 A2 0.011628f
C109 select2 x1.nSEL1 0.164995f
C110 select1 x1.gno0 0.312176f
C111 A6 x1.gpo3 1.72e-19
C112 x1.nSEL1 select0 0.169954f
C113 select2 x1.gpo1 4.34e-19
C114 x1.gpo1 select0 4.71e-19
C115 x1.gno0 VPWR 0.889132f
C116 select1 a_5645_5909# 0.03417f
C117 a_5671_6037# VPWR 4.32e-19
C118 a_5645_5493# a_5699_5631# 0.006584f
C119 a_5645_5909# VPWR 0.162117f
C120 x1.nSEL2 A1 0.566094f
C121 x1.gpo3 A4 3.96247f
C122 A5 x1.gpo3 0.098584f
C123 x1.gno3 A7 0.180503f
C124 x5.A x1.gpo0 0.35382f
C125 a_5645_6085# select2 1.67e-19
C126 select2 x1.nSEL2 4.00521f
C127 a_5645_6085# select0 0.143958f
C128 select1 x1.nSEL1 0.275603f
C129 x1.nSEL2 select0 0.131913f
C130 x1.gpo0 x3.Z3 0.354991f
C131 A3 x1.gpo3 0.00162f
C132 x1.nSEL1 VPWR 0.472688f
C133 select1 x1.gpo1 3.1e-20
C134 A6 x1.gno3 1.76e-19
C135 x1.gpo1 VPWR 3.26715f
C136 a_5645_5493# x1.nSEL0 0.081627f
C137 a_5671_6589# select0 0.001558f
C138 m2_5776_5494# x1.gno0 0.06935f
C139 x1.gpo3 A2 1.55e-19
C140 x1.gno3 A4 3.82666f
C141 A5 x1.gno3 0.005885f
C142 a_5645_6085# select1 0.254026f
C143 x1.gno0 x3.Z3 0.428132f
C144 select1 x1.nSEL2 0.140519f
C145 a_5645_6085# VPWR 0.193284f
C146 x5.A x1.gno0 0.430802f
C147 A3 x1.gno3 0.16467f
C148 x1.nSEL2 VPWR 3.6311f
C149 x1.nSEL0 x1.gpo0 6.21e-20
C150 a_5645_6461# select0 0.086353f
C151 x1.gpo3 A1 1.62e-19
C152 a_5645_6461# select2 0.009143f
C153 x1.gno0 a_5699_5631# 0.001144f
C154 m2_5776_5494# x1.nSEL1 0.00815f
C155 a_5671_6589# VPWR 0.001496f
C156 x1.gpo3 select0 0.001185f
C157 x1.gpo1 x3.Z3 0.350405f
C158 select2 x1.gpo3 0.006992f
C159 A2 x1.gno3 1.76e-19
C160 x5.A x1.gpo1 0.350703f
C161 a_5699_5631# x1.nSEL1 0.00175f
C162 x1.gno0 x1.nSEL0 0.002613f
C163 a_5645_5493# x1.gno0 0.128677f
C164 select1 a_5645_6461# 0.261734f
C165 a_5645_5493# a_5645_5909# 0.002207f
C166 a_5671_6037# x1.nSEL0 2.51e-19
C167 a_5645_5909# x1.nSEL0 0.03096f
C168 m2_5776_5494# x1.nSEL2 4e-19
C169 x1.gno3 A1 1.72e-19
C170 a_5645_6461# VPWR 0.171399f
C171 select1 x1.gpo3 3.7e-19
C172 x1.nSEL2 x3.Z3 4.15404f
C173 x5.A x1.nSEL2 4.05923f
C174 x1.gno3 select0 0.218342f
C175 a_5645_6637# select0 0.279858f
C176 x1.nSEL0 x1.nSEL1 0.352716f
C177 select2 x1.gno3 5.71e-20
C178 a_5645_5493# x1.nSEL1 0.193944f
C179 x1.gno0 x1.gpo0 2.99937f
C180 x1.gpo3 VPWR 2.92994f
C181 x1.nSEL2 a_5699_5631# 1.95e-19
C182 a_5645_5909# x1.gpo0 9.98e-19
C183 select1 x1.gno3 0.059776f
C184 select1 a_5645_6637# 0.127717f
C185 x1.nSEL1 x1.gpo0 1.17e-19
C186 x1.gpo1 x1.gpo0 0.101838f
C187 a_5645_6085# x1.nSEL0 0.001174f
C188 x1.nSEL2 x1.nSEL0 0.043717f
C189 a_5645_5493# x1.nSEL2 0.001336f
C190 a_5699_7287# select0 1.4e-19
C191 a_5645_7149# select0 0.220366f
C192 x1.gno3 VPWR 1.35568f
C193 a_5645_6637# VPWR 0.262163f
C194 a_5671_6037# x1.gno0 1.22e-20
C195 a_5671_6037# a_5645_5909# 0.004764f
C196 a_5645_5909# x1.gno0 0.012357f
C197 x1.gpo3 x3.Z3 0.3315f
C198 x5.A x1.gpo3 0.278763f
C199 a_5671_6037# x1.nSEL1 9.57e-19
C200 x1.gno0 x1.nSEL1 0.034871f
C201 x1.nSEL2 x1.gpo0 0.045168f
C202 select1 a_5699_7287# 8.84e-19
C203 x1.gno0 x1.gpo1 0.069439f
C204 select1 a_5645_7149# 0.125445f
C205 a_5645_5909# x1.nSEL1 0.073392f
C206 a_5645_7149# VPWR 0.217381f
C207 a_5645_6461# x1.nSEL0 1.91e-20
C208 a_5699_7287# VPWR 8.97e-19
C209 x1.gno3 x3.Z3 0.446539f
C210 x5.A x1.gno3 0.446599f
C211 a_5645_6085# x1.gno0 1.45e-19
C212 x1.gno0 x1.nSEL2 0.645006f
C213 a_5671_6037# x1.nSEL2 1.08e-19
C214 a_5645_6085# a_5645_5909# 0.185422f
C215 a_5645_5909# x1.nSEL2 3.56e-19
C216 a_5645_6461# x1.gpo0 1.19e-20
C217 a_5645_6085# x1.nSEL1 0.041068f
C218 x1.nSEL2 x1.nSEL1 0.10521f
C219 x1.gpo3 x1.gpo0 0.080341f
C220 x1.nSEL0 x1.gno3 2.26e-20
C221 x1.nSEL2 x1.gpo1 1.7e-20
C222 a_5645_6637# x1.nSEL0 1.21e-20
C223 a_5671_6589# x1.nSEL1 4.08e-19
C224 a_5645_6461# x1.gno0 7.95e-20
C225 a_5645_6085# x1.nSEL2 3.26e-19
C226 x1.gno0 x1.gpo3 0.848624f
C227 x1.gno3 x1.gpo0 0.066343f
C228 a_5645_6461# x1.nSEL1 7.84e-19
C229 a_5645_6461# x1.gpo1 2.46e-19
C230 a_5671_6589# x1.nSEL2 9.76e-20
C231 x1.gpo3 x1.gpo1 0.069892f
C232 a_5645_6637# x1.gno0 1.69e-20
C233 x1.gno0 x1.gno3 0.145529f
C234 a_5645_6461# x1.nSEL2 3.51e-19
C235 a_5645_6085# a_5645_6461# 3.02e-19
C236 x1.nSEL2 x1.gpo3 1.12e-19
C237 a_5645_6637# x1.nSEL1 1.59e-19
C238 x1.gpo1 x1.gno3 0.062916f
C239 a_5645_6637# x1.gpo1 2.95e-20
C240 a_5645_6461# a_5671_6589# 0.004764f
C241 x1.nSEL2 x1.gno3 9.02e-19
C242 a_5645_6637# x1.nSEL2 2.27e-19
C243 a_5671_6589# x1.gno3 3.22e-19
C244 a_5645_7149# x1.nSEL2 1.19e-19
C245 a_5645_6461# x1.gno3 6.84e-19
C246 a_5645_6461# a_5645_6637# 0.185422f
C247 x1.gpo3 x1.gno3 5.58658f
C248 a_5645_6637# x1.gpo3 4.96e-19
C249 a_5645_6637# x1.gno3 0.003645f
C250 a_5699_7287# x1.gpo3 1e-19
C251 a_5645_7149# x1.gpo3 2.98e-19
C252 a_5699_7287# x1.gno3 0.001562f
C253 a_5645_7149# x1.gno3 0.134079f
C254 a_5699_7287# a_5645_7149# 0.006584f
C255 x1.gno2 A8 0.006957f
C256 x1.gno2 A7 3.80762f
C257 x1.gno2 A6 0.156179f
C258 x1.gno2 A4 0.007342f
C259 x1.gno2 A5 2.86e-19
C260 x1.gno2 A3 3.78522f
C261 x1.gno2 A2 0.137879f
C262 x1.gno2 A1 2.84e-19
C263 x1.gno2 select2 0.00233f
C264 x1.gno2 select0 0.254198f
C265 select1 x1.gno2 0.272271f
C266 x1.gno2 VPWR 0.767412f
C267 x1.gno2 x5.A 0.429924f
C268 x1.gno2 x3.Z3 0.429865f
C269 x1.gno2 x1.nSEL0 4.01e-20
C270 x1.gno2 x1.gpo0 0.056456f
C271 x1.gno2 x1.gno0 0.089083f
C272 x1.gno2 a_5671_6037# 5.17e-20
C273 x1.gno2 a_5645_5909# 6.68e-19
C274 x1.gno2 x1.nSEL1 0.012418f
C275 x1.gno2 x1.gpo1 4.59188f
C276 a_5645_6085# x1.gno2 0.048646f
C277 x1.gno2 x1.nSEL2 1.63e-19
C278 x1.gno2 a_5671_6589# 0.001073f
C279 a_5645_6461# x1.gno2 0.104374f
C280 x1.gno2 x1.gpo3 0.072782f
C281 x1.gno2 x1.gno3 0.195239f
C282 x1.gno2 a_5645_6637# 0.004289f
C283 x1.gno2 a_5699_7287# 1.07e-20
C284 x1.gno2 a_5645_7149# 1.07e-20
C285 x1.gno1 Z 9.36e-20
C286 x1.gpo2 Z 2.44e-19
C287 A8 x1.gpo2 0.161339f
C288 x1.gno1 A7 0.006482f
C289 x1.gno1 A6 3.81297f
C290 x1.gpo2 A7 4.00999f
C291 x1.gno1 A4 6.05e-19
C292 x1.gno1 A5 0.145599f
C293 x1.gpo2 A6 0.001573f
C294 x1.gno1 A3 0.007138f
C295 x1.gpo2 A4 0.162086f
C296 A5 x1.gpo2 2.05e-19
C297 x1.gpo2 A3 3.96087f
C298 x1.gno1 A2 3.7791f
C299 x1.gpo2 A2 0.001569f
C300 x1.gno1 A1 0.13437f
C301 x1.gno1 select2 0.001516f
C302 x1.gno1 select0 0.114399f
C303 x1.gpo2 A1 1.96e-19
C304 select2 x1.gpo2 1.6e-19
C305 x1.gpo2 select0 2.74e-19
C306 x1.gno1 select1 0.108644f
C307 x1.gno1 VPWR 0.699246f
C308 select1 x1.gpo2 0.003325f
C309 x1.gpo2 VPWR 3.24607f
C310 x1.gno1 x3.Z3 0.429208f
C311 x1.gno1 x5.A 0.429382f
C312 x1.gno1 a_5699_5631# 8.86e-19
C313 x1.gpo2 x3.Z3 0.358391f
C314 x5.A x1.gpo2 0.358718f
C315 x1.gno1 x1.nSEL0 0.154394f
C316 x1.gno1 a_5645_5493# 0.039612f
C317 x1.gno1 x1.gpo0 4.59887f
C318 x1.gpo2 x1.gpo0 0.062293f
C319 x1.gno1 x1.gno0 0.146872f
C320 x1.gno1 a_5671_6037# 0.002395f
C321 x1.gno1 a_5645_5909# 0.106139f
C322 x1.gno0 x1.gpo2 0.076333f
C323 x1.gno1 x1.nSEL1 0.209954f
C324 x1.gno1 x1.gpo1 3.78638f
C325 x1.gpo2 x1.gpo1 0.096269f
C326 a_5645_6085# x1.gno1 0.016995f
C327 x1.gno1 x1.nSEL2 0.019435f
C328 x1.gno1 a_5671_6589# 3.11e-20
C329 x1.gpo2 x1.nSEL2 3.82e-20
C330 a_5671_6589# x1.gpo2 4.39e-19
C331 x1.gno1 a_5645_6461# 1.61e-19
C332 x1.gno1 x1.gpo3 0.068595f
C333 a_5645_6461# x1.gpo2 0.001353f
C334 x1.gpo2 x1.gpo3 0.109471f
C335 x1.gno1 x1.gno3 0.061048f
C336 x1.gno1 a_5645_6637# 1.03e-19
C337 x1.gpo2 x1.gno3 5.65242f
C338 a_5645_6637# x1.gpo2 4.69e-19
C339 x1.gno1 a_5699_7287# 8.14e-21
C340 x1.gno1 a_5645_7149# 7.58e-21
C341 Z VGND 6.578722f
C342 A8 VGND 3.687544f
C343 A7 VGND 3.163578f
C344 A6 VGND 3.279698f
C345 A5 VGND 3.5005f
C346 A4 VGND 3.017403f
C347 A3 VGND 3.186499f
C348 A2 VGND 3.320398f
C349 A1 VGND 4.042872f
C350 select2 VGND 6.567346f
C351 select0 VGND 1.45124f
C352 select1 VGND 1.80202f
C353 VPWR VGND 0.117673p
C354 m2_5776_5494# VGND 0.065655f $ **FLOATING
C355 x3.Z3 VGND 16.058199f
C356 x5.A VGND 12.524099f
C357 a_5699_5631# VGND 0.006505f
C358 a_5645_5493# VGND 0.266782f
C359 x1.nSEL0 VGND 0.650696f
C360 x1.gpo0 VGND 10.456742f
C361 x1.gno0 VGND 11.723553f
C362 a_5671_6037# VGND 0.004461f
C363 a_5645_5909# VGND 0.220868f
C364 x1.nSEL1 VGND 0.682637f
C365 x1.gpo1 VGND 10.05377f
C366 x1.gno1 VGND 7.03383f
C367 a_5645_6085# VGND 0.23458f
C368 x1.nSEL2 VGND 5.45531f
C369 x1.gpo2 VGND 3.19357f
C370 a_5671_6589# VGND 0.006801f
C371 x1.gno2 VGND 6.82653f
C372 a_5645_6461# VGND 0.232731f
C373 x1.gpo3 VGND 12.517524f
C374 a_5645_6637# VGND 0.249604f
C375 x1.gno3 VGND 13.497057f
C376 a_5699_7287# VGND 0.006583f
C377 a_5645_7149# VGND 0.307391f
C378 x1.gpo1.t3 VGND 0.018013f
C379 x1.gpo1.t2 VGND 0.018013f
C380 x1.gpo1.n0 VGND 0.042951f
C381 x1.gpo1.n1 VGND 0.084381f
C382 x1.gpo1.n2 VGND 0.026255f
C383 x1.gpo1.t5 VGND 0.911601f
C384 x1.gpo1.t7 VGND 0.937021f
C385 x1.gpo1.n3 VGND 3.3244f
C386 x1.gpo1.t4 VGND 0.911601f
C387 x1.gpo1.t6 VGND 0.937021f
C388 x1.gpo1.n4 VGND 3.3244f
C389 x1.gpo1.n5 VGND 1.96615f
C390 x1.gpo1.t1 VGND 0.027712f
C391 x1.gpo1.t0 VGND 0.027712f
C392 x1.gpo1.n6 VGND 0.057149f
C393 x1.gpo1.n7 VGND 0.119653f
C394 A8.t1 VGND 0.893325f
C395 A8.t0 VGND 0.512841f
C396 A8.n0 VGND 4.96695f
C397 A8.t3 VGND 0.924602f
C398 A8.t2 VGND 0.65407f
C399 A8.n1 VGND 5.0783f
C400 A8.n2 VGND 0.803255f
C401 A8.n3 VGND 0.258761f
C402 A6.t3 VGND 0.763965f
C403 A6.t2 VGND 0.438578f
C404 A6.n0 VGND 4.2477f
C405 A6.t0 VGND 0.790712f
C406 A6.t1 VGND 0.559356f
C407 A6.n1 VGND 4.34292f
C408 A6.n2 VGND 0.686937f
C409 A6.n3 VGND 0.222065f
C410 A3.t1 VGND 0.893857f
C411 A3.t0 VGND 0.513146f
C412 A3.n0 VGND 4.9699f
C413 A3.t3 VGND 0.925152f
C414 A3.t2 VGND 0.654459f
C415 A3.n1 VGND 5.08132f
C416 A3.n2 VGND 0.803733f
C417 A3.n3 VGND 0.264783f
C418 A7.t1 VGND 0.893857f
C419 A7.t0 VGND 0.513146f
C420 A7.n0 VGND 4.9699f
C421 A7.t2 VGND 0.925152f
C422 A7.t3 VGND 0.654459f
C423 A7.n1 VGND 5.08132f
C424 A7.n2 VGND 0.803733f
C425 A7.n3 VGND 0.264783f
C426 A4.t1 VGND 0.893325f
C427 A4.t0 VGND 0.512841f
C428 A4.n0 VGND 4.96695f
C429 A4.t2 VGND 0.924602f
C430 A4.t3 VGND 0.65407f
C431 A4.n1 VGND 5.0783f
C432 A4.n2 VGND 0.803255f
C433 A4.n3 VGND 0.258761f
C434 A2.t1 VGND 0.763965f
C435 A2.t2 VGND 0.438578f
C436 A2.n0 VGND 4.2477f
C437 A2.t0 VGND 0.790712f
C438 A2.t3 VGND 0.559356f
C439 A2.n1 VGND 4.34292f
C440 A2.n2 VGND 0.686937f
C441 A2.n3 VGND 0.222065f
C442 A1.t2 VGND 0.795131f
C443 A1.t3 VGND 0.45647f
C444 A1.n0 VGND 4.42098f
C445 A1.t0 VGND 0.82297f
C446 A1.t1 VGND 0.582175f
C447 A1.n1 VGND 4.52009f
C448 A1.n2 VGND 0.714961f
C449 A1.n3 VGND 0.223162f
C450 x1.gpo0.t3 VGND 0.01774f
C451 x1.gpo0.t2 VGND 0.01774f
C452 x1.gpo0.n0 VGND 0.0423f
C453 x1.gpo0.n1 VGND 0.083102f
C454 x1.gpo0.n2 VGND 0.025857f
C455 x1.gpo0.t6 VGND 0.897787f
C456 x1.gpo0.t7 VGND 0.922822f
C457 x1.gpo0.n3 VGND 3.26002f
C458 x1.gpo0.t4 VGND 0.897787f
C459 x1.gpo0.t5 VGND 0.922822f
C460 x1.gpo0.n4 VGND 3.29215f
C461 x1.gpo0.n5 VGND 1.7367f
C462 x1.gpo0.t1 VGND 0.027292f
C463 x1.gpo0.t0 VGND 0.027292f
C464 x1.gpo0.n6 VGND 0.056236f
C465 x1.gpo0.n7 VGND 0.120059f
C466 x1.gpo3.t2 VGND 0.01237f
C467 x1.gpo3.t3 VGND 0.01237f
C468 x1.gpo3.n0 VGND 0.029497f
C469 x1.gpo3.n1 VGND 0.056891f
C470 x1.gpo3.t6 VGND 0.626043f
C471 x1.gpo3.t4 VGND 0.643501f
C472 x1.gpo3.n2 VGND 2.2877f
C473 x1.gpo3.t5 VGND 0.626043f
C474 x1.gpo3.t7 VGND 0.643501f
C475 x1.gpo3.n3 VGND 2.2877f
C476 x1.gpo3.n4 VGND 2.68712f
C477 x1.gpo3.n5 VGND 0.0412f
C478 x1.gpo3.n6 VGND 0.01803f
C479 x1.gpo3.t0 VGND 0.019031f
C480 x1.gpo3.t1 VGND 0.019031f
C481 x1.gpo3.n7 VGND 0.041797f
C482 x1.gno3.t1 VGND 0.053338f
C483 x1.gno3.n0 VGND 0.061486f
C484 x1.gno3.t6 VGND 0.60277f
C485 x1.gno3.t9 VGND 0.588227f
C486 x1.gno3.n1 VGND 2.63915f
C487 x1.gno3.n2 VGND 1.63117f
C488 x1.gno3.t3 VGND 0.60277f
C489 x1.gno3.t5 VGND 0.588227f
C490 x1.gno3.n3 VGND 2.63915f
C491 x1.gno3.n4 VGND 2.31307f
C492 x1.gno3.t4 VGND 0.033483f
C493 x1.gno3.t2 VGND 0.019731f
C494 x1.gno3.t8 VGND 0.033483f
C495 x1.gno3.t7 VGND 0.019731f
C496 x1.gno3.n5 VGND 0.05618f
C497 x1.gno3.n6 VGND 0.083224f
C498 x1.gno3.n7 VGND 0.037258f
C499 x1.gno3.n8 VGND 0.301796f
C500 x1.gno3.t0 VGND 0.13622f
C501 x1.gno3.n9 VGND 0.024501f
C502 x1.gno3.n10 VGND 0.027448f
C503 A5.t3 VGND 0.770284f
C504 A5.t2 VGND 0.442205f
C505 A5.n0 VGND 4.28283f
C506 A5.t0 VGND 0.797252f
C507 A5.t1 VGND 0.563982f
C508 A5.n1 VGND 4.37884f
C509 A5.n2 VGND 0.692619f
C510 A5.n3 VGND 0.216188f
C511 x1.gno0.n0 VGND 1.21068f
C512 x1.gno0.t1 VGND 0.038064f
C513 x1.gno0.n1 VGND 0.043923f
C514 x1.gno0.t9 VGND 0.430161f
C515 x1.gno0.t7 VGND 0.419783f
C516 x1.gno0.n2 VGND 1.8834f
C517 x1.gno0.t2 VGND 0.430161f
C518 x1.gno0.t3 VGND 0.419783f
C519 x1.gno0.n3 VGND 1.8834f
C520 x1.gno0.n4 VGND 0.892351f
C521 x1.gno0.n5 VGND 0.304041f
C522 x1.gno0.t8 VGND 0.023895f
C523 x1.gno0.t5 VGND 0.014081f
C524 x1.gno0.t6 VGND 0.023895f
C525 x1.gno0.t4 VGND 0.014081f
C526 x1.gno0.n6 VGND 0.040092f
C527 x1.gno0.n7 VGND 0.059217f
C528 x1.gno0.n8 VGND 0.057595f
C529 x1.gno0.n9 VGND 0.1251f
C530 x1.gno0.t0 VGND 0.097212f
C531 x1.gno0.n10 VGND 0.017485f
C532 x1.gno0.n11 VGND 0.019588f
C533 VPWR.n0 VGND 0.078152f
C534 VPWR.n1 VGND 0.253693f
C535 VPWR.n2 VGND 0.122926f
C536 VPWR.n3 VGND 0.122926f
C537 VPWR.n4 VGND 0.122525f
C538 VPWR.n5 VGND 0.169863f
C539 VPWR.n6 VGND 0.547624f
C540 VPWR.t1 VGND 0.790353f
C541 VPWR.n7 VGND 0.763087f
C542 VPWR.t0 VGND 0.790353f
C543 VPWR.n8 VGND 0.547624f
C544 VPWR.n9 VGND 0.004814f
C545 VPWR.n10 VGND 0.134493f
C546 VPWR.n11 VGND 0.040318f
C547 VPWR.n12 VGND 0.138067f
C548 VPWR.n13 VGND 0.057005f
C549 VPWR.n14 VGND 0.253704f
C550 VPWR.n15 VGND 0.122531f
C551 VPWR.n16 VGND 1.03197f
C552 VPWR.n17 VGND 1.03197f
C553 VPWR.n18 VGND 0.169845f
C554 VPWR.n19 VGND 0.124397f
C555 VPWR.t7 VGND 1.37216f
C556 VPWR.n22 VGND 0.124397f
C557 VPWR.n23 VGND 5.27e-19
C558 VPWR.n24 VGND 0.07554f
C559 VPWR.n25 VGND 0.013735f
C560 VPWR.n26 VGND 0.149327f
C561 VPWR.n27 VGND 0.079843f
C562 VPWR.n28 VGND 0.162134f
C563 VPWR.n29 VGND 0.188097f
C564 VPWR.n30 VGND 0.253704f
C565 VPWR.n31 VGND 0.004119f
C566 VPWR.n32 VGND 0.169845f
C567 VPWR.n33 VGND 0.124397f
C568 VPWR.t77 VGND 1.37216f
C569 VPWR.n35 VGND 1.03197f
C570 VPWR.n36 VGND 0.124397f
C571 VPWR.n38 VGND 1.03197f
C572 VPWR.n39 VGND 0.122531f
C573 VPWR.n40 VGND 0.009862f
C574 VPWR.n41 VGND 0.075465f
C575 VPWR.n42 VGND 0.013861f
C576 VPWR.n43 VGND 0.149327f
C577 VPWR.n44 VGND 0.079211f
C578 VPWR.n45 VGND 0.128376f
C579 VPWR.n46 VGND 0.184404f
C580 VPWR.n47 VGND 0.253704f
C581 VPWR.n48 VGND 0.00437f
C582 VPWR.n49 VGND 0.169845f
C583 VPWR.n50 VGND 0.124397f
C584 VPWR.t6 VGND 1.37216f
C585 VPWR.n52 VGND 1.03197f
C586 VPWR.n53 VGND 0.124397f
C587 VPWR.n55 VGND 1.03197f
C588 VPWR.n56 VGND 0.122531f
C589 VPWR.n57 VGND 0.009878f
C590 VPWR.n58 VGND 0.075214f
C591 VPWR.n59 VGND 0.013861f
C592 VPWR.n60 VGND 0.149327f
C593 VPWR.n61 VGND 0.079211f
C594 VPWR.n62 VGND 0.125941f
C595 VPWR.n63 VGND 0.167914f
C596 VPWR.n64 VGND 0.010164f
C597 VPWR.n65 VGND 0.00773f
C598 VPWR.t39 VGND 0.015599f
C599 VPWR.n66 VGND 0.015344f
C600 VPWR.t13 VGND 0.001675f
C601 VPWR.t55 VGND 0.002544f
C602 VPWR.n67 VGND 0.004395f
C603 VPWR.t37 VGND 0.015899f
C604 VPWR.t76 VGND 0.015599f
C605 VPWR.n68 VGND 0.014858f
C606 VPWR.n69 VGND 0.00773f
C607 VPWR.n70 VGND 0.006997f
C608 VPWR.t43 VGND 0.002296f
C609 VPWR.n71 VGND 0.006515f
C610 VPWR.t35 VGND 0.009437f
C611 VPWR.n72 VGND 0.008687f
C612 VPWR.n73 VGND 0.007753f
C613 VPWR.t9 VGND 0.015603f
C614 VPWR.n74 VGND 0.001276f
C615 VPWR.t51 VGND 0.00669f
C616 VPWR.t64 VGND 0.011043f
C617 VPWR.n75 VGND 0.010887f
C618 VPWR.n76 VGND 0.013048f
C619 VPWR.t79 VGND 0.046088f
C620 VPWR.n77 VGND 0.041686f
C621 VPWR.t41 VGND 0.00125f
C622 VPWR.t47 VGND 0.003352f
C623 VPWR.n78 VGND 0.0153f
C624 VPWR.t65 VGND 0.011043f
C625 VPWR.n79 VGND 0.008081f
C626 VPWR.n80 VGND 0.030158f
C627 VPWR.n81 VGND 0.023827f
C628 VPWR.n82 VGND 0.030949f
C629 VPWR.n83 VGND 0.01787f
C630 VPWR.n84 VGND 0.013048f
C631 VPWR.n85 VGND 0.009786f
C632 VPWR.n86 VGND 0.006143f
C633 VPWR.n87 VGND 0.019352f
C634 VPWR.n88 VGND 0.030339f
C635 VPWR.t44 VGND 0.031357f
C636 VPWR.n89 VGND 0.002361f
C637 VPWR.n90 VGND 0.002411f
C638 VPWR.n91 VGND 0.009786f
C639 VPWR.n92 VGND 0.003014f
C640 VPWR.t33 VGND 0.015814f
C641 VPWR.n93 VGND 0.012977f
C642 VPWR.n94 VGND 0.00773f
C643 VPWR.t80 VGND 0.046088f
C644 VPWR.n95 VGND 0.011488f
C645 VPWR.n96 VGND 0.00773f
C646 VPWR.t3 VGND 0.00125f
C647 VPWR.t62 VGND 0.003352f
C648 VPWR.n97 VGND 0.0153f
C649 VPWR.t82 VGND 0.046088f
C650 VPWR.t17 VGND 0.00669f
C651 VPWR.n98 VGND 0.020658f
C652 VPWR.n99 VGND 0.011843f
C653 VPWR.n100 VGND 0.006143f
C654 VPWR.t67 VGND 0.011043f
C655 VPWR.n101 VGND 0.010887f
C656 VPWR.n102 VGND 0.041686f
C657 VPWR.n103 VGND 0.01787f
C658 VPWR.n104 VGND 0.030949f
C659 VPWR.t68 VGND 0.011043f
C660 VPWR.t49 VGND 0.015815f
C661 VPWR.n105 VGND 0.004468f
C662 VPWR.n106 VGND 0.005319f
C663 VPWR.t16 VGND 0.063133f
C664 VPWR.t61 VGND 0.061042f
C665 VPWR.t66 VGND 0.045154f
C666 VPWR.t2 VGND 0.064805f
C667 VPWR.t23 VGND 0.063133f
C668 VPWR.t10 VGND 0.071913f
C669 VPWR.t56 VGND 0.052262f
C670 VPWR.t20 VGND 0.028013f
C671 VPWR.t32 VGND 0.012961f
C672 VPWR.t48 VGND 0.045572f
C673 VPWR.n107 VGND 0.059469f
C674 VPWR.n108 VGND 0.041241f
C675 VPWR.n109 VGND 0.012122f
C676 VPWR.n110 VGND 0.01945f
C677 VPWR.n111 VGND 0.023827f
C678 VPWR.n112 VGND 0.008084f
C679 VPWR.n113 VGND 0.064395f
C680 VPWR.n114 VGND 0.087594f
C681 VPWR.t73 VGND 0.011043f
C682 VPWR.n115 VGND 0.021596f
C683 VPWR.n116 VGND 0.041686f
C684 VPWR.n117 VGND 0.025689f
C685 VPWR.t74 VGND 0.011043f
C686 VPWR.t27 VGND 0.015891f
C687 VPWR.n118 VGND 0.018568f
C688 VPWR.t72 VGND 0.142033f
C689 VPWR.t69 VGND 0.087258f
C690 VPWR.t52 VGND 0.035804f
C691 VPWR.t58 VGND 0.049557f
C692 VPWR.t14 VGND 0.035804f
C693 VPWR.t18 VGND 0.049557f
C694 VPWR.t29 VGND 0.035804f
C695 VPWR.t26 VGND 0.053589f
C696 VPWR.n119 VGND 0.058661f
C697 VPWR.n120 VGND 0.00773f
C698 VPWR.n121 VGND 0.003365f
C699 VPWR.t19 VGND 0.015891f
C700 VPWR.n122 VGND 0.003365f
C701 VPWR.t59 VGND 0.015891f
C702 VPWR.n123 VGND 0.227132f
C703 VPWR.n124 VGND 0.013294f
C704 VPWR.n125 VGND 0.008081f
C705 VPWR.t81 VGND 0.046809f
C706 VPWR.t70 VGND 0.011043f
C707 VPWR.n126 VGND 0.04634f
C708 VPWR.n127 VGND 0.023029f
C709 VPWR.t71 VGND 0.011043f
C710 VPWR.n128 VGND 0.030158f
C711 VPWR.n129 VGND 0.027736f
C712 VPWR.n130 VGND 0.017403f
C713 VPWR.n131 VGND 0.013581f
C714 VPWR.n132 VGND 0.013243f
C715 VPWR.t53 VGND 0.015899f
C716 VPWR.n133 VGND 0.020008f
C717 VPWR.n134 VGND 0.00773f
C718 VPWR.n135 VGND 0.013048f
C719 VPWR.n136 VGND 0.009786f
C720 VPWR.n137 VGND 0.018769f
C721 VPWR.t15 VGND 0.015899f
C722 VPWR.n138 VGND 0.02031f
C723 VPWR.n139 VGND 0.00773f
C724 VPWR.n140 VGND 0.013048f
C725 VPWR.n141 VGND 0.009786f
C726 VPWR.n142 VGND 0.018769f
C727 VPWR.t30 VGND 0.015899f
C728 VPWR.n143 VGND 0.02031f
C729 VPWR.n144 VGND 0.003365f
C730 VPWR.n145 VGND 0.013048f
C731 VPWR.n146 VGND 0.009786f
C732 VPWR.n147 VGND 0.004964f
C733 VPWR.n148 VGND 0.027117f
C734 VPWR.n149 VGND 0.012122f
C735 VPWR.n150 VGND 0.01945f
C736 VPWR.n151 VGND 0.033134f
C737 VPWR.n152 VGND 0.006595f
C738 VPWR.n153 VGND 0.059927f
C739 VPWR.n154 VGND 0.058109f
C740 VPWR.n155 VGND 0.001347f
C741 VPWR.t21 VGND 0.001675f
C742 VPWR.t57 VGND 0.002544f
C743 VPWR.n156 VGND 0.004395f
C744 VPWR.n157 VGND 0.029498f
C745 VPWR.t25 VGND 0.015891f
C746 VPWR.n158 VGND 0.018518f
C747 VPWR.t11 VGND 0.005236f
C748 VPWR.t45 VGND 0.013917f
C749 VPWR.n159 VGND 0.007895f
C750 VPWR.t24 VGND 0.015603f
C751 VPWR.n160 VGND 0.016462f
C752 VPWR.n161 VGND 0.021174f
C753 VPWR.n162 VGND 0.002788f
C754 VPWR.n163 VGND 0.013048f
C755 VPWR.n164 VGND 0.00773f
C756 VPWR.n165 VGND 0.004468f
C757 VPWR.n166 VGND 0.004964f
C758 VPWR.n167 VGND 0.026569f
C759 VPWR.n168 VGND 0.072449f
C760 VPWR.t12 VGND 0.013797f
C761 VPWR.t38 VGND 0.035956f
C762 VPWR.t36 VGND 0.040137f
C763 VPWR.t54 VGND 0.028013f
C764 VPWR.t42 VGND 0.052262f
C765 VPWR.t75 VGND 0.073585f
C766 VPWR.t8 VGND 0.035956f
C767 VPWR.t34 VGND 0.028013f
C768 VPWR.t40 VGND 0.064805f
C769 VPWR.t63 VGND 0.045154f
C770 VPWR.t46 VGND 0.061042f
C771 VPWR.t50 VGND 0.063133f
C772 VPWR.n169 VGND 0.042993f
C773 VPWR.n170 VGND 0.01249f
C774 VPWR.n171 VGND 0.008891f
C775 VPWR.n172 VGND 0.002361f
C776 VPWR.n173 VGND 0.017322f
C777 VPWR.n174 VGND 0.006606f
C778 VPWR.n175 VGND 0.013048f
C779 VPWR.n176 VGND 0.009786f
C780 VPWR.n177 VGND 0.005817f
C781 VPWR.n178 VGND 0.019774f
C782 VPWR.n179 VGND 0.014151f
C783 VPWR.n180 VGND 0.009006f
C784 VPWR.n181 VGND 0.025467f
C785 VPWR.n182 VGND 0.279991f
C786 VPWR.n183 VGND 0.651519f
C787 VPWR.n184 VGND 0.253704f
C788 VPWR.n185 VGND 0.051921f
C789 VPWR.n186 VGND 0.122531f
C790 VPWR.n187 VGND 1.03197f
C791 VPWR.n188 VGND 1.03197f
C792 VPWR.n189 VGND 0.169845f
C793 VPWR.n190 VGND 0.124397f
C794 VPWR.t60 VGND 1.37216f
C795 VPWR.n193 VGND 0.124397f
C796 VPWR.n194 VGND 4.77e-19
C797 VPWR.n195 VGND 0.07554f
C798 VPWR.n196 VGND 0.013785f
C799 VPWR.n197 VGND 0.149327f
C800 VPWR.n198 VGND 0.079793f
C801 VPWR.n199 VGND 0.15219f
C802 VPWR.n200 VGND 0.253704f
C803 VPWR.n201 VGND 0.00437f
C804 VPWR.n202 VGND 0.169845f
C805 VPWR.n203 VGND 0.124397f
C806 VPWR.t5 VGND 1.37216f
C807 VPWR.n205 VGND 1.03197f
C808 VPWR.n206 VGND 0.124397f
C809 VPWR.n208 VGND 1.03197f
C810 VPWR.n209 VGND 0.122531f
C811 VPWR.n210 VGND 0.075214f
C812 VPWR.n211 VGND 0.013861f
C813 VPWR.n212 VGND 0.149327f
C814 VPWR.n213 VGND 0.079211f
C815 VPWR.n214 VGND 0.153404f
C816 VPWR.n215 VGND 0.196603f
C817 VPWR.n216 VGND 0.116414f
C818 VPWR.n217 VGND 0.075465f
C819 VPWR.n218 VGND 0.013861f
C820 VPWR.n219 VGND 1.03197f
C821 VPWR.n220 VGND 1.03197f
C822 VPWR.n221 VGND 0.122531f
C823 VPWR.n222 VGND 0.079211f
C824 VPWR.n223 VGND 0.149327f
C825 VPWR.n224 VGND 0.253704f
C826 VPWR.n225 VGND 0.169845f
C827 VPWR.n226 VGND 0.124397f
C828 VPWR.t78 VGND 1.37216f
C829 VPWR.n229 VGND 0.124397f
C830 VPWR.n230 VGND 0.004119f
C831 VPWR.n231 VGND 0.009862f
C832 VPWR.n232 VGND 0.235683f
C833 VPWR.n233 VGND 0.097082f
C834 VPWR.n234 VGND 5.27e-19
C835 VPWR.n235 VGND 0.079843f
C836 VPWR.n236 VGND 0.149327f
C837 VPWR.n237 VGND 0.169845f
C838 VPWR.n238 VGND 0.124397f
C839 VPWR.t22 VGND 1.37216f
C840 VPWR.n239 VGND 0.253704f
C841 VPWR.n241 VGND 1.03197f
C842 VPWR.n242 VGND 0.124397f
C843 VPWR.n244 VGND 1.03197f
C844 VPWR.n245 VGND 0.122531f
C845 VPWR.n246 VGND 0.07554f
C846 VPWR.n247 VGND 0.013735f
C847 VPWR.n248 VGND 0.013528f
C848 VPWR.n249 VGND 0.191035f
C849 VPWR.n250 VGND 0.253704f
C850 VPWR.n251 VGND 0.07554f
C851 VPWR.n252 VGND 1.03197f
C852 VPWR.n253 VGND 1.03197f
C853 VPWR.n254 VGND 0.122531f
C854 VPWR.n255 VGND 0.169845f
C855 VPWR.n256 VGND 0.124397f
C856 VPWR.t4 VGND 1.37216f
C857 VPWR.n259 VGND 0.124397f
C858 VPWR.n260 VGND 4.77e-19
C859 VPWR.n261 VGND 0.013492f
C860 VPWR.n262 VGND 0.013785f
C861 VPWR.n263 VGND 0.149327f
C862 VPWR.n264 VGND 0.079793f
C863 VPWR.n265 VGND 0.142932f
C864 VPWR.n266 VGND 0.154755f
C865 VPWR.n267 VGND 0.390936f
C866 VPWR.n268 VGND 0.078152f
C867 VPWR.n269 VGND 0.253693f
C868 VPWR.n270 VGND 0.122926f
C869 VPWR.n271 VGND 0.122926f
C870 VPWR.n272 VGND 0.122525f
C871 VPWR.n273 VGND 0.169863f
C872 VPWR.n274 VGND 0.547624f
C873 VPWR.t28 VGND 0.790353f
C874 VPWR.n275 VGND 0.763087f
C875 VPWR.t31 VGND 0.790353f
C876 VPWR.n276 VGND 0.547624f
C877 VPWR.n277 VGND 0.004814f
C878 VPWR.n278 VGND 0.134493f
C879 VPWR.n279 VGND 0.040288f
C880 VPWR.n280 VGND 0.072753f
C881 Z.t5 VGND 0.434416f
C882 Z.n0 VGND 0.540283f
C883 Z.t4 VGND 0.446377f
C884 Z.t1 VGND 0.336375f
C885 Z.n1 VGND 2.25255f
C886 Z.n2 VGND 0.762169f
C887 Z.t0 VGND 0.329756f
C888 Z.n3 VGND 0.492384f
C889 Z.n4 VGND 0.648657f
C890 Z.n5 VGND 0.805956f
C891 Z.t2 VGND 0.434416f
C892 Z.n6 VGND 0.540283f
C893 Z.t3 VGND 0.446377f
C894 Z.t6 VGND 0.336375f
C895 Z.n7 VGND 2.25255f
C896 Z.n8 VGND 0.762169f
C897 Z.t7 VGND 0.329756f
C898 Z.n9 VGND 0.492384f
C899 Z.n10 VGND 0.664311f
C900 Z.n11 VGND 0.690962f
C901 select2.t3 VGND 0.587307f
C902 select2.t4 VGND 0.573137f
C903 select2.n0 VGND 2.59595f
C904 select2.t1 VGND 0.032624f
C905 select2.t7 VGND 0.019225f
C906 select2.t6 VGND 0.032624f
C907 select2.t5 VGND 0.019225f
C908 select2.n1 VGND 0.054739f
C909 select2.n2 VGND 0.080926f
C910 select2.n3 VGND 0.080283f
C911 select2.n4 VGND 1.30573f
C912 select2.t2 VGND 0.689904f
C913 select2.t0 VGND 0.709143f
C914 select2.n5 VGND 2.58376f
C915 select2.n6 VGND 1.7346f
C916 select2.n7 VGND 4.54427f
C917 select2.n8 VGND 1.56778f
C918 select2.n9 VGND 0.081638f
C919 select1.t6 VGND 0.031316f
C920 select1.t5 VGND 0.018454f
C921 select1.t3 VGND 0.031316f
C922 select1.t1 VGND 0.018454f
C923 select1.n0 VGND 0.052544f
C924 select1.n1 VGND 0.077632f
C925 select1.n2 VGND 0.047269f
C926 select1.t9 VGND 0.014491f
C927 select1.t7 VGND 0.03056f
C928 select1.n3 VGND 0.109737f
C929 select1.n4 VGND 0.021277f
C930 select1.n5 VGND 0.018327f
C931 select1.t4 VGND 0.022078f
C932 select1.t2 VGND 0.015172f
C933 select1.n6 VGND 0.064155f
C934 select1.n7 VGND 0.014778f
C935 select1.n8 VGND 0.105859f
C936 select1.n9 VGND 0.383423f
C937 select1.t8 VGND 0.026898f
C938 select1.t0 VGND 0.018264f
C939 select1.n10 VGND 0.063549f
C940 select1.n11 VGND 0.015211f
C941 select1.n12 VGND 0.098666f
C942 select1.n13 VGND 0.442567f
C943 select1.n14 VGND 0.578172f
.ends

