VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_patdeegan_anamux
  CLASS BLOCK ;
  FOREIGN tt_um_patdeegan_anamux ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 20.879999 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.759998 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.759998 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 31.320000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.873000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.873000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.094999 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.746000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.746000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 143.192490 ;
    ANTENNADIFFAREA 298.813782 ;
    PORT
      LAYER met4 ;
        RECT 26.400 3.740 31.500 216.500 ;
    END
  END VDPWR
  PIN VSS
    ANTENNAGATEAREA 224.938492 ;
    ANTENNADIFFAREA 237.083939 ;
    PORT
      LAYER met4 ;
        RECT 148.900 7.040 153.990 222.340 ;
    END
  END VSS
  OBS
      LAYER nwell ;
        RECT 92.685 163.695 101.345 165.300 ;
      LAYER pwell ;
        RECT 92.880 162.495 94.710 163.305 ;
        RECT 94.730 162.495 96.080 163.405 ;
        RECT 96.110 162.495 97.460 163.405 ;
        RECT 97.490 162.495 98.840 163.405 ;
        RECT 98.870 162.580 99.300 163.365 ;
        RECT 99.320 162.495 101.150 163.305 ;
        RECT 93.020 162.305 93.190 162.495 ;
        RECT 94.860 162.305 95.030 162.495 ;
        RECT 96.240 162.305 96.410 162.495 ;
        RECT 94.860 162.285 95.010 162.305 ;
        RECT 97.620 162.285 97.790 162.495 ;
        RECT 99.460 162.305 99.630 162.495 ;
        RECT 100.380 162.285 100.550 162.475 ;
        RECT 103.140 162.305 103.310 162.475 ;
        RECT 103.140 162.285 103.290 162.305 ;
        RECT 93.080 161.465 95.010 162.285 ;
        RECT 95.180 161.605 97.930 162.285 ;
        RECT 97.940 161.605 100.690 162.285 ;
        RECT 93.080 161.375 94.030 161.465 ;
        RECT 95.180 161.375 96.110 161.605 ;
        RECT 97.940 161.375 98.870 161.605 ;
        RECT 100.710 161.415 101.140 162.200 ;
        RECT 101.360 161.465 103.290 162.285 ;
        RECT 101.360 161.375 102.310 161.465 ;
      LAYER nwell ;
        RECT 92.685 159.480 103.645 161.085 ;
        RECT 92.685 158.255 103.185 159.480 ;
      LAYER pwell ;
        RECT 92.880 157.055 94.710 157.865 ;
        RECT 94.730 157.140 95.160 157.925 ;
        RECT 95.190 157.055 96.540 157.965 ;
        RECT 96.570 157.055 97.920 157.965 ;
        RECT 97.950 157.140 98.380 157.925 ;
        RECT 98.410 157.055 99.760 157.965 ;
        RECT 99.790 157.055 101.140 157.965 ;
        RECT 101.160 157.055 102.990 157.865 ;
        RECT 93.020 156.865 93.190 157.055 ;
        RECT 95.320 156.865 95.490 157.055 ;
        RECT 96.700 156.865 96.870 157.055 ;
        RECT 98.540 156.865 98.710 157.055 ;
        RECT 99.920 156.865 100.090 157.055 ;
        RECT 101.300 156.865 101.470 157.055 ;
        RECT 61.475 130.460 63.785 149.650 ;
      LAYER nwell ;
        RECT 63.795 128.790 66.105 152.160 ;
      LAYER pwell ;
        RECT 66.765 130.650 69.075 149.840 ;
      LAYER nwell ;
        RECT 69.085 128.980 71.395 152.350 ;
      LAYER pwell ;
        RECT 74.825 149.920 94.015 152.230 ;
      LAYER nwell ;
        RECT 73.155 147.600 96.525 149.910 ;
      LAYER pwell ;
        RECT 107.920 147.525 110.990 151.825 ;
        RECT 74.835 144.570 94.025 146.880 ;
      LAYER nwell ;
        RECT 73.165 142.250 96.535 144.560 ;
      LAYER pwell ;
        RECT 104.930 144.255 110.990 147.525 ;
        RECT 74.805 139.220 93.995 141.530 ;
        RECT 104.930 139.955 108.000 144.255 ;
      LAYER nwell ;
        RECT 73.135 136.900 96.505 139.210 ;
      LAYER pwell ;
        RECT 74.845 133.940 94.035 136.250 ;
      LAYER nwell ;
        RECT 73.175 131.620 96.545 133.930 ;
      LAYER pwell ;
        RECT 74.835 128.350 94.025 130.660 ;
        RECT 104.930 130.045 108.000 137.615 ;
        RECT 108.040 134.645 111.110 142.215 ;
      LAYER nwell ;
        RECT 73.165 126.030 96.535 128.340 ;
        RECT 58.600 122.160 67.260 123.765 ;
      LAYER pwell ;
        RECT 74.845 123.000 94.035 125.310 ;
        RECT 58.795 120.960 60.625 121.770 ;
        RECT 60.645 120.960 61.995 121.870 ;
        RECT 62.025 120.960 63.375 121.870 ;
        RECT 63.405 120.960 64.755 121.870 ;
        RECT 64.785 121.045 65.215 121.830 ;
        RECT 65.235 120.960 67.065 121.770 ;
        RECT 58.935 120.770 59.105 120.960 ;
        RECT 60.775 120.770 60.945 120.960 ;
        RECT 62.155 120.770 62.325 120.960 ;
        RECT 60.775 120.750 60.925 120.770 ;
        RECT 63.535 120.750 63.705 120.960 ;
        RECT 65.375 120.770 65.545 120.960 ;
        RECT 66.295 120.750 66.465 120.940 ;
        RECT 69.055 120.770 69.225 120.940 ;
        RECT 69.055 120.750 69.205 120.770 ;
        RECT 58.995 119.930 60.925 120.750 ;
        RECT 61.095 120.070 63.845 120.750 ;
        RECT 63.855 120.070 66.605 120.750 ;
        RECT 58.995 119.840 59.945 119.930 ;
        RECT 61.095 119.840 62.025 120.070 ;
        RECT 63.855 119.840 64.785 120.070 ;
        RECT 66.625 119.880 67.055 120.665 ;
        RECT 67.275 119.930 69.205 120.750 ;
      LAYER nwell ;
        RECT 73.175 120.680 96.545 122.990 ;
      LAYER pwell ;
        RECT 104.930 121.885 108.000 127.275 ;
        RECT 108.040 124.655 111.110 132.225 ;
        RECT 67.275 119.840 68.225 119.930 ;
      LAYER nwell ;
        RECT 58.600 117.945 69.560 119.550 ;
        RECT 58.600 116.720 69.100 117.945 ;
      LAYER pwell ;
        RECT 74.815 117.650 94.005 119.960 ;
        RECT 104.930 119.705 111.050 121.885 ;
        RECT 58.795 115.520 60.625 116.330 ;
        RECT 60.645 115.605 61.075 116.390 ;
        RECT 61.105 115.520 62.455 116.430 ;
        RECT 62.485 115.520 63.835 116.430 ;
        RECT 63.865 115.605 64.295 116.390 ;
        RECT 64.325 115.520 65.675 116.430 ;
        RECT 65.705 115.520 67.055 116.430 ;
        RECT 67.075 115.520 68.905 116.330 ;
        RECT 58.935 115.330 59.105 115.520 ;
        RECT 61.235 115.330 61.405 115.520 ;
        RECT 62.615 115.330 62.785 115.520 ;
        RECT 64.455 115.330 64.625 115.520 ;
        RECT 65.835 115.330 66.005 115.520 ;
        RECT 67.215 115.330 67.385 115.520 ;
      LAYER nwell ;
        RECT 73.145 115.330 96.515 117.640 ;
      LAYER pwell ;
        RECT 107.980 117.095 111.050 119.705 ;
        RECT 74.855 112.370 94.045 114.680 ;
        RECT 104.920 114.315 111.050 117.095 ;
        RECT 44.590 109.305 63.780 111.615 ;
      LAYER nwell ;
        RECT 73.185 110.050 96.555 112.360 ;
      LAYER pwell ;
        RECT 104.920 109.525 107.990 114.315 ;
      LAYER nwell ;
        RECT 42.920 106.985 66.290 109.295 ;
      LAYER pwell ;
        RECT 44.600 103.955 63.790 106.265 ;
      LAYER nwell ;
        RECT 42.930 101.635 66.300 103.945 ;
      LAYER pwell ;
        RECT 44.570 98.605 63.760 100.915 ;
      LAYER nwell ;
        RECT 42.900 96.285 66.270 98.595 ;
      LAYER pwell ;
        RECT 44.610 93.325 63.800 95.635 ;
      LAYER nwell ;
        RECT 42.940 91.005 66.310 93.315 ;
        RECT 83.200 73.245 84.720 73.255 ;
        RECT 71.840 71.640 89.240 73.245 ;
      LAYER pwell ;
        RECT 72.045 70.525 72.475 71.310 ;
        RECT 72.505 70.440 73.855 71.350 ;
        RECT 73.885 70.440 75.235 71.350 ;
        RECT 75.265 70.440 76.615 71.350 ;
        RECT 76.645 70.440 77.995 71.350 ;
        RECT 78.025 70.440 79.375 71.350 ;
        RECT 79.405 70.440 80.755 71.350 ;
        RECT 80.785 70.440 82.135 71.350 ;
        RECT 82.165 70.440 83.515 71.350 ;
        RECT 83.545 70.440 84.895 71.350 ;
        RECT 84.925 70.525 85.355 71.310 ;
        RECT 85.385 70.525 85.815 71.310 ;
        RECT 85.845 70.525 86.275 71.310 ;
        RECT 86.305 70.525 86.735 71.310 ;
        RECT 86.755 70.440 88.945 71.350 ;
      LAYER nwell ;
        RECT 95.315 70.855 97.425 82.045 ;
        RECT 98.815 70.855 104.325 82.045 ;
      LAYER pwell ;
        RECT 72.635 70.250 72.805 70.440 ;
        RECT 73.555 70.230 73.725 70.420 ;
        RECT 74.015 70.250 74.185 70.440 ;
        RECT 74.935 70.230 75.105 70.420 ;
        RECT 75.395 70.250 75.565 70.440 ;
        RECT 76.315 70.230 76.485 70.420 ;
        RECT 76.775 70.250 76.945 70.440 ;
        RECT 77.695 70.230 77.865 70.420 ;
        RECT 78.155 70.250 78.325 70.440 ;
        RECT 79.075 70.230 79.245 70.420 ;
        RECT 79.535 70.250 79.705 70.440 ;
        RECT 80.455 70.230 80.625 70.420 ;
        RECT 80.915 70.250 81.085 70.440 ;
        RECT 81.835 70.230 82.005 70.420 ;
        RECT 82.295 70.250 82.465 70.440 ;
        RECT 83.215 70.230 83.385 70.420 ;
        RECT 83.675 70.250 83.845 70.440 ;
        RECT 84.595 70.230 84.765 70.420 ;
        RECT 86.900 70.250 87.070 70.440 ;
        RECT 72.045 69.360 72.475 70.145 ;
        RECT 72.505 69.320 73.855 70.230 ;
        RECT 73.885 69.320 75.235 70.230 ;
        RECT 75.265 69.320 76.615 70.230 ;
        RECT 76.645 69.320 77.995 70.230 ;
        RECT 78.025 69.320 79.375 70.230 ;
        RECT 79.405 69.320 80.755 70.230 ;
        RECT 80.785 69.320 82.135 70.230 ;
        RECT 82.165 69.320 83.515 70.230 ;
        RECT 83.545 69.320 84.895 70.230 ;
        RECT 84.925 69.360 85.355 70.145 ;
      LAYER nwell ;
        RECT 71.840 67.425 85.560 69.030 ;
      LAYER pwell ;
        RECT 95.315 64.355 97.425 69.455 ;
        RECT 98.815 64.355 104.325 69.455 ;
      LAYER nwell ;
        RECT 77.250 62.715 85.910 64.320 ;
      LAYER pwell ;
        RECT 77.445 61.515 79.275 62.325 ;
        RECT 79.295 61.515 80.645 62.425 ;
        RECT 80.675 61.515 82.025 62.425 ;
        RECT 82.055 61.515 83.405 62.425 ;
        RECT 83.435 61.600 83.865 62.385 ;
        RECT 83.885 61.515 85.715 62.325 ;
        RECT 77.585 61.325 77.755 61.515 ;
        RECT 79.425 61.325 79.595 61.515 ;
        RECT 80.805 61.325 80.975 61.515 ;
        RECT 79.425 61.305 79.575 61.325 ;
        RECT 82.185 61.305 82.355 61.515 ;
        RECT 84.025 61.325 84.195 61.515 ;
        RECT 84.945 61.305 85.115 61.495 ;
        RECT 87.705 61.325 87.875 61.495 ;
        RECT 87.705 61.305 87.855 61.325 ;
        RECT 77.645 60.485 79.575 61.305 ;
        RECT 79.745 60.625 82.495 61.305 ;
        RECT 82.505 60.625 85.255 61.305 ;
        RECT 77.645 60.395 78.595 60.485 ;
        RECT 79.745 60.395 80.675 60.625 ;
        RECT 82.505 60.395 83.435 60.625 ;
        RECT 85.275 60.435 85.705 61.220 ;
        RECT 85.925 60.485 87.855 61.305 ;
        RECT 85.925 60.395 86.875 60.485 ;
      LAYER nwell ;
        RECT 77.250 58.500 88.210 60.105 ;
        RECT 77.250 57.275 87.750 58.500 ;
      LAYER pwell ;
        RECT 77.445 56.075 79.275 56.885 ;
        RECT 79.295 56.160 79.725 56.945 ;
        RECT 79.755 56.075 81.105 56.985 ;
        RECT 81.135 56.075 82.485 56.985 ;
        RECT 82.515 56.160 82.945 56.945 ;
        RECT 82.975 56.075 84.325 56.985 ;
        RECT 84.355 56.075 85.705 56.985 ;
        RECT 85.725 56.075 87.555 56.885 ;
        RECT 103.415 56.250 103.585 56.440 ;
        RECT 104.795 56.250 104.965 56.440 ;
        RECT 111.225 56.250 111.395 56.440 ;
        RECT 111.695 56.250 111.865 56.440 ;
        RECT 115.385 56.295 115.545 56.405 ;
        RECT 116.755 56.250 116.925 56.440 ;
        RECT 122.275 56.250 122.445 56.440 ;
        RECT 127.795 56.250 127.965 56.440 ;
        RECT 129.635 56.250 129.805 56.440 ;
        RECT 135.155 56.250 135.325 56.440 ;
        RECT 138.835 56.250 139.005 56.440 ;
        RECT 141.135 56.250 141.305 56.440 ;
        RECT 77.585 55.885 77.755 56.075 ;
        RECT 79.885 55.885 80.055 56.075 ;
        RECT 81.265 55.885 81.435 56.075 ;
        RECT 83.105 55.885 83.275 56.075 ;
        RECT 84.485 55.885 84.655 56.075 ;
        RECT 85.865 55.885 86.035 56.075 ;
        RECT 103.275 55.440 104.645 56.250 ;
        RECT 104.655 55.440 110.165 56.250 ;
        RECT 110.175 55.470 111.545 56.250 ;
        RECT 111.555 55.440 115.225 56.250 ;
        RECT 116.165 55.380 116.595 56.165 ;
        RECT 116.615 55.440 122.125 56.250 ;
        RECT 122.135 55.440 127.645 56.250 ;
        RECT 127.655 55.440 129.025 56.250 ;
        RECT 129.045 55.380 129.475 56.165 ;
        RECT 129.495 55.440 135.005 56.250 ;
        RECT 135.015 55.440 138.685 56.250 ;
        RECT 138.695 55.440 140.065 56.250 ;
        RECT 140.075 55.440 141.445 56.250 ;
      LAYER nwell ;
        RECT 103.080 52.220 141.640 55.050 ;
      LAYER pwell ;
        RECT 63.240 49.860 82.430 52.170 ;
        RECT 103.275 51.020 104.645 51.830 ;
        RECT 104.655 51.020 110.165 51.830 ;
        RECT 110.175 51.020 115.685 51.830 ;
        RECT 116.165 51.105 116.595 51.890 ;
        RECT 116.615 51.020 122.125 51.830 ;
        RECT 122.135 51.020 127.645 51.830 ;
        RECT 127.655 51.020 133.165 51.830 ;
        RECT 133.175 51.020 138.685 51.830 ;
        RECT 138.695 51.020 140.065 51.830 ;
        RECT 140.075 51.020 141.445 51.830 ;
        RECT 103.415 50.810 103.585 51.020 ;
        RECT 104.795 50.810 104.965 51.020 ;
        RECT 106.630 50.860 106.750 50.970 ;
        RECT 107.095 50.810 107.265 51.000 ;
        RECT 110.315 50.810 110.485 51.020 ;
        RECT 115.835 50.970 116.005 51.000 ;
        RECT 115.830 50.860 116.005 50.970 ;
        RECT 115.835 50.810 116.005 50.860 ;
        RECT 116.755 50.830 116.925 51.020 ;
        RECT 121.355 50.810 121.525 51.000 ;
        RECT 122.275 50.830 122.445 51.020 ;
        RECT 126.875 50.810 127.045 51.000 ;
        RECT 127.795 50.830 127.965 51.020 ;
        RECT 128.710 50.860 128.830 50.970 ;
        RECT 129.635 50.810 129.805 51.000 ;
        RECT 133.315 50.830 133.485 51.020 ;
        RECT 135.155 50.810 135.325 51.000 ;
        RECT 138.835 50.810 139.005 51.020 ;
        RECT 141.135 50.810 141.305 51.020 ;
        RECT 103.275 50.000 104.645 50.810 ;
        RECT 104.655 50.000 106.485 50.810 ;
        RECT 106.995 49.900 110.165 50.810 ;
        RECT 110.175 50.000 115.685 50.810 ;
        RECT 115.695 50.000 121.205 50.810 ;
        RECT 121.215 50.000 126.725 50.810 ;
        RECT 126.735 50.000 128.565 50.810 ;
        RECT 129.045 49.940 129.475 50.725 ;
        RECT 129.495 50.000 135.005 50.810 ;
        RECT 135.015 50.000 138.685 50.810 ;
        RECT 138.695 50.000 140.065 50.810 ;
        RECT 140.075 50.000 141.445 50.810 ;
      LAYER nwell ;
        RECT 61.570 47.540 84.940 49.850 ;
      LAYER pwell ;
        RECT 63.250 44.510 82.440 46.820 ;
      LAYER nwell ;
        RECT 103.080 46.780 141.640 49.610 ;
      LAYER pwell ;
        RECT 103.275 45.580 104.645 46.390 ;
        RECT 104.655 45.580 106.485 46.390 ;
        RECT 106.995 46.260 108.345 46.490 ;
        RECT 109.880 46.260 110.790 46.480 ;
        RECT 106.995 45.580 114.305 46.260 ;
        RECT 114.315 45.580 116.145 46.390 ;
        RECT 116.165 45.665 116.595 46.450 ;
        RECT 116.615 45.580 122.125 46.390 ;
        RECT 122.135 45.580 127.645 46.390 ;
        RECT 127.655 45.580 133.165 46.390 ;
        RECT 133.175 45.580 138.685 46.390 ;
        RECT 138.695 45.580 140.065 46.390 ;
        RECT 140.075 45.580 141.445 46.390 ;
        RECT 103.415 45.370 103.585 45.580 ;
        RECT 104.795 45.530 104.965 45.580 ;
        RECT 106.635 45.530 106.805 45.560 ;
        RECT 104.790 45.420 104.965 45.530 ;
        RECT 106.630 45.420 106.805 45.530 ;
        RECT 104.795 45.390 104.965 45.420 ;
        RECT 106.635 45.370 106.805 45.420 ;
        RECT 113.995 45.370 114.165 45.580 ;
        RECT 114.455 45.370 114.625 45.580 ;
        RECT 116.755 45.390 116.925 45.580 ;
        RECT 119.975 45.370 120.145 45.560 ;
        RECT 122.275 45.390 122.445 45.580 ;
        RECT 125.495 45.370 125.665 45.560 ;
        RECT 127.795 45.390 127.965 45.580 ;
        RECT 129.635 45.370 129.805 45.560 ;
        RECT 133.315 45.390 133.485 45.580 ;
        RECT 135.155 45.370 135.325 45.560 ;
        RECT 138.835 45.370 139.005 45.580 ;
        RECT 141.135 45.370 141.305 45.580 ;
        RECT 103.275 44.560 104.645 45.370 ;
      LAYER nwell ;
        RECT 61.580 42.190 84.950 44.500 ;
      LAYER pwell ;
        RECT 105.115 44.460 106.930 45.370 ;
        RECT 106.995 44.690 114.305 45.370 ;
        RECT 106.995 44.460 108.345 44.690 ;
        RECT 109.880 44.470 110.790 44.690 ;
        RECT 114.315 44.560 119.825 45.370 ;
        RECT 119.835 44.560 125.345 45.370 ;
        RECT 125.355 44.560 129.025 45.370 ;
        RECT 129.045 44.500 129.475 45.285 ;
        RECT 129.495 44.560 135.005 45.370 ;
        RECT 135.015 44.560 138.685 45.370 ;
        RECT 138.695 44.560 140.065 45.370 ;
        RECT 140.075 44.560 141.445 45.370 ;
        RECT 63.220 39.160 82.410 41.470 ;
      LAYER nwell ;
        RECT 103.080 41.340 141.640 44.170 ;
      LAYER pwell ;
        RECT 103.275 40.140 104.645 40.950 ;
        RECT 104.655 40.140 108.325 40.950 ;
        RECT 110.165 40.820 111.085 41.050 ;
        RECT 108.795 40.140 111.085 40.820 ;
        RECT 111.095 40.140 112.925 40.820 ;
        RECT 112.935 40.140 114.285 41.050 ;
        RECT 114.315 40.140 116.145 40.950 ;
        RECT 116.165 40.225 116.595 41.010 ;
        RECT 116.615 40.140 122.125 40.950 ;
        RECT 122.135 40.140 127.645 40.950 ;
        RECT 127.655 40.140 133.165 40.950 ;
        RECT 133.175 40.140 138.685 40.950 ;
        RECT 138.695 40.140 140.065 40.950 ;
        RECT 140.075 40.140 141.445 40.950 ;
        RECT 103.415 39.930 103.585 40.140 ;
        RECT 104.795 39.930 104.965 40.140 ;
        RECT 108.470 39.980 108.590 40.090 ;
        RECT 108.935 39.950 109.105 40.140 ;
        RECT 110.315 39.930 110.485 40.120 ;
        RECT 111.235 39.950 111.405 40.140 ;
        RECT 113.080 39.950 113.250 40.140 ;
        RECT 114.455 39.950 114.625 40.140 ;
        RECT 115.835 39.930 116.005 40.120 ;
        RECT 116.755 39.950 116.925 40.140 ;
        RECT 121.355 39.930 121.525 40.120 ;
        RECT 122.275 39.950 122.445 40.140 ;
        RECT 126.875 39.930 127.045 40.120 ;
        RECT 127.795 39.950 127.965 40.140 ;
        RECT 128.710 39.980 128.830 40.090 ;
        RECT 129.635 39.930 129.805 40.120 ;
        RECT 133.315 39.950 133.485 40.140 ;
        RECT 135.155 39.930 135.325 40.120 ;
        RECT 138.835 39.930 139.005 40.140 ;
        RECT 141.135 39.930 141.305 40.140 ;
      LAYER nwell ;
        RECT 61.550 36.840 84.920 39.150 ;
      LAYER pwell ;
        RECT 103.275 39.120 104.645 39.930 ;
        RECT 104.655 39.120 110.165 39.930 ;
        RECT 110.175 39.120 115.685 39.930 ;
        RECT 115.695 39.120 121.205 39.930 ;
        RECT 121.215 39.120 126.725 39.930 ;
        RECT 126.735 39.120 128.565 39.930 ;
        RECT 129.045 39.060 129.475 39.845 ;
        RECT 129.495 39.120 135.005 39.930 ;
        RECT 135.015 39.120 138.685 39.930 ;
        RECT 138.695 39.120 140.065 39.930 ;
        RECT 140.075 39.120 141.445 39.930 ;
        RECT 63.260 33.880 82.450 36.190 ;
      LAYER nwell ;
        RECT 103.080 35.900 141.640 38.730 ;
      LAYER pwell ;
        RECT 103.275 34.700 104.645 35.510 ;
        RECT 104.655 34.700 106.485 35.510 ;
        RECT 106.580 34.700 115.685 35.380 ;
        RECT 116.165 34.785 116.595 35.570 ;
        RECT 116.615 34.700 118.445 35.510 ;
        RECT 119.000 34.700 128.105 35.380 ;
        RECT 128.115 34.700 133.625 35.510 ;
        RECT 133.635 34.700 139.145 35.510 ;
        RECT 140.075 34.700 141.445 35.510 ;
        RECT 103.415 34.490 103.585 34.700 ;
        RECT 104.795 34.490 104.965 34.700 ;
        RECT 110.315 34.490 110.485 34.680 ;
        RECT 115.375 34.510 115.545 34.700 ;
        RECT 115.830 34.645 115.950 34.650 ;
        RECT 115.830 34.540 116.005 34.645 ;
        RECT 115.845 34.535 116.005 34.540 ;
        RECT 116.755 34.490 116.925 34.700 ;
        RECT 118.590 34.540 118.710 34.650 ;
        RECT 126.415 34.490 126.585 34.680 ;
        RECT 127.795 34.490 127.965 34.700 ;
        RECT 128.255 34.510 128.425 34.700 ;
        RECT 129.635 34.490 129.805 34.680 ;
        RECT 132.855 34.490 133.025 34.680 ;
        RECT 133.775 34.510 133.945 34.700 ;
        RECT 136.535 34.490 136.705 34.680 ;
        RECT 136.995 34.490 137.165 34.680 ;
        RECT 139.305 34.545 139.465 34.655 ;
        RECT 139.750 34.540 139.870 34.650 ;
        RECT 141.135 34.490 141.305 34.700 ;
      LAYER nwell ;
        RECT 61.590 31.560 84.960 33.870 ;
      LAYER pwell ;
        RECT 103.275 33.680 104.645 34.490 ;
        RECT 104.655 33.680 110.165 34.490 ;
        RECT 110.175 33.680 115.685 34.490 ;
        RECT 116.615 33.810 119.365 34.490 ;
        RECT 118.435 33.580 119.365 33.810 ;
        RECT 119.415 33.810 126.725 34.490 ;
        RECT 119.415 33.580 120.765 33.810 ;
        RECT 122.300 33.590 123.210 33.810 ;
        RECT 126.735 33.710 128.105 34.490 ;
        RECT 129.045 33.620 129.475 34.405 ;
        RECT 129.495 33.810 132.705 34.490 ;
        RECT 132.715 33.810 135.465 34.490 ;
        RECT 131.570 33.580 132.705 33.810 ;
        RECT 134.535 33.580 135.465 33.810 ;
        RECT 135.475 33.710 136.845 34.490 ;
        RECT 136.855 33.680 139.605 34.490 ;
        RECT 140.075 33.680 141.445 34.490 ;
      LAYER nwell ;
        RECT 103.080 30.460 141.640 33.290 ;
      LAYER pwell ;
        RECT 103.275 29.260 104.645 30.070 ;
        RECT 104.655 29.260 107.405 30.070 ;
        RECT 107.415 29.260 108.765 30.170 ;
        RECT 112.310 29.940 113.220 30.160 ;
        RECT 114.755 29.940 116.105 30.170 ;
        RECT 108.795 29.260 116.105 29.940 ;
        RECT 116.165 29.345 116.595 30.130 ;
        RECT 116.615 29.260 118.445 30.070 ;
        RECT 119.055 29.260 122.505 30.170 ;
        RECT 125.340 29.940 126.265 30.170 ;
        RECT 122.595 29.260 126.265 29.940 ;
        RECT 126.275 29.260 135.380 29.940 ;
        RECT 135.475 29.260 139.145 30.070 ;
        RECT 140.075 29.260 141.445 30.070 ;
        RECT 103.415 29.050 103.585 29.260 ;
        RECT 104.795 29.070 104.965 29.260 ;
        RECT 105.710 29.050 105.880 29.240 ;
        RECT 106.175 29.050 106.345 29.240 ;
        RECT 107.560 29.070 107.730 29.260 ;
        RECT 108.935 29.070 109.105 29.260 ;
        RECT 116.295 29.050 116.465 29.240 ;
        RECT 116.755 29.050 116.925 29.260 ;
        RECT 118.600 29.210 118.770 29.240 ;
        RECT 118.590 29.100 118.770 29.210 ;
        RECT 118.600 29.050 118.770 29.100 ;
        RECT 121.815 29.050 121.985 29.240 ;
        RECT 122.275 29.070 122.445 29.260 ;
        RECT 125.950 29.070 126.120 29.260 ;
        RECT 126.415 29.070 126.585 29.260 ;
        RECT 129.635 29.050 129.805 29.240 ;
        RECT 131.015 29.050 131.185 29.240 ;
        RECT 135.615 29.070 135.785 29.260 ;
        RECT 138.375 29.050 138.545 29.240 ;
        RECT 139.305 29.105 139.465 29.215 ;
        RECT 141.135 29.050 141.305 29.260 ;
        RECT 103.275 28.240 104.645 29.050 ;
        RECT 104.675 28.140 106.025 29.050 ;
        RECT 106.035 28.370 113.345 29.050 ;
        RECT 109.550 28.150 110.460 28.370 ;
        RECT 111.995 28.140 113.345 28.370 ;
        RECT 113.395 28.140 116.565 29.050 ;
        RECT 116.615 28.240 118.445 29.050 ;
        RECT 118.455 28.140 121.375 29.050 ;
        RECT 121.675 28.370 128.985 29.050 ;
        RECT 125.190 28.150 126.100 28.370 ;
        RECT 127.635 28.140 128.985 28.370 ;
        RECT 129.045 28.180 129.475 28.965 ;
        RECT 129.495 28.240 130.865 29.050 ;
        RECT 130.875 28.370 138.185 29.050 ;
        RECT 134.390 28.150 135.300 28.370 ;
        RECT 136.835 28.140 138.185 28.370 ;
        RECT 138.235 28.240 140.065 29.050 ;
        RECT 140.075 28.240 141.445 29.050 ;
      LAYER nwell ;
        RECT 103.080 25.020 141.640 27.850 ;
      LAYER pwell ;
        RECT 103.275 23.820 104.645 24.630 ;
        RECT 104.655 23.820 107.405 24.630 ;
        RECT 110.930 24.500 111.840 24.720 ;
        RECT 113.375 24.500 114.725 24.730 ;
        RECT 107.415 23.820 114.725 24.500 ;
        RECT 114.775 23.820 116.145 24.630 ;
        RECT 116.165 23.905 116.595 24.690 ;
        RECT 117.755 24.640 118.705 24.730 ;
        RECT 116.775 23.820 118.705 24.640 ;
        RECT 120.285 24.500 121.205 24.730 ;
        RECT 118.915 23.820 121.205 24.500 ;
        RECT 121.215 24.500 122.135 24.730 ;
        RECT 127.030 24.500 127.940 24.720 ;
        RECT 129.475 24.500 130.825 24.730 ;
        RECT 134.390 24.500 135.300 24.720 ;
        RECT 136.835 24.500 138.185 24.730 ;
        RECT 121.215 23.820 123.505 24.500 ;
        RECT 123.515 23.820 130.825 24.500 ;
        RECT 130.875 23.820 138.185 24.500 ;
        RECT 138.235 23.820 140.065 24.630 ;
        RECT 140.075 23.820 141.445 24.630 ;
        RECT 103.415 23.610 103.585 23.820 ;
        RECT 104.795 23.610 104.965 23.820 ;
        RECT 107.555 23.630 107.725 23.820 ;
        RECT 108.475 23.610 108.645 23.800 ;
        RECT 109.855 23.610 110.025 23.800 ;
        RECT 114.915 23.630 115.085 23.820 ;
        RECT 116.775 23.800 116.925 23.820 ;
        RECT 115.375 23.630 115.545 23.800 ;
        RECT 115.845 23.655 116.005 23.765 ;
        RECT 116.755 23.630 116.925 23.800 ;
        RECT 115.375 23.610 115.525 23.630 ;
        RECT 103.275 22.800 104.645 23.610 ;
        RECT 104.655 22.800 108.325 23.610 ;
        RECT 108.335 22.800 109.705 23.610 ;
        RECT 109.795 22.700 113.245 23.610 ;
        RECT 113.595 22.790 115.525 23.610 ;
        RECT 116.775 23.610 116.925 23.630 ;
        RECT 119.055 23.610 119.225 23.820 ;
        RECT 123.195 23.630 123.365 23.820 ;
        RECT 123.655 23.630 123.825 23.820 ;
        RECT 124.585 23.655 124.745 23.765 ;
        RECT 128.255 23.610 128.425 23.800 ;
        RECT 128.710 23.660 128.830 23.770 ;
        RECT 131.015 23.630 131.185 23.820 ;
        RECT 132.395 23.610 132.565 23.800 ;
        RECT 135.610 23.610 135.780 23.800 ;
        RECT 138.375 23.630 138.545 23.820 ;
        RECT 138.835 23.610 139.005 23.800 ;
        RECT 139.305 23.655 139.465 23.765 ;
        RECT 141.135 23.610 141.305 23.820 ;
        RECT 116.775 22.790 118.705 23.610 ;
        RECT 118.915 22.800 124.425 23.610 ;
        RECT 125.355 22.930 128.565 23.610 ;
        RECT 113.595 22.700 114.545 22.790 ;
        RECT 117.755 22.700 118.705 22.790 ;
        RECT 125.355 22.700 126.490 22.930 ;
        RECT 129.045 22.740 129.475 23.525 ;
        RECT 129.495 22.930 132.705 23.610 ;
        RECT 129.495 22.700 130.630 22.930 ;
        RECT 133.005 22.700 135.925 23.610 ;
        RECT 135.935 22.700 139.105 23.610 ;
        RECT 140.075 22.800 141.445 23.610 ;
      LAYER nwell ;
        RECT 103.080 19.580 141.640 22.410 ;
      LAYER pwell ;
        RECT 103.275 18.380 104.645 19.190 ;
        RECT 104.655 18.380 106.025 19.160 ;
        RECT 106.495 18.380 107.865 19.160 ;
        RECT 107.875 18.380 110.625 19.190 ;
        RECT 111.095 18.380 112.465 19.160 ;
        RECT 112.475 18.380 116.145 19.190 ;
        RECT 116.165 18.465 116.595 19.250 ;
        RECT 116.615 18.380 117.985 19.160 ;
        RECT 117.995 18.380 119.825 19.190 ;
        RECT 120.295 18.380 121.665 19.160 ;
        RECT 121.675 18.380 124.425 19.190 ;
        RECT 124.895 18.380 126.265 19.160 ;
        RECT 126.275 18.380 129.025 19.190 ;
        RECT 129.045 18.465 129.475 19.250 ;
        RECT 129.495 18.380 130.865 19.160 ;
        RECT 130.875 18.380 133.625 19.190 ;
        RECT 134.095 18.380 135.465 19.160 ;
        RECT 135.475 18.380 137.305 19.190 ;
        RECT 137.315 18.380 138.685 19.160 ;
        RECT 138.695 18.380 140.065 19.160 ;
        RECT 140.075 18.380 141.445 19.190 ;
        RECT 103.415 18.190 103.585 18.380 ;
        RECT 105.705 18.190 105.875 18.380 ;
        RECT 106.170 18.220 106.290 18.330 ;
        RECT 107.545 18.190 107.715 18.380 ;
        RECT 108.015 18.190 108.185 18.380 ;
        RECT 110.770 18.220 110.890 18.330 ;
        RECT 112.145 18.190 112.315 18.380 ;
        RECT 112.615 18.190 112.785 18.380 ;
        RECT 117.665 18.190 117.835 18.380 ;
        RECT 118.135 18.190 118.305 18.380 ;
        RECT 119.970 18.220 120.090 18.330 ;
        RECT 121.345 18.190 121.515 18.380 ;
        RECT 121.815 18.190 121.985 18.380 ;
        RECT 124.570 18.220 124.690 18.330 ;
        RECT 125.945 18.190 126.115 18.380 ;
        RECT 126.415 18.190 126.585 18.380 ;
        RECT 130.545 18.190 130.715 18.380 ;
        RECT 131.015 18.190 131.185 18.380 ;
        RECT 133.770 18.220 133.890 18.330 ;
        RECT 135.145 18.190 135.315 18.380 ;
        RECT 135.615 18.190 135.785 18.380 ;
        RECT 137.465 18.190 137.635 18.380 ;
        RECT 139.745 18.190 139.915 18.380 ;
        RECT 141.135 18.190 141.305 18.380 ;
      LAYER li1 ;
        RECT 92.875 165.025 101.155 165.195 ;
        RECT 92.960 163.935 94.630 165.025 ;
        RECT 92.960 163.245 93.710 163.765 ;
        RECT 93.880 163.415 94.630 163.935 ;
        RECT 94.840 163.885 95.070 165.025 ;
        RECT 95.240 163.875 95.570 164.855 ;
        RECT 95.740 163.885 95.950 165.025 ;
        RECT 96.220 163.885 96.450 165.025 ;
        RECT 96.620 163.875 96.950 164.855 ;
        RECT 97.120 163.885 97.330 165.025 ;
        RECT 97.600 163.885 97.830 165.025 ;
        RECT 98.000 163.875 98.330 164.855 ;
        RECT 98.500 163.885 98.710 165.025 ;
        RECT 95.320 163.760 95.570 163.875 ;
        RECT 94.820 163.700 95.150 163.715 ;
        RECT 94.815 163.480 95.150 163.700 ;
        RECT 94.820 163.465 95.150 163.480 ;
        RECT 95.320 163.460 95.595 163.760 ;
        RECT 96.200 163.465 96.530 163.715 ;
        RECT 92.960 162.475 94.630 163.245 ;
        RECT 94.840 162.475 95.070 163.295 ;
        RECT 95.320 163.275 95.570 163.460 ;
        RECT 95.240 162.645 95.570 163.275 ;
        RECT 95.740 162.475 95.950 163.295 ;
        RECT 96.220 162.475 96.450 163.295 ;
        RECT 96.700 163.275 96.950 163.875 ;
        RECT 97.580 163.710 97.910 163.715 ;
        RECT 97.565 163.470 97.910 163.710 ;
        RECT 97.580 163.465 97.910 163.470 ;
        RECT 98.080 163.710 98.330 163.875 ;
        RECT 98.940 163.860 99.230 165.025 ;
        RECT 99.400 163.935 101.070 165.025 ;
        RECT 98.080 163.470 98.425 163.710 ;
        RECT 96.620 162.645 96.950 163.275 ;
        RECT 97.120 162.475 97.330 163.295 ;
        RECT 97.600 162.475 97.830 163.295 ;
        RECT 98.080 163.275 98.330 163.470 ;
        RECT 98.000 162.645 98.330 163.275 ;
        RECT 98.500 162.475 98.710 163.295 ;
        RECT 99.400 163.245 100.150 163.765 ;
        RECT 100.320 163.415 101.070 163.935 ;
        RECT 98.940 162.475 99.230 163.200 ;
        RECT 99.400 162.475 101.070 163.245 ;
        RECT 92.875 162.305 103.455 162.475 ;
        RECT 92.960 161.845 93.520 162.135 ;
        RECT 93.690 161.845 93.940 162.305 ;
        RECT 92.960 161.790 93.210 161.845 ;
        RECT 92.955 160.650 93.210 161.790 ;
        RECT 94.560 161.675 94.890 162.035 ;
        RECT 93.500 161.485 94.890 161.675 ;
        RECT 95.280 161.615 95.520 162.135 ;
        RECT 95.690 161.810 96.085 162.305 ;
        RECT 96.650 161.975 96.820 162.120 ;
        RECT 96.445 161.780 96.820 161.975 ;
        RECT 93.500 161.395 93.670 161.485 ;
        RECT 93.380 161.065 93.670 161.395 ;
        RECT 93.840 161.065 94.180 161.315 ;
        RECT 94.400 161.065 95.075 161.315 ;
        RECT 92.960 160.475 93.210 160.650 ;
        RECT 93.500 160.815 93.670 161.065 ;
        RECT 93.500 160.645 94.440 160.815 ;
        RECT 94.810 160.705 95.075 161.065 ;
        RECT 95.280 160.810 95.455 161.615 ;
        RECT 96.445 161.445 96.615 161.780 ;
        RECT 97.100 161.735 97.340 162.110 ;
        RECT 97.510 161.800 97.845 162.305 ;
        RECT 97.100 161.585 97.320 161.735 ;
        RECT 95.630 161.085 96.615 161.445 ;
        RECT 96.785 161.255 97.320 161.585 ;
        RECT 95.630 161.065 96.915 161.085 ;
        RECT 96.055 160.915 96.915 161.065 ;
        RECT 92.960 159.925 93.420 160.475 ;
        RECT 93.610 159.755 93.940 160.475 ;
        RECT 94.140 160.095 94.440 160.645 ;
        RECT 94.610 159.755 94.890 160.425 ;
        RECT 95.280 160.025 95.585 160.810 ;
        RECT 95.760 160.435 96.455 160.745 ;
        RECT 95.765 159.755 96.450 160.225 ;
        RECT 96.630 159.970 96.915 160.915 ;
        RECT 97.085 160.605 97.320 161.255 ;
        RECT 97.490 160.775 97.790 161.625 ;
        RECT 98.040 161.615 98.280 162.135 ;
        RECT 98.450 161.810 98.845 162.305 ;
        RECT 99.410 161.975 99.580 162.120 ;
        RECT 99.205 161.780 99.580 161.975 ;
        RECT 98.040 160.810 98.215 161.615 ;
        RECT 99.205 161.445 99.375 161.780 ;
        RECT 99.860 161.735 100.100 162.110 ;
        RECT 100.270 161.800 100.605 162.305 ;
        RECT 99.860 161.585 100.080 161.735 ;
        RECT 98.390 161.085 99.375 161.445 ;
        RECT 99.545 161.255 100.080 161.585 ;
        RECT 98.390 161.065 99.675 161.085 ;
        RECT 98.815 160.915 99.675 161.065 ;
        RECT 97.085 160.375 97.760 160.605 ;
        RECT 97.090 159.755 97.420 160.205 ;
        RECT 97.590 159.945 97.760 160.375 ;
        RECT 98.040 160.025 98.345 160.810 ;
        RECT 98.520 160.435 99.215 160.745 ;
        RECT 98.525 159.755 99.210 160.225 ;
        RECT 99.390 159.970 99.675 160.915 ;
        RECT 99.845 160.605 100.080 161.255 ;
        RECT 100.250 160.775 100.550 161.625 ;
        RECT 100.780 161.580 101.070 162.305 ;
        RECT 101.240 161.845 101.800 162.135 ;
        RECT 101.970 161.845 102.220 162.305 ;
        RECT 99.845 160.375 100.520 160.605 ;
        RECT 99.850 159.755 100.180 160.205 ;
        RECT 100.350 159.945 100.520 160.375 ;
        RECT 100.780 159.755 101.070 160.920 ;
        RECT 101.240 160.475 101.490 161.845 ;
        RECT 102.840 161.675 103.170 162.035 ;
        RECT 101.780 161.485 103.170 161.675 ;
        RECT 101.780 161.395 101.950 161.485 ;
        RECT 101.660 161.065 101.950 161.395 ;
        RECT 102.120 161.065 102.460 161.315 ;
        RECT 102.680 161.065 103.355 161.315 ;
        RECT 101.780 160.815 101.950 161.065 ;
        RECT 102.735 160.990 103.355 161.065 ;
        RECT 101.780 160.645 102.720 160.815 ;
        RECT 103.090 160.705 103.355 160.990 ;
        RECT 101.240 159.925 101.700 160.475 ;
        RECT 101.890 159.755 102.220 160.475 ;
        RECT 102.420 160.095 102.720 160.645 ;
        RECT 102.890 159.755 103.170 160.425 ;
        RECT 92.875 159.585 103.455 159.755 ;
        RECT 92.960 158.495 94.630 159.585 ;
        RECT 92.960 157.805 93.710 158.325 ;
        RECT 93.880 157.975 94.630 158.495 ;
        RECT 94.800 158.420 95.090 159.585 ;
        RECT 95.300 158.445 95.530 159.585 ;
        RECT 95.700 158.435 96.030 159.415 ;
        RECT 96.200 158.445 96.410 159.585 ;
        RECT 96.680 158.445 96.910 159.585 ;
        RECT 97.080 158.435 97.410 159.415 ;
        RECT 97.580 158.445 97.790 159.585 ;
        RECT 95.280 158.025 95.610 158.275 ;
        RECT 92.960 157.035 94.630 157.805 ;
        RECT 94.800 157.035 95.090 157.760 ;
        RECT 95.300 157.035 95.530 157.855 ;
        RECT 95.780 157.835 96.030 158.435 ;
        RECT 96.660 158.025 96.990 158.275 ;
        RECT 95.700 157.205 96.030 157.835 ;
        RECT 96.200 157.035 96.410 157.855 ;
        RECT 96.680 157.035 96.910 157.855 ;
        RECT 97.160 157.835 97.410 158.435 ;
        RECT 98.020 158.420 98.310 159.585 ;
        RECT 98.520 158.445 98.750 159.585 ;
        RECT 98.920 158.435 99.250 159.415 ;
        RECT 99.420 158.445 99.630 159.585 ;
        RECT 99.900 158.445 100.130 159.585 ;
        RECT 100.300 158.435 100.630 159.415 ;
        RECT 100.800 158.445 101.010 159.585 ;
        RECT 101.240 158.495 102.910 159.585 ;
        RECT 98.500 158.025 98.830 158.275 ;
        RECT 97.080 157.205 97.410 157.835 ;
        RECT 97.580 157.035 97.790 157.855 ;
        RECT 98.020 157.035 98.310 157.760 ;
        RECT 98.520 157.035 98.750 157.855 ;
        RECT 99.000 157.835 99.250 158.435 ;
        RECT 99.880 158.270 100.210 158.275 ;
        RECT 99.855 158.030 100.210 158.270 ;
        RECT 99.880 158.025 100.210 158.030 ;
        RECT 98.920 157.205 99.250 157.835 ;
        RECT 99.420 157.035 99.630 157.855 ;
        RECT 99.900 157.035 100.130 157.855 ;
        RECT 100.380 157.835 100.630 158.435 ;
        RECT 100.300 157.205 100.630 157.835 ;
        RECT 100.800 157.035 101.010 157.855 ;
        RECT 101.240 157.805 101.990 158.325 ;
        RECT 102.160 157.975 102.910 158.495 ;
        RECT 101.240 157.035 102.910 157.805 ;
        RECT 92.875 156.865 102.995 157.035 ;
        RECT 69.265 152.000 71.215 152.170 ;
        RECT 75.015 152.050 95.005 152.370 ;
        RECT 63.975 151.810 65.925 151.980 ;
        RECT 63.975 151.540 64.145 151.810 ;
        RECT 61.335 150.150 62.485 150.640 ;
        RECT 61.335 149.470 63.595 150.150 ;
        RECT 61.335 149.300 63.605 149.470 ;
        RECT 61.335 130.810 61.825 149.300 ;
        RECT 62.455 148.790 62.805 148.960 ;
        RECT 62.225 140.580 62.395 148.620 ;
        RECT 62.865 140.580 63.035 148.620 ;
        RECT 62.455 140.240 62.805 140.410 ;
        RECT 62.455 139.700 62.805 139.870 ;
        RECT 62.225 131.490 62.395 139.530 ;
        RECT 62.865 131.490 63.035 139.530 ;
        RECT 62.455 131.150 62.805 131.320 ;
        RECT 63.435 130.810 63.605 149.300 ;
        RECT 61.335 130.650 63.605 130.810 ;
        RECT 61.655 130.640 63.605 130.650 ;
        RECT 63.785 129.810 64.145 151.540 ;
        RECT 64.775 151.300 65.125 151.470 ;
        RECT 64.545 141.045 64.715 151.085 ;
        RECT 65.185 141.045 65.355 151.085 ;
        RECT 64.775 140.660 65.125 140.830 ;
        RECT 64.775 140.120 65.125 140.290 ;
        RECT 64.545 129.865 64.715 139.905 ;
        RECT 65.185 129.865 65.355 139.905 ;
        RECT 63.105 129.760 64.145 129.810 ;
        RECT 62.835 129.140 64.145 129.760 ;
        RECT 64.775 129.480 65.125 129.650 ;
        RECT 65.755 129.140 65.925 151.810 ;
        RECT 69.265 151.730 69.435 152.000 ;
        RECT 66.625 150.340 67.775 150.830 ;
        RECT 66.625 149.660 68.885 150.340 ;
        RECT 66.625 149.490 68.895 149.660 ;
        RECT 66.625 131.000 67.115 149.490 ;
        RECT 67.745 148.980 68.095 149.150 ;
        RECT 67.515 140.770 67.685 148.810 ;
        RECT 68.155 140.770 68.325 148.810 ;
        RECT 67.745 140.430 68.095 140.600 ;
        RECT 67.745 139.890 68.095 140.060 ;
        RECT 67.515 131.680 67.685 139.720 ;
        RECT 68.155 131.680 68.325 139.720 ;
        RECT 67.745 131.340 68.095 131.510 ;
        RECT 68.725 131.000 68.895 149.490 ;
        RECT 66.625 130.840 68.895 131.000 ;
        RECT 66.945 130.830 68.895 130.840 ;
        RECT 69.075 130.000 69.435 151.730 ;
        RECT 70.065 151.490 70.415 151.660 ;
        RECT 69.835 141.235 70.005 151.275 ;
        RECT 70.475 141.235 70.645 151.275 ;
        RECT 70.065 140.850 70.415 141.020 ;
        RECT 70.065 140.310 70.415 140.480 ;
        RECT 69.835 130.055 70.005 140.095 ;
        RECT 70.475 130.055 70.645 140.095 ;
        RECT 68.395 129.950 69.435 130.000 ;
        RECT 62.835 128.970 65.925 129.140 ;
        RECT 68.125 129.330 69.435 129.950 ;
        RECT 70.065 129.670 70.415 129.840 ;
        RECT 71.045 129.330 71.215 152.000 ;
        RECT 75.005 151.880 95.005 152.050 ;
        RECT 73.265 150.860 74.125 150.870 ;
        RECT 73.165 150.600 74.125 150.860 ;
        RECT 73.165 149.920 74.175 150.600 ;
        RECT 75.005 150.270 75.175 151.880 ;
        RECT 75.855 151.310 83.895 151.480 ;
        RECT 84.945 151.310 92.985 151.480 ;
        RECT 75.515 150.900 75.685 151.250 ;
        RECT 84.065 150.900 84.235 151.250 ;
        RECT 84.605 150.900 84.775 151.250 ;
        RECT 93.155 150.900 93.325 151.250 ;
        RECT 93.665 151.220 95.005 151.880 ;
        RECT 108.030 151.645 111.700 154.055 ;
        RECT 108.030 151.475 111.710 151.645 ;
        RECT 75.855 150.670 83.895 150.840 ;
        RECT 84.945 150.670 92.985 150.840 ;
        RECT 93.665 150.270 94.515 151.220 ;
        RECT 75.005 150.110 94.515 150.270 ;
        RECT 75.005 150.100 93.835 150.110 ;
        RECT 73.165 149.730 95.905 149.920 ;
        RECT 73.165 149.560 96.345 149.730 ;
        RECT 73.165 147.950 73.505 149.560 ;
        RECT 74.230 148.990 84.270 149.160 ;
        RECT 85.410 148.990 95.450 149.160 ;
        RECT 73.845 148.580 74.015 148.930 ;
        RECT 84.485 148.580 84.655 148.930 ;
        RECT 85.025 148.580 85.195 148.930 ;
        RECT 95.665 148.580 95.835 148.930 ;
        RECT 74.230 148.350 84.270 148.520 ;
        RECT 85.410 148.350 95.450 148.520 ;
        RECT 96.175 147.950 96.345 149.560 ;
        RECT 73.165 147.790 96.345 147.950 ;
        RECT 73.335 147.780 96.345 147.790 ;
        RECT 103.980 147.345 105.280 147.435 ;
        RECT 103.980 147.175 107.820 147.345 ;
        RECT 75.025 146.700 95.015 147.020 ;
        RECT 75.015 146.530 95.015 146.700 ;
        RECT 73.275 145.510 74.135 145.520 ;
        RECT 73.175 145.250 74.135 145.510 ;
        RECT 73.175 144.570 74.185 145.250 ;
        RECT 75.015 144.920 75.185 146.530 ;
        RECT 75.865 145.960 83.905 146.130 ;
        RECT 84.955 145.960 92.995 146.130 ;
        RECT 75.525 145.550 75.695 145.900 ;
        RECT 84.075 145.550 84.245 145.900 ;
        RECT 84.615 145.550 84.785 145.900 ;
        RECT 93.165 145.550 93.335 145.900 ;
        RECT 93.675 145.870 95.015 146.530 ;
        RECT 75.865 145.320 83.905 145.490 ;
        RECT 84.955 145.320 92.995 145.490 ;
        RECT 93.675 144.920 94.525 145.870 ;
        RECT 75.015 144.760 94.525 144.920 ;
        RECT 75.015 144.750 93.845 144.760 ;
        RECT 73.175 144.380 95.915 144.570 ;
        RECT 73.175 144.210 96.355 144.380 ;
        RECT 73.175 142.600 73.515 144.210 ;
        RECT 74.240 143.640 84.280 143.810 ;
        RECT 85.420 143.640 95.460 143.810 ;
        RECT 73.855 143.230 74.025 143.580 ;
        RECT 84.495 143.230 84.665 143.580 ;
        RECT 85.035 143.230 85.205 143.580 ;
        RECT 95.675 143.230 95.845 143.580 ;
        RECT 74.240 143.000 84.280 143.170 ;
        RECT 85.420 143.000 95.460 143.170 ;
        RECT 96.185 142.600 96.355 144.210 ;
        RECT 73.175 142.440 96.355 142.600 ;
        RECT 73.345 142.430 96.355 142.440 ;
        RECT 74.995 141.350 94.985 141.670 ;
        RECT 74.985 141.180 94.985 141.350 ;
        RECT 73.245 140.160 74.105 140.170 ;
        RECT 73.145 139.900 74.105 140.160 ;
        RECT 73.145 139.220 74.155 139.900 ;
        RECT 74.985 139.570 75.155 141.180 ;
        RECT 75.835 140.610 83.875 140.780 ;
        RECT 84.925 140.610 92.965 140.780 ;
        RECT 75.495 140.200 75.665 140.550 ;
        RECT 84.045 140.200 84.215 140.550 ;
        RECT 84.585 140.200 84.755 140.550 ;
        RECT 93.135 140.200 93.305 140.550 ;
        RECT 93.645 140.520 94.985 141.180 ;
        RECT 75.835 139.970 83.875 140.140 ;
        RECT 84.925 139.970 92.965 140.140 ;
        RECT 93.645 139.570 94.495 140.520 ;
        RECT 74.985 139.410 94.495 139.570 ;
        RECT 103.980 140.305 105.280 147.175 ;
        RECT 105.760 144.535 107.170 146.695 ;
        RECT 105.760 140.785 107.170 142.945 ;
        RECT 107.650 140.305 107.820 147.175 ;
        RECT 108.100 144.605 108.270 151.475 ;
        RECT 108.750 148.835 110.160 150.995 ;
        RECT 108.750 145.085 110.160 147.245 ;
        RECT 110.640 144.605 111.710 151.475 ;
        RECT 108.100 144.435 111.710 144.605 ;
        RECT 110.640 142.035 111.710 144.435 ;
        RECT 103.980 140.135 107.820 140.305 ;
        RECT 108.220 141.865 111.710 142.035 ;
        RECT 74.985 139.400 93.815 139.410 ;
        RECT 73.145 139.030 95.885 139.220 ;
        RECT 73.145 138.860 96.325 139.030 ;
        RECT 73.145 137.250 73.485 138.860 ;
        RECT 74.210 138.290 84.250 138.460 ;
        RECT 85.390 138.290 95.430 138.460 ;
        RECT 73.825 137.880 73.995 138.230 ;
        RECT 84.465 137.880 84.635 138.230 ;
        RECT 85.005 137.880 85.175 138.230 ;
        RECT 95.645 137.880 95.815 138.230 ;
        RECT 74.210 137.650 84.250 137.820 ;
        RECT 85.390 137.650 95.430 137.820 ;
        RECT 96.155 137.250 96.325 138.860 ;
        RECT 73.145 137.090 96.325 137.250 ;
        RECT 73.315 137.080 96.325 137.090 ;
        RECT 103.980 137.435 105.280 140.135 ;
        RECT 103.980 137.265 107.820 137.435 ;
        RECT 75.035 136.070 95.025 136.390 ;
        RECT 75.025 135.900 95.025 136.070 ;
        RECT 73.285 134.880 74.145 134.890 ;
        RECT 73.185 134.620 74.145 134.880 ;
        RECT 73.185 133.940 74.195 134.620 ;
        RECT 75.025 134.290 75.195 135.900 ;
        RECT 75.875 135.330 83.915 135.500 ;
        RECT 84.965 135.330 93.005 135.500 ;
        RECT 75.535 134.920 75.705 135.270 ;
        RECT 84.085 134.920 84.255 135.270 ;
        RECT 84.625 134.920 84.795 135.270 ;
        RECT 93.175 134.920 93.345 135.270 ;
        RECT 93.685 135.240 95.025 135.900 ;
        RECT 75.875 134.690 83.915 134.860 ;
        RECT 84.965 134.690 93.005 134.860 ;
        RECT 93.685 134.290 94.535 135.240 ;
        RECT 75.025 134.130 94.535 134.290 ;
        RECT 75.025 134.120 93.855 134.130 ;
        RECT 73.185 133.750 95.925 133.940 ;
        RECT 73.185 133.580 96.365 133.750 ;
        RECT 73.185 131.970 73.525 133.580 ;
        RECT 74.250 133.010 84.290 133.180 ;
        RECT 85.430 133.010 95.470 133.180 ;
        RECT 73.865 132.600 74.035 132.950 ;
        RECT 84.505 132.600 84.675 132.950 ;
        RECT 85.045 132.600 85.215 132.950 ;
        RECT 95.685 132.600 95.855 132.950 ;
        RECT 74.250 132.370 84.290 132.540 ;
        RECT 85.430 132.370 95.470 132.540 ;
        RECT 96.195 131.970 96.365 133.580 ;
        RECT 73.185 131.810 96.365 131.970 ;
        RECT 73.355 131.800 96.365 131.810 ;
        RECT 75.025 130.480 95.015 130.800 ;
        RECT 68.125 129.160 71.215 129.330 ;
        RECT 75.015 130.310 95.015 130.480 ;
        RECT 73.275 129.290 74.135 129.300 ;
        RECT 68.125 129.090 71.205 129.160 ;
        RECT 68.135 128.990 71.205 129.090 ;
        RECT 73.175 129.030 74.135 129.290 ;
        RECT 62.835 128.900 65.915 128.970 ;
        RECT 62.845 128.800 65.915 128.900 ;
        RECT 73.175 128.350 74.185 129.030 ;
        RECT 75.015 128.700 75.185 130.310 ;
        RECT 75.865 129.740 83.905 129.910 ;
        RECT 84.955 129.740 92.995 129.910 ;
        RECT 75.525 129.330 75.695 129.680 ;
        RECT 84.075 129.330 84.245 129.680 ;
        RECT 84.615 129.330 84.785 129.680 ;
        RECT 93.165 129.330 93.335 129.680 ;
        RECT 93.675 129.650 95.015 130.310 ;
        RECT 103.980 130.395 105.280 137.265 ;
        RECT 105.760 134.625 107.170 136.785 ;
        RECT 105.760 130.875 107.170 133.035 ;
        RECT 107.650 130.395 107.820 137.265 ;
        RECT 108.220 134.995 108.390 141.865 ;
        RECT 108.870 139.225 110.280 141.385 ;
        RECT 108.870 135.475 110.280 137.635 ;
        RECT 110.640 134.995 111.710 141.865 ;
        RECT 108.220 134.825 111.710 134.995 ;
        RECT 110.640 132.045 111.710 134.825 ;
        RECT 103.980 130.225 107.820 130.395 ;
        RECT 108.220 131.875 111.710 132.045 ;
        RECT 75.865 129.100 83.905 129.270 ;
        RECT 84.955 129.100 92.995 129.270 ;
        RECT 93.675 128.700 94.525 129.650 ;
        RECT 75.015 128.540 94.525 128.700 ;
        RECT 75.015 128.530 93.845 128.540 ;
        RECT 73.175 128.160 95.915 128.350 ;
        RECT 73.175 127.990 96.355 128.160 ;
        RECT 73.175 126.380 73.515 127.990 ;
        RECT 74.240 127.420 84.280 127.590 ;
        RECT 85.420 127.420 95.460 127.590 ;
        RECT 73.855 127.010 74.025 127.360 ;
        RECT 84.495 127.010 84.665 127.360 ;
        RECT 85.035 127.010 85.205 127.360 ;
        RECT 95.675 127.010 95.845 127.360 ;
        RECT 74.240 126.780 84.280 126.950 ;
        RECT 85.420 126.780 95.460 126.950 ;
        RECT 96.185 126.380 96.355 127.990 ;
        RECT 73.175 126.220 96.355 126.380 ;
        RECT 73.345 126.210 96.355 126.220 ;
        RECT 103.980 127.095 105.280 130.225 ;
        RECT 103.980 126.925 107.820 127.095 ;
        RECT 75.035 125.130 95.025 125.450 ;
        RECT 75.025 124.960 95.025 125.130 ;
        RECT 73.285 123.940 74.145 123.950 ;
        RECT 73.185 123.680 74.145 123.940 ;
        RECT 58.790 123.490 67.070 123.660 ;
        RECT 58.875 122.400 60.545 123.490 ;
        RECT 58.875 121.710 59.625 122.230 ;
        RECT 59.795 121.880 60.545 122.400 ;
        RECT 60.755 122.350 60.985 123.490 ;
        RECT 61.155 122.340 61.485 123.320 ;
        RECT 61.655 122.350 61.865 123.490 ;
        RECT 62.135 122.350 62.365 123.490 ;
        RECT 62.535 122.340 62.865 123.320 ;
        RECT 63.035 122.350 63.245 123.490 ;
        RECT 63.515 122.350 63.745 123.490 ;
        RECT 63.915 122.340 64.245 123.320 ;
        RECT 64.415 122.350 64.625 123.490 ;
        RECT 61.235 122.225 61.485 122.340 ;
        RECT 60.735 122.165 61.065 122.180 ;
        RECT 60.730 121.945 61.065 122.165 ;
        RECT 60.735 121.930 61.065 121.945 ;
        RECT 61.235 121.925 61.510 122.225 ;
        RECT 62.115 121.930 62.445 122.180 ;
        RECT 58.875 120.940 60.545 121.710 ;
        RECT 60.755 120.940 60.985 121.760 ;
        RECT 61.235 121.740 61.485 121.925 ;
        RECT 61.155 121.110 61.485 121.740 ;
        RECT 61.655 120.940 61.865 121.760 ;
        RECT 62.135 120.940 62.365 121.760 ;
        RECT 62.615 121.740 62.865 122.340 ;
        RECT 63.495 122.175 63.825 122.180 ;
        RECT 63.480 121.935 63.825 122.175 ;
        RECT 63.495 121.930 63.825 121.935 ;
        RECT 63.995 122.175 64.245 122.340 ;
        RECT 64.855 122.325 65.145 123.490 ;
        RECT 65.315 122.400 66.985 123.490 ;
        RECT 63.995 121.935 64.340 122.175 ;
        RECT 62.535 121.110 62.865 121.740 ;
        RECT 63.035 120.940 63.245 121.760 ;
        RECT 63.515 120.940 63.745 121.760 ;
        RECT 63.995 121.740 64.245 121.935 ;
        RECT 63.915 121.110 64.245 121.740 ;
        RECT 64.415 120.940 64.625 121.760 ;
        RECT 65.315 121.710 66.065 122.230 ;
        RECT 66.235 121.880 66.985 122.400 ;
        RECT 73.185 123.000 74.195 123.680 ;
        RECT 75.025 123.350 75.195 124.960 ;
        RECT 75.875 124.390 83.915 124.560 ;
        RECT 84.965 124.390 93.005 124.560 ;
        RECT 75.535 123.980 75.705 124.330 ;
        RECT 84.085 123.980 84.255 124.330 ;
        RECT 84.625 123.980 84.795 124.330 ;
        RECT 93.175 123.980 93.345 124.330 ;
        RECT 93.685 124.300 95.025 124.960 ;
        RECT 75.875 123.750 83.915 123.920 ;
        RECT 84.965 123.750 93.005 123.920 ;
        RECT 93.685 123.350 94.535 124.300 ;
        RECT 75.025 123.190 94.535 123.350 ;
        RECT 75.025 123.180 93.855 123.190 ;
        RECT 73.185 122.810 95.925 123.000 ;
        RECT 73.185 122.640 96.365 122.810 ;
        RECT 64.855 120.940 65.145 121.665 ;
        RECT 65.315 120.940 66.985 121.710 ;
        RECT 73.185 121.030 73.525 122.640 ;
        RECT 74.250 122.070 84.290 122.240 ;
        RECT 85.430 122.070 95.470 122.240 ;
        RECT 73.865 121.660 74.035 122.010 ;
        RECT 84.505 121.660 84.675 122.010 ;
        RECT 85.045 121.660 85.215 122.010 ;
        RECT 95.685 121.660 95.855 122.010 ;
        RECT 74.250 121.430 84.290 121.600 ;
        RECT 85.430 121.430 95.470 121.600 ;
        RECT 96.195 121.030 96.365 122.640 ;
        RECT 58.790 120.770 69.370 120.940 ;
        RECT 73.185 120.870 96.365 121.030 ;
        RECT 73.355 120.860 96.365 120.870 ;
        RECT 58.875 120.310 59.435 120.600 ;
        RECT 59.605 120.310 59.855 120.770 ;
        RECT 58.875 120.255 59.125 120.310 ;
        RECT 58.870 119.115 59.125 120.255 ;
        RECT 60.475 120.140 60.805 120.500 ;
        RECT 59.415 119.950 60.805 120.140 ;
        RECT 61.195 120.080 61.435 120.600 ;
        RECT 61.605 120.275 62.000 120.770 ;
        RECT 62.565 120.440 62.735 120.585 ;
        RECT 62.360 120.245 62.735 120.440 ;
        RECT 59.415 119.860 59.585 119.950 ;
        RECT 59.295 119.530 59.585 119.860 ;
        RECT 59.755 119.530 60.095 119.780 ;
        RECT 60.315 119.530 60.990 119.780 ;
        RECT 58.875 118.940 59.125 119.115 ;
        RECT 59.415 119.280 59.585 119.530 ;
        RECT 59.415 119.110 60.355 119.280 ;
        RECT 60.725 119.170 60.990 119.530 ;
        RECT 61.195 119.275 61.370 120.080 ;
        RECT 62.360 119.910 62.530 120.245 ;
        RECT 63.015 120.200 63.255 120.575 ;
        RECT 63.425 120.265 63.760 120.770 ;
        RECT 63.015 120.050 63.235 120.200 ;
        RECT 61.545 119.550 62.530 119.910 ;
        RECT 62.700 119.720 63.235 120.050 ;
        RECT 61.545 119.530 62.830 119.550 ;
        RECT 61.970 119.380 62.830 119.530 ;
        RECT 58.875 118.390 59.335 118.940 ;
        RECT 59.525 118.220 59.855 118.940 ;
        RECT 60.055 118.560 60.355 119.110 ;
        RECT 60.525 118.220 60.805 118.890 ;
        RECT 61.195 118.490 61.500 119.275 ;
        RECT 61.675 118.900 62.370 119.210 ;
        RECT 61.680 118.220 62.365 118.690 ;
        RECT 62.545 118.435 62.830 119.380 ;
        RECT 63.000 119.070 63.235 119.720 ;
        RECT 63.405 119.240 63.705 120.090 ;
        RECT 63.955 120.080 64.195 120.600 ;
        RECT 64.365 120.275 64.760 120.770 ;
        RECT 65.325 120.440 65.495 120.585 ;
        RECT 65.120 120.245 65.495 120.440 ;
        RECT 63.955 119.275 64.130 120.080 ;
        RECT 65.120 119.910 65.290 120.245 ;
        RECT 65.775 120.200 66.015 120.575 ;
        RECT 66.185 120.265 66.520 120.770 ;
        RECT 65.775 120.050 65.995 120.200 ;
        RECT 64.305 119.550 65.290 119.910 ;
        RECT 65.460 119.720 65.995 120.050 ;
        RECT 64.305 119.530 65.590 119.550 ;
        RECT 64.730 119.380 65.590 119.530 ;
        RECT 63.000 118.840 63.675 119.070 ;
        RECT 63.005 118.220 63.335 118.670 ;
        RECT 63.505 118.410 63.675 118.840 ;
        RECT 63.955 118.490 64.260 119.275 ;
        RECT 64.435 118.900 65.130 119.210 ;
        RECT 64.440 118.220 65.125 118.690 ;
        RECT 65.305 118.435 65.590 119.380 ;
        RECT 65.760 119.070 65.995 119.720 ;
        RECT 66.165 119.240 66.465 120.090 ;
        RECT 66.695 120.045 66.985 120.770 ;
        RECT 67.155 120.310 67.715 120.600 ;
        RECT 67.885 120.310 68.135 120.770 ;
        RECT 65.760 118.840 66.435 119.070 ;
        RECT 65.765 118.220 66.095 118.670 ;
        RECT 66.265 118.410 66.435 118.840 ;
        RECT 66.695 118.220 66.985 119.385 ;
        RECT 67.155 118.940 67.405 120.310 ;
        RECT 68.755 120.140 69.085 120.500 ;
        RECT 67.695 119.950 69.085 120.140 ;
        RECT 67.695 119.860 67.865 119.950 ;
        RECT 67.575 119.530 67.865 119.860 ;
        RECT 75.005 119.780 94.995 120.100 ;
        RECT 68.035 119.530 68.375 119.780 ;
        RECT 68.595 119.530 69.270 119.780 ;
        RECT 67.695 119.280 67.865 119.530 ;
        RECT 68.650 119.455 69.270 119.530 ;
        RECT 67.695 119.110 68.635 119.280 ;
        RECT 69.005 119.170 69.270 119.455 ;
        RECT 74.995 119.610 94.995 119.780 ;
        RECT 67.155 118.390 67.615 118.940 ;
        RECT 67.805 118.220 68.135 118.940 ;
        RECT 68.335 118.560 68.635 119.110 ;
        RECT 68.805 118.220 69.085 118.890 ;
        RECT 73.255 118.590 74.115 118.600 ;
        RECT 73.155 118.330 74.115 118.590 ;
        RECT 58.790 118.050 69.370 118.220 ;
        RECT 58.875 116.960 60.545 118.050 ;
        RECT 58.875 116.270 59.625 116.790 ;
        RECT 59.795 116.440 60.545 116.960 ;
        RECT 60.715 116.885 61.005 118.050 ;
        RECT 61.215 116.910 61.445 118.050 ;
        RECT 61.615 116.900 61.945 117.880 ;
        RECT 62.115 116.910 62.325 118.050 ;
        RECT 62.595 116.910 62.825 118.050 ;
        RECT 62.995 116.900 63.325 117.880 ;
        RECT 63.495 116.910 63.705 118.050 ;
        RECT 61.195 116.490 61.525 116.740 ;
        RECT 58.875 115.500 60.545 116.270 ;
        RECT 60.715 115.500 61.005 116.225 ;
        RECT 61.215 115.500 61.445 116.320 ;
        RECT 61.695 116.300 61.945 116.900 ;
        RECT 62.575 116.490 62.905 116.740 ;
        RECT 61.615 115.670 61.945 116.300 ;
        RECT 62.115 115.500 62.325 116.320 ;
        RECT 62.595 115.500 62.825 116.320 ;
        RECT 63.075 116.300 63.325 116.900 ;
        RECT 63.935 116.885 64.225 118.050 ;
        RECT 64.435 116.910 64.665 118.050 ;
        RECT 64.835 116.900 65.165 117.880 ;
        RECT 65.335 116.910 65.545 118.050 ;
        RECT 65.815 116.910 66.045 118.050 ;
        RECT 66.215 116.900 66.545 117.880 ;
        RECT 66.715 116.910 66.925 118.050 ;
        RECT 67.155 116.960 68.825 118.050 ;
        RECT 64.415 116.490 64.745 116.740 ;
        RECT 62.995 115.670 63.325 116.300 ;
        RECT 63.495 115.500 63.705 116.320 ;
        RECT 63.935 115.500 64.225 116.225 ;
        RECT 64.435 115.500 64.665 116.320 ;
        RECT 64.915 116.300 65.165 116.900 ;
        RECT 65.795 116.735 66.125 116.740 ;
        RECT 65.770 116.495 66.125 116.735 ;
        RECT 65.795 116.490 66.125 116.495 ;
        RECT 64.835 115.670 65.165 116.300 ;
        RECT 65.335 115.500 65.545 116.320 ;
        RECT 65.815 115.500 66.045 116.320 ;
        RECT 66.295 116.300 66.545 116.900 ;
        RECT 66.215 115.670 66.545 116.300 ;
        RECT 66.715 115.500 66.925 116.320 ;
        RECT 67.155 116.270 67.905 116.790 ;
        RECT 68.075 116.440 68.825 116.960 ;
        RECT 73.155 117.650 74.165 118.330 ;
        RECT 74.995 118.000 75.165 119.610 ;
        RECT 75.845 119.040 83.885 119.210 ;
        RECT 84.935 119.040 92.975 119.210 ;
        RECT 75.505 118.630 75.675 118.980 ;
        RECT 84.055 118.630 84.225 118.980 ;
        RECT 84.595 118.630 84.765 118.980 ;
        RECT 93.145 118.630 93.315 118.980 ;
        RECT 93.655 118.950 94.995 119.610 ;
        RECT 103.980 120.055 105.280 126.925 ;
        RECT 105.760 124.285 107.170 126.445 ;
        RECT 105.760 120.535 107.170 122.695 ;
        RECT 107.650 120.055 107.820 126.925 ;
        RECT 108.220 125.005 108.390 131.875 ;
        RECT 108.870 129.235 110.280 131.395 ;
        RECT 108.870 125.485 110.280 127.645 ;
        RECT 110.640 125.005 111.710 131.875 ;
        RECT 108.220 124.835 111.710 125.005 ;
        RECT 110.640 121.705 111.710 124.835 ;
        RECT 103.980 119.885 107.820 120.055 ;
        RECT 108.160 121.535 111.710 121.705 ;
        RECT 75.845 118.400 83.885 118.570 ;
        RECT 84.935 118.400 92.975 118.570 ;
        RECT 93.655 118.000 94.505 118.950 ;
        RECT 74.995 117.840 94.505 118.000 ;
        RECT 74.995 117.830 93.825 117.840 ;
        RECT 73.155 117.460 95.895 117.650 ;
        RECT 73.155 117.290 96.335 117.460 ;
        RECT 67.155 115.500 68.825 116.270 ;
        RECT 73.155 115.680 73.495 117.290 ;
        RECT 74.220 116.720 84.260 116.890 ;
        RECT 85.400 116.720 95.440 116.890 ;
        RECT 73.835 116.310 74.005 116.660 ;
        RECT 84.475 116.310 84.645 116.660 ;
        RECT 85.015 116.310 85.185 116.660 ;
        RECT 95.655 116.310 95.825 116.660 ;
        RECT 74.220 116.080 84.260 116.250 ;
        RECT 85.400 116.080 95.440 116.250 ;
        RECT 96.165 115.680 96.335 117.290 ;
        RECT 73.155 115.520 96.335 115.680 ;
        RECT 73.325 115.510 96.335 115.520 ;
        RECT 103.980 116.915 105.280 119.885 ;
        RECT 103.980 116.745 107.810 116.915 ;
        RECT 58.790 115.330 68.910 115.500 ;
        RECT 75.045 114.500 95.035 114.820 ;
        RECT 75.035 114.330 95.035 114.500 ;
        RECT 73.295 113.310 74.155 113.320 ;
        RECT 73.195 113.050 74.155 113.310 ;
        RECT 73.195 112.370 74.205 113.050 ;
        RECT 75.035 112.720 75.205 114.330 ;
        RECT 75.885 113.760 83.925 113.930 ;
        RECT 84.975 113.760 93.015 113.930 ;
        RECT 75.545 113.350 75.715 113.700 ;
        RECT 84.095 113.350 84.265 113.700 ;
        RECT 84.635 113.350 84.805 113.700 ;
        RECT 93.185 113.350 93.355 113.700 ;
        RECT 93.695 113.670 95.035 114.330 ;
        RECT 75.885 113.120 83.925 113.290 ;
        RECT 84.975 113.120 93.015 113.290 ;
        RECT 93.695 112.720 94.545 113.670 ;
        RECT 75.035 112.560 94.545 112.720 ;
        RECT 75.035 112.550 93.865 112.560 ;
        RECT 73.195 112.180 95.935 112.370 ;
        RECT 73.195 112.010 96.375 112.180 ;
        RECT 44.780 111.435 64.770 111.755 ;
        RECT 44.770 111.265 64.770 111.435 ;
        RECT 43.030 110.245 43.890 110.255 ;
        RECT 42.930 109.985 43.890 110.245 ;
        RECT 42.930 109.305 43.940 109.985 ;
        RECT 44.770 109.655 44.940 111.265 ;
        RECT 45.620 110.695 53.660 110.865 ;
        RECT 54.710 110.695 62.750 110.865 ;
        RECT 45.280 110.285 45.450 110.635 ;
        RECT 53.830 110.285 54.000 110.635 ;
        RECT 54.370 110.285 54.540 110.635 ;
        RECT 62.920 110.285 63.090 110.635 ;
        RECT 63.430 110.605 64.770 111.265 ;
        RECT 45.620 110.055 53.660 110.225 ;
        RECT 54.710 110.055 62.750 110.225 ;
        RECT 63.430 109.655 64.280 110.605 ;
        RECT 73.195 110.400 73.535 112.010 ;
        RECT 74.260 111.440 84.300 111.610 ;
        RECT 85.440 111.440 95.480 111.610 ;
        RECT 73.875 111.030 74.045 111.380 ;
        RECT 84.515 111.030 84.685 111.380 ;
        RECT 85.055 111.030 85.225 111.380 ;
        RECT 95.695 111.030 95.865 111.380 ;
        RECT 74.260 110.800 84.300 110.970 ;
        RECT 85.440 110.800 95.480 110.970 ;
        RECT 96.205 110.400 96.375 112.010 ;
        RECT 73.195 110.240 96.375 110.400 ;
        RECT 73.365 110.230 96.375 110.240 ;
        RECT 44.770 109.495 64.280 109.655 ;
        RECT 103.980 109.875 105.280 116.745 ;
        RECT 105.750 114.105 107.160 116.265 ;
        RECT 107.640 114.735 107.810 116.745 ;
        RECT 108.160 114.735 108.330 121.535 ;
        RECT 108.810 118.895 110.220 121.055 ;
        RECT 108.810 115.145 110.220 117.305 ;
        RECT 110.640 114.735 111.710 121.535 ;
        RECT 107.640 113.985 111.830 114.735 ;
        RECT 107.610 113.045 111.830 113.985 ;
        RECT 105.750 110.355 107.160 112.515 ;
        RECT 107.610 109.875 111.690 113.045 ;
        RECT 44.770 109.485 63.600 109.495 ;
        RECT 42.930 109.115 65.670 109.305 ;
        RECT 42.930 108.945 66.110 109.115 ;
        RECT 42.930 107.335 43.270 108.945 ;
        RECT 43.995 108.375 54.035 108.545 ;
        RECT 55.175 108.375 65.215 108.545 ;
        RECT 43.610 107.965 43.780 108.315 ;
        RECT 54.250 107.965 54.420 108.315 ;
        RECT 54.790 107.965 54.960 108.315 ;
        RECT 65.430 107.965 65.600 108.315 ;
        RECT 43.995 107.735 54.035 107.905 ;
        RECT 55.175 107.735 65.215 107.905 ;
        RECT 65.940 107.335 66.110 108.945 ;
        RECT 103.980 108.615 111.690 109.875 ;
        RECT 103.980 108.565 108.910 108.615 ;
        RECT 42.930 107.175 66.110 107.335 ;
        RECT 43.100 107.165 66.110 107.175 ;
        RECT 44.790 106.085 64.780 106.405 ;
        RECT 44.780 105.915 64.780 106.085 ;
        RECT 43.040 104.895 43.900 104.905 ;
        RECT 42.940 104.635 43.900 104.895 ;
        RECT 42.940 103.955 43.950 104.635 ;
        RECT 44.780 104.305 44.950 105.915 ;
        RECT 45.630 105.345 53.670 105.515 ;
        RECT 54.720 105.345 62.760 105.515 ;
        RECT 45.290 104.935 45.460 105.285 ;
        RECT 53.840 104.935 54.010 105.285 ;
        RECT 54.380 104.935 54.550 105.285 ;
        RECT 62.930 104.935 63.100 105.285 ;
        RECT 63.440 105.255 64.780 105.915 ;
        RECT 45.630 104.705 53.670 104.875 ;
        RECT 54.720 104.705 62.760 104.875 ;
        RECT 63.440 104.305 64.290 105.255 ;
        RECT 44.780 104.145 64.290 104.305 ;
        RECT 44.780 104.135 63.610 104.145 ;
        RECT 42.940 103.765 65.680 103.955 ;
        RECT 42.940 103.595 66.120 103.765 ;
        RECT 42.940 101.985 43.280 103.595 ;
        RECT 44.005 103.025 54.045 103.195 ;
        RECT 55.185 103.025 65.225 103.195 ;
        RECT 43.620 102.615 43.790 102.965 ;
        RECT 54.260 102.615 54.430 102.965 ;
        RECT 54.800 102.615 54.970 102.965 ;
        RECT 65.440 102.615 65.610 102.965 ;
        RECT 44.005 102.385 54.045 102.555 ;
        RECT 55.185 102.385 65.225 102.555 ;
        RECT 65.950 101.985 66.120 103.595 ;
        RECT 42.940 101.825 66.120 101.985 ;
        RECT 43.110 101.815 66.120 101.825 ;
        RECT 44.760 100.735 64.750 101.055 ;
        RECT 44.750 100.565 64.750 100.735 ;
        RECT 43.010 99.545 43.870 99.555 ;
        RECT 42.910 99.285 43.870 99.545 ;
        RECT 42.910 98.605 43.920 99.285 ;
        RECT 44.750 98.955 44.920 100.565 ;
        RECT 45.600 99.995 53.640 100.165 ;
        RECT 54.690 99.995 62.730 100.165 ;
        RECT 45.260 99.585 45.430 99.935 ;
        RECT 53.810 99.585 53.980 99.935 ;
        RECT 54.350 99.585 54.520 99.935 ;
        RECT 62.900 99.585 63.070 99.935 ;
        RECT 63.410 99.905 64.750 100.565 ;
        RECT 45.600 99.355 53.640 99.525 ;
        RECT 54.690 99.355 62.730 99.525 ;
        RECT 63.410 98.955 64.260 99.905 ;
        RECT 44.750 98.795 64.260 98.955 ;
        RECT 44.750 98.785 63.580 98.795 ;
        RECT 42.910 98.415 65.650 98.605 ;
        RECT 42.910 98.245 66.090 98.415 ;
        RECT 42.910 96.635 43.250 98.245 ;
        RECT 43.975 97.675 54.015 97.845 ;
        RECT 55.155 97.675 65.195 97.845 ;
        RECT 43.590 97.265 43.760 97.615 ;
        RECT 54.230 97.265 54.400 97.615 ;
        RECT 54.770 97.265 54.940 97.615 ;
        RECT 65.410 97.265 65.580 97.615 ;
        RECT 43.975 97.035 54.015 97.205 ;
        RECT 55.155 97.035 65.195 97.205 ;
        RECT 65.920 96.635 66.090 98.245 ;
        RECT 42.910 96.475 66.090 96.635 ;
        RECT 43.080 96.465 66.090 96.475 ;
        RECT 44.800 95.455 64.790 95.775 ;
        RECT 44.790 95.285 64.790 95.455 ;
        RECT 43.050 94.265 43.910 94.275 ;
        RECT 42.950 94.005 43.910 94.265 ;
        RECT 42.950 93.325 43.960 94.005 ;
        RECT 44.790 93.675 44.960 95.285 ;
        RECT 45.640 94.715 53.680 94.885 ;
        RECT 54.730 94.715 62.770 94.885 ;
        RECT 45.300 94.305 45.470 94.655 ;
        RECT 53.850 94.305 54.020 94.655 ;
        RECT 54.390 94.305 54.560 94.655 ;
        RECT 62.940 94.305 63.110 94.655 ;
        RECT 63.450 94.625 64.790 95.285 ;
        RECT 45.640 94.075 53.680 94.245 ;
        RECT 54.730 94.075 62.770 94.245 ;
        RECT 63.450 93.675 64.300 94.625 ;
        RECT 44.790 93.515 64.300 93.675 ;
        RECT 44.790 93.505 63.620 93.515 ;
        RECT 42.950 93.135 65.690 93.325 ;
        RECT 42.950 92.965 66.130 93.135 ;
        RECT 42.950 91.355 43.290 92.965 ;
        RECT 44.015 92.395 54.055 92.565 ;
        RECT 55.195 92.395 65.235 92.565 ;
        RECT 43.630 91.985 43.800 92.335 ;
        RECT 54.270 91.985 54.440 92.335 ;
        RECT 54.810 91.985 54.980 92.335 ;
        RECT 65.450 91.985 65.620 92.335 ;
        RECT 44.015 91.755 54.055 91.925 ;
        RECT 55.195 91.755 65.235 91.925 ;
        RECT 65.960 91.355 66.130 92.965 ;
        RECT 42.950 91.195 66.130 91.355 ;
        RECT 43.120 91.185 66.130 91.195 ;
        RECT 95.965 81.865 96.765 81.905 ;
        RECT 99.465 81.865 103.665 81.905 ;
        RECT 95.495 81.695 97.245 81.865 ;
        RECT 72.030 72.970 89.050 73.140 ;
        RECT 72.115 71.805 72.405 72.970 ;
        RECT 72.615 71.830 72.845 72.970 ;
        RECT 73.015 71.820 73.345 72.800 ;
        RECT 73.515 71.830 73.725 72.970 ;
        RECT 73.995 71.830 74.225 72.970 ;
        RECT 74.395 71.820 74.725 72.800 ;
        RECT 74.895 71.830 75.105 72.970 ;
        RECT 75.375 71.830 75.605 72.970 ;
        RECT 75.775 71.820 76.105 72.800 ;
        RECT 76.275 71.830 76.485 72.970 ;
        RECT 76.755 71.830 76.985 72.970 ;
        RECT 77.155 71.820 77.485 72.800 ;
        RECT 77.655 71.830 77.865 72.970 ;
        RECT 78.135 71.830 78.365 72.970 ;
        RECT 78.535 71.820 78.865 72.800 ;
        RECT 79.035 71.830 79.245 72.970 ;
        RECT 79.515 71.830 79.745 72.970 ;
        RECT 79.915 71.820 80.245 72.800 ;
        RECT 80.415 71.830 80.625 72.970 ;
        RECT 80.895 71.830 81.125 72.970 ;
        RECT 81.295 71.820 81.625 72.800 ;
        RECT 81.795 71.830 82.005 72.970 ;
        RECT 82.275 71.830 82.505 72.970 ;
        RECT 82.675 71.820 83.005 72.800 ;
        RECT 83.175 71.830 83.385 72.970 ;
        RECT 83.655 71.830 83.885 72.970 ;
        RECT 84.055 71.820 84.385 72.800 ;
        RECT 84.555 71.830 84.765 72.970 ;
        RECT 72.595 71.410 72.925 71.660 ;
        RECT 72.115 70.420 72.405 71.145 ;
        RECT 72.615 70.420 72.845 71.240 ;
        RECT 73.095 71.220 73.345 71.820 ;
        RECT 73.975 71.410 74.305 71.660 ;
        RECT 73.015 70.590 73.345 71.220 ;
        RECT 73.515 70.420 73.725 71.240 ;
        RECT 73.995 70.420 74.225 71.240 ;
        RECT 74.475 71.220 74.725 71.820 ;
        RECT 75.355 71.410 75.685 71.660 ;
        RECT 74.395 70.590 74.725 71.220 ;
        RECT 74.895 70.420 75.105 71.240 ;
        RECT 75.375 70.420 75.605 71.240 ;
        RECT 75.855 71.220 76.105 71.820 ;
        RECT 76.735 71.410 77.065 71.660 ;
        RECT 75.775 70.590 76.105 71.220 ;
        RECT 76.275 70.420 76.485 71.240 ;
        RECT 76.755 70.420 76.985 71.240 ;
        RECT 77.235 71.220 77.485 71.820 ;
        RECT 78.115 71.410 78.445 71.660 ;
        RECT 77.155 70.590 77.485 71.220 ;
        RECT 77.655 70.420 77.865 71.240 ;
        RECT 78.135 70.420 78.365 71.240 ;
        RECT 78.615 71.220 78.865 71.820 ;
        RECT 79.495 71.410 79.825 71.660 ;
        RECT 78.535 70.590 78.865 71.220 ;
        RECT 79.035 70.420 79.245 71.240 ;
        RECT 79.515 70.420 79.745 71.240 ;
        RECT 79.995 71.220 80.245 71.820 ;
        RECT 80.875 71.410 81.205 71.660 ;
        RECT 79.915 70.590 80.245 71.220 ;
        RECT 80.415 70.420 80.625 71.240 ;
        RECT 80.895 70.420 81.125 71.240 ;
        RECT 81.375 71.220 81.625 71.820 ;
        RECT 82.255 71.410 82.585 71.660 ;
        RECT 81.295 70.590 81.625 71.220 ;
        RECT 81.795 70.420 82.005 71.240 ;
        RECT 82.275 70.420 82.505 71.240 ;
        RECT 82.755 71.220 83.005 71.820 ;
        RECT 83.635 71.410 83.965 71.660 ;
        RECT 82.675 70.590 83.005 71.220 ;
        RECT 83.175 70.420 83.385 71.240 ;
        RECT 83.655 70.420 83.885 71.240 ;
        RECT 84.135 71.220 84.385 71.820 ;
        RECT 84.995 71.805 85.285 72.970 ;
        RECT 85.455 71.805 85.745 72.970 ;
        RECT 85.915 71.805 86.205 72.970 ;
        RECT 86.375 71.805 86.665 72.970 ;
        RECT 86.835 71.830 87.095 72.970 ;
        RECT 87.265 72.000 87.595 72.800 ;
        RECT 87.765 72.170 87.935 72.970 ;
        RECT 88.105 72.000 88.435 72.800 ;
        RECT 88.605 72.170 88.860 72.970 ;
        RECT 87.265 71.830 88.965 72.000 ;
        RECT 86.835 71.410 87.595 71.660 ;
        RECT 87.765 71.410 88.515 71.660 ;
        RECT 88.685 71.625 88.965 71.830 ;
        RECT 88.685 71.455 88.970 71.625 ;
        RECT 88.685 71.240 88.965 71.455 ;
        RECT 84.055 70.590 84.385 71.220 ;
        RECT 84.555 70.420 84.765 71.240 ;
        RECT 84.995 70.420 85.285 71.145 ;
        RECT 85.455 70.420 85.745 71.145 ;
        RECT 85.915 70.420 86.205 71.145 ;
        RECT 86.375 70.420 86.665 71.145 ;
        RECT 86.835 71.050 87.935 71.220 ;
        RECT 86.835 70.590 87.175 71.050 ;
        RECT 87.345 70.420 87.515 70.880 ;
        RECT 87.685 70.800 87.935 71.050 ;
        RECT 88.105 70.990 88.965 71.240 ;
        RECT 95.495 71.205 95.665 81.695 ;
        RECT 96.205 81.185 96.535 81.355 ;
        RECT 96.065 71.930 96.235 80.970 ;
        RECT 96.505 71.930 96.675 80.970 ;
        RECT 96.205 71.545 96.535 71.715 ;
        RECT 97.075 71.205 97.245 81.695 ;
        RECT 95.495 71.035 97.245 71.205 ;
        RECT 98.995 81.695 104.145 81.865 ;
        RECT 98.995 71.205 99.165 81.695 ;
        RECT 99.465 81.655 103.665 81.695 ;
        RECT 100.205 81.185 100.535 81.355 ;
        RECT 101.165 81.185 101.495 81.355 ;
        RECT 102.125 81.185 102.455 81.355 ;
        RECT 103.085 81.185 103.415 81.355 ;
        RECT 99.565 71.930 99.735 80.970 ;
        RECT 100.045 71.930 100.215 80.970 ;
        RECT 100.525 71.930 100.695 80.970 ;
        RECT 101.005 71.930 101.175 80.970 ;
        RECT 101.485 71.930 101.655 80.970 ;
        RECT 101.965 71.930 102.135 80.970 ;
        RECT 102.445 71.930 102.615 80.970 ;
        RECT 102.925 71.930 103.095 80.970 ;
        RECT 103.405 71.930 103.575 80.970 ;
        RECT 99.725 71.545 100.055 71.715 ;
        RECT 100.685 71.545 101.015 71.715 ;
        RECT 101.645 71.545 101.975 71.715 ;
        RECT 102.605 71.545 102.935 71.715 ;
        RECT 103.975 71.205 104.145 81.695 ;
        RECT 98.995 71.035 104.145 71.205 ;
        RECT 88.525 70.800 88.855 70.820 ;
        RECT 87.685 70.590 88.855 70.800 ;
        RECT 72.030 70.250 89.050 70.420 ;
        RECT 72.115 69.525 72.405 70.250 ;
        RECT 72.635 69.430 72.845 70.250 ;
        RECT 73.015 69.450 73.345 70.080 ;
        RECT 72.115 67.700 72.405 68.865 ;
        RECT 73.015 68.850 73.265 69.450 ;
        RECT 73.515 69.430 73.745 70.250 ;
        RECT 74.015 69.430 74.225 70.250 ;
        RECT 74.395 69.450 74.725 70.080 ;
        RECT 73.435 69.010 73.765 69.260 ;
        RECT 74.395 68.850 74.645 69.450 ;
        RECT 74.895 69.430 75.125 70.250 ;
        RECT 75.395 69.430 75.605 70.250 ;
        RECT 75.775 69.450 76.105 70.080 ;
        RECT 74.815 69.010 75.145 69.260 ;
        RECT 75.775 68.850 76.025 69.450 ;
        RECT 76.275 69.430 76.505 70.250 ;
        RECT 76.775 69.430 76.985 70.250 ;
        RECT 77.155 69.450 77.485 70.080 ;
        RECT 76.195 69.010 76.525 69.260 ;
        RECT 77.155 68.850 77.405 69.450 ;
        RECT 77.655 69.430 77.885 70.250 ;
        RECT 78.155 69.430 78.365 70.250 ;
        RECT 78.535 69.450 78.865 70.080 ;
        RECT 77.575 69.010 77.905 69.260 ;
        RECT 78.535 68.850 78.785 69.450 ;
        RECT 79.035 69.430 79.265 70.250 ;
        RECT 79.535 69.430 79.745 70.250 ;
        RECT 79.915 69.450 80.245 70.080 ;
        RECT 78.955 69.010 79.285 69.260 ;
        RECT 79.915 68.850 80.165 69.450 ;
        RECT 80.415 69.430 80.645 70.250 ;
        RECT 80.915 69.430 81.125 70.250 ;
        RECT 81.295 69.450 81.625 70.080 ;
        RECT 80.335 69.010 80.665 69.260 ;
        RECT 81.295 68.850 81.545 69.450 ;
        RECT 81.795 69.430 82.025 70.250 ;
        RECT 82.295 69.430 82.505 70.250 ;
        RECT 82.675 69.450 83.005 70.080 ;
        RECT 81.715 69.010 82.045 69.260 ;
        RECT 82.675 68.850 82.925 69.450 ;
        RECT 83.175 69.430 83.405 70.250 ;
        RECT 83.675 69.430 83.885 70.250 ;
        RECT 84.055 69.450 84.385 70.080 ;
        RECT 83.095 69.010 83.425 69.260 ;
        RECT 84.055 68.850 84.305 69.450 ;
        RECT 84.555 69.430 84.785 70.250 ;
        RECT 84.995 69.525 85.285 70.250 ;
        RECT 84.475 69.010 84.805 69.260 ;
        RECT 95.495 69.105 97.245 69.275 ;
        RECT 72.635 67.700 72.845 68.840 ;
        RECT 73.015 67.870 73.345 68.850 ;
        RECT 73.515 67.700 73.745 68.840 ;
        RECT 74.015 67.700 74.225 68.840 ;
        RECT 74.395 67.870 74.725 68.850 ;
        RECT 74.895 67.700 75.125 68.840 ;
        RECT 75.395 67.700 75.605 68.840 ;
        RECT 75.775 67.870 76.105 68.850 ;
        RECT 76.275 67.700 76.505 68.840 ;
        RECT 76.775 67.700 76.985 68.840 ;
        RECT 77.155 67.870 77.485 68.850 ;
        RECT 77.655 67.700 77.885 68.840 ;
        RECT 78.155 67.700 78.365 68.840 ;
        RECT 78.535 67.870 78.865 68.850 ;
        RECT 79.035 67.700 79.265 68.840 ;
        RECT 79.535 67.700 79.745 68.840 ;
        RECT 79.915 67.870 80.245 68.850 ;
        RECT 80.415 67.700 80.645 68.840 ;
        RECT 80.915 67.700 81.125 68.840 ;
        RECT 81.295 67.870 81.625 68.850 ;
        RECT 81.795 67.700 82.025 68.840 ;
        RECT 82.295 67.700 82.505 68.840 ;
        RECT 82.675 67.870 83.005 68.850 ;
        RECT 83.175 67.700 83.405 68.840 ;
        RECT 83.675 67.700 83.885 68.840 ;
        RECT 84.055 67.870 84.385 68.850 ;
        RECT 84.555 67.700 84.785 68.840 ;
        RECT 84.995 67.700 85.285 68.865 ;
        RECT 72.030 67.530 85.370 67.700 ;
        RECT 95.495 64.705 95.665 69.105 ;
        RECT 96.205 68.595 96.535 68.765 ;
        RECT 96.065 65.385 96.235 68.425 ;
        RECT 96.505 65.385 96.675 68.425 ;
        RECT 96.205 65.045 96.535 65.215 ;
        RECT 97.075 64.705 97.245 69.105 ;
        RECT 95.495 64.535 97.245 64.705 ;
        RECT 98.995 69.105 104.145 69.275 ;
        RECT 98.995 64.705 99.165 69.105 ;
        RECT 100.205 68.595 100.535 68.765 ;
        RECT 101.165 68.595 101.495 68.765 ;
        RECT 102.125 68.595 102.455 68.765 ;
        RECT 103.085 68.595 103.415 68.765 ;
        RECT 99.565 65.385 99.735 68.425 ;
        RECT 100.045 65.385 100.215 68.425 ;
        RECT 100.525 65.385 100.695 68.425 ;
        RECT 101.005 65.385 101.175 68.425 ;
        RECT 101.485 65.385 101.655 68.425 ;
        RECT 101.965 65.385 102.135 68.425 ;
        RECT 102.445 65.385 102.615 68.425 ;
        RECT 102.925 65.385 103.095 68.425 ;
        RECT 103.405 65.385 103.575 68.425 ;
        RECT 99.725 65.045 100.055 65.215 ;
        RECT 100.685 65.045 101.015 65.215 ;
        RECT 101.645 65.045 101.975 65.215 ;
        RECT 102.605 65.045 102.935 65.215 ;
        RECT 103.975 64.705 104.145 69.105 ;
        RECT 98.995 64.535 104.145 64.705 ;
        RECT 95.915 64.455 96.815 64.535 ;
        RECT 99.565 64.505 103.715 64.535 ;
        RECT 77.440 64.045 85.720 64.215 ;
        RECT 77.525 62.955 79.195 64.045 ;
        RECT 77.525 62.265 78.275 62.785 ;
        RECT 78.445 62.435 79.195 62.955 ;
        RECT 79.405 62.905 79.635 64.045 ;
        RECT 79.805 62.895 80.135 63.875 ;
        RECT 80.305 62.905 80.515 64.045 ;
        RECT 80.785 62.905 81.015 64.045 ;
        RECT 81.185 62.895 81.515 63.875 ;
        RECT 81.685 62.905 81.895 64.045 ;
        RECT 82.165 62.905 82.395 64.045 ;
        RECT 82.565 62.895 82.895 63.875 ;
        RECT 83.065 62.905 83.275 64.045 ;
        RECT 79.885 62.780 80.135 62.895 ;
        RECT 79.385 62.720 79.715 62.735 ;
        RECT 79.380 62.500 79.715 62.720 ;
        RECT 79.385 62.485 79.715 62.500 ;
        RECT 79.885 62.480 80.160 62.780 ;
        RECT 80.765 62.485 81.095 62.735 ;
        RECT 77.525 61.495 79.195 62.265 ;
        RECT 79.405 61.495 79.635 62.315 ;
        RECT 79.885 62.295 80.135 62.480 ;
        RECT 79.805 61.665 80.135 62.295 ;
        RECT 80.305 61.495 80.515 62.315 ;
        RECT 80.785 61.495 81.015 62.315 ;
        RECT 81.265 62.295 81.515 62.895 ;
        RECT 82.145 62.730 82.475 62.735 ;
        RECT 82.130 62.490 82.475 62.730 ;
        RECT 82.145 62.485 82.475 62.490 ;
        RECT 82.645 62.730 82.895 62.895 ;
        RECT 83.505 62.880 83.795 64.045 ;
        RECT 83.965 62.955 85.635 64.045 ;
        RECT 82.645 62.490 82.990 62.730 ;
        RECT 81.185 61.665 81.515 62.295 ;
        RECT 81.685 61.495 81.895 62.315 ;
        RECT 82.165 61.495 82.395 62.315 ;
        RECT 82.645 62.295 82.895 62.490 ;
        RECT 82.565 61.665 82.895 62.295 ;
        RECT 83.065 61.495 83.275 62.315 ;
        RECT 83.965 62.265 84.715 62.785 ;
        RECT 84.885 62.435 85.635 62.955 ;
        RECT 83.505 61.495 83.795 62.220 ;
        RECT 83.965 61.495 85.635 62.265 ;
        RECT 77.440 61.325 88.020 61.495 ;
        RECT 77.525 60.865 78.085 61.155 ;
        RECT 78.255 60.865 78.505 61.325 ;
        RECT 77.525 60.810 77.775 60.865 ;
        RECT 77.520 59.670 77.775 60.810 ;
        RECT 79.125 60.695 79.455 61.055 ;
        RECT 78.065 60.505 79.455 60.695 ;
        RECT 79.845 60.635 80.085 61.155 ;
        RECT 80.255 60.830 80.650 61.325 ;
        RECT 81.215 60.995 81.385 61.140 ;
        RECT 81.010 60.800 81.385 60.995 ;
        RECT 78.065 60.415 78.235 60.505 ;
        RECT 77.945 60.085 78.235 60.415 ;
        RECT 78.405 60.085 78.745 60.335 ;
        RECT 78.965 60.085 79.640 60.335 ;
        RECT 77.525 59.495 77.775 59.670 ;
        RECT 78.065 59.835 78.235 60.085 ;
        RECT 78.065 59.665 79.005 59.835 ;
        RECT 79.375 59.725 79.640 60.085 ;
        RECT 79.845 59.830 80.020 60.635 ;
        RECT 81.010 60.465 81.180 60.800 ;
        RECT 81.665 60.755 81.905 61.130 ;
        RECT 82.075 60.820 82.410 61.325 ;
        RECT 81.665 60.605 81.885 60.755 ;
        RECT 80.195 60.105 81.180 60.465 ;
        RECT 81.350 60.275 81.885 60.605 ;
        RECT 80.195 60.085 81.480 60.105 ;
        RECT 80.620 59.935 81.480 60.085 ;
        RECT 77.525 58.945 77.985 59.495 ;
        RECT 78.175 58.775 78.505 59.495 ;
        RECT 78.705 59.115 79.005 59.665 ;
        RECT 79.175 58.775 79.455 59.445 ;
        RECT 79.845 59.045 80.150 59.830 ;
        RECT 80.325 59.455 81.020 59.765 ;
        RECT 80.330 58.775 81.015 59.245 ;
        RECT 81.195 58.990 81.480 59.935 ;
        RECT 81.650 59.625 81.885 60.275 ;
        RECT 82.055 59.795 82.355 60.645 ;
        RECT 82.605 60.635 82.845 61.155 ;
        RECT 83.015 60.830 83.410 61.325 ;
        RECT 83.975 60.995 84.145 61.140 ;
        RECT 83.770 60.800 84.145 60.995 ;
        RECT 82.605 59.830 82.780 60.635 ;
        RECT 83.770 60.465 83.940 60.800 ;
        RECT 84.425 60.755 84.665 61.130 ;
        RECT 84.835 60.820 85.170 61.325 ;
        RECT 84.425 60.605 84.645 60.755 ;
        RECT 82.955 60.105 83.940 60.465 ;
        RECT 84.110 60.275 84.645 60.605 ;
        RECT 82.955 60.085 84.240 60.105 ;
        RECT 83.380 59.935 84.240 60.085 ;
        RECT 81.650 59.395 82.325 59.625 ;
        RECT 81.655 58.775 81.985 59.225 ;
        RECT 82.155 58.965 82.325 59.395 ;
        RECT 82.605 59.045 82.910 59.830 ;
        RECT 83.085 59.455 83.780 59.765 ;
        RECT 83.090 58.775 83.775 59.245 ;
        RECT 83.955 58.990 84.240 59.935 ;
        RECT 84.410 59.625 84.645 60.275 ;
        RECT 84.815 59.795 85.115 60.645 ;
        RECT 85.345 60.600 85.635 61.325 ;
        RECT 85.805 60.865 86.365 61.155 ;
        RECT 86.535 60.865 86.785 61.325 ;
        RECT 84.410 59.395 85.085 59.625 ;
        RECT 84.415 58.775 84.745 59.225 ;
        RECT 84.915 58.965 85.085 59.395 ;
        RECT 85.345 58.775 85.635 59.940 ;
        RECT 85.805 59.495 86.055 60.865 ;
        RECT 87.405 60.695 87.735 61.055 ;
        RECT 86.345 60.505 87.735 60.695 ;
        RECT 86.345 60.415 86.515 60.505 ;
        RECT 86.225 60.085 86.515 60.415 ;
        RECT 86.685 60.085 87.025 60.335 ;
        RECT 87.245 60.085 87.920 60.335 ;
        RECT 86.345 59.835 86.515 60.085 ;
        RECT 87.300 60.010 87.920 60.085 ;
        RECT 86.345 59.665 87.285 59.835 ;
        RECT 87.655 59.725 87.920 60.010 ;
        RECT 85.805 58.945 86.265 59.495 ;
        RECT 86.455 58.775 86.785 59.495 ;
        RECT 86.985 59.115 87.285 59.665 ;
        RECT 87.455 58.775 87.735 59.445 ;
        RECT 77.440 58.605 88.020 58.775 ;
        RECT 77.525 57.515 79.195 58.605 ;
        RECT 77.525 56.825 78.275 57.345 ;
        RECT 78.445 56.995 79.195 57.515 ;
        RECT 79.365 57.440 79.655 58.605 ;
        RECT 79.865 57.465 80.095 58.605 ;
        RECT 80.265 57.455 80.595 58.435 ;
        RECT 80.765 57.465 80.975 58.605 ;
        RECT 81.245 57.465 81.475 58.605 ;
        RECT 81.645 57.455 81.975 58.435 ;
        RECT 82.145 57.465 82.355 58.605 ;
        RECT 79.845 57.045 80.175 57.295 ;
        RECT 77.525 56.055 79.195 56.825 ;
        RECT 79.365 56.055 79.655 56.780 ;
        RECT 79.865 56.055 80.095 56.875 ;
        RECT 80.345 56.855 80.595 57.455 ;
        RECT 81.225 57.045 81.555 57.295 ;
        RECT 80.265 56.225 80.595 56.855 ;
        RECT 80.765 56.055 80.975 56.875 ;
        RECT 81.245 56.055 81.475 56.875 ;
        RECT 81.725 56.855 81.975 57.455 ;
        RECT 82.585 57.440 82.875 58.605 ;
        RECT 83.085 57.465 83.315 58.605 ;
        RECT 83.485 57.455 83.815 58.435 ;
        RECT 83.985 57.465 84.195 58.605 ;
        RECT 84.465 57.465 84.695 58.605 ;
        RECT 84.865 57.455 85.195 58.435 ;
        RECT 85.365 57.465 85.575 58.605 ;
        RECT 85.805 57.515 87.475 58.605 ;
        RECT 83.065 57.045 83.395 57.295 ;
        RECT 81.645 56.225 81.975 56.855 ;
        RECT 82.145 56.055 82.355 56.875 ;
        RECT 82.585 56.055 82.875 56.780 ;
        RECT 83.085 56.055 83.315 56.875 ;
        RECT 83.565 56.855 83.815 57.455 ;
        RECT 84.445 57.290 84.775 57.295 ;
        RECT 84.420 57.050 84.775 57.290 ;
        RECT 84.445 57.045 84.775 57.050 ;
        RECT 83.485 56.225 83.815 56.855 ;
        RECT 83.985 56.055 84.195 56.875 ;
        RECT 84.465 56.055 84.695 56.875 ;
        RECT 84.945 56.855 85.195 57.455 ;
        RECT 84.865 56.225 85.195 56.855 ;
        RECT 85.365 56.055 85.575 56.875 ;
        RECT 85.805 56.825 86.555 57.345 ;
        RECT 86.725 56.995 87.475 57.515 ;
        RECT 85.805 56.055 87.475 56.825 ;
        RECT 103.270 56.270 141.450 56.440 ;
        RECT 77.440 55.885 87.560 56.055 ;
        RECT 103.355 55.520 104.565 56.270 ;
        RECT 104.735 55.725 110.080 56.270 ;
        RECT 103.355 54.980 103.875 55.520 ;
        RECT 104.045 54.810 104.565 55.350 ;
        RECT 106.320 54.895 106.660 55.725 ;
        RECT 110.255 55.595 110.515 56.100 ;
        RECT 110.695 55.890 111.025 56.270 ;
        RECT 111.205 55.720 111.375 56.100 ;
        RECT 103.355 53.720 104.565 54.810 ;
        RECT 108.140 54.155 108.490 55.405 ;
        RECT 110.255 54.795 110.435 55.595 ;
        RECT 110.710 55.550 111.375 55.720 ;
        RECT 110.710 55.295 110.880 55.550 ;
        RECT 111.635 55.500 115.145 56.270 ;
        RECT 116.235 55.545 116.525 56.270 ;
        RECT 116.695 55.725 122.040 56.270 ;
        RECT 122.215 55.725 127.560 56.270 ;
        RECT 110.605 54.965 110.880 55.295 ;
        RECT 111.105 55.000 111.445 55.370 ;
        RECT 111.635 54.980 113.285 55.500 ;
        RECT 110.710 54.820 110.880 54.965 ;
        RECT 104.735 53.720 110.080 54.155 ;
        RECT 110.255 53.890 110.525 54.795 ;
        RECT 110.710 54.650 111.385 54.820 ;
        RECT 113.455 54.810 115.145 55.330 ;
        RECT 118.280 54.895 118.620 55.725 ;
        RECT 110.695 53.720 111.025 54.480 ;
        RECT 111.205 53.890 111.385 54.650 ;
        RECT 111.635 53.720 115.145 54.810 ;
        RECT 116.235 53.720 116.525 54.885 ;
        RECT 120.100 54.155 120.450 55.405 ;
        RECT 123.800 54.895 124.140 55.725 ;
        RECT 127.735 55.520 128.945 56.270 ;
        RECT 129.115 55.545 129.405 56.270 ;
        RECT 129.575 55.725 134.920 56.270 ;
        RECT 125.620 54.155 125.970 55.405 ;
        RECT 127.735 54.980 128.255 55.520 ;
        RECT 128.425 54.810 128.945 55.350 ;
        RECT 131.160 54.895 131.500 55.725 ;
        RECT 135.095 55.500 138.605 56.270 ;
        RECT 138.775 55.520 139.985 56.270 ;
        RECT 140.155 55.520 141.365 56.270 ;
        RECT 116.695 53.720 122.040 54.155 ;
        RECT 122.215 53.720 127.560 54.155 ;
        RECT 127.735 53.720 128.945 54.810 ;
        RECT 129.115 53.720 129.405 54.885 ;
        RECT 132.980 54.155 133.330 55.405 ;
        RECT 135.095 54.980 136.745 55.500 ;
        RECT 136.915 54.810 138.605 55.330 ;
        RECT 138.775 54.980 139.295 55.520 ;
        RECT 139.465 54.810 139.985 55.350 ;
        RECT 129.575 53.720 134.920 54.155 ;
        RECT 135.095 53.720 138.605 54.810 ;
        RECT 138.775 53.720 139.985 54.810 ;
        RECT 140.155 54.810 140.675 55.350 ;
        RECT 140.845 54.980 141.365 55.520 ;
        RECT 140.155 53.720 141.365 54.810 ;
        RECT 103.270 53.550 141.450 53.720 ;
        RECT 103.355 52.460 104.565 53.550 ;
        RECT 104.735 53.115 110.080 53.550 ;
        RECT 110.255 53.115 115.600 53.550 ;
        RECT 63.430 51.990 83.420 52.310 ;
        RECT 63.420 51.820 83.420 51.990 ;
        RECT 61.680 50.800 62.540 50.810 ;
        RECT 61.580 50.540 62.540 50.800 ;
        RECT 61.580 49.860 62.590 50.540 ;
        RECT 63.420 50.210 63.590 51.820 ;
        RECT 64.270 51.250 72.310 51.420 ;
        RECT 73.360 51.250 81.400 51.420 ;
        RECT 63.930 50.840 64.100 51.190 ;
        RECT 72.480 50.840 72.650 51.190 ;
        RECT 73.020 50.840 73.190 51.190 ;
        RECT 81.570 50.840 81.740 51.190 ;
        RECT 82.080 51.160 83.420 51.820 ;
        RECT 103.355 51.750 103.875 52.290 ;
        RECT 104.045 51.920 104.565 52.460 ;
        RECT 64.270 50.610 72.310 50.780 ;
        RECT 73.360 50.610 81.400 50.780 ;
        RECT 82.080 50.210 82.930 51.160 ;
        RECT 103.355 51.000 104.565 51.750 ;
        RECT 106.320 51.545 106.660 52.375 ;
        RECT 108.140 51.865 108.490 53.115 ;
        RECT 111.840 51.545 112.180 52.375 ;
        RECT 113.660 51.865 114.010 53.115 ;
        RECT 116.235 52.385 116.525 53.550 ;
        RECT 116.695 53.115 122.040 53.550 ;
        RECT 122.215 53.115 127.560 53.550 ;
        RECT 127.735 53.115 133.080 53.550 ;
        RECT 133.255 53.115 138.600 53.550 ;
        RECT 104.735 51.000 110.080 51.545 ;
        RECT 110.255 51.000 115.600 51.545 ;
        RECT 116.235 51.000 116.525 51.725 ;
        RECT 118.280 51.545 118.620 52.375 ;
        RECT 120.100 51.865 120.450 53.115 ;
        RECT 123.800 51.545 124.140 52.375 ;
        RECT 125.620 51.865 125.970 53.115 ;
        RECT 129.320 51.545 129.660 52.375 ;
        RECT 131.140 51.865 131.490 53.115 ;
        RECT 134.840 51.545 135.180 52.375 ;
        RECT 136.660 51.865 137.010 53.115 ;
        RECT 138.775 52.460 139.985 53.550 ;
        RECT 138.775 51.750 139.295 52.290 ;
        RECT 139.465 51.920 139.985 52.460 ;
        RECT 140.155 52.460 141.365 53.550 ;
        RECT 140.155 51.920 140.675 52.460 ;
        RECT 140.845 51.750 141.365 52.290 ;
        RECT 116.695 51.000 122.040 51.545 ;
        RECT 122.215 51.000 127.560 51.545 ;
        RECT 127.735 51.000 133.080 51.545 ;
        RECT 133.255 51.000 138.600 51.545 ;
        RECT 138.775 51.000 139.985 51.750 ;
        RECT 140.155 51.000 141.365 51.750 ;
        RECT 103.270 50.830 141.450 51.000 ;
        RECT 63.420 50.050 82.930 50.210 ;
        RECT 103.355 50.080 104.565 50.830 ;
        RECT 63.420 50.040 82.250 50.050 ;
        RECT 61.580 49.670 84.320 49.860 ;
        RECT 61.580 49.500 84.760 49.670 ;
        RECT 103.355 49.540 103.875 50.080 ;
        RECT 104.735 50.060 106.405 50.830 ;
        RECT 107.085 50.440 107.415 50.830 ;
        RECT 107.585 50.260 107.755 50.580 ;
        RECT 107.925 50.440 108.255 50.830 ;
        RECT 108.670 50.430 109.625 50.600 ;
        RECT 107.035 50.090 109.285 50.260 ;
        RECT 61.580 47.890 61.920 49.500 ;
        RECT 62.645 48.930 72.685 49.100 ;
        RECT 73.825 48.930 83.865 49.100 ;
        RECT 62.260 48.520 62.430 48.870 ;
        RECT 72.900 48.520 73.070 48.870 ;
        RECT 73.440 48.520 73.610 48.870 ;
        RECT 84.080 48.520 84.250 48.870 ;
        RECT 62.645 48.290 72.685 48.460 ;
        RECT 73.825 48.290 83.865 48.460 ;
        RECT 84.590 47.890 84.760 49.500 ;
        RECT 104.045 49.370 104.565 49.910 ;
        RECT 104.735 49.540 105.485 50.060 ;
        RECT 105.655 49.370 106.405 49.890 ;
        RECT 103.355 48.280 104.565 49.370 ;
        RECT 104.735 48.280 106.405 49.370 ;
        RECT 107.035 49.130 107.205 50.090 ;
        RECT 107.375 49.470 107.620 49.920 ;
        RECT 107.790 49.640 108.340 49.840 ;
        RECT 108.510 49.670 108.885 49.840 ;
        RECT 108.510 49.470 108.680 49.670 ;
        RECT 109.055 49.590 109.285 50.090 ;
        RECT 107.375 49.300 108.680 49.470 ;
        RECT 109.455 49.550 109.625 50.430 ;
        RECT 109.795 49.995 110.085 50.830 ;
        RECT 110.255 50.285 115.600 50.830 ;
        RECT 115.775 50.285 121.120 50.830 ;
        RECT 121.295 50.285 126.640 50.830 ;
        RECT 109.455 49.380 110.085 49.550 ;
        RECT 111.840 49.455 112.180 50.285 ;
        RECT 107.035 48.450 107.415 49.130 ;
        RECT 108.005 48.280 108.175 49.130 ;
        RECT 108.345 48.960 109.585 49.130 ;
        RECT 108.345 48.450 108.675 48.960 ;
        RECT 108.845 48.280 109.015 48.790 ;
        RECT 109.185 48.450 109.585 48.960 ;
        RECT 109.765 48.450 110.085 49.380 ;
        RECT 113.660 48.715 114.010 49.965 ;
        RECT 117.360 49.455 117.700 50.285 ;
        RECT 119.180 48.715 119.530 49.965 ;
        RECT 122.880 49.455 123.220 50.285 ;
        RECT 126.815 50.060 128.485 50.830 ;
        RECT 129.115 50.105 129.405 50.830 ;
        RECT 129.575 50.285 134.920 50.830 ;
        RECT 124.700 48.715 125.050 49.965 ;
        RECT 126.815 49.540 127.565 50.060 ;
        RECT 127.735 49.370 128.485 49.890 ;
        RECT 131.160 49.455 131.500 50.285 ;
        RECT 135.095 50.060 138.605 50.830 ;
        RECT 138.775 50.080 139.985 50.830 ;
        RECT 140.155 50.080 141.365 50.830 ;
        RECT 110.255 48.280 115.600 48.715 ;
        RECT 115.775 48.280 121.120 48.715 ;
        RECT 121.295 48.280 126.640 48.715 ;
        RECT 126.815 48.280 128.485 49.370 ;
        RECT 129.115 48.280 129.405 49.445 ;
        RECT 132.980 48.715 133.330 49.965 ;
        RECT 135.095 49.540 136.745 50.060 ;
        RECT 136.915 49.370 138.605 49.890 ;
        RECT 138.775 49.540 139.295 50.080 ;
        RECT 139.465 49.370 139.985 49.910 ;
        RECT 129.575 48.280 134.920 48.715 ;
        RECT 135.095 48.280 138.605 49.370 ;
        RECT 138.775 48.280 139.985 49.370 ;
        RECT 140.155 49.370 140.675 49.910 ;
        RECT 140.845 49.540 141.365 50.080 ;
        RECT 140.155 48.280 141.365 49.370 ;
        RECT 103.270 48.110 141.450 48.280 ;
        RECT 61.580 47.730 84.760 47.890 ;
        RECT 61.750 47.720 84.760 47.730 ;
        RECT 103.355 47.020 104.565 48.110 ;
        RECT 104.735 47.020 106.405 48.110 ;
        RECT 107.095 47.050 107.425 47.895 ;
        RECT 107.595 47.100 107.765 48.110 ;
        RECT 107.935 47.380 108.275 47.940 ;
        RECT 108.505 47.610 108.820 48.110 ;
        RECT 109.000 47.640 109.885 47.810 ;
        RECT 63.440 46.640 83.430 46.960 ;
        RECT 63.430 46.470 83.430 46.640 ;
        RECT 61.690 45.450 62.550 45.460 ;
        RECT 61.590 45.190 62.550 45.450 ;
        RECT 61.590 44.510 62.600 45.190 ;
        RECT 63.430 44.860 63.600 46.470 ;
        RECT 64.280 45.900 72.320 46.070 ;
        RECT 73.370 45.900 81.410 46.070 ;
        RECT 63.940 45.490 64.110 45.840 ;
        RECT 72.490 45.490 72.660 45.840 ;
        RECT 73.030 45.490 73.200 45.840 ;
        RECT 81.580 45.490 81.750 45.840 ;
        RECT 82.090 45.810 83.430 46.470 ;
        RECT 103.355 46.310 103.875 46.850 ;
        RECT 104.045 46.480 104.565 47.020 ;
        RECT 104.735 46.330 105.485 46.850 ;
        RECT 105.655 46.500 106.405 47.020 ;
        RECT 107.035 46.970 107.425 47.050 ;
        RECT 107.935 47.005 108.830 47.380 ;
        RECT 107.035 46.920 107.250 46.970 ;
        RECT 107.035 46.340 107.205 46.920 ;
        RECT 107.935 46.800 108.125 47.005 ;
        RECT 109.000 46.800 109.170 47.640 ;
        RECT 110.110 47.610 110.360 47.940 ;
        RECT 107.375 46.470 108.125 46.800 ;
        RECT 108.295 46.470 109.170 46.800 ;
        RECT 64.280 45.260 72.320 45.430 ;
        RECT 73.370 45.260 81.410 45.430 ;
        RECT 82.090 44.860 82.940 45.810 ;
        RECT 103.355 45.560 104.565 46.310 ;
        RECT 104.735 45.560 106.405 46.330 ;
        RECT 107.035 46.300 107.260 46.340 ;
        RECT 107.925 46.300 108.125 46.470 ;
        RECT 107.035 46.215 107.415 46.300 ;
        RECT 107.085 45.780 107.415 46.215 ;
        RECT 107.585 45.560 107.755 46.170 ;
        RECT 107.925 45.775 108.255 46.300 ;
        RECT 108.515 45.560 108.725 46.090 ;
        RECT 109.000 46.010 109.170 46.470 ;
        RECT 109.340 46.510 109.660 47.470 ;
        RECT 109.830 46.720 110.020 47.440 ;
        RECT 110.190 46.540 110.360 47.610 ;
        RECT 110.530 47.310 110.700 48.110 ;
        RECT 110.870 47.665 111.975 47.835 ;
        RECT 110.870 47.050 111.040 47.665 ;
        RECT 112.185 47.515 112.435 47.940 ;
        RECT 112.605 47.650 112.870 48.110 ;
        RECT 111.210 47.130 111.740 47.495 ;
        RECT 112.185 47.385 112.490 47.515 ;
        RECT 110.530 46.960 111.040 47.050 ;
        RECT 110.530 46.790 111.400 46.960 ;
        RECT 110.530 46.720 110.700 46.790 ;
        RECT 110.820 46.540 111.020 46.570 ;
        RECT 109.340 46.180 109.805 46.510 ;
        RECT 110.190 46.240 111.020 46.540 ;
        RECT 110.190 46.010 110.360 46.240 ;
        RECT 109.000 45.840 109.785 46.010 ;
        RECT 109.955 45.840 110.360 46.010 ;
        RECT 110.540 45.560 110.910 46.060 ;
        RECT 111.230 46.010 111.400 46.790 ;
        RECT 111.570 46.430 111.740 47.130 ;
        RECT 111.910 46.600 112.150 47.195 ;
        RECT 111.570 46.210 112.095 46.430 ;
        RECT 112.320 46.280 112.490 47.385 ;
        RECT 112.265 46.150 112.490 46.280 ;
        RECT 112.660 46.190 112.940 47.140 ;
        RECT 112.265 46.010 112.435 46.150 ;
        RECT 111.230 45.840 111.905 46.010 ;
        RECT 112.100 45.840 112.435 46.010 ;
        RECT 112.605 45.560 112.855 46.020 ;
        RECT 113.110 45.820 113.295 47.940 ;
        RECT 113.465 47.610 113.795 48.110 ;
        RECT 113.965 47.440 114.135 47.940 ;
        RECT 113.470 47.270 114.135 47.440 ;
        RECT 113.470 46.280 113.700 47.270 ;
        RECT 113.870 46.450 114.220 47.100 ;
        RECT 114.395 47.020 116.065 48.110 ;
        RECT 114.395 46.330 115.145 46.850 ;
        RECT 115.315 46.500 116.065 47.020 ;
        RECT 116.235 46.945 116.525 48.110 ;
        RECT 116.695 47.675 122.040 48.110 ;
        RECT 122.215 47.675 127.560 48.110 ;
        RECT 127.735 47.675 133.080 48.110 ;
        RECT 133.255 47.675 138.600 48.110 ;
        RECT 113.470 46.110 114.135 46.280 ;
        RECT 113.465 45.560 113.795 45.940 ;
        RECT 113.965 45.820 114.135 46.110 ;
        RECT 114.395 45.560 116.065 46.330 ;
        RECT 116.235 45.560 116.525 46.285 ;
        RECT 118.280 46.105 118.620 46.935 ;
        RECT 120.100 46.425 120.450 47.675 ;
        RECT 123.800 46.105 124.140 46.935 ;
        RECT 125.620 46.425 125.970 47.675 ;
        RECT 129.320 46.105 129.660 46.935 ;
        RECT 131.140 46.425 131.490 47.675 ;
        RECT 134.840 46.105 135.180 46.935 ;
        RECT 136.660 46.425 137.010 47.675 ;
        RECT 138.775 47.020 139.985 48.110 ;
        RECT 138.775 46.310 139.295 46.850 ;
        RECT 139.465 46.480 139.985 47.020 ;
        RECT 140.155 47.020 141.365 48.110 ;
        RECT 140.155 46.480 140.675 47.020 ;
        RECT 140.845 46.310 141.365 46.850 ;
        RECT 116.695 45.560 122.040 46.105 ;
        RECT 122.215 45.560 127.560 46.105 ;
        RECT 127.735 45.560 133.080 46.105 ;
        RECT 133.255 45.560 138.600 46.105 ;
        RECT 138.775 45.560 139.985 46.310 ;
        RECT 140.155 45.560 141.365 46.310 ;
        RECT 103.270 45.390 141.450 45.560 ;
        RECT 63.430 44.700 82.940 44.860 ;
        RECT 63.430 44.690 82.260 44.700 ;
        RECT 103.355 44.640 104.565 45.390 ;
        RECT 105.205 44.660 105.505 45.390 ;
        RECT 61.590 44.320 84.330 44.510 ;
        RECT 61.590 44.150 84.770 44.320 ;
        RECT 61.590 42.540 61.930 44.150 ;
        RECT 62.655 43.580 72.695 43.750 ;
        RECT 73.835 43.580 83.875 43.750 ;
        RECT 62.270 43.170 62.440 43.520 ;
        RECT 72.910 43.170 73.080 43.520 ;
        RECT 73.450 43.170 73.620 43.520 ;
        RECT 84.090 43.170 84.260 43.520 ;
        RECT 62.655 42.940 72.695 43.110 ;
        RECT 73.835 42.940 83.875 43.110 ;
        RECT 84.600 42.540 84.770 44.150 ;
        RECT 103.355 44.100 103.875 44.640 ;
        RECT 105.685 44.480 105.915 45.100 ;
        RECT 106.115 44.830 106.340 45.210 ;
        RECT 106.510 45.000 106.840 45.390 ;
        RECT 106.115 44.650 106.445 44.830 ;
        RECT 104.045 43.930 104.565 44.470 ;
        RECT 105.210 44.150 105.505 44.480 ;
        RECT 105.685 44.150 106.100 44.480 ;
        RECT 106.270 43.980 106.445 44.650 ;
        RECT 106.615 44.150 106.855 44.800 ;
        RECT 107.085 44.735 107.415 45.170 ;
        RECT 107.585 44.780 107.755 45.390 ;
        RECT 107.035 44.650 107.415 44.735 ;
        RECT 107.925 44.650 108.255 45.175 ;
        RECT 108.515 44.860 108.725 45.390 ;
        RECT 109.000 44.940 109.785 45.110 ;
        RECT 109.955 44.940 110.360 45.110 ;
        RECT 107.035 44.610 107.260 44.650 ;
        RECT 107.035 44.030 107.205 44.610 ;
        RECT 107.925 44.480 108.125 44.650 ;
        RECT 109.000 44.480 109.170 44.940 ;
        RECT 107.375 44.150 108.125 44.480 ;
        RECT 108.295 44.150 109.170 44.480 ;
        RECT 107.035 43.980 107.250 44.030 ;
        RECT 103.355 42.840 104.565 43.930 ;
        RECT 105.205 43.620 106.100 43.950 ;
        RECT 106.270 43.790 106.855 43.980 ;
        RECT 107.035 43.900 107.425 43.980 ;
        RECT 105.205 43.450 106.410 43.620 ;
        RECT 105.205 43.020 105.535 43.450 ;
        RECT 105.715 42.840 105.910 43.280 ;
        RECT 106.080 43.020 106.410 43.450 ;
        RECT 106.580 43.020 106.855 43.790 ;
        RECT 107.095 43.055 107.425 43.900 ;
        RECT 107.935 43.945 108.125 44.150 ;
        RECT 107.595 42.840 107.765 43.850 ;
        RECT 107.935 43.570 108.830 43.945 ;
        RECT 107.935 43.010 108.275 43.570 ;
        RECT 108.505 42.840 108.820 43.340 ;
        RECT 109.000 43.310 109.170 44.150 ;
        RECT 109.340 44.440 109.805 44.770 ;
        RECT 110.190 44.710 110.360 44.940 ;
        RECT 110.540 44.890 110.910 45.390 ;
        RECT 111.230 44.940 111.905 45.110 ;
        RECT 112.100 44.940 112.435 45.110 ;
        RECT 109.340 43.480 109.660 44.440 ;
        RECT 110.190 44.410 111.020 44.710 ;
        RECT 109.830 43.510 110.020 44.230 ;
        RECT 110.190 43.340 110.360 44.410 ;
        RECT 110.820 44.380 111.020 44.410 ;
        RECT 110.530 44.160 110.700 44.230 ;
        RECT 111.230 44.160 111.400 44.940 ;
        RECT 112.265 44.800 112.435 44.940 ;
        RECT 112.605 44.930 112.855 45.390 ;
        RECT 110.530 43.990 111.400 44.160 ;
        RECT 111.570 44.520 112.095 44.740 ;
        RECT 112.265 44.670 112.490 44.800 ;
        RECT 110.530 43.900 111.040 43.990 ;
        RECT 109.000 43.140 109.885 43.310 ;
        RECT 110.110 43.010 110.360 43.340 ;
        RECT 110.530 42.840 110.700 43.640 ;
        RECT 110.870 43.285 111.040 43.900 ;
        RECT 111.570 43.820 111.740 44.520 ;
        RECT 111.210 43.455 111.740 43.820 ;
        RECT 111.910 43.755 112.150 44.350 ;
        RECT 112.320 43.565 112.490 44.670 ;
        RECT 112.660 43.810 112.940 44.760 ;
        RECT 112.185 43.435 112.490 43.565 ;
        RECT 110.870 43.115 111.975 43.285 ;
        RECT 112.185 43.010 112.435 43.435 ;
        RECT 112.605 42.840 112.870 43.300 ;
        RECT 113.110 43.010 113.295 45.130 ;
        RECT 113.465 45.010 113.795 45.390 ;
        RECT 113.965 44.840 114.135 45.130 ;
        RECT 114.395 44.845 119.740 45.390 ;
        RECT 119.915 44.845 125.260 45.390 ;
        RECT 113.470 44.670 114.135 44.840 ;
        RECT 113.470 43.680 113.700 44.670 ;
        RECT 113.870 43.850 114.220 44.500 ;
        RECT 115.980 44.015 116.320 44.845 ;
        RECT 113.470 43.510 114.135 43.680 ;
        RECT 113.465 42.840 113.795 43.340 ;
        RECT 113.965 43.010 114.135 43.510 ;
        RECT 117.800 43.275 118.150 44.525 ;
        RECT 121.500 44.015 121.840 44.845 ;
        RECT 125.435 44.620 128.945 45.390 ;
        RECT 129.115 44.665 129.405 45.390 ;
        RECT 129.575 44.845 134.920 45.390 ;
        RECT 123.320 43.275 123.670 44.525 ;
        RECT 125.435 44.100 127.085 44.620 ;
        RECT 127.255 43.930 128.945 44.450 ;
        RECT 131.160 44.015 131.500 44.845 ;
        RECT 135.095 44.620 138.605 45.390 ;
        RECT 138.775 44.640 139.985 45.390 ;
        RECT 140.155 44.640 141.365 45.390 ;
        RECT 114.395 42.840 119.740 43.275 ;
        RECT 119.915 42.840 125.260 43.275 ;
        RECT 125.435 42.840 128.945 43.930 ;
        RECT 129.115 42.840 129.405 44.005 ;
        RECT 132.980 43.275 133.330 44.525 ;
        RECT 135.095 44.100 136.745 44.620 ;
        RECT 136.915 43.930 138.605 44.450 ;
        RECT 138.775 44.100 139.295 44.640 ;
        RECT 139.465 43.930 139.985 44.470 ;
        RECT 129.575 42.840 134.920 43.275 ;
        RECT 135.095 42.840 138.605 43.930 ;
        RECT 138.775 42.840 139.985 43.930 ;
        RECT 140.155 43.930 140.675 44.470 ;
        RECT 140.845 44.100 141.365 44.640 ;
        RECT 140.155 42.840 141.365 43.930 ;
        RECT 103.270 42.670 141.450 42.840 ;
        RECT 61.590 42.380 84.770 42.540 ;
        RECT 61.760 42.370 84.770 42.380 ;
        RECT 63.410 41.290 83.400 41.610 ;
        RECT 103.355 41.580 104.565 42.670 ;
        RECT 104.735 41.580 108.245 42.670 ;
        RECT 108.875 42.115 109.480 42.670 ;
        RECT 109.655 42.160 110.135 42.500 ;
        RECT 110.305 42.125 110.560 42.670 ;
        RECT 108.875 42.015 109.490 42.115 ;
        RECT 109.305 41.990 109.490 42.015 ;
        RECT 63.400 41.120 83.400 41.290 ;
        RECT 61.660 40.100 62.520 40.110 ;
        RECT 61.560 39.840 62.520 40.100 ;
        RECT 61.560 39.160 62.570 39.840 ;
        RECT 63.400 39.510 63.570 41.120 ;
        RECT 64.250 40.550 72.290 40.720 ;
        RECT 73.340 40.550 81.380 40.720 ;
        RECT 63.910 40.140 64.080 40.490 ;
        RECT 72.460 40.140 72.630 40.490 ;
        RECT 73.000 40.140 73.170 40.490 ;
        RECT 81.550 40.140 81.720 40.490 ;
        RECT 82.060 40.460 83.400 41.120 ;
        RECT 103.355 40.870 103.875 41.410 ;
        RECT 104.045 41.040 104.565 41.580 ;
        RECT 104.735 40.890 106.385 41.410 ;
        RECT 106.555 41.060 108.245 41.580 ;
        RECT 108.875 41.395 109.135 41.845 ;
        RECT 109.305 41.745 109.635 41.990 ;
        RECT 109.805 41.670 110.560 41.920 ;
        RECT 110.730 41.800 111.005 42.500 ;
        RECT 109.790 41.635 110.560 41.670 ;
        RECT 109.775 41.625 110.560 41.635 ;
        RECT 109.770 41.610 110.665 41.625 ;
        RECT 109.750 41.595 110.665 41.610 ;
        RECT 109.730 41.585 110.665 41.595 ;
        RECT 109.705 41.575 110.665 41.585 ;
        RECT 109.635 41.545 110.665 41.575 ;
        RECT 109.615 41.515 110.665 41.545 ;
        RECT 109.595 41.485 110.665 41.515 ;
        RECT 109.565 41.460 110.665 41.485 ;
        RECT 109.530 41.425 110.665 41.460 ;
        RECT 109.500 41.420 110.665 41.425 ;
        RECT 109.500 41.415 109.890 41.420 ;
        RECT 109.500 41.405 109.865 41.415 ;
        RECT 109.500 41.400 109.850 41.405 ;
        RECT 109.500 41.395 109.835 41.400 ;
        RECT 108.875 41.390 109.835 41.395 ;
        RECT 108.875 41.380 109.825 41.390 ;
        RECT 108.875 41.375 109.815 41.380 ;
        RECT 108.875 41.365 109.805 41.375 ;
        RECT 108.875 41.355 109.800 41.365 ;
        RECT 108.875 41.350 109.795 41.355 ;
        RECT 108.875 41.335 109.785 41.350 ;
        RECT 108.875 41.320 109.780 41.335 ;
        RECT 108.875 41.295 109.770 41.320 ;
        RECT 108.875 41.225 109.765 41.295 ;
        RECT 64.250 39.910 72.290 40.080 ;
        RECT 73.340 39.910 81.380 40.080 ;
        RECT 82.060 39.510 82.910 40.460 ;
        RECT 103.355 40.120 104.565 40.870 ;
        RECT 104.735 40.120 108.245 40.890 ;
        RECT 108.875 40.670 109.425 41.055 ;
        RECT 109.595 40.500 109.765 41.225 ;
        RECT 108.875 40.330 109.765 40.500 ;
        RECT 109.935 40.825 110.265 41.250 ;
        RECT 110.435 41.025 110.665 41.420 ;
        RECT 109.935 40.340 110.155 40.825 ;
        RECT 110.835 40.770 111.005 41.800 ;
        RECT 110.325 40.120 110.575 40.660 ;
        RECT 110.745 40.290 111.005 40.770 ;
        RECT 111.175 41.700 111.445 42.470 ;
        RECT 111.615 41.890 111.945 42.670 ;
        RECT 112.150 42.065 112.335 42.470 ;
        RECT 112.505 42.245 112.840 42.670 ;
        RECT 112.150 41.890 112.815 42.065 ;
        RECT 111.175 41.530 112.305 41.700 ;
        RECT 111.175 40.620 111.345 41.530 ;
        RECT 111.515 40.780 111.875 41.360 ;
        RECT 112.055 41.030 112.305 41.530 ;
        RECT 112.475 40.860 112.815 41.890 ;
        RECT 113.025 41.700 113.355 42.485 ;
        RECT 113.025 41.530 113.705 41.700 ;
        RECT 113.885 41.530 114.215 42.670 ;
        RECT 114.395 41.580 116.065 42.670 ;
        RECT 113.015 41.110 113.365 41.360 ;
        RECT 113.535 40.930 113.705 41.530 ;
        RECT 113.875 41.110 114.225 41.360 ;
        RECT 112.130 40.690 112.815 40.860 ;
        RECT 111.175 40.290 111.435 40.620 ;
        RECT 111.645 40.120 111.920 40.600 ;
        RECT 112.130 40.290 112.335 40.690 ;
        RECT 112.505 40.120 112.840 40.520 ;
        RECT 113.035 40.120 113.275 40.930 ;
        RECT 113.445 40.290 113.775 40.930 ;
        RECT 113.945 40.120 114.215 40.930 ;
        RECT 114.395 40.890 115.145 41.410 ;
        RECT 115.315 41.060 116.065 41.580 ;
        RECT 116.235 41.505 116.525 42.670 ;
        RECT 116.695 42.235 122.040 42.670 ;
        RECT 122.215 42.235 127.560 42.670 ;
        RECT 127.735 42.235 133.080 42.670 ;
        RECT 133.255 42.235 138.600 42.670 ;
        RECT 114.395 40.120 116.065 40.890 ;
        RECT 116.235 40.120 116.525 40.845 ;
        RECT 118.280 40.665 118.620 41.495 ;
        RECT 120.100 40.985 120.450 42.235 ;
        RECT 123.800 40.665 124.140 41.495 ;
        RECT 125.620 40.985 125.970 42.235 ;
        RECT 129.320 40.665 129.660 41.495 ;
        RECT 131.140 40.985 131.490 42.235 ;
        RECT 134.840 40.665 135.180 41.495 ;
        RECT 136.660 40.985 137.010 42.235 ;
        RECT 138.775 41.580 139.985 42.670 ;
        RECT 138.775 40.870 139.295 41.410 ;
        RECT 139.465 41.040 139.985 41.580 ;
        RECT 140.155 41.580 141.365 42.670 ;
        RECT 140.155 41.040 140.675 41.580 ;
        RECT 140.845 40.870 141.365 41.410 ;
        RECT 116.695 40.120 122.040 40.665 ;
        RECT 122.215 40.120 127.560 40.665 ;
        RECT 127.735 40.120 133.080 40.665 ;
        RECT 133.255 40.120 138.600 40.665 ;
        RECT 138.775 40.120 139.985 40.870 ;
        RECT 140.155 40.120 141.365 40.870 ;
        RECT 103.270 39.950 141.450 40.120 ;
        RECT 63.400 39.350 82.910 39.510 ;
        RECT 63.400 39.340 82.230 39.350 ;
        RECT 103.355 39.200 104.565 39.950 ;
        RECT 104.735 39.405 110.080 39.950 ;
        RECT 110.255 39.405 115.600 39.950 ;
        RECT 115.775 39.405 121.120 39.950 ;
        RECT 121.295 39.405 126.640 39.950 ;
        RECT 61.560 38.970 84.300 39.160 ;
        RECT 61.560 38.800 84.740 38.970 ;
        RECT 61.560 37.190 61.900 38.800 ;
        RECT 62.625 38.230 72.665 38.400 ;
        RECT 73.805 38.230 83.845 38.400 ;
        RECT 62.240 37.820 62.410 38.170 ;
        RECT 72.880 37.820 73.050 38.170 ;
        RECT 73.420 37.820 73.590 38.170 ;
        RECT 84.060 37.820 84.230 38.170 ;
        RECT 62.625 37.590 72.665 37.760 ;
        RECT 73.805 37.590 83.845 37.760 ;
        RECT 84.570 37.190 84.740 38.800 ;
        RECT 103.355 38.660 103.875 39.200 ;
        RECT 104.045 38.490 104.565 39.030 ;
        RECT 106.320 38.575 106.660 39.405 ;
        RECT 103.355 37.400 104.565 38.490 ;
        RECT 108.140 37.835 108.490 39.085 ;
        RECT 111.840 38.575 112.180 39.405 ;
        RECT 113.660 37.835 114.010 39.085 ;
        RECT 117.360 38.575 117.700 39.405 ;
        RECT 119.180 37.835 119.530 39.085 ;
        RECT 122.880 38.575 123.220 39.405 ;
        RECT 126.815 39.180 128.485 39.950 ;
        RECT 129.115 39.225 129.405 39.950 ;
        RECT 129.575 39.405 134.920 39.950 ;
        RECT 124.700 37.835 125.050 39.085 ;
        RECT 126.815 38.660 127.565 39.180 ;
        RECT 127.735 38.490 128.485 39.010 ;
        RECT 131.160 38.575 131.500 39.405 ;
        RECT 135.095 39.180 138.605 39.950 ;
        RECT 138.775 39.200 139.985 39.950 ;
        RECT 140.155 39.200 141.365 39.950 ;
        RECT 104.735 37.400 110.080 37.835 ;
        RECT 110.255 37.400 115.600 37.835 ;
        RECT 115.775 37.400 121.120 37.835 ;
        RECT 121.295 37.400 126.640 37.835 ;
        RECT 126.815 37.400 128.485 38.490 ;
        RECT 129.115 37.400 129.405 38.565 ;
        RECT 132.980 37.835 133.330 39.085 ;
        RECT 135.095 38.660 136.745 39.180 ;
        RECT 136.915 38.490 138.605 39.010 ;
        RECT 138.775 38.660 139.295 39.200 ;
        RECT 139.465 38.490 139.985 39.030 ;
        RECT 129.575 37.400 134.920 37.835 ;
        RECT 135.095 37.400 138.605 38.490 ;
        RECT 138.775 37.400 139.985 38.490 ;
        RECT 140.155 38.490 140.675 39.030 ;
        RECT 140.845 38.660 141.365 39.200 ;
        RECT 140.155 37.400 141.365 38.490 ;
        RECT 103.270 37.230 141.450 37.400 ;
        RECT 61.560 37.030 84.740 37.190 ;
        RECT 61.730 37.020 84.740 37.030 ;
        RECT 63.450 36.010 83.440 36.330 ;
        RECT 103.355 36.140 104.565 37.230 ;
        RECT 104.735 36.140 106.405 37.230 ;
        RECT 106.665 36.485 106.935 37.230 ;
        RECT 107.565 37.225 113.840 37.230 ;
        RECT 107.105 36.315 107.395 37.055 ;
        RECT 107.565 36.500 107.820 37.225 ;
        RECT 108.005 36.330 108.265 37.055 ;
        RECT 108.435 36.500 108.680 37.225 ;
        RECT 108.865 36.330 109.125 37.055 ;
        RECT 109.295 36.500 109.540 37.225 ;
        RECT 109.725 36.330 109.985 37.055 ;
        RECT 110.155 36.500 110.400 37.225 ;
        RECT 110.570 36.330 110.830 37.055 ;
        RECT 111.000 36.500 111.260 37.225 ;
        RECT 111.430 36.330 111.690 37.055 ;
        RECT 111.860 36.500 112.120 37.225 ;
        RECT 112.290 36.330 112.550 37.055 ;
        RECT 112.720 36.500 112.980 37.225 ;
        RECT 113.150 36.330 113.410 37.055 ;
        RECT 113.580 36.430 113.840 37.225 ;
        RECT 108.005 36.315 113.410 36.330 ;
        RECT 63.440 35.840 83.440 36.010 ;
        RECT 61.700 34.820 62.560 34.830 ;
        RECT 61.600 34.560 62.560 34.820 ;
        RECT 61.600 33.880 62.610 34.560 ;
        RECT 63.440 34.230 63.610 35.840 ;
        RECT 64.290 35.270 72.330 35.440 ;
        RECT 73.380 35.270 81.420 35.440 ;
        RECT 63.950 34.860 64.120 35.210 ;
        RECT 72.500 34.860 72.670 35.210 ;
        RECT 73.040 34.860 73.210 35.210 ;
        RECT 81.590 34.860 81.760 35.210 ;
        RECT 82.100 35.180 83.440 35.840 ;
        RECT 103.355 35.430 103.875 35.970 ;
        RECT 104.045 35.600 104.565 36.140 ;
        RECT 104.735 35.450 105.485 35.970 ;
        RECT 105.655 35.620 106.405 36.140 ;
        RECT 106.665 36.090 113.410 36.315 ;
        RECT 106.665 35.500 107.830 36.090 ;
        RECT 114.010 35.920 114.260 37.055 ;
        RECT 114.440 36.420 114.700 37.230 ;
        RECT 114.875 35.920 115.120 37.060 ;
        RECT 115.300 36.420 115.595 37.230 ;
        RECT 116.235 36.065 116.525 37.230 ;
        RECT 116.695 36.140 118.365 37.230 ;
        RECT 119.085 36.485 119.355 37.230 ;
        RECT 119.985 37.225 126.260 37.230 ;
        RECT 119.525 36.315 119.815 37.055 ;
        RECT 119.985 36.500 120.240 37.225 ;
        RECT 120.425 36.330 120.685 37.055 ;
        RECT 120.855 36.500 121.100 37.225 ;
        RECT 121.285 36.330 121.545 37.055 ;
        RECT 121.715 36.500 121.960 37.225 ;
        RECT 122.145 36.330 122.405 37.055 ;
        RECT 122.575 36.500 122.820 37.225 ;
        RECT 122.990 36.330 123.250 37.055 ;
        RECT 123.420 36.500 123.680 37.225 ;
        RECT 123.850 36.330 124.110 37.055 ;
        RECT 124.280 36.500 124.540 37.225 ;
        RECT 124.710 36.330 124.970 37.055 ;
        RECT 125.140 36.500 125.400 37.225 ;
        RECT 125.570 36.330 125.830 37.055 ;
        RECT 126.000 36.430 126.260 37.225 ;
        RECT 120.425 36.315 125.830 36.330 ;
        RECT 108.000 35.670 115.120 35.920 ;
        RECT 64.290 34.630 72.330 34.800 ;
        RECT 73.380 34.630 81.420 34.800 ;
        RECT 82.100 34.230 82.950 35.180 ;
        RECT 103.355 34.680 104.565 35.430 ;
        RECT 104.735 34.680 106.405 35.450 ;
        RECT 106.665 35.330 113.410 35.500 ;
        RECT 106.665 34.680 106.965 35.160 ;
        RECT 107.135 34.875 107.395 35.330 ;
        RECT 107.565 34.680 107.825 35.160 ;
        RECT 108.005 34.875 108.265 35.330 ;
        RECT 108.435 34.680 108.685 35.160 ;
        RECT 108.865 34.875 109.125 35.330 ;
        RECT 109.295 34.680 109.545 35.160 ;
        RECT 109.725 34.875 109.985 35.330 ;
        RECT 110.155 34.680 110.400 35.160 ;
        RECT 110.570 34.875 110.845 35.330 ;
        RECT 111.015 34.680 111.260 35.160 ;
        RECT 111.430 34.875 111.690 35.330 ;
        RECT 111.860 34.680 112.120 35.160 ;
        RECT 112.290 34.875 112.550 35.330 ;
        RECT 112.720 34.680 112.980 35.160 ;
        RECT 113.150 34.875 113.410 35.330 ;
        RECT 113.580 34.680 113.840 35.240 ;
        RECT 114.010 34.860 114.260 35.670 ;
        RECT 114.440 34.680 114.700 35.205 ;
        RECT 114.870 34.860 115.120 35.670 ;
        RECT 115.290 35.360 115.605 35.920 ;
        RECT 116.695 35.450 117.445 35.970 ;
        RECT 117.615 35.620 118.365 36.140 ;
        RECT 119.085 36.090 125.830 36.315 ;
        RECT 119.085 35.500 120.250 36.090 ;
        RECT 126.430 35.920 126.680 37.055 ;
        RECT 126.860 36.420 127.120 37.230 ;
        RECT 127.295 35.920 127.540 37.060 ;
        RECT 127.720 36.420 128.015 37.230 ;
        RECT 128.195 36.795 133.540 37.230 ;
        RECT 133.715 36.795 139.060 37.230 ;
        RECT 120.420 35.670 127.540 35.920 ;
        RECT 115.300 34.680 115.605 35.190 ;
        RECT 116.235 34.680 116.525 35.405 ;
        RECT 116.695 34.680 118.365 35.450 ;
        RECT 119.085 35.330 125.830 35.500 ;
        RECT 119.085 34.680 119.385 35.160 ;
        RECT 119.555 34.875 119.815 35.330 ;
        RECT 119.985 34.680 120.245 35.160 ;
        RECT 120.425 34.875 120.685 35.330 ;
        RECT 120.855 34.680 121.105 35.160 ;
        RECT 121.285 34.875 121.545 35.330 ;
        RECT 121.715 34.680 121.965 35.160 ;
        RECT 122.145 34.875 122.405 35.330 ;
        RECT 122.575 34.680 122.820 35.160 ;
        RECT 122.990 34.875 123.265 35.330 ;
        RECT 123.435 34.680 123.680 35.160 ;
        RECT 123.850 34.875 124.110 35.330 ;
        RECT 124.280 34.680 124.540 35.160 ;
        RECT 124.710 34.875 124.970 35.330 ;
        RECT 125.140 34.680 125.400 35.160 ;
        RECT 125.570 34.875 125.830 35.330 ;
        RECT 126.000 34.680 126.260 35.240 ;
        RECT 126.430 34.860 126.680 35.670 ;
        RECT 126.860 34.680 127.120 35.205 ;
        RECT 127.290 34.860 127.540 35.670 ;
        RECT 127.710 35.360 128.025 35.920 ;
        RECT 129.780 35.225 130.120 36.055 ;
        RECT 131.600 35.545 131.950 36.795 ;
        RECT 135.300 35.225 135.640 36.055 ;
        RECT 137.120 35.545 137.470 36.795 ;
        RECT 140.155 36.140 141.365 37.230 ;
        RECT 140.155 35.600 140.675 36.140 ;
        RECT 140.845 35.430 141.365 35.970 ;
        RECT 127.720 34.680 128.025 35.190 ;
        RECT 128.195 34.680 133.540 35.225 ;
        RECT 133.715 34.680 139.060 35.225 ;
        RECT 140.155 34.680 141.365 35.430 ;
        RECT 103.270 34.510 141.450 34.680 ;
        RECT 63.440 34.070 82.950 34.230 ;
        RECT 63.440 34.060 82.270 34.070 ;
        RECT 61.600 33.690 84.340 33.880 ;
        RECT 103.355 33.760 104.565 34.510 ;
        RECT 104.735 33.965 110.080 34.510 ;
        RECT 110.255 33.965 115.600 34.510 ;
        RECT 116.700 34.005 117.035 34.510 ;
        RECT 61.600 33.520 84.780 33.690 ;
        RECT 61.600 31.910 61.940 33.520 ;
        RECT 62.665 32.950 72.705 33.120 ;
        RECT 73.845 32.950 83.885 33.120 ;
        RECT 62.280 32.540 62.450 32.890 ;
        RECT 72.920 32.540 73.090 32.890 ;
        RECT 73.460 32.540 73.630 32.890 ;
        RECT 84.100 32.540 84.270 32.890 ;
        RECT 62.665 32.310 72.705 32.480 ;
        RECT 73.845 32.310 83.885 32.480 ;
        RECT 84.610 31.910 84.780 33.520 ;
        RECT 103.355 33.220 103.875 33.760 ;
        RECT 104.045 33.050 104.565 33.590 ;
        RECT 106.320 33.135 106.660 33.965 ;
        RECT 103.355 31.960 104.565 33.050 ;
        RECT 108.140 32.395 108.490 33.645 ;
        RECT 111.840 33.135 112.180 33.965 ;
        RECT 117.205 33.940 117.445 34.315 ;
        RECT 117.725 34.180 117.895 34.325 ;
        RECT 117.725 33.985 118.100 34.180 ;
        RECT 118.460 34.015 118.855 34.510 ;
        RECT 113.660 32.395 114.010 33.645 ;
        RECT 116.755 32.980 117.055 33.830 ;
        RECT 117.225 33.790 117.445 33.940 ;
        RECT 117.225 33.460 117.760 33.790 ;
        RECT 117.930 33.650 118.100 33.985 ;
        RECT 119.025 33.820 119.265 34.340 ;
        RECT 119.505 33.855 119.835 34.290 ;
        RECT 120.005 33.900 120.175 34.510 ;
        RECT 117.225 32.810 117.460 33.460 ;
        RECT 117.930 33.290 118.915 33.650 ;
        RECT 116.785 32.580 117.460 32.810 ;
        RECT 117.630 33.270 118.915 33.290 ;
        RECT 117.630 33.120 118.490 33.270 ;
        RECT 119.090 33.150 119.265 33.820 ;
        RECT 104.735 31.960 110.080 32.395 ;
        RECT 110.255 31.960 115.600 32.395 ;
        RECT 116.785 32.150 116.955 32.580 ;
        RECT 117.125 31.960 117.455 32.410 ;
        RECT 117.630 32.175 117.915 33.120 ;
        RECT 119.055 33.015 119.265 33.150 ;
        RECT 119.455 33.770 119.835 33.855 ;
        RECT 120.345 33.770 120.675 34.295 ;
        RECT 120.935 33.980 121.145 34.510 ;
        RECT 121.420 34.060 122.205 34.230 ;
        RECT 122.375 34.060 122.780 34.230 ;
        RECT 119.455 33.730 119.680 33.770 ;
        RECT 119.455 33.150 119.625 33.730 ;
        RECT 120.345 33.600 120.545 33.770 ;
        RECT 121.420 33.600 121.590 34.060 ;
        RECT 119.795 33.270 120.545 33.600 ;
        RECT 120.715 33.270 121.590 33.600 ;
        RECT 119.455 33.100 119.670 33.150 ;
        RECT 119.455 33.020 119.845 33.100 ;
        RECT 118.090 32.640 118.785 32.950 ;
        RECT 118.095 31.960 118.780 32.430 ;
        RECT 118.960 32.230 119.265 33.015 ;
        RECT 119.515 32.175 119.845 33.020 ;
        RECT 120.355 33.065 120.545 33.270 ;
        RECT 120.015 31.960 120.185 32.970 ;
        RECT 120.355 32.690 121.250 33.065 ;
        RECT 120.355 32.130 120.695 32.690 ;
        RECT 120.925 31.960 121.240 32.460 ;
        RECT 121.420 32.430 121.590 33.270 ;
        RECT 121.760 33.560 122.225 33.890 ;
        RECT 122.610 33.830 122.780 34.060 ;
        RECT 122.960 34.010 123.330 34.510 ;
        RECT 123.650 34.060 124.325 34.230 ;
        RECT 124.520 34.060 124.855 34.230 ;
        RECT 121.760 32.600 122.080 33.560 ;
        RECT 122.610 33.530 123.440 33.830 ;
        RECT 122.250 32.630 122.440 33.350 ;
        RECT 122.610 32.460 122.780 33.530 ;
        RECT 123.240 33.500 123.440 33.530 ;
        RECT 122.950 33.280 123.120 33.350 ;
        RECT 123.650 33.280 123.820 34.060 ;
        RECT 124.685 33.920 124.855 34.060 ;
        RECT 125.025 34.050 125.275 34.510 ;
        RECT 122.950 33.110 123.820 33.280 ;
        RECT 123.990 33.640 124.515 33.860 ;
        RECT 124.685 33.790 124.910 33.920 ;
        RECT 122.950 33.020 123.460 33.110 ;
        RECT 121.420 32.260 122.305 32.430 ;
        RECT 122.530 32.130 122.780 32.460 ;
        RECT 122.950 31.960 123.120 32.760 ;
        RECT 123.290 32.405 123.460 33.020 ;
        RECT 123.990 32.940 124.160 33.640 ;
        RECT 123.630 32.575 124.160 32.940 ;
        RECT 124.330 32.875 124.570 33.470 ;
        RECT 124.740 32.685 124.910 33.790 ;
        RECT 125.080 32.930 125.360 33.880 ;
        RECT 124.605 32.555 124.910 32.685 ;
        RECT 123.290 32.235 124.395 32.405 ;
        RECT 124.605 32.130 124.855 32.555 ;
        RECT 125.025 31.960 125.290 32.420 ;
        RECT 125.530 32.130 125.715 34.250 ;
        RECT 125.885 34.130 126.215 34.510 ;
        RECT 126.385 33.960 126.555 34.250 ;
        RECT 125.890 33.790 126.555 33.960 ;
        RECT 126.815 33.835 127.075 34.340 ;
        RECT 127.255 34.130 127.585 34.510 ;
        RECT 127.765 33.960 127.935 34.340 ;
        RECT 125.890 32.800 126.120 33.790 ;
        RECT 126.290 32.970 126.640 33.620 ;
        RECT 126.815 33.035 126.985 33.835 ;
        RECT 127.270 33.790 127.935 33.960 ;
        RECT 127.270 33.535 127.440 33.790 ;
        RECT 129.115 33.785 129.405 34.510 ;
        RECT 129.660 34.010 130.155 34.340 ;
        RECT 127.155 33.205 127.440 33.535 ;
        RECT 127.675 33.240 128.005 33.610 ;
        RECT 127.270 33.060 127.440 33.205 ;
        RECT 125.890 32.630 126.555 32.800 ;
        RECT 125.885 31.960 126.215 32.460 ;
        RECT 126.385 32.130 126.555 32.630 ;
        RECT 126.815 32.130 127.085 33.035 ;
        RECT 127.270 32.890 127.935 33.060 ;
        RECT 127.255 31.960 127.585 32.720 ;
        RECT 127.765 32.130 127.935 32.890 ;
        RECT 129.115 31.960 129.405 33.125 ;
        RECT 129.575 32.520 129.815 33.830 ;
        RECT 129.985 33.100 130.155 34.010 ;
        RECT 130.375 33.270 130.725 34.235 ;
        RECT 130.905 33.270 131.205 34.240 ;
        RECT 131.385 33.270 131.665 34.240 ;
        RECT 131.845 33.710 132.115 34.510 ;
        RECT 132.285 33.790 132.625 34.300 ;
        RECT 132.800 34.005 133.135 34.510 ;
        RECT 133.305 33.940 133.545 34.315 ;
        RECT 133.825 34.180 133.995 34.325 ;
        RECT 133.825 33.985 134.200 34.180 ;
        RECT 134.560 34.015 134.955 34.510 ;
        RECT 131.860 33.270 132.190 33.520 ;
        RECT 131.860 33.100 132.175 33.270 ;
        RECT 129.985 32.930 132.175 33.100 ;
        RECT 129.580 31.960 129.915 32.340 ;
        RECT 130.085 32.130 130.335 32.930 ;
        RECT 130.555 31.960 130.885 32.680 ;
        RECT 131.070 32.130 131.320 32.930 ;
        RECT 131.785 31.960 132.115 32.760 ;
        RECT 132.365 32.390 132.625 33.790 ;
        RECT 132.855 32.980 133.155 33.830 ;
        RECT 133.325 33.790 133.545 33.940 ;
        RECT 133.325 33.460 133.860 33.790 ;
        RECT 134.030 33.650 134.200 33.985 ;
        RECT 135.125 33.820 135.365 34.340 ;
        RECT 133.325 32.810 133.560 33.460 ;
        RECT 134.030 33.290 135.015 33.650 ;
        RECT 132.285 32.130 132.625 32.390 ;
        RECT 132.885 32.580 133.560 32.810 ;
        RECT 133.730 33.270 135.015 33.290 ;
        RECT 133.730 33.120 134.590 33.270 ;
        RECT 135.190 33.150 135.365 33.820 ;
        RECT 132.885 32.150 133.055 32.580 ;
        RECT 133.225 31.960 133.555 32.410 ;
        RECT 133.730 32.175 134.015 33.120 ;
        RECT 135.155 33.015 135.365 33.150 ;
        RECT 134.190 32.640 134.885 32.950 ;
        RECT 134.195 31.960 134.880 32.430 ;
        RECT 135.060 32.230 135.365 33.015 ;
        RECT 135.555 33.835 135.815 34.340 ;
        RECT 135.995 34.130 136.325 34.510 ;
        RECT 136.505 33.960 136.675 34.340 ;
        RECT 135.555 33.035 135.725 33.835 ;
        RECT 136.010 33.790 136.675 33.960 ;
        RECT 136.010 33.535 136.180 33.790 ;
        RECT 136.935 33.740 139.525 34.510 ;
        RECT 140.155 33.760 141.365 34.510 ;
        RECT 135.895 33.205 136.180 33.535 ;
        RECT 136.415 33.240 136.745 33.610 ;
        RECT 136.935 33.220 138.145 33.740 ;
        RECT 136.010 33.060 136.180 33.205 ;
        RECT 135.555 32.130 135.825 33.035 ;
        RECT 136.010 32.890 136.675 33.060 ;
        RECT 138.315 33.050 139.525 33.570 ;
        RECT 135.995 31.960 136.325 32.720 ;
        RECT 136.505 32.130 136.675 32.890 ;
        RECT 136.935 31.960 139.525 33.050 ;
        RECT 140.155 33.050 140.675 33.590 ;
        RECT 140.845 33.220 141.365 33.760 ;
        RECT 140.155 31.960 141.365 33.050 ;
        RECT 61.600 31.750 84.780 31.910 ;
        RECT 103.270 31.790 141.450 31.960 ;
        RECT 61.770 31.740 84.780 31.750 ;
        RECT 103.355 30.700 104.565 31.790 ;
        RECT 104.735 30.700 107.325 31.790 ;
        RECT 103.355 29.990 103.875 30.530 ;
        RECT 104.045 30.160 104.565 30.700 ;
        RECT 104.735 30.010 105.945 30.530 ;
        RECT 106.115 30.180 107.325 30.700 ;
        RECT 107.505 30.820 107.835 31.605 ;
        RECT 107.505 30.650 108.185 30.820 ;
        RECT 108.365 30.650 108.695 31.790 ;
        RECT 108.965 31.120 109.135 31.620 ;
        RECT 109.305 31.290 109.635 31.790 ;
        RECT 108.965 30.950 109.630 31.120 ;
        RECT 107.495 30.230 107.845 30.480 ;
        RECT 108.015 30.050 108.185 30.650 ;
        RECT 108.355 30.230 108.705 30.480 ;
        RECT 108.880 30.130 109.230 30.780 ;
        RECT 103.355 29.240 104.565 29.990 ;
        RECT 104.735 29.240 107.325 30.010 ;
        RECT 107.515 29.240 107.755 30.050 ;
        RECT 107.925 29.410 108.255 30.050 ;
        RECT 108.425 29.240 108.695 30.050 ;
        RECT 109.400 29.960 109.630 30.950 ;
        RECT 108.965 29.790 109.630 29.960 ;
        RECT 108.965 29.500 109.135 29.790 ;
        RECT 109.305 29.240 109.635 29.620 ;
        RECT 109.805 29.500 109.990 31.620 ;
        RECT 110.230 31.330 110.495 31.790 ;
        RECT 110.665 31.195 110.915 31.620 ;
        RECT 111.125 31.345 112.230 31.515 ;
        RECT 110.610 31.065 110.915 31.195 ;
        RECT 110.160 29.870 110.440 30.820 ;
        RECT 110.610 29.960 110.780 31.065 ;
        RECT 110.950 30.280 111.190 30.875 ;
        RECT 111.360 30.810 111.890 31.175 ;
        RECT 111.360 30.110 111.530 30.810 ;
        RECT 112.060 30.730 112.230 31.345 ;
        RECT 112.400 30.990 112.570 31.790 ;
        RECT 112.740 31.290 112.990 31.620 ;
        RECT 113.215 31.320 114.100 31.490 ;
        RECT 112.060 30.640 112.570 30.730 ;
        RECT 110.610 29.830 110.835 29.960 ;
        RECT 111.005 29.890 111.530 30.110 ;
        RECT 111.700 30.470 112.570 30.640 ;
        RECT 110.245 29.240 110.495 29.700 ;
        RECT 110.665 29.690 110.835 29.830 ;
        RECT 111.700 29.690 111.870 30.470 ;
        RECT 112.400 30.400 112.570 30.470 ;
        RECT 112.080 30.220 112.280 30.250 ;
        RECT 112.740 30.220 112.910 31.290 ;
        RECT 113.080 30.400 113.270 31.120 ;
        RECT 112.080 29.920 112.910 30.220 ;
        RECT 113.440 30.190 113.760 31.150 ;
        RECT 110.665 29.520 111.000 29.690 ;
        RECT 111.195 29.520 111.870 29.690 ;
        RECT 112.190 29.240 112.560 29.740 ;
        RECT 112.740 29.690 112.910 29.920 ;
        RECT 113.295 29.860 113.760 30.190 ;
        RECT 113.930 30.480 114.100 31.320 ;
        RECT 114.280 31.290 114.595 31.790 ;
        RECT 114.825 31.060 115.165 31.620 ;
        RECT 114.270 30.685 115.165 31.060 ;
        RECT 115.335 30.780 115.505 31.790 ;
        RECT 114.975 30.480 115.165 30.685 ;
        RECT 115.675 30.730 116.005 31.575 ;
        RECT 115.675 30.650 116.065 30.730 ;
        RECT 115.850 30.600 116.065 30.650 ;
        RECT 116.235 30.625 116.525 31.790 ;
        RECT 116.695 30.700 118.365 31.790 ;
        RECT 113.930 30.150 114.805 30.480 ;
        RECT 114.975 30.150 115.725 30.480 ;
        RECT 113.930 29.690 114.100 30.150 ;
        RECT 114.975 29.980 115.175 30.150 ;
        RECT 115.895 30.020 116.065 30.600 ;
        RECT 115.840 29.980 116.065 30.020 ;
        RECT 112.740 29.520 113.145 29.690 ;
        RECT 113.315 29.520 114.100 29.690 ;
        RECT 114.375 29.240 114.585 29.770 ;
        RECT 114.845 29.455 115.175 29.980 ;
        RECT 115.685 29.895 116.065 29.980 ;
        RECT 116.695 30.010 117.445 30.530 ;
        RECT 117.615 30.180 118.365 30.700 ;
        RECT 119.210 30.690 119.540 31.790 ;
        RECT 120.015 31.190 120.340 31.620 ;
        RECT 120.510 31.370 120.840 31.790 ;
        RECT 121.585 31.360 121.995 31.790 ;
        RECT 120.015 31.020 121.995 31.190 ;
        RECT 120.015 30.610 120.720 31.020 ;
        RECT 118.995 30.230 119.640 30.440 ;
        RECT 119.810 30.230 120.380 30.440 ;
        RECT 115.345 29.240 115.515 29.850 ;
        RECT 115.685 29.460 116.015 29.895 ;
        RECT 116.235 29.240 116.525 29.965 ;
        RECT 116.695 29.240 118.365 30.010 ;
        RECT 119.150 29.890 120.320 30.060 ;
        RECT 119.150 29.425 119.480 29.890 ;
        RECT 119.650 29.240 119.820 29.710 ;
        RECT 119.990 29.410 120.320 29.890 ;
        RECT 120.550 29.410 120.720 30.610 ;
        RECT 120.890 30.680 121.515 30.850 ;
        RECT 120.890 29.980 121.060 30.680 ;
        RECT 121.730 30.480 121.995 31.020 ;
        RECT 122.165 30.635 122.505 31.620 ;
        RECT 122.675 30.970 123.020 31.790 ;
        RECT 121.230 30.150 121.560 30.480 ;
        RECT 121.730 30.150 122.080 30.480 ;
        RECT 122.250 29.980 122.505 30.635 ;
        RECT 122.675 30.230 123.020 30.800 ;
        RECT 123.190 30.480 123.365 31.580 ;
        RECT 123.535 31.210 123.865 31.445 ;
        RECT 124.155 31.390 124.555 31.790 ;
        RECT 125.425 31.390 125.755 31.790 ;
        RECT 123.535 31.040 125.615 31.210 ;
        RECT 123.535 30.650 124.090 31.040 ;
        RECT 123.190 30.230 123.750 30.480 ;
        RECT 123.920 30.400 124.090 30.650 ;
        RECT 124.260 30.650 125.275 30.870 ;
        RECT 125.445 30.770 125.615 31.040 ;
        RECT 125.925 30.950 126.185 31.620 ;
        RECT 126.365 30.980 126.660 31.790 ;
        RECT 124.260 30.510 124.535 30.650 ;
        RECT 125.445 30.600 125.840 30.770 ;
        RECT 123.920 30.230 124.115 30.400 ;
        RECT 120.890 29.810 121.430 29.980 ;
        RECT 121.260 29.605 121.430 29.810 ;
        RECT 121.710 29.240 121.880 29.980 ;
        RECT 122.145 29.605 122.505 29.980 ;
        RECT 122.675 29.880 123.775 30.060 ;
        RECT 122.275 29.580 122.445 29.605 ;
        RECT 122.675 29.475 123.015 29.880 ;
        RECT 123.185 29.240 123.355 29.710 ;
        RECT 123.525 29.475 123.775 29.880 ;
        RECT 123.945 29.845 124.115 30.230 ;
        RECT 123.945 29.475 124.195 29.845 ;
        RECT 124.365 29.720 124.535 30.510 ;
        RECT 124.705 30.060 124.880 30.255 ;
        RECT 125.050 30.230 125.500 30.430 ;
        RECT 125.670 30.150 125.840 30.600 ;
        RECT 124.705 29.890 125.200 30.060 ;
        RECT 126.010 29.980 126.185 30.950 ;
        RECT 126.840 30.480 127.085 31.620 ;
        RECT 127.260 30.980 127.520 31.790 ;
        RECT 128.120 31.785 134.395 31.790 ;
        RECT 127.700 30.480 127.950 31.615 ;
        RECT 128.120 30.990 128.380 31.785 ;
        RECT 128.550 30.890 128.810 31.615 ;
        RECT 128.980 31.060 129.240 31.785 ;
        RECT 129.410 30.890 129.670 31.615 ;
        RECT 129.840 31.060 130.100 31.785 ;
        RECT 130.270 30.890 130.530 31.615 ;
        RECT 130.700 31.060 130.960 31.785 ;
        RECT 131.130 30.890 131.390 31.615 ;
        RECT 131.560 31.060 131.805 31.785 ;
        RECT 131.975 30.890 132.235 31.615 ;
        RECT 132.420 31.060 132.665 31.785 ;
        RECT 132.835 30.890 133.095 31.615 ;
        RECT 133.280 31.060 133.525 31.785 ;
        RECT 133.695 30.890 133.955 31.615 ;
        RECT 134.140 31.060 134.395 31.785 ;
        RECT 128.550 30.875 133.955 30.890 ;
        RECT 134.565 30.875 134.855 31.615 ;
        RECT 135.025 31.045 135.295 31.790 ;
        RECT 128.550 30.650 135.295 30.875 ;
        RECT 135.555 30.700 139.065 31.790 ;
        RECT 124.980 29.750 125.200 29.890 ;
        RECT 124.365 29.550 124.810 29.720 ;
        RECT 124.980 29.580 125.205 29.750 ;
        RECT 124.980 29.535 125.200 29.580 ;
        RECT 125.480 29.240 125.650 29.905 ;
        RECT 125.845 29.410 126.185 29.980 ;
        RECT 126.355 29.920 126.670 30.480 ;
        RECT 126.840 30.230 133.960 30.480 ;
        RECT 126.355 29.240 126.660 29.750 ;
        RECT 126.840 29.420 127.090 30.230 ;
        RECT 127.260 29.240 127.520 29.765 ;
        RECT 127.700 29.420 127.950 30.230 ;
        RECT 134.130 30.060 135.295 30.650 ;
        RECT 128.550 29.890 135.295 30.060 ;
        RECT 135.555 30.010 137.205 30.530 ;
        RECT 137.375 30.180 139.065 30.700 ;
        RECT 140.155 30.700 141.365 31.790 ;
        RECT 140.155 30.160 140.675 30.700 ;
        RECT 128.120 29.240 128.380 29.800 ;
        RECT 128.550 29.435 128.810 29.890 ;
        RECT 128.980 29.240 129.240 29.720 ;
        RECT 129.410 29.435 129.670 29.890 ;
        RECT 129.840 29.240 130.100 29.720 ;
        RECT 130.270 29.435 130.530 29.890 ;
        RECT 130.700 29.240 130.945 29.720 ;
        RECT 131.115 29.435 131.390 29.890 ;
        RECT 131.560 29.240 131.805 29.720 ;
        RECT 131.975 29.435 132.235 29.890 ;
        RECT 132.415 29.240 132.665 29.720 ;
        RECT 132.835 29.435 133.095 29.890 ;
        RECT 133.275 29.240 133.525 29.720 ;
        RECT 133.695 29.435 133.955 29.890 ;
        RECT 134.135 29.240 134.395 29.720 ;
        RECT 134.565 29.435 134.825 29.890 ;
        RECT 134.995 29.240 135.295 29.720 ;
        RECT 135.555 29.240 139.065 30.010 ;
        RECT 140.845 29.990 141.365 30.530 ;
        RECT 140.155 29.240 141.365 29.990 ;
        RECT 103.270 29.070 141.450 29.240 ;
        RECT 103.355 28.320 104.565 29.070 ;
        RECT 103.355 27.780 103.875 28.320 ;
        RECT 104.745 28.260 105.015 29.070 ;
        RECT 105.185 28.260 105.515 28.900 ;
        RECT 105.685 28.260 105.925 29.070 ;
        RECT 106.205 28.520 106.375 28.810 ;
        RECT 106.545 28.690 106.875 29.070 ;
        RECT 106.205 28.350 106.870 28.520 ;
        RECT 104.045 27.610 104.565 28.150 ;
        RECT 104.735 27.830 105.085 28.080 ;
        RECT 105.255 27.660 105.425 28.260 ;
        RECT 105.595 27.830 105.945 28.080 ;
        RECT 103.355 26.520 104.565 27.610 ;
        RECT 104.745 26.520 105.075 27.660 ;
        RECT 105.255 27.490 105.935 27.660 ;
        RECT 106.120 27.530 106.470 28.180 ;
        RECT 105.605 26.705 105.935 27.490 ;
        RECT 106.640 27.360 106.870 28.350 ;
        RECT 106.205 27.190 106.870 27.360 ;
        RECT 106.205 26.690 106.375 27.190 ;
        RECT 106.545 26.520 106.875 27.020 ;
        RECT 107.045 26.690 107.230 28.810 ;
        RECT 107.485 28.610 107.735 29.070 ;
        RECT 107.905 28.620 108.240 28.790 ;
        RECT 108.435 28.620 109.110 28.790 ;
        RECT 107.905 28.480 108.075 28.620 ;
        RECT 107.400 27.490 107.680 28.440 ;
        RECT 107.850 28.350 108.075 28.480 ;
        RECT 107.850 27.245 108.020 28.350 ;
        RECT 108.245 28.200 108.770 28.420 ;
        RECT 108.190 27.435 108.430 28.030 ;
        RECT 108.600 27.500 108.770 28.200 ;
        RECT 108.940 27.840 109.110 28.620 ;
        RECT 109.430 28.570 109.800 29.070 ;
        RECT 109.980 28.620 110.385 28.790 ;
        RECT 110.555 28.620 111.340 28.790 ;
        RECT 109.980 28.390 110.150 28.620 ;
        RECT 109.320 28.090 110.150 28.390 ;
        RECT 110.535 28.120 111.000 28.450 ;
        RECT 109.320 28.060 109.520 28.090 ;
        RECT 109.640 27.840 109.810 27.910 ;
        RECT 108.940 27.670 109.810 27.840 ;
        RECT 109.300 27.580 109.810 27.670 ;
        RECT 107.850 27.115 108.155 27.245 ;
        RECT 108.600 27.135 109.130 27.500 ;
        RECT 107.470 26.520 107.735 26.980 ;
        RECT 107.905 26.690 108.155 27.115 ;
        RECT 109.300 26.965 109.470 27.580 ;
        RECT 108.365 26.795 109.470 26.965 ;
        RECT 109.640 26.520 109.810 27.320 ;
        RECT 109.980 27.020 110.150 28.090 ;
        RECT 110.320 27.190 110.510 27.910 ;
        RECT 110.680 27.160 111.000 28.120 ;
        RECT 111.170 28.160 111.340 28.620 ;
        RECT 111.615 28.540 111.825 29.070 ;
        RECT 112.085 28.330 112.415 28.855 ;
        RECT 112.585 28.460 112.755 29.070 ;
        RECT 112.925 28.415 113.255 28.850 ;
        RECT 112.925 28.330 113.305 28.415 ;
        RECT 112.215 28.160 112.415 28.330 ;
        RECT 113.080 28.290 113.305 28.330 ;
        RECT 111.170 27.830 112.045 28.160 ;
        RECT 112.215 27.830 112.965 28.160 ;
        RECT 109.980 26.690 110.230 27.020 ;
        RECT 111.170 26.990 111.340 27.830 ;
        RECT 112.215 27.625 112.405 27.830 ;
        RECT 113.135 27.710 113.305 28.290 ;
        RECT 113.475 28.235 113.765 29.070 ;
        RECT 113.935 28.670 114.890 28.840 ;
        RECT 115.305 28.680 115.635 29.070 ;
        RECT 113.935 27.790 114.105 28.670 ;
        RECT 115.805 28.500 115.975 28.820 ;
        RECT 116.145 28.680 116.475 29.070 ;
        RECT 114.275 28.330 116.525 28.500 ;
        RECT 114.275 27.830 114.505 28.330 ;
        RECT 114.675 27.910 115.050 28.080 ;
        RECT 113.090 27.660 113.305 27.710 ;
        RECT 111.510 27.250 112.405 27.625 ;
        RECT 112.915 27.580 113.305 27.660 ;
        RECT 113.475 27.620 114.105 27.790 ;
        RECT 114.880 27.710 115.050 27.910 ;
        RECT 115.220 27.880 115.770 28.080 ;
        RECT 115.940 27.710 116.185 28.160 ;
        RECT 110.455 26.820 111.340 26.990 ;
        RECT 111.520 26.520 111.835 27.020 ;
        RECT 112.065 26.690 112.405 27.250 ;
        RECT 112.575 26.520 112.745 27.530 ;
        RECT 112.915 26.735 113.245 27.580 ;
        RECT 113.475 26.690 113.795 27.620 ;
        RECT 114.880 27.540 116.185 27.710 ;
        RECT 116.355 27.370 116.525 28.330 ;
        RECT 116.695 28.300 118.365 29.070 ;
        RECT 118.545 28.345 118.875 28.855 ;
        RECT 119.045 28.670 119.375 29.070 ;
        RECT 120.425 28.500 120.755 28.840 ;
        RECT 120.925 28.670 121.255 29.070 ;
        RECT 121.845 28.520 122.015 28.810 ;
        RECT 122.185 28.690 122.515 29.070 ;
        RECT 116.695 27.780 117.445 28.300 ;
        RECT 117.615 27.610 118.365 28.130 ;
        RECT 113.975 27.200 115.215 27.370 ;
        RECT 113.975 26.690 114.375 27.200 ;
        RECT 114.545 26.520 114.715 27.030 ;
        RECT 114.885 26.690 115.215 27.200 ;
        RECT 115.385 26.520 115.555 27.370 ;
        RECT 116.145 26.690 116.525 27.370 ;
        RECT 116.695 26.520 118.365 27.610 ;
        RECT 118.545 27.710 118.735 28.345 ;
        RECT 119.045 28.330 121.410 28.500 ;
        RECT 121.845 28.350 122.510 28.520 ;
        RECT 119.045 28.160 119.215 28.330 ;
        RECT 118.905 27.830 119.215 28.160 ;
        RECT 119.385 27.830 119.690 28.160 ;
        RECT 118.545 27.580 118.765 27.710 ;
        RECT 118.545 26.730 118.875 27.580 ;
        RECT 119.045 26.520 119.295 27.660 ;
        RECT 119.475 27.500 119.690 27.830 ;
        RECT 119.865 27.500 120.150 28.160 ;
        RECT 120.345 27.500 120.610 28.160 ;
        RECT 120.825 27.500 121.070 28.160 ;
        RECT 121.240 27.330 121.410 28.330 ;
        RECT 121.760 27.530 122.110 28.180 ;
        RECT 122.280 27.360 122.510 28.350 ;
        RECT 119.485 27.160 120.775 27.330 ;
        RECT 119.485 26.740 119.735 27.160 ;
        RECT 119.965 26.520 120.295 26.990 ;
        RECT 120.525 26.740 120.775 27.160 ;
        RECT 120.955 27.160 121.410 27.330 ;
        RECT 121.845 27.190 122.510 27.360 ;
        RECT 120.955 26.730 121.285 27.160 ;
        RECT 121.845 26.690 122.015 27.190 ;
        RECT 122.185 26.520 122.515 27.020 ;
        RECT 122.685 26.690 122.870 28.810 ;
        RECT 123.125 28.610 123.375 29.070 ;
        RECT 123.545 28.620 123.880 28.790 ;
        RECT 124.075 28.620 124.750 28.790 ;
        RECT 123.545 28.480 123.715 28.620 ;
        RECT 123.040 27.490 123.320 28.440 ;
        RECT 123.490 28.350 123.715 28.480 ;
        RECT 123.490 27.245 123.660 28.350 ;
        RECT 123.885 28.200 124.410 28.420 ;
        RECT 123.830 27.435 124.070 28.030 ;
        RECT 124.240 27.500 124.410 28.200 ;
        RECT 124.580 27.840 124.750 28.620 ;
        RECT 125.070 28.570 125.440 29.070 ;
        RECT 125.620 28.620 126.025 28.790 ;
        RECT 126.195 28.620 126.980 28.790 ;
        RECT 125.620 28.390 125.790 28.620 ;
        RECT 124.960 28.090 125.790 28.390 ;
        RECT 126.175 28.120 126.640 28.450 ;
        RECT 124.960 28.060 125.160 28.090 ;
        RECT 125.280 27.840 125.450 27.910 ;
        RECT 124.580 27.670 125.450 27.840 ;
        RECT 124.940 27.580 125.450 27.670 ;
        RECT 123.490 27.115 123.795 27.245 ;
        RECT 124.240 27.135 124.770 27.500 ;
        RECT 123.110 26.520 123.375 26.980 ;
        RECT 123.545 26.690 123.795 27.115 ;
        RECT 124.940 26.965 125.110 27.580 ;
        RECT 124.005 26.795 125.110 26.965 ;
        RECT 125.280 26.520 125.450 27.320 ;
        RECT 125.620 27.020 125.790 28.090 ;
        RECT 125.960 27.190 126.150 27.910 ;
        RECT 126.320 27.160 126.640 28.120 ;
        RECT 126.810 28.160 126.980 28.620 ;
        RECT 127.255 28.540 127.465 29.070 ;
        RECT 127.725 28.330 128.055 28.855 ;
        RECT 128.225 28.460 128.395 29.070 ;
        RECT 128.565 28.415 128.895 28.850 ;
        RECT 128.565 28.330 128.945 28.415 ;
        RECT 129.115 28.345 129.405 29.070 ;
        RECT 127.855 28.160 128.055 28.330 ;
        RECT 128.720 28.290 128.945 28.330 ;
        RECT 126.810 27.830 127.685 28.160 ;
        RECT 127.855 27.830 128.605 28.160 ;
        RECT 125.620 26.690 125.870 27.020 ;
        RECT 126.810 26.990 126.980 27.830 ;
        RECT 127.855 27.625 128.045 27.830 ;
        RECT 128.775 27.710 128.945 28.290 ;
        RECT 129.575 28.320 130.785 29.070 ;
        RECT 131.045 28.520 131.215 28.810 ;
        RECT 131.385 28.690 131.715 29.070 ;
        RECT 131.045 28.350 131.710 28.520 ;
        RECT 129.575 27.780 130.095 28.320 ;
        RECT 128.730 27.660 128.945 27.710 ;
        RECT 127.150 27.250 128.045 27.625 ;
        RECT 128.555 27.580 128.945 27.660 ;
        RECT 126.095 26.820 126.980 26.990 ;
        RECT 127.160 26.520 127.475 27.020 ;
        RECT 127.705 26.690 128.045 27.250 ;
        RECT 128.215 26.520 128.385 27.530 ;
        RECT 128.555 26.735 128.885 27.580 ;
        RECT 129.115 26.520 129.405 27.685 ;
        RECT 130.265 27.610 130.785 28.150 ;
        RECT 129.575 26.520 130.785 27.610 ;
        RECT 130.960 27.530 131.310 28.180 ;
        RECT 131.480 27.360 131.710 28.350 ;
        RECT 131.045 27.190 131.710 27.360 ;
        RECT 131.045 26.690 131.215 27.190 ;
        RECT 131.385 26.520 131.715 27.020 ;
        RECT 131.885 26.690 132.070 28.810 ;
        RECT 132.325 28.610 132.575 29.070 ;
        RECT 132.745 28.620 133.080 28.790 ;
        RECT 133.275 28.620 133.950 28.790 ;
        RECT 132.745 28.480 132.915 28.620 ;
        RECT 132.240 27.490 132.520 28.440 ;
        RECT 132.690 28.350 132.915 28.480 ;
        RECT 132.690 27.245 132.860 28.350 ;
        RECT 133.085 28.200 133.610 28.420 ;
        RECT 133.030 27.435 133.270 28.030 ;
        RECT 133.440 27.500 133.610 28.200 ;
        RECT 133.780 27.840 133.950 28.620 ;
        RECT 134.270 28.570 134.640 29.070 ;
        RECT 134.820 28.620 135.225 28.790 ;
        RECT 135.395 28.620 136.180 28.790 ;
        RECT 134.820 28.390 134.990 28.620 ;
        RECT 134.160 28.090 134.990 28.390 ;
        RECT 135.375 28.120 135.840 28.450 ;
        RECT 134.160 28.060 134.360 28.090 ;
        RECT 134.480 27.840 134.650 27.910 ;
        RECT 133.780 27.670 134.650 27.840 ;
        RECT 134.140 27.580 134.650 27.670 ;
        RECT 132.690 27.115 132.995 27.245 ;
        RECT 133.440 27.135 133.970 27.500 ;
        RECT 132.310 26.520 132.575 26.980 ;
        RECT 132.745 26.690 132.995 27.115 ;
        RECT 134.140 26.965 134.310 27.580 ;
        RECT 133.205 26.795 134.310 26.965 ;
        RECT 134.480 26.520 134.650 27.320 ;
        RECT 134.820 27.020 134.990 28.090 ;
        RECT 135.160 27.190 135.350 27.910 ;
        RECT 135.520 27.160 135.840 28.120 ;
        RECT 136.010 28.160 136.180 28.620 ;
        RECT 136.455 28.540 136.665 29.070 ;
        RECT 136.925 28.330 137.255 28.855 ;
        RECT 137.425 28.460 137.595 29.070 ;
        RECT 137.765 28.415 138.095 28.850 ;
        RECT 137.765 28.330 138.145 28.415 ;
        RECT 137.055 28.160 137.255 28.330 ;
        RECT 137.920 28.290 138.145 28.330 ;
        RECT 136.010 27.830 136.885 28.160 ;
        RECT 137.055 27.830 137.805 28.160 ;
        RECT 134.820 26.690 135.070 27.020 ;
        RECT 136.010 26.990 136.180 27.830 ;
        RECT 137.055 27.625 137.245 27.830 ;
        RECT 137.975 27.710 138.145 28.290 ;
        RECT 138.315 28.300 139.985 29.070 ;
        RECT 140.155 28.320 141.365 29.070 ;
        RECT 138.315 27.780 139.065 28.300 ;
        RECT 137.930 27.660 138.145 27.710 ;
        RECT 136.350 27.250 137.245 27.625 ;
        RECT 137.755 27.580 138.145 27.660 ;
        RECT 139.235 27.610 139.985 28.130 ;
        RECT 135.295 26.820 136.180 26.990 ;
        RECT 136.360 26.520 136.675 27.020 ;
        RECT 136.905 26.690 137.245 27.250 ;
        RECT 137.415 26.520 137.585 27.530 ;
        RECT 137.755 26.735 138.085 27.580 ;
        RECT 138.315 26.520 139.985 27.610 ;
        RECT 140.155 27.610 140.675 28.150 ;
        RECT 140.845 27.780 141.365 28.320 ;
        RECT 140.155 26.520 141.365 27.610 ;
        RECT 103.270 26.350 141.450 26.520 ;
        RECT 103.355 25.260 104.565 26.350 ;
        RECT 104.735 25.260 107.325 26.350 ;
        RECT 107.585 25.680 107.755 26.180 ;
        RECT 107.925 25.850 108.255 26.350 ;
        RECT 107.585 25.510 108.250 25.680 ;
        RECT 103.355 24.550 103.875 25.090 ;
        RECT 104.045 24.720 104.565 25.260 ;
        RECT 104.735 24.570 105.945 25.090 ;
        RECT 106.115 24.740 107.325 25.260 ;
        RECT 107.500 24.690 107.850 25.340 ;
        RECT 103.355 23.800 104.565 24.550 ;
        RECT 104.735 23.800 107.325 24.570 ;
        RECT 108.020 24.520 108.250 25.510 ;
        RECT 107.585 24.350 108.250 24.520 ;
        RECT 107.585 24.060 107.755 24.350 ;
        RECT 107.925 23.800 108.255 24.180 ;
        RECT 108.425 24.060 108.610 26.180 ;
        RECT 108.850 25.890 109.115 26.350 ;
        RECT 109.285 25.755 109.535 26.180 ;
        RECT 109.745 25.905 110.850 26.075 ;
        RECT 109.230 25.625 109.535 25.755 ;
        RECT 108.780 24.430 109.060 25.380 ;
        RECT 109.230 24.520 109.400 25.625 ;
        RECT 109.570 24.840 109.810 25.435 ;
        RECT 109.980 25.370 110.510 25.735 ;
        RECT 109.980 24.670 110.150 25.370 ;
        RECT 110.680 25.290 110.850 25.905 ;
        RECT 111.020 25.550 111.190 26.350 ;
        RECT 111.360 25.850 111.610 26.180 ;
        RECT 111.835 25.880 112.720 26.050 ;
        RECT 110.680 25.200 111.190 25.290 ;
        RECT 109.230 24.390 109.455 24.520 ;
        RECT 109.625 24.450 110.150 24.670 ;
        RECT 110.320 25.030 111.190 25.200 ;
        RECT 108.865 23.800 109.115 24.260 ;
        RECT 109.285 24.250 109.455 24.390 ;
        RECT 110.320 24.250 110.490 25.030 ;
        RECT 111.020 24.960 111.190 25.030 ;
        RECT 110.700 24.780 110.900 24.810 ;
        RECT 111.360 24.780 111.530 25.850 ;
        RECT 111.700 24.960 111.890 25.680 ;
        RECT 110.700 24.480 111.530 24.780 ;
        RECT 112.060 24.750 112.380 25.710 ;
        RECT 109.285 24.080 109.620 24.250 ;
        RECT 109.815 24.080 110.490 24.250 ;
        RECT 110.810 23.800 111.180 24.300 ;
        RECT 111.360 24.250 111.530 24.480 ;
        RECT 111.915 24.420 112.380 24.750 ;
        RECT 112.550 25.040 112.720 25.880 ;
        RECT 112.900 25.850 113.215 26.350 ;
        RECT 113.445 25.620 113.785 26.180 ;
        RECT 112.890 25.245 113.785 25.620 ;
        RECT 113.955 25.340 114.125 26.350 ;
        RECT 113.595 25.040 113.785 25.245 ;
        RECT 114.295 25.290 114.625 26.135 ;
        RECT 114.295 25.210 114.685 25.290 ;
        RECT 114.855 25.260 116.065 26.350 ;
        RECT 114.470 25.160 114.685 25.210 ;
        RECT 112.550 24.710 113.425 25.040 ;
        RECT 113.595 24.710 114.345 25.040 ;
        RECT 112.550 24.250 112.720 24.710 ;
        RECT 113.595 24.540 113.795 24.710 ;
        RECT 114.515 24.580 114.685 25.160 ;
        RECT 114.460 24.540 114.685 24.580 ;
        RECT 111.360 24.080 111.765 24.250 ;
        RECT 111.935 24.080 112.720 24.250 ;
        RECT 112.995 23.800 113.205 24.330 ;
        RECT 113.465 24.015 113.795 24.540 ;
        RECT 114.305 24.455 114.685 24.540 ;
        RECT 114.855 24.550 115.375 25.090 ;
        RECT 115.545 24.720 116.065 25.260 ;
        RECT 116.235 25.185 116.525 26.350 ;
        RECT 116.895 25.680 117.175 26.350 ;
        RECT 117.345 25.460 117.645 26.010 ;
        RECT 117.845 25.630 118.175 26.350 ;
        RECT 118.365 25.630 118.825 26.180 ;
        RECT 118.995 25.795 119.600 26.350 ;
        RECT 119.775 25.840 120.255 26.180 ;
        RECT 120.425 25.805 120.680 26.350 ;
        RECT 118.995 25.695 119.610 25.795 ;
        RECT 116.710 25.040 116.975 25.400 ;
        RECT 117.345 25.290 118.285 25.460 ;
        RECT 118.115 25.040 118.285 25.290 ;
        RECT 116.710 24.790 117.385 25.040 ;
        RECT 117.605 24.790 117.945 25.040 ;
        RECT 118.115 24.710 118.405 25.040 ;
        RECT 118.115 24.620 118.285 24.710 ;
        RECT 113.965 23.800 114.135 24.410 ;
        RECT 114.305 24.020 114.635 24.455 ;
        RECT 114.855 23.800 116.065 24.550 ;
        RECT 116.235 23.800 116.525 24.525 ;
        RECT 116.895 24.430 118.285 24.620 ;
        RECT 116.895 24.070 117.225 24.430 ;
        RECT 118.575 24.260 118.825 25.630 ;
        RECT 119.425 25.670 119.610 25.695 ;
        RECT 118.995 25.075 119.255 25.525 ;
        RECT 119.425 25.425 119.755 25.670 ;
        RECT 119.925 25.350 120.680 25.600 ;
        RECT 120.850 25.480 121.125 26.180 ;
        RECT 119.910 25.315 120.680 25.350 ;
        RECT 119.895 25.305 120.680 25.315 ;
        RECT 119.890 25.290 120.785 25.305 ;
        RECT 119.870 25.275 120.785 25.290 ;
        RECT 119.850 25.265 120.785 25.275 ;
        RECT 119.825 25.255 120.785 25.265 ;
        RECT 119.755 25.225 120.785 25.255 ;
        RECT 119.735 25.195 120.785 25.225 ;
        RECT 119.715 25.165 120.785 25.195 ;
        RECT 119.685 25.140 120.785 25.165 ;
        RECT 119.650 25.105 120.785 25.140 ;
        RECT 119.620 25.100 120.785 25.105 ;
        RECT 119.620 25.095 120.010 25.100 ;
        RECT 119.620 25.085 119.985 25.095 ;
        RECT 119.620 25.080 119.970 25.085 ;
        RECT 119.620 25.075 119.955 25.080 ;
        RECT 118.995 25.070 119.955 25.075 ;
        RECT 118.995 25.060 119.945 25.070 ;
        RECT 118.995 25.055 119.935 25.060 ;
        RECT 118.995 25.045 119.925 25.055 ;
        RECT 118.995 25.035 119.920 25.045 ;
        RECT 118.995 25.030 119.915 25.035 ;
        RECT 118.995 25.015 119.905 25.030 ;
        RECT 118.995 25.000 119.900 25.015 ;
        RECT 118.995 24.975 119.890 25.000 ;
        RECT 118.995 24.905 119.885 24.975 ;
        RECT 118.995 24.350 119.545 24.735 ;
        RECT 117.845 23.800 118.095 24.260 ;
        RECT 118.265 23.970 118.825 24.260 ;
        RECT 119.715 24.180 119.885 24.905 ;
        RECT 118.995 24.010 119.885 24.180 ;
        RECT 120.055 24.505 120.385 24.930 ;
        RECT 120.555 24.705 120.785 25.100 ;
        RECT 120.055 24.020 120.275 24.505 ;
        RECT 120.955 24.450 121.125 25.480 ;
        RECT 120.445 23.800 120.695 24.340 ;
        RECT 120.865 23.970 121.125 24.450 ;
        RECT 121.295 25.480 121.570 26.180 ;
        RECT 121.740 25.805 121.995 26.350 ;
        RECT 122.165 25.840 122.645 26.180 ;
        RECT 122.820 25.795 123.425 26.350 ;
        RECT 122.810 25.695 123.425 25.795 ;
        RECT 122.810 25.670 122.995 25.695 ;
        RECT 121.295 24.450 121.465 25.480 ;
        RECT 121.740 25.350 122.495 25.600 ;
        RECT 122.665 25.425 122.995 25.670 ;
        RECT 123.685 25.680 123.855 26.180 ;
        RECT 124.025 25.850 124.355 26.350 ;
        RECT 121.740 25.315 122.510 25.350 ;
        RECT 121.740 25.305 122.525 25.315 ;
        RECT 121.635 25.290 122.530 25.305 ;
        RECT 121.635 25.275 122.550 25.290 ;
        RECT 121.635 25.265 122.570 25.275 ;
        RECT 121.635 25.255 122.595 25.265 ;
        RECT 121.635 25.225 122.665 25.255 ;
        RECT 121.635 25.195 122.685 25.225 ;
        RECT 121.635 25.165 122.705 25.195 ;
        RECT 121.635 25.140 122.735 25.165 ;
        RECT 121.635 25.105 122.770 25.140 ;
        RECT 121.635 25.100 122.800 25.105 ;
        RECT 121.635 24.705 121.865 25.100 ;
        RECT 122.410 25.095 122.800 25.100 ;
        RECT 122.435 25.085 122.800 25.095 ;
        RECT 122.450 25.080 122.800 25.085 ;
        RECT 122.465 25.075 122.800 25.080 ;
        RECT 123.165 25.075 123.425 25.525 ;
        RECT 123.685 25.510 124.350 25.680 ;
        RECT 122.465 25.070 123.425 25.075 ;
        RECT 122.475 25.060 123.425 25.070 ;
        RECT 122.485 25.055 123.425 25.060 ;
        RECT 122.495 25.045 123.425 25.055 ;
        RECT 122.500 25.035 123.425 25.045 ;
        RECT 122.505 25.030 123.425 25.035 ;
        RECT 122.515 25.015 123.425 25.030 ;
        RECT 122.520 25.000 123.425 25.015 ;
        RECT 122.530 24.975 123.425 25.000 ;
        RECT 122.035 24.505 122.365 24.930 ;
        RECT 121.295 23.970 121.555 24.450 ;
        RECT 121.725 23.800 121.975 24.340 ;
        RECT 122.145 24.020 122.365 24.505 ;
        RECT 122.535 24.905 123.425 24.975 ;
        RECT 122.535 24.180 122.705 24.905 ;
        RECT 122.875 24.350 123.425 24.735 ;
        RECT 123.600 24.690 123.950 25.340 ;
        RECT 124.120 24.520 124.350 25.510 ;
        RECT 123.685 24.350 124.350 24.520 ;
        RECT 122.535 24.010 123.425 24.180 ;
        RECT 123.685 24.060 123.855 24.350 ;
        RECT 124.025 23.800 124.355 24.180 ;
        RECT 124.525 24.060 124.710 26.180 ;
        RECT 124.950 25.890 125.215 26.350 ;
        RECT 125.385 25.755 125.635 26.180 ;
        RECT 125.845 25.905 126.950 26.075 ;
        RECT 125.330 25.625 125.635 25.755 ;
        RECT 124.880 24.430 125.160 25.380 ;
        RECT 125.330 24.520 125.500 25.625 ;
        RECT 125.670 24.840 125.910 25.435 ;
        RECT 126.080 25.370 126.610 25.735 ;
        RECT 126.080 24.670 126.250 25.370 ;
        RECT 126.780 25.290 126.950 25.905 ;
        RECT 127.120 25.550 127.290 26.350 ;
        RECT 127.460 25.850 127.710 26.180 ;
        RECT 127.935 25.880 128.820 26.050 ;
        RECT 126.780 25.200 127.290 25.290 ;
        RECT 125.330 24.390 125.555 24.520 ;
        RECT 125.725 24.450 126.250 24.670 ;
        RECT 126.420 25.030 127.290 25.200 ;
        RECT 124.965 23.800 125.215 24.260 ;
        RECT 125.385 24.250 125.555 24.390 ;
        RECT 126.420 24.250 126.590 25.030 ;
        RECT 127.120 24.960 127.290 25.030 ;
        RECT 126.800 24.780 127.000 24.810 ;
        RECT 127.460 24.780 127.630 25.850 ;
        RECT 127.800 24.960 127.990 25.680 ;
        RECT 126.800 24.480 127.630 24.780 ;
        RECT 128.160 24.750 128.480 25.710 ;
        RECT 125.385 24.080 125.720 24.250 ;
        RECT 125.915 24.080 126.590 24.250 ;
        RECT 126.910 23.800 127.280 24.300 ;
        RECT 127.460 24.250 127.630 24.480 ;
        RECT 128.015 24.420 128.480 24.750 ;
        RECT 128.650 25.040 128.820 25.880 ;
        RECT 129.000 25.850 129.315 26.350 ;
        RECT 129.545 25.620 129.885 26.180 ;
        RECT 128.990 25.245 129.885 25.620 ;
        RECT 130.055 25.340 130.225 26.350 ;
        RECT 129.695 25.040 129.885 25.245 ;
        RECT 130.395 25.290 130.725 26.135 ;
        RECT 131.045 25.680 131.215 26.180 ;
        RECT 131.385 25.850 131.715 26.350 ;
        RECT 131.045 25.510 131.710 25.680 ;
        RECT 130.395 25.210 130.785 25.290 ;
        RECT 130.570 25.160 130.785 25.210 ;
        RECT 128.650 24.710 129.525 25.040 ;
        RECT 129.695 24.710 130.445 25.040 ;
        RECT 128.650 24.250 128.820 24.710 ;
        RECT 129.695 24.540 129.895 24.710 ;
        RECT 130.615 24.580 130.785 25.160 ;
        RECT 130.960 24.690 131.310 25.340 ;
        RECT 130.560 24.540 130.785 24.580 ;
        RECT 127.460 24.080 127.865 24.250 ;
        RECT 128.035 24.080 128.820 24.250 ;
        RECT 129.095 23.800 129.305 24.330 ;
        RECT 129.565 24.015 129.895 24.540 ;
        RECT 130.405 24.455 130.785 24.540 ;
        RECT 131.480 24.520 131.710 25.510 ;
        RECT 130.065 23.800 130.235 24.410 ;
        RECT 130.405 24.020 130.735 24.455 ;
        RECT 131.045 24.350 131.710 24.520 ;
        RECT 131.045 24.060 131.215 24.350 ;
        RECT 131.385 23.800 131.715 24.180 ;
        RECT 131.885 24.060 132.070 26.180 ;
        RECT 132.310 25.890 132.575 26.350 ;
        RECT 132.745 25.755 132.995 26.180 ;
        RECT 133.205 25.905 134.310 26.075 ;
        RECT 132.690 25.625 132.995 25.755 ;
        RECT 132.240 24.430 132.520 25.380 ;
        RECT 132.690 24.520 132.860 25.625 ;
        RECT 133.030 24.840 133.270 25.435 ;
        RECT 133.440 25.370 133.970 25.735 ;
        RECT 133.440 24.670 133.610 25.370 ;
        RECT 134.140 25.290 134.310 25.905 ;
        RECT 134.480 25.550 134.650 26.350 ;
        RECT 134.820 25.850 135.070 26.180 ;
        RECT 135.295 25.880 136.180 26.050 ;
        RECT 134.140 25.200 134.650 25.290 ;
        RECT 132.690 24.390 132.915 24.520 ;
        RECT 133.085 24.450 133.610 24.670 ;
        RECT 133.780 25.030 134.650 25.200 ;
        RECT 132.325 23.800 132.575 24.260 ;
        RECT 132.745 24.250 132.915 24.390 ;
        RECT 133.780 24.250 133.950 25.030 ;
        RECT 134.480 24.960 134.650 25.030 ;
        RECT 134.160 24.780 134.360 24.810 ;
        RECT 134.820 24.780 134.990 25.850 ;
        RECT 135.160 24.960 135.350 25.680 ;
        RECT 134.160 24.480 134.990 24.780 ;
        RECT 135.520 24.750 135.840 25.710 ;
        RECT 132.745 24.080 133.080 24.250 ;
        RECT 133.275 24.080 133.950 24.250 ;
        RECT 134.270 23.800 134.640 24.300 ;
        RECT 134.820 24.250 134.990 24.480 ;
        RECT 135.375 24.420 135.840 24.750 ;
        RECT 136.010 25.040 136.180 25.880 ;
        RECT 136.360 25.850 136.675 26.350 ;
        RECT 136.905 25.620 137.245 26.180 ;
        RECT 136.350 25.245 137.245 25.620 ;
        RECT 137.415 25.340 137.585 26.350 ;
        RECT 137.055 25.040 137.245 25.245 ;
        RECT 137.755 25.290 138.085 26.135 ;
        RECT 137.755 25.210 138.145 25.290 ;
        RECT 138.315 25.260 139.985 26.350 ;
        RECT 137.930 25.160 138.145 25.210 ;
        RECT 136.010 24.710 136.885 25.040 ;
        RECT 137.055 24.710 137.805 25.040 ;
        RECT 136.010 24.250 136.180 24.710 ;
        RECT 137.055 24.540 137.255 24.710 ;
        RECT 137.975 24.580 138.145 25.160 ;
        RECT 137.920 24.540 138.145 24.580 ;
        RECT 134.820 24.080 135.225 24.250 ;
        RECT 135.395 24.080 136.180 24.250 ;
        RECT 136.455 23.800 136.665 24.330 ;
        RECT 136.925 24.015 137.255 24.540 ;
        RECT 137.765 24.455 138.145 24.540 ;
        RECT 138.315 24.570 139.065 25.090 ;
        RECT 139.235 24.740 139.985 25.260 ;
        RECT 140.155 25.260 141.365 26.350 ;
        RECT 140.155 24.720 140.675 25.260 ;
        RECT 137.425 23.800 137.595 24.410 ;
        RECT 137.765 24.020 138.095 24.455 ;
        RECT 138.315 23.800 139.985 24.570 ;
        RECT 140.845 24.550 141.365 25.090 ;
        RECT 140.155 23.800 141.365 24.550 ;
        RECT 103.270 23.630 141.450 23.800 ;
        RECT 103.355 22.880 104.565 23.630 ;
        RECT 103.355 22.340 103.875 22.880 ;
        RECT 104.735 22.860 108.245 23.630 ;
        RECT 108.415 22.880 109.625 23.630 ;
        RECT 109.855 23.265 110.025 23.290 ;
        RECT 109.795 22.890 110.155 23.265 ;
        RECT 110.420 22.890 110.590 23.630 ;
        RECT 110.870 23.060 111.040 23.265 ;
        RECT 110.870 22.890 111.410 23.060 ;
        RECT 104.045 22.170 104.565 22.710 ;
        RECT 104.735 22.340 106.385 22.860 ;
        RECT 106.555 22.170 108.245 22.690 ;
        RECT 108.415 22.340 108.935 22.880 ;
        RECT 109.105 22.170 109.625 22.710 ;
        RECT 103.355 21.080 104.565 22.170 ;
        RECT 104.735 21.080 108.245 22.170 ;
        RECT 108.415 21.080 109.625 22.170 ;
        RECT 109.795 22.235 110.050 22.890 ;
        RECT 110.220 22.390 110.570 22.720 ;
        RECT 110.740 22.390 111.070 22.720 ;
        RECT 109.795 21.250 110.135 22.235 ;
        RECT 110.305 21.850 110.570 22.390 ;
        RECT 111.240 22.190 111.410 22.890 ;
        RECT 110.785 22.020 111.410 22.190 ;
        RECT 111.580 22.260 111.750 23.460 ;
        RECT 111.980 22.980 112.310 23.460 ;
        RECT 112.480 23.160 112.650 23.630 ;
        RECT 112.820 22.980 113.150 23.445 ;
        RECT 111.980 22.810 113.150 22.980 ;
        RECT 113.475 23.170 114.035 23.460 ;
        RECT 114.205 23.170 114.455 23.630 ;
        RECT 111.920 22.430 112.490 22.640 ;
        RECT 112.660 22.430 113.305 22.640 ;
        RECT 111.580 21.850 112.285 22.260 ;
        RECT 110.305 21.680 112.285 21.850 ;
        RECT 110.305 21.080 110.715 21.510 ;
        RECT 111.460 21.080 111.790 21.500 ;
        RECT 111.960 21.250 112.285 21.680 ;
        RECT 112.760 21.080 113.090 22.180 ;
        RECT 113.475 21.800 113.725 23.170 ;
        RECT 115.075 23.000 115.405 23.360 ;
        RECT 114.015 22.810 115.405 23.000 ;
        RECT 116.895 23.000 117.225 23.360 ;
        RECT 117.845 23.170 118.095 23.630 ;
        RECT 118.265 23.170 118.825 23.460 ;
        RECT 116.895 22.810 118.285 23.000 ;
        RECT 114.015 22.720 114.185 22.810 ;
        RECT 113.895 22.390 114.185 22.720 ;
        RECT 118.115 22.720 118.285 22.810 ;
        RECT 114.355 22.390 114.695 22.640 ;
        RECT 114.915 22.390 115.590 22.640 ;
        RECT 114.015 22.140 114.185 22.390 ;
        RECT 114.015 21.970 114.955 22.140 ;
        RECT 115.325 22.030 115.590 22.390 ;
        RECT 116.710 22.390 117.385 22.640 ;
        RECT 117.605 22.390 117.945 22.640 ;
        RECT 118.115 22.390 118.405 22.720 ;
        RECT 116.710 22.030 116.975 22.390 ;
        RECT 118.115 22.140 118.285 22.390 ;
        RECT 113.475 21.250 113.935 21.800 ;
        RECT 114.125 21.080 114.455 21.800 ;
        RECT 114.655 21.420 114.955 21.970 ;
        RECT 117.345 21.970 118.285 22.140 ;
        RECT 115.125 21.080 115.405 21.750 ;
        RECT 116.895 21.080 117.175 21.750 ;
        RECT 117.345 21.420 117.645 21.970 ;
        RECT 118.575 21.800 118.825 23.170 ;
        RECT 118.995 23.085 124.340 23.630 ;
        RECT 120.580 22.255 120.920 23.085 ;
        RECT 125.435 22.910 125.775 23.420 ;
        RECT 117.845 21.080 118.175 21.800 ;
        RECT 118.365 21.250 118.825 21.800 ;
        RECT 122.400 21.515 122.750 22.765 ;
        RECT 118.995 21.080 124.340 21.515 ;
        RECT 125.435 21.510 125.695 22.910 ;
        RECT 125.945 22.830 126.215 23.630 ;
        RECT 125.870 22.390 126.200 22.640 ;
        RECT 126.395 22.390 126.675 23.360 ;
        RECT 126.855 22.390 127.155 23.360 ;
        RECT 127.335 22.390 127.685 23.355 ;
        RECT 127.905 23.130 128.400 23.460 ;
        RECT 125.885 22.220 126.200 22.390 ;
        RECT 127.905 22.220 128.075 23.130 ;
        RECT 125.885 22.050 128.075 22.220 ;
        RECT 125.435 21.250 125.775 21.510 ;
        RECT 125.945 21.080 126.275 21.880 ;
        RECT 126.740 21.250 126.990 22.050 ;
        RECT 127.175 21.080 127.505 21.800 ;
        RECT 127.725 21.250 127.975 22.050 ;
        RECT 128.245 21.640 128.485 22.950 ;
        RECT 129.115 22.905 129.405 23.630 ;
        RECT 129.575 22.910 129.915 23.420 ;
        RECT 128.145 21.080 128.480 21.460 ;
        RECT 129.115 21.080 129.405 22.245 ;
        RECT 129.575 21.510 129.835 22.910 ;
        RECT 130.085 22.830 130.355 23.630 ;
        RECT 130.010 22.390 130.340 22.640 ;
        RECT 130.535 22.390 130.815 23.360 ;
        RECT 130.995 22.390 131.295 23.360 ;
        RECT 131.475 22.390 131.825 23.355 ;
        RECT 132.045 23.130 132.540 23.460 ;
        RECT 133.125 23.230 133.455 23.630 ;
        RECT 130.025 22.220 130.340 22.390 ;
        RECT 132.045 22.220 132.215 23.130 ;
        RECT 133.625 23.060 133.955 23.400 ;
        RECT 135.005 23.230 135.335 23.630 ;
        RECT 130.025 22.050 132.215 22.220 ;
        RECT 129.575 21.250 129.915 21.510 ;
        RECT 130.085 21.080 130.415 21.880 ;
        RECT 130.880 21.250 131.130 22.050 ;
        RECT 131.315 21.080 131.645 21.800 ;
        RECT 131.865 21.250 132.115 22.050 ;
        RECT 132.385 21.640 132.625 22.950 ;
        RECT 132.970 22.890 135.335 23.060 ;
        RECT 135.505 22.905 135.835 23.415 ;
        RECT 132.970 21.890 133.140 22.890 ;
        RECT 135.165 22.720 135.335 22.890 ;
        RECT 133.310 22.060 133.555 22.720 ;
        RECT 133.770 22.060 134.035 22.720 ;
        RECT 134.230 22.060 134.515 22.720 ;
        RECT 134.690 22.390 134.995 22.720 ;
        RECT 135.165 22.390 135.475 22.720 ;
        RECT 134.690 22.060 134.905 22.390 ;
        RECT 132.970 21.720 133.425 21.890 ;
        RECT 132.285 21.080 132.620 21.460 ;
        RECT 133.095 21.290 133.425 21.720 ;
        RECT 133.605 21.720 134.895 21.890 ;
        RECT 133.605 21.300 133.855 21.720 ;
        RECT 134.085 21.080 134.415 21.550 ;
        RECT 134.645 21.300 134.895 21.720 ;
        RECT 135.085 21.080 135.335 22.220 ;
        RECT 135.645 22.140 135.835 22.905 ;
        RECT 136.015 22.795 136.305 23.630 ;
        RECT 136.475 23.230 137.430 23.400 ;
        RECT 137.845 23.240 138.175 23.630 ;
        RECT 136.475 22.350 136.645 23.230 ;
        RECT 138.345 23.060 138.515 23.380 ;
        RECT 138.685 23.240 139.015 23.630 ;
        RECT 136.815 22.890 139.065 23.060 ;
        RECT 136.815 22.390 137.045 22.890 ;
        RECT 137.215 22.470 137.590 22.640 ;
        RECT 135.505 21.290 135.835 22.140 ;
        RECT 136.015 22.180 136.645 22.350 ;
        RECT 137.420 22.270 137.590 22.470 ;
        RECT 137.760 22.440 138.310 22.640 ;
        RECT 138.480 22.270 138.725 22.720 ;
        RECT 136.015 21.250 136.335 22.180 ;
        RECT 137.420 22.100 138.725 22.270 ;
        RECT 138.895 21.930 139.065 22.890 ;
        RECT 140.155 22.880 141.365 23.630 ;
        RECT 136.515 21.760 137.755 21.930 ;
        RECT 136.515 21.250 136.915 21.760 ;
        RECT 137.085 21.080 137.255 21.590 ;
        RECT 137.425 21.250 137.755 21.760 ;
        RECT 137.925 21.080 138.095 21.930 ;
        RECT 138.685 21.250 139.065 21.930 ;
        RECT 140.155 22.170 140.675 22.710 ;
        RECT 140.845 22.340 141.365 22.880 ;
        RECT 140.155 21.080 141.365 22.170 ;
        RECT 103.270 20.910 141.450 21.080 ;
        RECT 103.355 19.820 104.565 20.910 ;
        RECT 103.355 19.110 103.875 19.650 ;
        RECT 104.045 19.280 104.565 19.820 ;
        RECT 104.735 19.835 105.005 20.740 ;
        RECT 105.175 20.150 105.505 20.910 ;
        RECT 105.685 19.980 105.865 20.740 ;
        RECT 103.355 18.360 104.565 19.110 ;
        RECT 104.735 19.035 104.915 19.835 ;
        RECT 105.190 19.810 105.865 19.980 ;
        RECT 106.575 19.835 106.845 20.740 ;
        RECT 107.015 20.150 107.345 20.910 ;
        RECT 107.525 19.980 107.705 20.740 ;
        RECT 105.190 19.665 105.360 19.810 ;
        RECT 105.085 19.335 105.360 19.665 ;
        RECT 105.190 19.080 105.360 19.335 ;
        RECT 105.585 19.260 105.925 19.630 ;
        RECT 104.735 18.530 104.995 19.035 ;
        RECT 105.190 18.910 105.855 19.080 ;
        RECT 105.175 18.360 105.505 18.740 ;
        RECT 105.685 18.530 105.855 18.910 ;
        RECT 106.575 19.035 106.755 19.835 ;
        RECT 107.030 19.810 107.705 19.980 ;
        RECT 107.955 19.820 110.545 20.910 ;
        RECT 107.030 19.665 107.200 19.810 ;
        RECT 106.925 19.335 107.200 19.665 ;
        RECT 107.030 19.080 107.200 19.335 ;
        RECT 107.425 19.260 107.765 19.630 ;
        RECT 107.955 19.130 109.165 19.650 ;
        RECT 109.335 19.300 110.545 19.820 ;
        RECT 111.175 19.835 111.445 20.740 ;
        RECT 111.615 20.150 111.945 20.910 ;
        RECT 112.125 19.980 112.305 20.740 ;
        RECT 106.575 18.530 106.835 19.035 ;
        RECT 107.030 18.910 107.695 19.080 ;
        RECT 107.015 18.360 107.345 18.740 ;
        RECT 107.525 18.530 107.695 18.910 ;
        RECT 107.955 18.360 110.545 19.130 ;
        RECT 111.175 19.035 111.355 19.835 ;
        RECT 111.630 19.810 112.305 19.980 ;
        RECT 112.555 19.820 116.065 20.910 ;
        RECT 111.630 19.665 111.800 19.810 ;
        RECT 111.525 19.335 111.800 19.665 ;
        RECT 111.630 19.080 111.800 19.335 ;
        RECT 112.025 19.260 112.365 19.630 ;
        RECT 112.555 19.130 114.205 19.650 ;
        RECT 114.375 19.300 116.065 19.820 ;
        RECT 116.235 19.745 116.525 20.910 ;
        RECT 116.695 19.835 116.965 20.740 ;
        RECT 117.135 20.150 117.465 20.910 ;
        RECT 117.645 19.980 117.825 20.740 ;
        RECT 111.175 18.530 111.435 19.035 ;
        RECT 111.630 18.910 112.295 19.080 ;
        RECT 111.615 18.360 111.945 18.740 ;
        RECT 112.125 18.530 112.295 18.910 ;
        RECT 112.555 18.360 116.065 19.130 ;
        RECT 116.235 18.360 116.525 19.085 ;
        RECT 116.695 19.035 116.875 19.835 ;
        RECT 117.150 19.810 117.825 19.980 ;
        RECT 118.075 19.820 119.745 20.910 ;
        RECT 117.150 19.665 117.320 19.810 ;
        RECT 117.045 19.335 117.320 19.665 ;
        RECT 117.150 19.080 117.320 19.335 ;
        RECT 117.545 19.260 117.885 19.630 ;
        RECT 118.075 19.130 118.825 19.650 ;
        RECT 118.995 19.300 119.745 19.820 ;
        RECT 120.375 19.835 120.645 20.740 ;
        RECT 120.815 20.150 121.145 20.910 ;
        RECT 121.325 19.980 121.505 20.740 ;
        RECT 116.695 18.530 116.955 19.035 ;
        RECT 117.150 18.910 117.815 19.080 ;
        RECT 117.135 18.360 117.465 18.740 ;
        RECT 117.645 18.530 117.815 18.910 ;
        RECT 118.075 18.360 119.745 19.130 ;
        RECT 120.375 19.035 120.555 19.835 ;
        RECT 120.830 19.810 121.505 19.980 ;
        RECT 121.755 19.820 124.345 20.910 ;
        RECT 120.830 19.665 121.000 19.810 ;
        RECT 120.725 19.335 121.000 19.665 ;
        RECT 120.830 19.080 121.000 19.335 ;
        RECT 121.225 19.260 121.565 19.630 ;
        RECT 121.755 19.130 122.965 19.650 ;
        RECT 123.135 19.300 124.345 19.820 ;
        RECT 124.975 19.835 125.245 20.740 ;
        RECT 125.415 20.150 125.745 20.910 ;
        RECT 125.925 19.980 126.105 20.740 ;
        RECT 120.375 18.530 120.635 19.035 ;
        RECT 120.830 18.910 121.495 19.080 ;
        RECT 120.815 18.360 121.145 18.740 ;
        RECT 121.325 18.530 121.495 18.910 ;
        RECT 121.755 18.360 124.345 19.130 ;
        RECT 124.975 19.035 125.155 19.835 ;
        RECT 125.430 19.810 126.105 19.980 ;
        RECT 126.355 19.820 128.945 20.910 ;
        RECT 125.430 19.665 125.600 19.810 ;
        RECT 125.325 19.335 125.600 19.665 ;
        RECT 125.430 19.080 125.600 19.335 ;
        RECT 125.825 19.260 126.165 19.630 ;
        RECT 126.355 19.130 127.565 19.650 ;
        RECT 127.735 19.300 128.945 19.820 ;
        RECT 129.115 19.745 129.405 20.910 ;
        RECT 129.575 19.835 129.845 20.740 ;
        RECT 130.015 20.150 130.345 20.910 ;
        RECT 130.525 19.980 130.705 20.740 ;
        RECT 124.975 18.530 125.235 19.035 ;
        RECT 125.430 18.910 126.095 19.080 ;
        RECT 125.415 18.360 125.745 18.740 ;
        RECT 125.925 18.530 126.095 18.910 ;
        RECT 126.355 18.360 128.945 19.130 ;
        RECT 129.115 18.360 129.405 19.085 ;
        RECT 129.575 19.035 129.755 19.835 ;
        RECT 130.030 19.810 130.705 19.980 ;
        RECT 130.955 19.820 133.545 20.910 ;
        RECT 130.030 19.665 130.200 19.810 ;
        RECT 129.925 19.335 130.200 19.665 ;
        RECT 130.030 19.080 130.200 19.335 ;
        RECT 130.425 19.260 130.765 19.630 ;
        RECT 130.955 19.130 132.165 19.650 ;
        RECT 132.335 19.300 133.545 19.820 ;
        RECT 134.175 19.835 134.445 20.740 ;
        RECT 134.615 20.150 134.945 20.910 ;
        RECT 135.125 19.980 135.305 20.740 ;
        RECT 129.575 18.530 129.835 19.035 ;
        RECT 130.030 18.910 130.695 19.080 ;
        RECT 130.015 18.360 130.345 18.740 ;
        RECT 130.525 18.530 130.695 18.910 ;
        RECT 130.955 18.360 133.545 19.130 ;
        RECT 134.175 19.035 134.355 19.835 ;
        RECT 134.630 19.810 135.305 19.980 ;
        RECT 135.555 19.820 137.225 20.910 ;
        RECT 134.630 19.665 134.800 19.810 ;
        RECT 134.525 19.335 134.800 19.665 ;
        RECT 134.630 19.080 134.800 19.335 ;
        RECT 135.025 19.260 135.365 19.630 ;
        RECT 135.555 19.130 136.305 19.650 ;
        RECT 136.475 19.300 137.225 19.820 ;
        RECT 137.475 19.980 137.655 20.740 ;
        RECT 137.835 20.150 138.165 20.910 ;
        RECT 137.475 19.810 138.150 19.980 ;
        RECT 138.335 19.835 138.605 20.740 ;
        RECT 137.980 19.665 138.150 19.810 ;
        RECT 137.415 19.260 137.755 19.630 ;
        RECT 137.980 19.335 138.255 19.665 ;
        RECT 134.175 18.530 134.435 19.035 ;
        RECT 134.630 18.910 135.295 19.080 ;
        RECT 134.615 18.360 134.945 18.740 ;
        RECT 135.125 18.530 135.295 18.910 ;
        RECT 135.555 18.360 137.225 19.130 ;
        RECT 137.980 19.080 138.150 19.335 ;
        RECT 137.485 18.910 138.150 19.080 ;
        RECT 138.425 19.035 138.605 19.835 ;
        RECT 137.485 18.530 137.655 18.910 ;
        RECT 137.835 18.360 138.165 18.740 ;
        RECT 138.345 18.530 138.605 19.035 ;
        RECT 138.775 19.835 139.045 20.740 ;
        RECT 139.215 20.150 139.545 20.910 ;
        RECT 139.725 19.980 139.905 20.740 ;
        RECT 138.775 19.035 138.955 19.835 ;
        RECT 139.230 19.810 139.905 19.980 ;
        RECT 140.155 19.820 141.365 20.910 ;
        RECT 139.230 19.665 139.400 19.810 ;
        RECT 139.125 19.335 139.400 19.665 ;
        RECT 139.230 19.080 139.400 19.335 ;
        RECT 139.625 19.260 139.965 19.630 ;
        RECT 140.155 19.280 140.675 19.820 ;
        RECT 140.845 19.110 141.365 19.650 ;
        RECT 138.775 18.530 139.035 19.035 ;
        RECT 139.230 18.910 139.895 19.080 ;
        RECT 139.215 18.360 139.545 18.740 ;
        RECT 139.725 18.530 139.895 18.910 ;
        RECT 140.155 18.360 141.365 19.110 ;
        RECT 103.270 18.190 141.450 18.360 ;
      LAYER met1 ;
        RECT 132.580 223.140 133.305 223.805 ;
        RECT 135.355 223.245 136.050 223.880 ;
        RECT 138.145 223.275 138.775 223.845 ;
        RECT 127.070 211.630 128.070 211.660 ;
        RECT 54.580 210.630 128.070 211.630 ;
        RECT 127.070 210.600 128.070 210.630 ;
        RECT 51.940 208.440 130.650 209.320 ;
        RECT 89.605 166.665 90.340 175.080 ;
        RECT 132.610 174.350 133.275 223.140 ;
        RECT 90.925 171.730 91.535 172.565 ;
        RECT 135.385 171.885 136.020 223.245 ;
        RECT 90.920 171.315 91.535 171.730 ;
        RECT 90.920 166.665 91.525 171.315 ;
        RECT 92.250 169.320 92.915 170.455 ;
        RECT 138.175 170.375 138.745 223.275 ;
        RECT 138.145 169.805 138.775 170.375 ;
        RECT 89.590 165.665 90.590 166.665 ;
        RECT 90.760 166.640 91.760 166.665 ;
        RECT 92.225 166.645 92.915 169.320 ;
        RECT 90.760 165.665 91.770 166.640 ;
        RECT 91.960 166.020 92.960 166.645 ;
        RECT 91.920 165.690 92.960 166.020 ;
        RECT 89.830 165.515 90.590 165.665 ;
        RECT 89.985 165.200 90.375 165.515 ;
        RECT 91.440 164.400 91.770 165.665 ;
        RECT 91.960 165.645 92.960 165.690 ;
        RECT 92.875 165.280 101.995 165.350 ;
        RECT 92.875 164.880 102.115 165.280 ;
        RECT 92.875 164.870 101.155 164.880 ;
        RECT 96.655 164.460 97.005 164.730 ;
        RECT 98.035 164.670 98.325 164.700 ;
        RECT 101.205 164.670 101.465 164.725 ;
        RECT 98.035 164.580 102.165 164.670 ;
        RECT 97.995 164.460 102.165 164.580 ;
        RECT 93.255 164.400 93.605 164.410 ;
        RECT 91.440 164.070 96.520 164.400 ;
        RECT 95.345 163.820 95.565 163.880 ;
        RECT 95.335 163.760 95.625 163.820 ;
        RECT 91.920 163.730 95.175 163.750 ;
        RECT 91.920 163.450 95.195 163.730 ;
        RECT 91.920 163.420 95.175 163.450 ;
        RECT 95.335 163.420 95.775 163.760 ;
        RECT 96.190 163.740 96.520 164.070 ;
        RECT 96.715 164.250 96.985 164.460 ;
        RECT 96.715 163.890 97.125 164.250 ;
        RECT 97.995 163.910 98.515 164.460 ;
        RECT 101.205 164.405 101.465 164.460 ;
        RECT 96.145 163.440 96.575 163.740 ;
        RECT 96.725 163.440 97.125 163.890 ;
        RECT 98.035 163.860 98.485 163.910 ;
        RECT 97.505 163.440 97.955 163.740 ;
        RECT 98.115 163.440 98.485 163.860 ;
        RECT 95.335 163.400 95.625 163.420 ;
        RECT 95.345 163.370 95.565 163.400 ;
        RECT 97.540 163.180 97.870 163.440 ;
        RECT 90.910 162.850 97.870 163.180 ;
        RECT 87.900 160.885 89.460 162.745 ;
        RECT 92.875 162.150 103.455 162.630 ;
        RECT 95.250 161.980 95.540 161.995 ;
        RECT 95.245 161.970 95.540 161.980 ;
        RECT 96.075 161.970 96.395 162.010 ;
        RECT 92.925 161.780 93.225 161.850 ;
        RECT 95.245 161.790 96.395 161.970 ;
        RECT 96.715 161.840 97.135 161.860 ;
        RECT 95.245 161.780 95.540 161.790 ;
        RECT 92.815 161.750 93.225 161.780 ;
        RECT 95.250 161.765 95.540 161.780 ;
        RECT 96.075 161.750 96.395 161.790 ;
        RECT 92.625 160.660 93.225 161.750 ;
        RECT 96.705 161.610 97.135 161.840 ;
        RECT 98.015 161.840 98.305 161.980 ;
        RECT 101.215 161.880 101.515 161.960 ;
        RECT 93.895 161.580 97.135 161.610 ;
        RECT 93.895 161.470 97.125 161.580 ;
        RECT 93.895 161.340 94.205 161.470 ;
        RECT 93.815 161.050 94.205 161.340 ;
        RECT 94.415 161.320 95.115 161.330 ;
        RECT 94.415 161.295 95.125 161.320 ;
        RECT 95.280 161.295 95.600 161.300 ;
        RECT 94.400 161.045 95.600 161.295 ;
        RECT 94.415 161.040 95.125 161.045 ;
        RECT 95.280 161.040 95.600 161.045 ;
        RECT 97.465 160.990 97.825 161.690 ;
        RECT 98.015 161.580 98.855 161.840 ;
        RECT 98.015 161.560 98.305 161.580 ;
        RECT 100.245 161.550 100.565 161.570 ;
        RECT 97.975 161.345 98.295 161.370 ;
        RECT 100.225 161.345 100.605 161.550 ;
        RECT 97.975 161.135 100.605 161.345 ;
        RECT 97.975 161.110 98.295 161.135 ;
        RECT 97.485 160.950 97.805 160.990 ;
        RECT 95.775 160.740 96.445 160.770 ;
        RECT 98.655 160.760 99.095 160.860 ;
        RECT 100.225 160.780 100.605 161.135 ;
        RECT 101.205 161.000 101.645 161.880 ;
        RECT 102.095 161.320 102.485 161.330 ;
        RECT 102.085 161.050 102.485 161.320 ;
        RECT 102.675 161.305 103.405 161.340 ;
        RECT 102.670 161.055 103.405 161.305 ;
        RECT 101.215 160.960 101.515 161.000 ;
        RECT 102.105 160.780 102.425 161.050 ;
        RECT 102.675 160.960 103.405 161.055 ;
        RECT 98.545 160.740 99.205 160.760 ;
        RECT 92.925 160.590 93.225 160.660 ;
        RECT 93.775 160.470 98.305 160.740 ;
        RECT 93.775 160.420 94.275 160.470 ;
        RECT 95.785 160.430 96.455 160.470 ;
        RECT 97.945 160.420 98.305 160.470 ;
        RECT 98.525 160.460 99.215 160.740 ;
        RECT 100.205 160.520 102.455 160.780 ;
        RECT 93.005 160.270 93.385 160.380 ;
        RECT 98.725 160.315 99.035 160.460 ;
        RECT 97.495 160.270 97.815 160.315 ;
        RECT 98.725 160.270 99.045 160.315 ;
        RECT 103.090 160.270 103.340 160.960 ;
        RECT 93.005 160.175 103.340 160.270 ;
        RECT 93.005 160.110 103.300 160.175 ;
        RECT 93.095 160.100 103.300 160.110 ;
        RECT 97.495 160.055 97.815 160.100 ;
        RECT 98.725 160.055 99.045 160.100 ;
        RECT 92.875 159.430 103.455 159.910 ;
        RECT 94.765 158.470 95.135 159.430 ;
        RECT 95.705 159.210 96.045 159.270 ;
        RECT 95.685 158.510 96.065 159.210 ;
        RECT 97.075 159.200 97.395 159.260 ;
        RECT 97.055 158.510 97.415 159.200 ;
        RECT 98.915 159.100 99.255 159.170 ;
        RECT 99.885 159.105 100.205 159.130 ;
        RECT 101.225 159.105 101.545 159.130 ;
        RECT 95.705 158.450 96.045 158.510 ;
        RECT 97.075 158.450 97.395 158.510 ;
        RECT 98.905 158.490 99.295 159.100 ;
        RECT 99.885 158.895 101.545 159.105 ;
        RECT 99.885 158.870 100.205 158.895 ;
        RECT 101.225 158.870 101.545 158.895 ;
        RECT 98.915 158.440 99.255 158.490 ;
        RECT 92.630 158.135 92.950 158.190 ;
        RECT 95.225 158.135 95.665 158.300 ;
        RECT 92.630 158.020 95.665 158.135 ;
        RECT 96.085 158.230 96.405 158.270 ;
        RECT 96.635 158.230 97.015 158.290 ;
        RECT 98.455 158.270 98.875 158.300 ;
        RECT 96.085 158.055 97.015 158.230 ;
        RECT 92.630 157.985 95.590 158.020 ;
        RECT 96.085 158.010 96.405 158.055 ;
        RECT 96.635 158.010 97.015 158.055 ;
        RECT 98.435 158.000 98.875 158.270 ;
        RECT 92.630 157.930 92.950 157.985 ;
        RECT 98.435 157.970 98.865 158.000 ;
        RECT 94.755 157.190 95.125 157.830 ;
        RECT 99.015 157.780 99.255 158.440 ;
        RECT 99.795 158.000 100.205 158.300 ;
        RECT 100.355 158.230 100.655 158.300 ;
        RECT 98.925 157.330 99.255 157.780 ;
        RECT 100.355 157.470 100.765 158.230 ;
        RECT 100.355 157.410 100.655 157.470 ;
        RECT 92.875 156.710 102.995 157.190 ;
        RECT 106.140 153.615 107.140 153.865 ;
        RECT 108.080 153.615 114.570 154.320 ;
        RECT 103.490 153.580 114.570 153.615 ;
        RECT 62.965 152.820 63.405 153.200 ;
        RECT 61.575 151.865 62.575 151.980 ;
        RECT 62.995 151.970 63.375 152.820 ;
        RECT 67.150 152.410 72.295 152.945 ;
        RECT 103.395 152.690 114.570 153.580 ;
        RECT 103.490 152.665 114.570 152.690 ;
        RECT 67.150 152.170 67.685 152.410 ;
        RECT 60.320 151.115 62.575 151.865 ;
        RECT 60.320 126.765 61.070 151.115 ;
        RECT 61.575 150.980 62.575 151.115 ;
        RECT 62.715 151.610 63.715 151.970 ;
        RECT 62.715 151.240 66.175 151.610 ;
        RECT 62.715 150.970 63.715 151.240 ;
        RECT 61.885 150.730 62.525 150.750 ;
        RECT 61.575 149.730 62.575 150.730 ;
        RECT 62.715 150.720 63.065 150.740 ;
        RECT 62.715 149.740 63.715 150.720 ;
        RECT 64.515 150.250 64.745 151.065 ;
        RECT 61.885 149.710 62.525 149.730 ;
        RECT 62.715 149.470 63.175 149.740 ;
        RECT 62.485 149.220 63.175 149.470 ;
        RECT 62.485 149.070 62.785 149.220 ;
        RECT 61.415 148.790 62.785 149.070 ;
        RECT 61.415 140.370 61.775 148.790 ;
        RECT 62.475 148.760 62.785 148.790 ;
        RECT 62.195 148.440 62.425 148.600 ;
        RECT 61.935 140.920 62.425 148.440 ;
        RECT 62.195 140.600 62.425 140.920 ;
        RECT 62.835 148.520 63.065 148.600 ;
        RECT 62.835 147.830 63.335 148.520 ;
        RECT 64.245 147.830 64.745 150.250 ;
        RECT 62.835 146.530 64.745 147.830 ;
        RECT 62.835 143.900 63.335 146.530 ;
        RECT 64.245 143.900 64.745 146.530 ;
        RECT 62.835 142.600 64.745 143.900 ;
        RECT 62.835 140.610 63.335 142.600 ;
        RECT 62.835 140.600 63.065 140.610 ;
        RECT 62.415 140.370 62.815 140.440 ;
        RECT 61.415 139.770 62.815 140.370 ;
        RECT 61.415 131.350 61.775 139.770 ;
        RECT 62.415 139.700 62.815 139.770 ;
        RECT 62.475 139.670 62.785 139.700 ;
        RECT 62.195 139.230 62.425 139.510 ;
        RECT 61.915 131.710 62.425 139.230 ;
        RECT 62.195 131.510 62.425 131.710 ;
        RECT 62.835 139.460 63.065 139.510 ;
        RECT 62.835 138.640 63.345 139.460 ;
        RECT 63.545 138.640 63.955 142.600 ;
        RECT 64.245 142.340 64.745 142.600 ;
        RECT 64.515 141.065 64.745 142.340 ;
        RECT 65.155 150.580 65.385 151.065 ;
        RECT 65.155 141.610 65.635 150.580 ;
        RECT 65.155 141.065 65.385 141.610 ;
        RECT 64.795 140.840 65.105 140.860 ;
        RECT 64.775 140.690 65.105 140.840 ;
        RECT 65.905 140.690 66.175 151.240 ;
        RECT 66.865 151.170 67.865 152.170 ;
        RECT 68.005 151.800 69.005 152.160 ;
        RECT 71.760 152.040 72.295 152.410 ;
        RECT 73.095 152.040 74.915 152.180 ;
        RECT 68.005 151.430 71.465 151.800 ;
        RECT 68.005 151.160 69.005 151.430 ;
        RECT 67.125 150.920 67.755 150.960 ;
        RECT 66.865 149.920 67.865 150.920 ;
        RECT 68.005 150.910 68.355 150.930 ;
        RECT 68.005 149.930 69.005 150.910 ;
        RECT 69.805 150.440 70.035 151.255 ;
        RECT 67.125 149.890 67.755 149.920 ;
        RECT 68.005 149.660 68.465 149.930 ;
        RECT 67.775 149.410 68.465 149.660 ;
        RECT 67.775 149.260 68.075 149.410 ;
        RECT 64.775 140.240 66.175 140.690 ;
        RECT 64.775 140.110 65.105 140.240 ;
        RECT 64.795 140.090 65.105 140.110 ;
        RECT 64.515 138.990 64.745 139.885 ;
        RECT 64.275 138.640 64.745 138.990 ;
        RECT 62.835 137.340 64.745 138.640 ;
        RECT 62.835 134.300 63.345 137.340 ;
        RECT 64.275 134.300 64.745 137.340 ;
        RECT 62.835 133.000 64.745 134.300 ;
        RECT 62.835 131.850 63.345 133.000 ;
        RECT 64.275 131.850 64.745 133.000 ;
        RECT 62.835 131.510 64.745 131.850 ;
        RECT 61.415 131.050 62.805 131.350 ;
        RECT 62.985 131.270 64.745 131.510 ;
        RECT 61.415 131.040 61.775 131.050 ;
        RECT 63.265 130.550 63.735 131.270 ;
        RECT 64.275 131.080 64.745 131.270 ;
        RECT 61.525 130.360 63.735 130.550 ;
        RECT 61.475 130.020 63.735 130.360 ;
        RECT 61.475 129.290 62.525 130.020 ;
        RECT 64.515 129.885 64.745 131.080 ;
        RECT 65.155 139.200 65.385 139.885 ;
        RECT 65.155 130.230 65.715 139.200 ;
        RECT 65.155 129.885 65.385 130.230 ;
        RECT 34.370 126.300 35.450 126.340 ;
        RECT 56.010 126.300 57.010 126.305 ;
        RECT 61.475 126.300 62.475 129.290 ;
        RECT 62.745 128.820 63.745 129.820 ;
        RECT 64.795 129.670 65.105 129.680 ;
        RECT 65.905 129.670 66.175 140.240 ;
        RECT 66.705 148.980 68.075 149.260 ;
        RECT 66.705 140.560 67.065 148.980 ;
        RECT 67.765 148.950 68.075 148.980 ;
        RECT 67.485 148.630 67.715 148.790 ;
        RECT 67.225 141.110 67.715 148.630 ;
        RECT 67.485 140.790 67.715 141.110 ;
        RECT 68.125 148.710 68.355 148.790 ;
        RECT 68.125 148.020 68.625 148.710 ;
        RECT 69.535 148.020 70.035 150.440 ;
        RECT 68.125 146.720 70.035 148.020 ;
        RECT 68.125 144.090 68.625 146.720 ;
        RECT 69.535 144.090 70.035 146.720 ;
        RECT 68.125 142.790 70.035 144.090 ;
        RECT 68.125 140.800 68.625 142.790 ;
        RECT 68.125 140.790 68.355 140.800 ;
        RECT 67.705 140.560 68.105 140.630 ;
        RECT 66.705 139.960 68.105 140.560 ;
        RECT 66.705 131.540 67.065 139.960 ;
        RECT 67.705 139.890 68.105 139.960 ;
        RECT 67.765 139.860 68.075 139.890 ;
        RECT 67.485 139.420 67.715 139.700 ;
        RECT 67.205 131.900 67.715 139.420 ;
        RECT 67.485 131.700 67.715 131.900 ;
        RECT 68.125 139.650 68.355 139.700 ;
        RECT 68.125 138.830 68.635 139.650 ;
        RECT 68.835 138.830 69.245 142.790 ;
        RECT 69.535 142.530 70.035 142.790 ;
        RECT 69.805 141.255 70.035 142.530 ;
        RECT 70.445 150.770 70.675 151.255 ;
        RECT 70.445 141.800 70.925 150.770 ;
        RECT 70.445 141.255 70.675 141.800 ;
        RECT 70.085 141.030 70.395 141.050 ;
        RECT 70.065 140.880 70.395 141.030 ;
        RECT 71.195 140.880 71.465 151.430 ;
        RECT 70.065 140.430 71.465 140.880 ;
        RECT 70.065 140.300 70.395 140.430 ;
        RECT 70.085 140.280 70.395 140.300 ;
        RECT 69.805 139.180 70.035 140.075 ;
        RECT 69.565 138.830 70.035 139.180 ;
        RECT 68.125 137.530 70.035 138.830 ;
        RECT 68.125 134.490 68.635 137.530 ;
        RECT 69.565 134.490 70.035 137.530 ;
        RECT 68.125 133.190 70.035 134.490 ;
        RECT 68.125 132.040 68.635 133.190 ;
        RECT 69.565 132.040 70.035 133.190 ;
        RECT 68.125 131.700 70.035 132.040 ;
        RECT 66.705 131.240 68.095 131.540 ;
        RECT 68.275 131.460 70.035 131.700 ;
        RECT 66.705 131.230 67.065 131.240 ;
        RECT 68.555 130.740 69.025 131.460 ;
        RECT 69.565 131.270 70.035 131.460 ;
        RECT 64.765 129.400 66.175 129.670 ;
        RECT 66.815 130.210 69.025 130.740 ;
        RECT 66.815 126.300 67.815 130.210 ;
        RECT 69.805 130.075 70.035 131.270 ;
        RECT 70.445 139.390 70.675 140.075 ;
        RECT 70.445 130.420 71.005 139.390 ;
        RECT 70.445 130.075 70.675 130.420 ;
        RECT 68.035 129.010 69.035 130.010 ;
        RECT 70.085 129.860 70.395 129.870 ;
        RECT 71.195 129.860 71.465 140.430 ;
        RECT 71.760 151.505 74.915 152.040 ;
        RECT 75.405 151.930 93.435 152.290 ;
        RECT 71.760 146.630 72.295 151.505 ;
        RECT 73.095 151.180 74.915 151.505 ;
        RECT 72.625 149.960 74.185 150.960 ;
        RECT 74.385 150.440 74.915 151.180 ;
        RECT 75.415 150.900 75.715 151.930 ;
        RECT 76.075 151.510 83.595 151.790 ;
        RECT 75.875 151.280 83.875 151.510 ;
        RECT 84.135 151.290 84.735 151.930 ;
        RECT 85.285 151.510 92.805 151.770 ;
        RECT 84.065 151.230 84.805 151.290 ;
        RECT 84.965 151.280 92.965 151.510 ;
        RECT 93.155 151.230 93.435 151.930 ;
        RECT 84.035 150.920 84.805 151.230 ;
        RECT 93.125 151.220 93.435 151.230 ;
        RECT 93.125 150.990 93.835 151.220 ;
        RECT 94.095 151.130 95.095 152.130 ;
        RECT 95.345 151.810 96.345 152.130 ;
        RECT 96.775 151.810 106.660 152.040 ;
        RECT 95.345 151.200 106.660 151.810 ;
        RECT 108.080 151.310 114.570 152.665 ;
        RECT 95.345 151.130 96.345 151.200 ;
        RECT 96.775 151.040 106.660 151.200 ;
        RECT 93.125 150.920 95.105 150.990 ;
        RECT 84.065 150.890 84.805 150.920 ;
        RECT 75.875 150.720 83.875 150.870 ;
        RECT 75.635 150.640 83.875 150.720 ;
        RECT 84.965 150.640 92.965 150.870 ;
        RECT 93.585 150.640 95.105 150.920 ;
        RECT 75.635 150.440 83.825 150.640 ;
        RECT 74.385 150.360 83.825 150.440 ;
        RECT 84.975 150.370 92.885 150.640 ;
        RECT 93.585 150.530 95.085 150.640 ;
        RECT 74.385 149.970 76.215 150.360 ;
        RECT 73.195 147.870 73.515 149.660 ;
        RECT 75.635 149.430 76.215 149.970 ;
        RECT 77.365 149.430 78.665 150.360 ;
        RECT 81.705 150.160 83.005 150.360 ;
        RECT 86.965 150.160 88.265 150.370 ;
        RECT 81.705 149.750 88.265 150.160 ;
        RECT 81.705 149.430 83.005 149.750 ;
        RECT 86.965 149.460 88.265 149.750 ;
        RECT 90.895 149.460 92.195 150.370 ;
        RECT 94.105 149.990 95.085 150.530 ;
        RECT 95.335 149.990 96.335 150.990 ;
        RECT 95.605 149.700 96.315 149.990 ;
        RECT 96.775 149.900 97.775 150.900 ;
        RECT 96.795 149.700 97.795 149.710 ;
        RECT 75.445 149.190 83.355 149.430 ;
        RECT 86.705 149.190 94.615 149.460 ;
        RECT 95.605 149.315 97.795 149.700 ;
        RECT 98.945 149.315 99.265 149.330 ;
        RECT 95.605 149.270 99.265 149.315 ;
        RECT 74.250 148.960 84.250 149.190 ;
        RECT 85.430 148.960 95.430 149.190 ;
        RECT 73.765 148.910 74.035 148.940 ;
        RECT 84.475 148.910 85.205 148.930 ;
        RECT 73.765 148.600 74.045 148.910 ;
        RECT 84.455 148.600 85.225 148.910 ;
        RECT 73.765 147.800 74.035 148.600 ;
        RECT 74.250 148.320 84.250 148.550 ;
        RECT 74.595 147.990 83.565 148.320 ;
        RECT 84.605 147.800 85.055 148.600 ;
        RECT 85.430 148.320 95.430 148.550 ;
        RECT 85.975 148.070 94.945 148.320 ;
        RECT 95.605 147.800 95.975 149.270 ;
        RECT 96.795 149.080 99.265 149.270 ;
        RECT 96.795 148.710 97.795 149.080 ;
        RECT 98.945 149.070 99.265 149.080 ;
        RECT 73.765 147.530 95.975 147.800 ;
        RECT 96.775 147.130 97.775 148.130 ;
        RECT 73.115 146.830 74.115 146.840 ;
        RECT 73.115 146.630 74.925 146.830 ;
        RECT 71.760 146.095 74.925 146.630 ;
        RECT 75.415 146.580 93.445 146.940 ;
        RECT 71.760 141.265 72.295 146.095 ;
        RECT 73.115 145.840 74.925 146.095 ;
        RECT 73.665 145.830 74.925 145.840 ;
        RECT 73.195 145.530 74.195 145.610 ;
        RECT 73.195 144.650 74.205 145.530 ;
        RECT 74.395 145.090 74.925 145.830 ;
        RECT 75.425 145.550 75.725 146.580 ;
        RECT 76.085 146.160 83.605 146.440 ;
        RECT 75.885 145.930 83.885 146.160 ;
        RECT 84.145 145.940 84.745 146.580 ;
        RECT 85.295 146.160 92.815 146.420 ;
        RECT 84.075 145.880 84.815 145.940 ;
        RECT 84.975 145.930 92.975 146.160 ;
        RECT 93.165 145.880 93.445 146.580 ;
        RECT 84.045 145.570 84.815 145.880 ;
        RECT 93.135 145.870 93.445 145.880 ;
        RECT 93.135 145.640 93.845 145.870 ;
        RECT 94.105 145.780 95.105 146.780 ;
        RECT 95.355 146.440 96.355 146.780 ;
        RECT 96.765 146.440 103.630 146.760 ;
        RECT 95.355 145.780 103.630 146.440 ;
        RECT 96.765 145.760 103.630 145.780 ;
        RECT 93.135 145.570 95.115 145.640 ;
        RECT 84.075 145.540 84.815 145.570 ;
        RECT 75.885 145.370 83.885 145.520 ;
        RECT 75.645 145.290 83.885 145.370 ;
        RECT 84.975 145.290 92.975 145.520 ;
        RECT 93.595 145.290 95.115 145.570 ;
        RECT 75.645 145.090 83.835 145.290 ;
        RECT 74.395 145.010 83.835 145.090 ;
        RECT 84.985 145.020 92.895 145.290 ;
        RECT 93.595 145.180 95.095 145.290 ;
        RECT 73.195 144.610 74.195 144.650 ;
        RECT 74.395 144.620 76.225 145.010 ;
        RECT 73.215 142.480 73.535 144.270 ;
        RECT 75.645 144.080 76.225 144.620 ;
        RECT 77.375 144.080 78.675 145.010 ;
        RECT 81.715 144.810 83.015 145.010 ;
        RECT 86.975 144.810 88.275 145.020 ;
        RECT 81.715 144.400 88.275 144.810 ;
        RECT 81.715 144.080 83.015 144.400 ;
        RECT 86.975 144.110 88.275 144.400 ;
        RECT 90.905 144.110 92.205 145.020 ;
        RECT 94.115 144.640 95.095 145.180 ;
        RECT 95.345 144.640 96.345 145.640 ;
        RECT 95.615 144.430 96.345 144.640 ;
        RECT 96.775 145.265 97.775 145.600 ;
        RECT 96.775 145.260 99.940 145.265 ;
        RECT 96.775 145.000 99.965 145.260 ;
        RECT 96.775 144.995 99.940 145.000 ;
        RECT 96.775 144.600 97.775 144.995 ;
        RECT 75.455 143.840 83.365 144.080 ;
        RECT 86.715 143.840 94.625 144.110 ;
        RECT 95.615 144.055 97.785 144.430 ;
        RECT 95.615 144.040 100.550 144.055 ;
        RECT 74.260 143.610 84.260 143.840 ;
        RECT 85.440 143.610 95.440 143.840 ;
        RECT 73.775 143.560 74.045 143.590 ;
        RECT 84.485 143.560 85.215 143.580 ;
        RECT 73.775 143.250 74.055 143.560 ;
        RECT 84.465 143.250 85.235 143.560 ;
        RECT 73.775 142.450 74.045 143.250 ;
        RECT 74.260 142.970 84.260 143.200 ;
        RECT 74.605 142.640 83.575 142.970 ;
        RECT 84.615 142.450 85.065 143.250 ;
        RECT 85.440 142.970 95.440 143.200 ;
        RECT 85.985 142.720 94.955 142.970 ;
        RECT 95.615 142.450 95.985 144.040 ;
        RECT 96.785 143.780 100.565 144.040 ;
        RECT 96.785 143.765 100.550 143.780 ;
        RECT 96.785 143.430 97.785 143.765 ;
        RECT 73.775 142.180 95.985 142.450 ;
        RECT 102.630 143.175 103.630 145.760 ;
        RECT 105.660 146.665 106.660 151.040 ;
        RECT 108.770 149.065 110.200 151.310 ;
        RECT 108.800 148.860 110.110 149.065 ;
        RECT 105.660 146.605 107.120 146.665 ;
        RECT 108.800 146.605 110.110 147.220 ;
        RECT 105.660 145.605 110.190 146.605 ;
        RECT 105.810 144.560 107.120 145.605 ;
        RECT 108.800 145.115 110.110 145.605 ;
        RECT 102.630 142.920 107.110 143.175 ;
        RECT 102.630 142.175 107.120 142.920 ;
        RECT 105.810 141.835 107.120 142.175 ;
        RECT 72.935 141.480 73.935 141.490 ;
        RECT 72.935 141.265 74.895 141.480 ;
        RECT 71.760 140.730 74.895 141.265 ;
        RECT 75.385 141.230 93.415 141.590 ;
        RECT 71.760 136.000 72.295 140.730 ;
        RECT 72.935 140.490 74.895 140.730 ;
        RECT 73.635 140.480 74.895 140.490 ;
        RECT 73.165 140.190 74.165 140.260 ;
        RECT 73.165 139.310 74.175 140.190 ;
        RECT 74.365 139.740 74.895 140.480 ;
        RECT 75.395 140.200 75.695 141.230 ;
        RECT 76.055 140.810 83.575 141.090 ;
        RECT 75.855 140.580 83.855 140.810 ;
        RECT 84.115 140.590 84.715 141.230 ;
        RECT 85.265 140.810 92.785 141.070 ;
        RECT 84.045 140.530 84.785 140.590 ;
        RECT 84.945 140.580 92.945 140.810 ;
        RECT 93.135 140.530 93.415 141.230 ;
        RECT 84.015 140.220 84.785 140.530 ;
        RECT 93.105 140.520 93.415 140.530 ;
        RECT 93.105 140.290 93.815 140.520 ;
        RECT 94.075 140.430 95.075 141.430 ;
        RECT 95.325 141.280 96.325 141.430 ;
        RECT 96.745 141.280 103.810 141.540 ;
        RECT 95.325 140.550 103.810 141.280 ;
        RECT 105.810 140.835 110.270 141.835 ;
        RECT 105.810 140.815 107.120 140.835 ;
        RECT 95.325 140.430 96.325 140.550 ;
        RECT 96.745 140.540 103.810 140.550 ;
        RECT 93.105 140.220 95.085 140.290 ;
        RECT 84.045 140.190 84.785 140.220 ;
        RECT 75.855 140.020 83.855 140.170 ;
        RECT 75.615 139.940 83.855 140.020 ;
        RECT 84.945 139.940 92.945 140.170 ;
        RECT 93.565 139.940 95.085 140.220 ;
        RECT 75.615 139.740 83.805 139.940 ;
        RECT 74.365 139.660 83.805 139.740 ;
        RECT 84.955 139.670 92.865 139.940 ;
        RECT 93.565 139.830 95.065 139.940 ;
        RECT 73.165 139.260 74.165 139.310 ;
        RECT 74.365 139.270 76.195 139.660 ;
        RECT 73.175 137.130 73.495 138.920 ;
        RECT 75.615 138.730 76.195 139.270 ;
        RECT 77.345 138.730 78.645 139.660 ;
        RECT 81.685 139.460 82.985 139.660 ;
        RECT 86.945 139.460 88.245 139.670 ;
        RECT 81.685 139.050 88.245 139.460 ;
        RECT 81.685 138.730 82.985 139.050 ;
        RECT 86.945 138.760 88.245 139.050 ;
        RECT 90.875 138.760 92.175 139.670 ;
        RECT 94.085 139.290 95.065 139.830 ;
        RECT 95.315 139.290 96.315 140.290 ;
        RECT 96.755 140.055 97.755 140.370 ;
        RECT 96.755 139.720 101.245 140.055 ;
        RECT 96.755 139.370 97.755 139.720 ;
        RECT 95.585 139.070 96.305 139.290 ;
        RECT 96.755 139.070 97.755 139.200 ;
        RECT 95.585 138.925 97.755 139.070 ;
        RECT 75.425 138.490 83.335 138.730 ;
        RECT 86.685 138.490 94.595 138.760 ;
        RECT 95.585 138.630 101.790 138.925 ;
        RECT 74.230 138.260 84.230 138.490 ;
        RECT 85.410 138.260 95.410 138.490 ;
        RECT 73.745 138.210 74.015 138.240 ;
        RECT 84.455 138.210 85.185 138.230 ;
        RECT 73.745 137.900 74.025 138.210 ;
        RECT 84.435 137.900 85.205 138.210 ;
        RECT 73.745 137.100 74.015 137.900 ;
        RECT 74.230 137.620 84.230 137.850 ;
        RECT 74.575 137.290 83.545 137.620 ;
        RECT 84.585 137.100 85.035 137.900 ;
        RECT 85.410 137.620 95.410 137.850 ;
        RECT 85.955 137.370 94.925 137.620 ;
        RECT 95.585 137.100 95.955 138.630 ;
        RECT 96.755 138.535 101.790 138.630 ;
        RECT 96.755 138.200 97.755 138.535 ;
        RECT 102.810 138.485 103.810 140.540 ;
        RECT 108.920 139.250 110.230 140.835 ;
        RECT 102.810 137.485 106.220 138.485 ;
        RECT 73.745 136.830 95.955 137.100 ;
        RECT 105.220 136.925 106.220 137.485 ;
        RECT 108.920 136.925 110.230 137.610 ;
        RECT 72.925 136.000 74.935 136.200 ;
        RECT 71.760 135.430 74.935 136.000 ;
        RECT 75.425 135.950 93.455 136.310 ;
        RECT 96.815 136.150 104.210 136.390 ;
        RECT 71.885 135.395 74.935 135.430 ;
        RECT 72.925 135.200 74.935 135.395 ;
        RECT 73.205 133.980 74.205 134.980 ;
        RECT 74.405 134.460 74.935 135.200 ;
        RECT 75.435 134.920 75.735 135.950 ;
        RECT 76.095 135.530 83.615 135.810 ;
        RECT 75.895 135.300 83.895 135.530 ;
        RECT 84.155 135.310 84.755 135.950 ;
        RECT 85.305 135.530 92.825 135.790 ;
        RECT 84.085 135.250 84.825 135.310 ;
        RECT 84.985 135.300 92.985 135.530 ;
        RECT 93.175 135.250 93.455 135.950 ;
        RECT 84.055 134.940 84.825 135.250 ;
        RECT 93.145 135.240 93.455 135.250 ;
        RECT 93.145 135.010 93.855 135.240 ;
        RECT 94.115 135.150 95.115 136.150 ;
        RECT 95.365 135.390 104.210 136.150 ;
        RECT 105.220 135.925 110.230 136.925 ;
        RECT 95.365 135.150 96.365 135.390 ;
        RECT 93.145 134.940 95.125 135.010 ;
        RECT 84.085 134.910 84.825 134.940 ;
        RECT 75.895 134.740 83.895 134.890 ;
        RECT 75.655 134.660 83.895 134.740 ;
        RECT 84.985 134.660 92.985 134.890 ;
        RECT 93.605 134.660 95.125 134.940 ;
        RECT 75.655 134.460 83.845 134.660 ;
        RECT 74.405 134.380 83.845 134.460 ;
        RECT 84.995 134.390 92.905 134.660 ;
        RECT 93.605 134.550 95.105 134.660 ;
        RECT 74.405 133.990 76.235 134.380 ;
        RECT 73.215 131.950 73.535 133.740 ;
        RECT 75.655 133.450 76.235 133.990 ;
        RECT 77.385 133.450 78.685 134.380 ;
        RECT 81.725 134.180 83.025 134.380 ;
        RECT 86.985 134.180 88.285 134.390 ;
        RECT 81.725 133.770 88.285 134.180 ;
        RECT 81.725 133.450 83.025 133.770 ;
        RECT 86.985 133.480 88.285 133.770 ;
        RECT 90.915 133.480 92.215 134.390 ;
        RECT 94.125 134.010 95.105 134.550 ;
        RECT 95.355 134.020 96.355 135.010 ;
        RECT 96.815 134.865 97.815 135.250 ;
        RECT 96.815 134.430 102.415 134.865 ;
        RECT 96.815 134.250 97.815 134.430 ;
        RECT 96.815 134.020 97.815 134.030 ;
        RECT 95.355 134.010 97.815 134.020 ;
        RECT 95.625 133.685 97.815 134.010 ;
        RECT 75.465 133.210 83.375 133.450 ;
        RECT 86.725 133.210 94.635 133.480 ;
        RECT 95.625 133.400 103.015 133.685 ;
        RECT 74.270 132.980 84.270 133.210 ;
        RECT 85.450 132.980 95.450 133.210 ;
        RECT 73.785 132.930 74.055 132.960 ;
        RECT 84.495 132.930 85.225 132.950 ;
        RECT 73.785 132.620 74.065 132.930 ;
        RECT 84.475 132.620 85.245 132.930 ;
        RECT 73.785 131.820 74.055 132.620 ;
        RECT 74.270 132.340 84.270 132.570 ;
        RECT 74.615 132.010 83.585 132.340 ;
        RECT 84.625 131.820 85.075 132.620 ;
        RECT 85.450 132.340 95.450 132.570 ;
        RECT 85.995 132.090 94.965 132.340 ;
        RECT 95.625 131.820 95.995 133.400 ;
        RECT 96.815 133.180 103.015 133.400 ;
        RECT 96.815 133.030 97.815 133.180 ;
        RECT 73.785 131.550 95.995 131.820 ;
        RECT 103.210 132.025 104.210 135.390 ;
        RECT 105.810 134.650 107.120 135.925 ;
        RECT 108.920 135.505 110.230 135.925 ;
        RECT 105.810 132.025 107.120 133.010 ;
        RECT 103.210 131.025 110.270 132.025 ;
        RECT 105.810 130.905 107.120 131.025 ;
        RECT 73.105 130.415 74.925 130.610 ;
        RECT 70.055 129.590 71.465 129.860 ;
        RECT 71.785 129.880 74.925 130.415 ;
        RECT 75.415 130.360 93.445 130.720 ;
        RECT 71.785 127.545 72.320 129.880 ;
        RECT 73.105 129.610 74.925 129.880 ;
        RECT 72.635 128.390 74.195 129.390 ;
        RECT 74.395 128.870 74.925 129.610 ;
        RECT 75.425 129.330 75.725 130.360 ;
        RECT 76.085 129.940 83.605 130.220 ;
        RECT 75.885 129.710 83.885 129.940 ;
        RECT 84.145 129.720 84.745 130.360 ;
        RECT 85.295 129.940 92.815 130.200 ;
        RECT 84.075 129.660 84.815 129.720 ;
        RECT 84.975 129.710 92.975 129.940 ;
        RECT 93.165 129.660 93.445 130.360 ;
        RECT 84.045 129.350 84.815 129.660 ;
        RECT 93.135 129.650 93.445 129.660 ;
        RECT 93.135 129.420 93.845 129.650 ;
        RECT 94.105 129.560 95.105 130.560 ;
        RECT 95.355 130.240 96.355 130.560 ;
        RECT 96.785 130.240 101.850 130.470 ;
        RECT 95.355 129.630 101.850 130.240 ;
        RECT 95.355 129.560 96.355 129.630 ;
        RECT 96.785 129.470 101.850 129.630 ;
        RECT 93.135 129.350 95.115 129.420 ;
        RECT 84.075 129.320 84.815 129.350 ;
        RECT 75.885 129.150 83.885 129.300 ;
        RECT 75.645 129.070 83.885 129.150 ;
        RECT 84.975 129.070 92.975 129.300 ;
        RECT 93.595 129.070 95.115 129.350 ;
        RECT 75.645 128.870 83.835 129.070 ;
        RECT 74.395 128.790 83.835 128.870 ;
        RECT 84.985 128.800 92.895 129.070 ;
        RECT 93.595 128.960 95.095 129.070 ;
        RECT 74.395 128.400 76.225 128.790 ;
        RECT 71.150 126.795 72.425 127.545 ;
        RECT 34.370 125.300 67.870 126.300 ;
        RECT 34.370 3.490 35.450 125.300 ;
        RECT 71.785 125.035 72.320 126.795 ;
        RECT 73.205 126.300 73.525 128.090 ;
        RECT 75.645 127.860 76.225 128.400 ;
        RECT 77.375 127.860 78.675 128.790 ;
        RECT 81.715 128.590 83.015 128.790 ;
        RECT 86.975 128.590 88.275 128.800 ;
        RECT 81.715 128.180 88.275 128.590 ;
        RECT 81.715 127.860 83.015 128.180 ;
        RECT 86.975 127.890 88.275 128.180 ;
        RECT 90.905 127.890 92.205 128.800 ;
        RECT 94.115 128.420 95.095 128.960 ;
        RECT 95.345 128.420 96.345 129.420 ;
        RECT 95.615 128.130 96.325 128.420 ;
        RECT 96.785 128.330 97.785 129.330 ;
        RECT 96.805 128.130 97.805 128.140 ;
        RECT 75.455 127.620 83.365 127.860 ;
        RECT 86.715 127.620 94.625 127.890 ;
        RECT 95.615 127.700 97.805 128.130 ;
        RECT 74.260 127.390 84.260 127.620 ;
        RECT 85.440 127.390 95.440 127.620 ;
        RECT 73.775 127.340 74.045 127.370 ;
        RECT 84.485 127.340 85.215 127.360 ;
        RECT 73.775 127.030 74.055 127.340 ;
        RECT 84.465 127.030 85.235 127.340 ;
        RECT 73.775 126.230 74.045 127.030 ;
        RECT 74.260 126.750 84.260 126.980 ;
        RECT 74.605 126.420 83.575 126.750 ;
        RECT 84.615 126.230 85.065 127.030 ;
        RECT 85.440 126.750 95.440 126.980 ;
        RECT 85.985 126.500 94.955 126.750 ;
        RECT 95.615 126.230 95.985 127.700 ;
        RECT 96.805 127.140 97.805 127.700 ;
        RECT 100.850 126.895 101.850 129.470 ;
        RECT 108.920 129.260 110.230 131.025 ;
        RECT 108.920 126.895 110.230 127.620 ;
        RECT 73.775 125.960 95.985 126.230 ;
        RECT 96.785 125.560 97.785 126.560 ;
        RECT 100.850 125.895 110.230 126.895 ;
        RECT 73.125 125.260 74.125 125.270 ;
        RECT 73.125 125.035 74.935 125.260 ;
        RECT 71.785 124.500 74.935 125.035 ;
        RECT 75.425 125.010 93.455 125.370 ;
        RECT 39.400 123.455 58.400 124.455 ;
        RECT 58.790 123.745 67.910 123.815 ;
        RECT 57.710 122.865 58.135 123.455 ;
        RECT 58.790 123.345 68.030 123.745 ;
        RECT 58.790 123.335 67.070 123.345 ;
        RECT 62.570 122.925 62.920 123.195 ;
        RECT 63.950 123.135 64.240 123.165 ;
        RECT 63.950 123.045 68.740 123.135 ;
        RECT 63.910 122.925 68.740 123.045 ;
        RECT 59.170 122.865 59.520 122.875 ;
        RECT 57.710 122.535 62.435 122.865 ;
        RECT 57.710 122.485 58.135 122.535 ;
        RECT 37.190 122.235 57.240 122.485 ;
        RECT 61.260 122.285 61.480 122.345 ;
        RECT 37.190 122.215 58.350 122.235 ;
        RECT 61.250 122.225 61.540 122.285 ;
        RECT 37.190 122.195 61.090 122.215 ;
        RECT 37.190 121.915 61.110 122.195 ;
        RECT 37.190 121.885 61.090 121.915 ;
        RECT 61.250 121.885 61.690 122.225 ;
        RECT 62.105 122.205 62.435 122.535 ;
        RECT 62.630 122.715 62.900 122.925 ;
        RECT 62.630 122.355 63.040 122.715 ;
        RECT 63.910 122.375 64.430 122.925 ;
        RECT 68.270 122.495 68.740 122.925 ;
        RECT 62.060 121.905 62.490 122.205 ;
        RECT 62.640 121.905 63.040 122.355 ;
        RECT 63.950 122.325 64.400 122.375 ;
        RECT 63.420 121.905 63.870 122.205 ;
        RECT 64.030 121.905 64.400 122.325 ;
        RECT 37.190 121.860 58.350 121.885 ;
        RECT 61.250 121.865 61.540 121.885 ;
        RECT 37.190 121.485 57.240 121.860 ;
        RECT 61.260 121.835 61.480 121.865 ;
        RECT 63.455 121.645 63.785 121.905 ;
        RECT 57.735 121.315 63.785 121.645 ;
        RECT 58.790 120.615 69.370 121.095 ;
        RECT 61.165 120.445 61.455 120.460 ;
        RECT 61.160 120.435 61.455 120.445 ;
        RECT 61.990 120.435 62.310 120.475 ;
        RECT 58.840 120.245 59.140 120.315 ;
        RECT 61.160 120.255 62.310 120.435 ;
        RECT 62.630 120.305 63.050 120.325 ;
        RECT 61.160 120.245 61.455 120.255 ;
        RECT 58.730 120.215 59.140 120.245 ;
        RECT 61.165 120.230 61.455 120.245 ;
        RECT 61.990 120.215 62.310 120.255 ;
        RECT 58.540 119.125 59.140 120.215 ;
        RECT 62.620 120.075 63.050 120.305 ;
        RECT 63.930 120.305 64.220 120.445 ;
        RECT 67.130 120.345 67.430 120.425 ;
        RECT 59.810 120.045 63.050 120.075 ;
        RECT 59.810 119.935 63.040 120.045 ;
        RECT 59.810 119.805 60.120 119.935 ;
        RECT 59.730 119.515 60.120 119.805 ;
        RECT 60.330 119.785 61.030 119.795 ;
        RECT 60.330 119.760 61.040 119.785 ;
        RECT 61.195 119.760 61.515 119.765 ;
        RECT 60.315 119.510 61.515 119.760 ;
        RECT 60.330 119.505 61.040 119.510 ;
        RECT 61.195 119.505 61.515 119.510 ;
        RECT 63.380 119.455 63.740 120.155 ;
        RECT 63.930 120.045 64.770 120.305 ;
        RECT 63.930 120.025 64.220 120.045 ;
        RECT 66.160 120.015 66.480 120.035 ;
        RECT 63.890 119.810 64.210 119.835 ;
        RECT 66.140 119.810 66.520 120.015 ;
        RECT 63.890 119.600 66.520 119.810 ;
        RECT 63.890 119.575 64.210 119.600 ;
        RECT 63.400 119.415 63.720 119.455 ;
        RECT 61.690 119.205 62.360 119.235 ;
        RECT 64.570 119.225 65.010 119.325 ;
        RECT 66.140 119.245 66.520 119.600 ;
        RECT 67.120 119.465 67.560 120.345 ;
        RECT 68.010 119.785 68.400 119.795 ;
        RECT 68.000 119.515 68.400 119.785 ;
        RECT 68.590 119.770 69.320 119.805 ;
        RECT 68.585 119.520 69.320 119.770 ;
        RECT 67.130 119.425 67.430 119.465 ;
        RECT 68.020 119.245 68.340 119.515 ;
        RECT 68.590 119.425 69.320 119.520 ;
        RECT 71.785 119.740 72.320 124.500 ;
        RECT 73.125 124.270 74.935 124.500 ;
        RECT 73.675 124.260 74.935 124.270 ;
        RECT 73.205 123.960 74.205 124.040 ;
        RECT 73.205 123.080 74.215 123.960 ;
        RECT 74.405 123.520 74.935 124.260 ;
        RECT 75.435 123.980 75.735 125.010 ;
        RECT 76.095 124.590 83.615 124.870 ;
        RECT 75.895 124.360 83.895 124.590 ;
        RECT 84.155 124.370 84.755 125.010 ;
        RECT 85.305 124.590 92.825 124.850 ;
        RECT 84.085 124.310 84.825 124.370 ;
        RECT 84.985 124.360 92.985 124.590 ;
        RECT 93.175 124.310 93.455 125.010 ;
        RECT 84.055 124.000 84.825 124.310 ;
        RECT 93.145 124.300 93.455 124.310 ;
        RECT 93.145 124.070 93.855 124.300 ;
        RECT 94.115 124.210 95.115 125.210 ;
        RECT 95.365 124.870 96.365 125.210 ;
        RECT 96.775 124.870 104.210 125.190 ;
        RECT 95.365 124.210 104.210 124.870 ;
        RECT 105.810 124.310 107.120 125.895 ;
        RECT 108.920 125.515 110.230 125.895 ;
        RECT 96.775 124.190 104.210 124.210 ;
        RECT 93.145 124.000 95.125 124.070 ;
        RECT 84.085 123.970 84.825 124.000 ;
        RECT 75.895 123.800 83.895 123.950 ;
        RECT 75.655 123.720 83.895 123.800 ;
        RECT 84.985 123.720 92.985 123.950 ;
        RECT 93.605 123.720 95.125 124.000 ;
        RECT 75.655 123.520 83.845 123.720 ;
        RECT 74.405 123.440 83.845 123.520 ;
        RECT 84.995 123.450 92.905 123.720 ;
        RECT 93.605 123.610 95.105 123.720 ;
        RECT 73.205 123.040 74.205 123.080 ;
        RECT 74.405 123.050 76.235 123.440 ;
        RECT 73.225 120.910 73.545 122.700 ;
        RECT 75.655 122.510 76.235 123.050 ;
        RECT 77.385 122.510 78.685 123.440 ;
        RECT 81.725 123.240 83.025 123.440 ;
        RECT 86.985 123.240 88.285 123.450 ;
        RECT 81.725 122.830 88.285 123.240 ;
        RECT 81.725 122.510 83.025 122.830 ;
        RECT 86.985 122.540 88.285 122.830 ;
        RECT 90.915 122.540 92.215 123.450 ;
        RECT 94.125 123.070 95.105 123.610 ;
        RECT 95.355 123.070 96.355 124.070 ;
        RECT 95.625 122.860 96.355 123.070 ;
        RECT 96.785 123.030 97.785 124.030 ;
        RECT 75.465 122.270 83.375 122.510 ;
        RECT 86.725 122.270 94.635 122.540 ;
        RECT 95.625 122.470 97.795 122.860 ;
        RECT 74.270 122.040 84.270 122.270 ;
        RECT 85.450 122.040 95.450 122.270 ;
        RECT 73.785 121.990 74.055 122.020 ;
        RECT 84.495 121.990 85.225 122.010 ;
        RECT 73.785 121.680 74.065 121.990 ;
        RECT 84.475 121.680 85.245 121.990 ;
        RECT 73.785 120.880 74.055 121.680 ;
        RECT 74.270 121.400 84.270 121.630 ;
        RECT 74.615 121.070 83.585 121.400 ;
        RECT 84.625 120.880 85.075 121.680 ;
        RECT 85.450 121.400 95.450 121.630 ;
        RECT 85.995 121.150 94.965 121.400 ;
        RECT 95.625 120.880 95.995 122.470 ;
        RECT 96.795 121.860 97.795 122.470 ;
        RECT 73.785 120.610 95.995 120.880 ;
        RECT 103.210 121.585 104.210 124.190 ;
        RECT 105.810 121.585 107.120 122.670 ;
        RECT 103.210 120.585 110.270 121.585 ;
        RECT 105.810 120.565 107.120 120.585 ;
        RECT 72.945 119.910 73.945 119.920 ;
        RECT 72.945 119.740 74.905 119.910 ;
        RECT 64.460 119.205 65.120 119.225 ;
        RECT 58.840 119.055 59.140 119.125 ;
        RECT 59.690 118.935 64.220 119.205 ;
        RECT 59.690 118.885 60.190 118.935 ;
        RECT 61.700 118.895 62.370 118.935 ;
        RECT 63.860 118.885 64.220 118.935 ;
        RECT 64.440 118.925 65.130 119.205 ;
        RECT 66.120 118.985 68.370 119.245 ;
        RECT 58.920 118.735 59.300 118.845 ;
        RECT 64.640 118.780 64.950 118.925 ;
        RECT 63.410 118.735 63.730 118.780 ;
        RECT 64.640 118.735 64.960 118.780 ;
        RECT 69.005 118.735 69.255 119.425 ;
        RECT 58.920 118.640 69.255 118.735 ;
        RECT 71.785 119.205 74.905 119.740 ;
        RECT 75.395 119.660 93.425 120.020 ;
        RECT 58.920 118.575 69.215 118.640 ;
        RECT 59.010 118.565 69.215 118.575 ;
        RECT 63.410 118.520 63.730 118.565 ;
        RECT 64.640 118.520 64.960 118.565 ;
        RECT 58.790 117.895 69.370 118.375 ;
        RECT 60.680 116.935 61.050 117.895 ;
        RECT 61.620 117.675 61.960 117.735 ;
        RECT 61.600 116.975 61.980 117.675 ;
        RECT 62.990 117.665 63.310 117.725 ;
        RECT 62.970 116.975 63.330 117.665 ;
        RECT 64.830 117.565 65.170 117.635 ;
        RECT 65.800 117.570 66.120 117.595 ;
        RECT 67.140 117.570 67.460 117.595 ;
        RECT 61.620 116.915 61.960 116.975 ;
        RECT 62.990 116.915 63.310 116.975 ;
        RECT 64.820 116.955 65.210 117.565 ;
        RECT 65.800 117.360 67.460 117.570 ;
        RECT 65.800 117.335 66.120 117.360 ;
        RECT 67.140 117.335 67.460 117.360 ;
        RECT 64.830 116.905 65.170 116.955 ;
        RECT 58.545 116.600 58.865 116.655 ;
        RECT 61.140 116.600 61.580 116.765 ;
        RECT 58.545 116.485 61.580 116.600 ;
        RECT 62.000 116.695 62.320 116.735 ;
        RECT 62.550 116.695 62.930 116.755 ;
        RECT 64.370 116.735 64.790 116.765 ;
        RECT 62.000 116.520 62.930 116.695 ;
        RECT 58.545 116.450 61.505 116.485 ;
        RECT 62.000 116.475 62.320 116.520 ;
        RECT 62.550 116.475 62.930 116.520 ;
        RECT 64.350 116.465 64.790 116.735 ;
        RECT 58.545 116.395 58.865 116.450 ;
        RECT 64.350 116.435 64.780 116.465 ;
        RECT 60.670 115.655 61.040 116.295 ;
        RECT 64.930 116.245 65.170 116.905 ;
        RECT 65.710 116.465 66.120 116.765 ;
        RECT 66.270 116.695 66.570 116.765 ;
        RECT 64.840 115.795 65.170 116.245 ;
        RECT 66.270 115.935 66.680 116.695 ;
        RECT 66.270 115.875 66.570 115.935 ;
        RECT 58.790 115.175 68.910 115.655 ;
        RECT 71.785 114.160 72.320 119.205 ;
        RECT 72.945 118.920 74.905 119.205 ;
        RECT 73.645 118.910 74.905 118.920 ;
        RECT 73.175 118.620 74.175 118.690 ;
        RECT 73.175 117.740 74.185 118.620 ;
        RECT 74.375 118.170 74.905 118.910 ;
        RECT 75.405 118.630 75.705 119.660 ;
        RECT 76.065 119.240 83.585 119.520 ;
        RECT 75.865 119.010 83.865 119.240 ;
        RECT 84.125 119.020 84.725 119.660 ;
        RECT 85.275 119.240 92.795 119.500 ;
        RECT 84.055 118.960 84.795 119.020 ;
        RECT 84.955 119.010 92.955 119.240 ;
        RECT 93.145 118.960 93.425 119.660 ;
        RECT 84.025 118.650 84.795 118.960 ;
        RECT 93.115 118.950 93.425 118.960 ;
        RECT 93.115 118.720 93.825 118.950 ;
        RECT 94.085 118.860 95.085 119.860 ;
        RECT 95.335 119.710 96.335 119.860 ;
        RECT 96.755 119.710 102.610 119.970 ;
        RECT 95.335 118.980 102.610 119.710 ;
        RECT 95.335 118.860 96.335 118.980 ;
        RECT 96.755 118.970 102.610 118.980 ;
        RECT 93.115 118.650 95.095 118.720 ;
        RECT 84.055 118.620 84.795 118.650 ;
        RECT 75.865 118.450 83.865 118.600 ;
        RECT 75.625 118.370 83.865 118.450 ;
        RECT 84.955 118.370 92.955 118.600 ;
        RECT 93.575 118.370 95.095 118.650 ;
        RECT 75.625 118.170 83.815 118.370 ;
        RECT 74.375 118.090 83.815 118.170 ;
        RECT 84.965 118.100 92.875 118.370 ;
        RECT 93.575 118.260 95.075 118.370 ;
        RECT 73.175 117.690 74.175 117.740 ;
        RECT 74.375 117.700 76.205 118.090 ;
        RECT 73.185 115.560 73.505 117.350 ;
        RECT 75.625 117.160 76.205 117.700 ;
        RECT 77.355 117.160 78.655 118.090 ;
        RECT 81.695 117.890 82.995 118.090 ;
        RECT 86.955 117.890 88.255 118.100 ;
        RECT 81.695 117.480 88.255 117.890 ;
        RECT 81.695 117.160 82.995 117.480 ;
        RECT 86.955 117.190 88.255 117.480 ;
        RECT 90.885 117.190 92.185 118.100 ;
        RECT 94.095 117.720 95.075 118.260 ;
        RECT 95.325 117.720 96.325 118.720 ;
        RECT 96.765 117.800 97.765 118.800 ;
        RECT 95.595 117.500 96.315 117.720 ;
        RECT 96.765 117.500 97.765 117.630 ;
        RECT 75.435 116.920 83.345 117.160 ;
        RECT 86.695 116.920 94.605 117.190 ;
        RECT 95.595 117.060 97.765 117.500 ;
        RECT 74.240 116.690 84.240 116.920 ;
        RECT 85.420 116.690 95.420 116.920 ;
        RECT 73.755 116.640 74.025 116.670 ;
        RECT 84.465 116.640 85.195 116.660 ;
        RECT 73.755 116.330 74.035 116.640 ;
        RECT 84.445 116.330 85.215 116.640 ;
        RECT 73.755 115.530 74.025 116.330 ;
        RECT 74.240 116.050 84.240 116.280 ;
        RECT 74.585 115.720 83.555 116.050 ;
        RECT 84.595 115.530 85.045 116.330 ;
        RECT 85.420 116.050 95.420 116.280 ;
        RECT 85.965 115.800 94.935 116.050 ;
        RECT 95.595 115.530 95.965 117.060 ;
        RECT 96.765 116.630 97.765 117.060 ;
        RECT 101.610 116.595 102.610 118.970 ;
        RECT 108.860 118.920 110.170 120.585 ;
        RECT 108.860 116.595 110.170 117.280 ;
        RECT 101.610 115.595 110.270 116.595 ;
        RECT 73.755 115.260 95.965 115.530 ;
        RECT 72.935 114.160 74.945 114.630 ;
        RECT 75.435 114.380 93.465 114.740 ;
        RECT 96.825 114.580 103.490 114.820 ;
        RECT 71.785 113.630 74.945 114.160 ;
        RECT 71.785 113.625 73.500 113.630 ;
        RECT 73.215 112.410 74.215 113.410 ;
        RECT 74.415 112.890 74.945 113.630 ;
        RECT 75.445 113.350 75.745 114.380 ;
        RECT 76.105 113.960 83.625 114.240 ;
        RECT 75.905 113.730 83.905 113.960 ;
        RECT 84.165 113.740 84.765 114.380 ;
        RECT 85.315 113.960 92.835 114.220 ;
        RECT 84.095 113.680 84.835 113.740 ;
        RECT 84.995 113.730 92.995 113.960 ;
        RECT 93.185 113.680 93.465 114.380 ;
        RECT 84.065 113.370 84.835 113.680 ;
        RECT 93.155 113.670 93.465 113.680 ;
        RECT 93.155 113.440 93.865 113.670 ;
        RECT 94.125 113.580 95.125 114.580 ;
        RECT 95.375 113.820 103.490 114.580 ;
        RECT 105.800 114.130 107.110 115.595 ;
        RECT 108.860 115.175 110.170 115.595 ;
        RECT 95.375 113.580 96.375 113.820 ;
        RECT 93.155 113.370 95.135 113.440 ;
        RECT 84.095 113.340 84.835 113.370 ;
        RECT 75.905 113.170 83.905 113.320 ;
        RECT 75.665 113.090 83.905 113.170 ;
        RECT 84.995 113.090 92.995 113.320 ;
        RECT 93.615 113.090 95.135 113.370 ;
        RECT 75.665 112.890 83.855 113.090 ;
        RECT 74.415 112.810 83.855 112.890 ;
        RECT 85.005 112.820 92.915 113.090 ;
        RECT 93.615 112.980 95.115 113.090 ;
        RECT 74.415 112.420 76.245 112.810 ;
        RECT 40.800 111.615 41.800 111.635 ;
        RECT 40.800 111.565 43.640 111.615 ;
        RECT 40.800 110.635 44.680 111.565 ;
        RECT 45.170 111.315 63.200 111.675 ;
        RECT 40.890 110.615 44.680 110.635 ;
        RECT 40.890 106.225 41.890 110.615 ;
        RECT 42.860 110.565 44.680 110.615 ;
        RECT 42.390 109.345 43.950 110.345 ;
        RECT 44.150 109.825 44.680 110.565 ;
        RECT 45.180 110.285 45.480 111.315 ;
        RECT 45.840 110.895 53.360 111.175 ;
        RECT 45.640 110.665 53.640 110.895 ;
        RECT 53.900 110.675 54.500 111.315 ;
        RECT 55.050 110.895 62.570 111.155 ;
        RECT 53.830 110.615 54.570 110.675 ;
        RECT 54.730 110.665 62.730 110.895 ;
        RECT 62.920 110.615 63.200 111.315 ;
        RECT 53.800 110.305 54.570 110.615 ;
        RECT 62.890 110.605 63.200 110.615 ;
        RECT 62.890 110.375 63.600 110.605 ;
        RECT 63.860 110.515 64.860 111.515 ;
        RECT 65.110 111.195 66.110 111.515 ;
        RECT 70.980 111.505 71.980 111.595 ;
        RECT 66.570 111.425 71.980 111.505 ;
        RECT 66.540 111.195 71.980 111.425 ;
        RECT 65.110 110.625 71.980 111.195 ;
        RECT 65.110 110.585 67.540 110.625 ;
        RECT 65.110 110.515 66.110 110.585 ;
        RECT 66.540 110.425 67.540 110.585 ;
        RECT 70.980 110.535 71.980 110.625 ;
        RECT 73.225 110.380 73.545 112.170 ;
        RECT 75.665 111.880 76.245 112.420 ;
        RECT 77.395 111.880 78.695 112.810 ;
        RECT 81.735 112.610 83.035 112.810 ;
        RECT 86.995 112.610 88.295 112.820 ;
        RECT 81.735 112.200 88.295 112.610 ;
        RECT 81.735 111.880 83.035 112.200 ;
        RECT 86.995 111.910 88.295 112.200 ;
        RECT 90.925 111.910 92.225 112.820 ;
        RECT 94.135 112.440 95.115 112.980 ;
        RECT 95.365 112.450 96.365 113.440 ;
        RECT 96.825 112.680 97.825 113.680 ;
        RECT 96.825 112.450 97.825 112.460 ;
        RECT 95.365 112.440 97.825 112.450 ;
        RECT 75.475 111.640 83.385 111.880 ;
        RECT 86.735 111.640 94.645 111.910 ;
        RECT 95.635 111.830 97.825 112.440 ;
        RECT 74.280 111.410 84.280 111.640 ;
        RECT 85.460 111.410 95.460 111.640 ;
        RECT 73.795 111.360 74.065 111.390 ;
        RECT 84.505 111.360 85.235 111.380 ;
        RECT 73.795 111.050 74.075 111.360 ;
        RECT 84.485 111.050 85.255 111.360 ;
        RECT 62.890 110.305 64.870 110.375 ;
        RECT 53.830 110.275 54.570 110.305 ;
        RECT 45.640 110.105 53.640 110.255 ;
        RECT 45.400 110.025 53.640 110.105 ;
        RECT 54.730 110.025 62.730 110.255 ;
        RECT 63.350 110.025 64.870 110.305 ;
        RECT 45.400 109.825 53.590 110.025 ;
        RECT 44.150 109.745 53.590 109.825 ;
        RECT 54.740 109.755 62.650 110.025 ;
        RECT 63.350 109.915 64.850 110.025 ;
        RECT 44.150 109.355 45.980 109.745 ;
        RECT 42.960 107.255 43.280 109.045 ;
        RECT 45.400 108.815 45.980 109.355 ;
        RECT 47.130 108.815 48.430 109.745 ;
        RECT 51.470 109.545 52.770 109.745 ;
        RECT 56.730 109.545 58.030 109.755 ;
        RECT 51.470 109.135 58.030 109.545 ;
        RECT 51.470 108.815 52.770 109.135 ;
        RECT 56.730 108.845 58.030 109.135 ;
        RECT 60.660 108.845 61.960 109.755 ;
        RECT 63.870 109.375 64.850 109.915 ;
        RECT 65.100 109.375 66.100 110.375 ;
        RECT 65.370 109.085 66.080 109.375 ;
        RECT 66.540 109.285 67.540 110.285 ;
        RECT 73.795 110.250 74.065 111.050 ;
        RECT 74.280 110.770 84.280 111.000 ;
        RECT 74.625 110.440 83.595 110.770 ;
        RECT 84.635 110.250 85.085 111.050 ;
        RECT 85.460 110.770 95.460 111.000 ;
        RECT 86.005 110.520 94.975 110.770 ;
        RECT 95.635 110.250 96.005 111.830 ;
        RECT 96.825 111.460 97.825 111.830 ;
        RECT 102.490 111.865 103.490 113.820 ;
        RECT 105.800 112.105 107.110 112.490 ;
        RECT 105.650 111.865 108.570 112.105 ;
        RECT 102.490 110.865 108.570 111.865 ;
        RECT 105.650 110.625 108.570 110.865 ;
        RECT 105.800 110.385 108.570 110.625 ;
        RECT 73.795 109.980 96.005 110.250 ;
        RECT 66.560 109.085 67.560 109.095 ;
        RECT 45.210 108.575 53.120 108.815 ;
        RECT 56.470 108.575 64.380 108.845 ;
        RECT 65.370 108.655 67.560 109.085 ;
        RECT 44.015 108.345 54.015 108.575 ;
        RECT 55.195 108.345 65.195 108.575 ;
        RECT 43.530 108.295 43.800 108.325 ;
        RECT 54.240 108.295 54.970 108.315 ;
        RECT 43.530 107.985 43.810 108.295 ;
        RECT 54.220 107.985 54.990 108.295 ;
        RECT 43.530 107.185 43.800 107.985 ;
        RECT 44.015 107.705 54.015 107.935 ;
        RECT 44.360 107.375 53.330 107.705 ;
        RECT 54.370 107.185 54.820 107.985 ;
        RECT 55.195 107.705 65.195 107.935 ;
        RECT 55.740 107.455 64.710 107.705 ;
        RECT 65.370 107.185 65.740 108.655 ;
        RECT 66.560 108.095 67.560 108.655 ;
        RECT 43.530 106.915 65.740 107.185 ;
        RECT 66.540 106.515 67.540 107.515 ;
        RECT 71.890 106.735 73.350 108.845 ;
        RECT 40.890 106.215 43.880 106.225 ;
        RECT 40.890 105.225 44.690 106.215 ;
        RECT 45.180 105.965 63.210 106.325 ;
        RECT 40.890 100.875 41.890 105.225 ;
        RECT 43.430 105.215 44.690 105.225 ;
        RECT 42.960 104.915 43.960 104.995 ;
        RECT 42.960 104.035 43.970 104.915 ;
        RECT 44.160 104.475 44.690 105.215 ;
        RECT 45.190 104.935 45.490 105.965 ;
        RECT 45.850 105.545 53.370 105.825 ;
        RECT 45.650 105.315 53.650 105.545 ;
        RECT 53.910 105.325 54.510 105.965 ;
        RECT 55.060 105.545 62.580 105.805 ;
        RECT 53.840 105.265 54.580 105.325 ;
        RECT 54.740 105.315 62.740 105.545 ;
        RECT 62.930 105.265 63.210 105.965 ;
        RECT 53.810 104.955 54.580 105.265 ;
        RECT 62.900 105.255 63.210 105.265 ;
        RECT 62.900 105.025 63.610 105.255 ;
        RECT 63.870 105.165 64.870 106.165 ;
        RECT 65.120 105.825 66.120 106.165 ;
        RECT 66.530 105.825 67.530 106.145 ;
        RECT 65.120 105.165 67.530 105.825 ;
        RECT 66.530 105.145 67.530 105.165 ;
        RECT 62.900 104.955 64.880 105.025 ;
        RECT 53.840 104.925 54.580 104.955 ;
        RECT 45.650 104.755 53.650 104.905 ;
        RECT 45.410 104.675 53.650 104.755 ;
        RECT 54.740 104.675 62.740 104.905 ;
        RECT 63.360 104.675 64.880 104.955 ;
        RECT 45.410 104.475 53.600 104.675 ;
        RECT 44.160 104.395 53.600 104.475 ;
        RECT 54.750 104.405 62.660 104.675 ;
        RECT 63.360 104.565 64.860 104.675 ;
        RECT 42.960 103.995 43.960 104.035 ;
        RECT 44.160 104.005 45.990 104.395 ;
        RECT 42.980 101.865 43.300 103.655 ;
        RECT 45.410 103.465 45.990 104.005 ;
        RECT 47.140 103.465 48.440 104.395 ;
        RECT 51.480 104.195 52.780 104.395 ;
        RECT 56.740 104.195 58.040 104.405 ;
        RECT 51.480 103.785 58.040 104.195 ;
        RECT 51.480 103.465 52.780 103.785 ;
        RECT 56.740 103.495 58.040 103.785 ;
        RECT 60.670 103.495 61.970 104.405 ;
        RECT 63.880 104.025 64.860 104.565 ;
        RECT 65.110 104.025 66.110 105.025 ;
        RECT 65.380 103.815 66.110 104.025 ;
        RECT 66.540 103.985 67.540 104.985 ;
        RECT 45.220 103.225 53.130 103.465 ;
        RECT 56.480 103.225 64.390 103.495 ;
        RECT 65.380 103.425 67.550 103.815 ;
        RECT 44.025 102.995 54.025 103.225 ;
        RECT 55.205 102.995 65.205 103.225 ;
        RECT 43.540 102.945 43.810 102.975 ;
        RECT 54.250 102.945 54.980 102.965 ;
        RECT 43.540 102.635 43.820 102.945 ;
        RECT 54.230 102.635 55.000 102.945 ;
        RECT 43.540 101.835 43.810 102.635 ;
        RECT 44.025 102.355 54.025 102.585 ;
        RECT 44.370 102.025 53.340 102.355 ;
        RECT 54.380 101.835 54.830 102.635 ;
        RECT 55.205 102.355 65.205 102.585 ;
        RECT 55.750 102.105 64.720 102.355 ;
        RECT 65.380 101.835 65.750 103.425 ;
        RECT 66.550 102.815 67.550 103.425 ;
        RECT 43.540 101.565 65.750 101.835 ;
        RECT 40.890 100.865 43.700 100.875 ;
        RECT 40.890 99.875 44.660 100.865 ;
        RECT 45.150 100.615 63.180 100.975 ;
        RECT 71.950 100.945 73.130 106.735 ;
        RECT 74.360 106.095 75.940 106.725 ;
        RECT 74.275 104.940 75.940 106.095 ;
        RECT 107.090 105.120 108.570 110.385 ;
        RECT 66.580 100.925 73.130 100.945 ;
        RECT 36.590 95.585 37.695 95.640 ;
        RECT 40.890 95.585 41.890 99.875 ;
        RECT 43.400 99.865 44.660 99.875 ;
        RECT 42.930 99.575 43.930 99.645 ;
        RECT 42.930 98.695 43.940 99.575 ;
        RECT 44.130 99.125 44.660 99.865 ;
        RECT 45.160 99.585 45.460 100.615 ;
        RECT 45.820 100.195 53.340 100.475 ;
        RECT 45.620 99.965 53.620 100.195 ;
        RECT 53.880 99.975 54.480 100.615 ;
        RECT 55.030 100.195 62.550 100.455 ;
        RECT 53.810 99.915 54.550 99.975 ;
        RECT 54.710 99.965 62.710 100.195 ;
        RECT 62.900 99.915 63.180 100.615 ;
        RECT 53.780 99.605 54.550 99.915 ;
        RECT 62.870 99.905 63.180 99.915 ;
        RECT 62.870 99.675 63.580 99.905 ;
        RECT 63.840 99.815 64.840 100.815 ;
        RECT 65.090 100.665 66.090 100.815 ;
        RECT 66.510 100.665 73.130 100.925 ;
        RECT 65.090 99.965 73.130 100.665 ;
        RECT 65.090 99.935 67.510 99.965 ;
        RECT 65.090 99.815 66.090 99.935 ;
        RECT 66.510 99.925 67.510 99.935 ;
        RECT 71.950 99.865 73.130 99.965 ;
        RECT 74.305 104.525 75.940 104.940 ;
        RECT 105.785 104.620 106.855 104.650 ;
        RECT 107.020 104.620 151.785 105.120 ;
        RECT 62.870 99.605 64.850 99.675 ;
        RECT 53.810 99.575 54.550 99.605 ;
        RECT 45.620 99.405 53.620 99.555 ;
        RECT 45.380 99.325 53.620 99.405 ;
        RECT 54.710 99.325 62.710 99.555 ;
        RECT 63.330 99.325 64.850 99.605 ;
        RECT 45.380 99.125 53.570 99.325 ;
        RECT 44.130 99.045 53.570 99.125 ;
        RECT 54.720 99.055 62.630 99.325 ;
        RECT 63.330 99.215 64.830 99.325 ;
        RECT 42.930 98.645 43.930 98.695 ;
        RECT 44.130 98.655 45.960 99.045 ;
        RECT 42.940 96.515 43.260 98.305 ;
        RECT 45.380 98.115 45.960 98.655 ;
        RECT 47.110 98.115 48.410 99.045 ;
        RECT 51.450 98.845 52.750 99.045 ;
        RECT 56.710 98.845 58.010 99.055 ;
        RECT 51.450 98.435 58.010 98.845 ;
        RECT 51.450 98.115 52.750 98.435 ;
        RECT 56.710 98.145 58.010 98.435 ;
        RECT 60.640 98.145 61.940 99.055 ;
        RECT 63.850 98.675 64.830 99.215 ;
        RECT 65.080 98.675 66.080 99.675 ;
        RECT 66.520 98.755 67.520 99.755 ;
        RECT 65.350 98.455 66.070 98.675 ;
        RECT 66.520 98.455 67.520 98.585 ;
        RECT 45.190 97.875 53.100 98.115 ;
        RECT 56.450 97.875 64.360 98.145 ;
        RECT 65.350 98.015 67.520 98.455 ;
        RECT 43.995 97.645 53.995 97.875 ;
        RECT 55.175 97.645 65.175 97.875 ;
        RECT 43.510 97.595 43.780 97.625 ;
        RECT 54.220 97.595 54.950 97.615 ;
        RECT 43.510 97.285 43.790 97.595 ;
        RECT 54.200 97.285 54.970 97.595 ;
        RECT 43.510 96.485 43.780 97.285 ;
        RECT 43.995 97.005 53.995 97.235 ;
        RECT 44.340 96.675 53.310 97.005 ;
        RECT 54.350 96.485 54.800 97.285 ;
        RECT 55.175 97.005 65.175 97.235 ;
        RECT 55.720 96.755 64.690 97.005 ;
        RECT 65.350 96.485 65.720 98.015 ;
        RECT 66.520 97.585 67.520 98.015 ;
        RECT 43.510 96.215 65.720 96.485 ;
        RECT 66.580 95.710 67.580 95.775 ;
        RECT 74.305 95.710 75.460 104.525 ;
        RECT 105.785 103.550 151.785 104.620 ;
        RECT 105.785 103.520 106.855 103.550 ;
        RECT 107.020 103.510 151.785 103.550 ;
        RECT 36.590 94.585 44.700 95.585 ;
        RECT 45.190 95.335 63.220 95.695 ;
        RECT 66.580 95.535 75.460 95.710 ;
        RECT 36.590 6.165 37.695 94.585 ;
        RECT 42.970 93.365 43.970 94.365 ;
        RECT 44.170 93.845 44.700 94.585 ;
        RECT 45.200 94.305 45.500 95.335 ;
        RECT 45.860 94.915 53.380 95.195 ;
        RECT 45.660 94.685 53.660 94.915 ;
        RECT 53.920 94.695 54.520 95.335 ;
        RECT 55.070 94.915 62.590 95.175 ;
        RECT 53.850 94.635 54.590 94.695 ;
        RECT 54.750 94.685 62.750 94.915 ;
        RECT 62.940 94.635 63.220 95.335 ;
        RECT 53.820 94.325 54.590 94.635 ;
        RECT 62.910 94.625 63.220 94.635 ;
        RECT 62.910 94.395 63.620 94.625 ;
        RECT 63.880 94.535 64.880 95.535 ;
        RECT 65.130 94.850 75.460 95.535 ;
        RECT 65.130 94.775 67.580 94.850 ;
        RECT 65.130 94.535 66.130 94.775 ;
        RECT 74.305 94.700 75.460 94.850 ;
        RECT 62.910 94.325 64.890 94.395 ;
        RECT 53.850 94.295 54.590 94.325 ;
        RECT 45.660 94.125 53.660 94.275 ;
        RECT 45.420 94.045 53.660 94.125 ;
        RECT 54.750 94.045 62.750 94.275 ;
        RECT 63.370 94.045 64.890 94.325 ;
        RECT 45.420 93.845 53.610 94.045 ;
        RECT 44.170 93.765 53.610 93.845 ;
        RECT 54.760 93.775 62.670 94.045 ;
        RECT 63.370 93.935 64.870 94.045 ;
        RECT 44.170 93.375 46.000 93.765 ;
        RECT 42.980 91.335 43.300 93.125 ;
        RECT 45.420 92.835 46.000 93.375 ;
        RECT 47.150 92.835 48.450 93.765 ;
        RECT 51.490 93.565 52.790 93.765 ;
        RECT 56.750 93.565 58.050 93.775 ;
        RECT 51.490 93.155 58.050 93.565 ;
        RECT 51.490 92.835 52.790 93.155 ;
        RECT 56.750 92.865 58.050 93.155 ;
        RECT 60.680 92.865 61.980 93.775 ;
        RECT 63.890 93.395 64.870 93.935 ;
        RECT 65.120 93.405 66.120 94.395 ;
        RECT 66.580 93.635 67.580 94.635 ;
        RECT 66.580 93.405 67.580 93.415 ;
        RECT 65.120 93.395 67.580 93.405 ;
        RECT 45.230 92.595 53.140 92.835 ;
        RECT 56.490 92.595 64.400 92.865 ;
        RECT 65.390 92.785 67.580 93.395 ;
        RECT 44.035 92.365 54.035 92.595 ;
        RECT 55.215 92.365 65.215 92.595 ;
        RECT 43.550 92.315 43.820 92.345 ;
        RECT 54.260 92.315 54.990 92.335 ;
        RECT 43.550 92.005 43.830 92.315 ;
        RECT 54.240 92.005 55.010 92.315 ;
        RECT 43.550 91.205 43.820 92.005 ;
        RECT 44.035 91.725 54.035 91.955 ;
        RECT 44.380 91.395 53.350 91.725 ;
        RECT 54.390 91.205 54.840 92.005 ;
        RECT 55.215 91.725 65.215 91.955 ;
        RECT 55.760 91.475 64.730 91.725 ;
        RECT 65.390 91.205 65.760 92.785 ;
        RECT 66.580 92.415 67.580 92.785 ;
        RECT 43.550 90.935 65.760 91.205 ;
        RECT 39.405 88.985 60.845 88.990 ;
        RECT 39.405 87.995 65.505 88.985 ;
        RECT 90.950 87.430 92.350 87.460 ;
        RECT 38.650 86.650 39.650 86.680 ;
        RECT 38.650 85.650 64.220 86.650 ;
        RECT 88.240 86.030 92.350 87.430 ;
        RECT 95.220 86.030 120.620 87.430 ;
        RECT 38.650 85.620 39.650 85.650 ;
        RECT 88.240 78.375 89.640 86.030 ;
        RECT 90.950 86.000 92.350 86.030 ;
        RECT 93.815 81.655 104.415 83.755 ;
        RECT 95.115 80.955 95.815 81.655 ;
        RECT 96.115 81.105 96.615 81.405 ;
        RECT 100.225 81.355 100.515 81.385 ;
        RECT 101.185 81.355 101.475 81.385 ;
        RECT 102.145 81.355 102.435 81.385 ;
        RECT 103.105 81.355 103.395 81.385 ;
        RECT 98.015 81.155 103.615 81.355 ;
        RECT 98.015 80.955 98.815 81.155 ;
        RECT 95.115 80.950 96.215 80.955 ;
        RECT 96.515 80.950 98.815 80.955 ;
        RECT 88.240 76.975 93.200 78.375 ;
        RECT 61.150 74.535 62.610 74.565 ;
        RECT 69.000 74.535 89.900 74.655 ;
        RECT 61.150 73.075 89.900 74.535 ;
        RECT 91.800 73.930 93.200 76.975 ;
        RECT 61.150 73.045 62.610 73.075 ;
        RECT 69.000 72.855 89.900 73.075 ;
        RECT 91.200 73.580 93.200 73.930 ;
        RECT 72.030 72.815 89.050 72.855 ;
        RECT 91.200 72.605 91.550 73.580 ;
        RECT 91.800 72.855 93.200 73.580 ;
        RECT 88.200 72.255 91.550 72.605 ;
        RECT 88.200 72.055 88.650 72.255 ;
        RECT 71.445 71.355 72.900 71.705 ;
        RECT 73.100 71.305 74.300 71.705 ;
        RECT 74.480 71.305 75.680 71.705 ;
        RECT 75.860 71.305 77.060 71.705 ;
        RECT 77.240 71.305 78.440 71.705 ;
        RECT 78.620 71.305 79.820 71.705 ;
        RECT 80.000 71.305 81.200 71.705 ;
        RECT 81.380 71.305 82.580 71.705 ;
        RECT 82.760 71.305 83.960 71.705 ;
        RECT 84.100 71.305 87.650 71.705 ;
        RECT 88.200 71.305 88.550 72.055 ;
        RECT 95.115 71.955 96.265 80.950 ;
        RECT 96.035 71.950 96.265 71.955 ;
        RECT 96.475 71.955 98.815 80.950 ;
        RECT 99.515 78.355 99.815 81.005 ;
        RECT 96.475 71.950 96.705 71.955 ;
        RECT 89.450 71.755 92.200 71.805 ;
        RECT 88.700 71.355 92.200 71.755 ;
        RECT 96.115 71.405 96.615 71.805 ;
        RECT 97.415 71.655 98.815 71.955 ;
        RECT 99.535 71.950 99.765 78.355 ;
        RECT 100.015 74.605 100.245 80.950 ;
        RECT 100.465 78.355 100.765 81.005 ;
        RECT 99.965 72.005 100.315 74.605 ;
        RECT 100.015 71.950 100.245 72.005 ;
        RECT 100.495 71.950 100.725 78.355 ;
        RECT 100.975 74.605 101.205 80.950 ;
        RECT 101.415 78.355 101.715 81.005 ;
        RECT 100.915 72.005 101.265 74.605 ;
        RECT 100.975 71.950 101.205 72.005 ;
        RECT 101.455 71.950 101.685 78.355 ;
        RECT 101.935 74.605 102.165 80.950 ;
        RECT 102.365 78.355 102.665 81.005 ;
        RECT 101.915 72.005 102.265 74.605 ;
        RECT 101.935 71.950 102.165 72.005 ;
        RECT 102.415 71.950 102.645 78.355 ;
        RECT 102.895 74.605 103.125 80.950 ;
        RECT 103.365 78.355 103.665 81.005 ;
        RECT 102.865 72.005 103.215 74.605 ;
        RECT 102.895 71.950 103.125 72.005 ;
        RECT 103.375 71.950 103.605 78.355 ;
        RECT 99.745 71.655 100.035 71.745 ;
        RECT 100.705 71.655 100.995 71.745 ;
        RECT 101.665 71.655 101.955 71.745 ;
        RECT 102.625 71.655 102.915 71.745 ;
        RECT 91.400 70.655 92.200 71.355 ;
        RECT 93.765 70.655 94.915 70.705 ;
        RECT 68.900 70.645 70.850 70.655 ;
        RECT 68.620 70.555 70.850 70.645 ;
        RECT 72.030 70.555 89.050 70.575 ;
        RECT 68.620 70.055 90.000 70.555 ;
        RECT 91.400 70.355 94.950 70.655 ;
        RECT 96.215 70.355 96.515 71.405 ;
        RECT 68.620 69.665 70.850 70.055 ;
        RECT 68.900 69.255 70.850 69.665 ;
        RECT 91.400 69.655 96.515 70.355 ;
        RECT 71.950 69.280 73.300 69.305 ;
        RECT 71.445 68.955 73.300 69.280 ;
        RECT 73.470 68.955 74.670 69.355 ;
        RECT 74.850 68.955 76.050 69.355 ;
        RECT 76.230 68.955 77.430 69.355 ;
        RECT 77.610 68.955 78.810 69.355 ;
        RECT 78.990 68.955 80.190 69.355 ;
        RECT 80.370 68.955 81.570 69.355 ;
        RECT 81.750 68.955 82.950 69.355 ;
        RECT 83.130 68.955 84.330 69.355 ;
        RECT 84.510 69.305 85.640 69.355 ;
        RECT 89.500 69.305 89.800 69.335 ;
        RECT 84.510 69.005 89.800 69.305 ;
        RECT 84.510 68.955 85.640 69.005 ;
        RECT 89.500 68.975 89.800 69.005 ;
        RECT 91.400 69.255 94.950 69.655 ;
        RECT 71.445 68.930 72.325 68.955 ;
        RECT 72.030 67.715 85.370 67.855 ;
        RECT 69.080 67.705 89.780 67.715 ;
        RECT 69.080 67.055 89.900 67.705 ;
        RECT 61.300 66.615 62.735 66.645 ;
        RECT 69.000 66.615 89.900 67.055 ;
        RECT 61.300 65.255 89.900 66.615 ;
        RECT 61.300 65.180 70.455 65.255 ;
        RECT 61.300 65.150 62.735 65.180 ;
        RECT 77.440 64.300 86.560 64.370 ;
        RECT 77.440 63.900 86.680 64.300 ;
        RECT 77.440 63.890 85.720 63.900 ;
        RECT 81.220 63.480 81.570 63.750 ;
        RECT 82.600 63.690 82.890 63.720 ;
        RECT 82.600 63.600 87.390 63.690 ;
        RECT 82.560 63.480 87.390 63.600 ;
        RECT 77.820 63.420 78.170 63.430 ;
        RECT 64.945 63.090 81.085 63.420 ;
        RECT 79.910 62.840 80.130 62.900 ;
        RECT 79.900 62.780 80.190 62.840 ;
        RECT 63.675 62.750 79.740 62.770 ;
        RECT 63.675 62.470 79.760 62.750 ;
        RECT 63.675 62.440 79.740 62.470 ;
        RECT 79.900 62.440 80.340 62.780 ;
        RECT 80.755 62.760 81.085 63.090 ;
        RECT 81.280 63.270 81.550 63.480 ;
        RECT 81.280 62.910 81.690 63.270 ;
        RECT 82.560 62.930 83.080 63.480 ;
        RECT 86.920 63.050 87.390 63.480 ;
        RECT 80.710 62.460 81.140 62.760 ;
        RECT 81.290 62.460 81.690 62.910 ;
        RECT 82.600 62.880 83.050 62.930 ;
        RECT 82.070 62.460 82.520 62.760 ;
        RECT 82.680 62.460 83.050 62.880 ;
        RECT 79.900 62.420 80.190 62.440 ;
        RECT 79.910 62.390 80.130 62.420 ;
        RECT 82.105 62.200 82.435 62.460 ;
        RECT 76.385 61.870 82.435 62.200 ;
        RECT 76.385 58.360 76.715 61.870 ;
        RECT 77.440 61.170 88.020 61.650 ;
        RECT 79.815 61.000 80.105 61.015 ;
        RECT 79.810 60.990 80.105 61.000 ;
        RECT 80.640 60.990 80.960 61.030 ;
        RECT 77.490 60.800 77.790 60.870 ;
        RECT 79.810 60.810 80.960 60.990 ;
        RECT 81.280 60.860 81.700 60.880 ;
        RECT 79.810 60.800 80.105 60.810 ;
        RECT 77.380 60.770 77.790 60.800 ;
        RECT 79.815 60.785 80.105 60.800 ;
        RECT 80.640 60.770 80.960 60.810 ;
        RECT 77.190 59.680 77.790 60.770 ;
        RECT 81.270 60.630 81.700 60.860 ;
        RECT 82.580 60.860 82.870 61.000 ;
        RECT 85.780 60.900 86.080 60.980 ;
        RECT 78.460 60.600 81.700 60.630 ;
        RECT 78.460 60.490 81.690 60.600 ;
        RECT 78.460 60.360 78.770 60.490 ;
        RECT 78.380 60.070 78.770 60.360 ;
        RECT 78.980 60.340 79.680 60.350 ;
        RECT 78.980 60.315 79.690 60.340 ;
        RECT 79.845 60.315 80.165 60.320 ;
        RECT 78.965 60.065 80.165 60.315 ;
        RECT 78.980 60.060 79.690 60.065 ;
        RECT 79.845 60.060 80.165 60.065 ;
        RECT 82.030 60.010 82.390 60.710 ;
        RECT 82.580 60.600 83.420 60.860 ;
        RECT 82.580 60.580 82.870 60.600 ;
        RECT 84.810 60.570 85.130 60.590 ;
        RECT 82.540 60.365 82.860 60.390 ;
        RECT 84.790 60.365 85.170 60.570 ;
        RECT 82.540 60.155 85.170 60.365 ;
        RECT 82.540 60.130 82.860 60.155 ;
        RECT 82.050 59.970 82.370 60.010 ;
        RECT 80.340 59.760 81.010 59.790 ;
        RECT 83.220 59.780 83.660 59.880 ;
        RECT 84.790 59.800 85.170 60.155 ;
        RECT 85.770 60.020 86.210 60.900 ;
        RECT 86.660 60.340 87.050 60.350 ;
        RECT 86.650 60.070 87.050 60.340 ;
        RECT 87.240 60.325 87.970 60.360 ;
        RECT 87.235 60.075 87.970 60.325 ;
        RECT 85.780 59.980 86.080 60.020 ;
        RECT 86.670 59.800 86.990 60.070 ;
        RECT 87.240 59.980 87.970 60.075 ;
        RECT 83.110 59.760 83.770 59.780 ;
        RECT 77.490 59.610 77.790 59.680 ;
        RECT 78.340 59.490 82.870 59.760 ;
        RECT 78.340 59.440 78.840 59.490 ;
        RECT 80.350 59.450 81.020 59.490 ;
        RECT 82.510 59.440 82.870 59.490 ;
        RECT 83.090 59.480 83.780 59.760 ;
        RECT 84.770 59.540 87.020 59.800 ;
        RECT 77.570 59.290 77.950 59.400 ;
        RECT 83.290 59.335 83.600 59.480 ;
        RECT 82.060 59.290 82.380 59.335 ;
        RECT 83.290 59.290 83.610 59.335 ;
        RECT 87.655 59.290 87.905 59.980 ;
        RECT 77.570 59.195 87.905 59.290 ;
        RECT 77.570 59.130 87.865 59.195 ;
        RECT 77.660 59.120 87.865 59.130 ;
        RECT 82.060 59.075 82.380 59.120 ;
        RECT 83.290 59.075 83.610 59.120 ;
        RECT 77.440 58.450 88.020 58.930 ;
        RECT 79.330 57.490 79.700 58.450 ;
        RECT 80.270 58.230 80.610 58.290 ;
        RECT 80.250 57.530 80.630 58.230 ;
        RECT 81.640 58.220 81.960 58.280 ;
        RECT 81.620 57.530 81.980 58.220 ;
        RECT 83.480 58.120 83.820 58.190 ;
        RECT 84.450 58.125 84.770 58.150 ;
        RECT 85.790 58.125 86.110 58.150 ;
        RECT 80.270 57.470 80.610 57.530 ;
        RECT 81.640 57.470 81.960 57.530 ;
        RECT 83.470 57.510 83.860 58.120 ;
        RECT 84.450 57.915 86.110 58.125 ;
        RECT 84.450 57.890 84.770 57.915 ;
        RECT 85.790 57.890 86.110 57.915 ;
        RECT 83.480 57.460 83.820 57.510 ;
        RECT 77.195 57.155 77.515 57.210 ;
        RECT 79.790 57.155 80.230 57.320 ;
        RECT 77.195 57.040 80.230 57.155 ;
        RECT 80.650 57.250 80.970 57.290 ;
        RECT 81.200 57.250 81.580 57.310 ;
        RECT 83.020 57.290 83.440 57.320 ;
        RECT 80.650 57.075 81.580 57.250 ;
        RECT 77.195 57.005 80.155 57.040 ;
        RECT 80.650 57.030 80.970 57.075 ;
        RECT 81.200 57.030 81.580 57.075 ;
        RECT 83.000 57.020 83.440 57.290 ;
        RECT 77.195 56.950 77.515 57.005 ;
        RECT 83.000 56.990 83.430 57.020 ;
        RECT 79.320 56.210 79.690 56.850 ;
        RECT 83.580 56.800 83.820 57.460 ;
        RECT 84.360 57.020 84.770 57.320 ;
        RECT 84.920 57.250 85.220 57.320 ;
        RECT 83.490 56.350 83.820 56.800 ;
        RECT 84.920 56.490 85.330 57.250 ;
        RECT 84.920 56.430 85.220 56.490 ;
        RECT 77.440 55.730 87.560 56.210 ;
        RECT 59.420 52.120 62.540 52.175 ;
        RECT 59.420 51.175 63.330 52.120 ;
        RECT 63.820 51.870 81.850 52.230 ;
        RECT 59.420 46.780 60.420 51.175 ;
        RECT 61.510 51.120 63.330 51.175 ;
        RECT 61.040 49.900 62.600 50.900 ;
        RECT 62.800 50.380 63.330 51.120 ;
        RECT 63.830 50.840 64.130 51.870 ;
        RECT 64.490 51.450 72.010 51.730 ;
        RECT 64.290 51.220 72.290 51.450 ;
        RECT 72.550 51.230 73.150 51.870 ;
        RECT 73.700 51.450 81.220 51.710 ;
        RECT 72.480 51.170 73.220 51.230 ;
        RECT 73.380 51.220 81.380 51.450 ;
        RECT 81.570 51.170 81.850 51.870 ;
        RECT 72.450 50.860 73.220 51.170 ;
        RECT 81.540 51.160 81.850 51.170 ;
        RECT 81.540 50.930 82.250 51.160 ;
        RECT 82.510 51.070 83.510 52.070 ;
        RECT 83.760 51.750 84.760 52.070 ;
        RECT 91.400 51.985 92.800 69.255 ;
        RECT 96.215 68.905 96.515 69.655 ;
        RECT 96.115 68.555 96.665 68.905 ;
        RECT 97.415 68.655 103.615 71.655 ;
        RECT 103.865 70.520 105.865 70.805 ;
        RECT 103.865 69.470 132.925 70.520 ;
        RECT 103.865 69.355 105.865 69.470 ;
        RECT 96.035 68.255 96.265 68.405 ;
        RECT 95.015 65.455 96.265 68.255 ;
        RECT 95.015 64.755 95.815 65.455 ;
        RECT 96.035 65.405 96.265 65.455 ;
        RECT 96.475 68.255 96.705 68.405 ;
        RECT 97.415 68.255 98.815 68.655 ;
        RECT 100.225 68.565 100.515 68.655 ;
        RECT 101.185 68.565 101.475 68.655 ;
        RECT 102.145 68.565 102.435 68.655 ;
        RECT 103.105 68.565 103.395 68.655 ;
        RECT 96.475 65.455 98.815 68.255 ;
        RECT 99.535 66.605 99.765 68.405 ;
        RECT 100.015 68.255 100.245 68.405 ;
        RECT 99.965 67.055 100.315 68.255 ;
        RECT 96.475 65.405 96.705 65.455 ;
        RECT 97.915 65.255 98.815 65.455 ;
        RECT 99.465 65.405 99.815 66.605 ;
        RECT 100.015 65.405 100.245 67.055 ;
        RECT 100.495 66.605 100.725 68.405 ;
        RECT 100.975 68.255 101.205 68.405 ;
        RECT 100.915 67.055 101.265 68.255 ;
        RECT 100.415 65.405 100.765 66.605 ;
        RECT 100.975 65.405 101.205 67.055 ;
        RECT 101.455 66.605 101.685 68.405 ;
        RECT 101.935 68.255 102.165 68.405 ;
        RECT 101.915 67.055 102.265 68.255 ;
        RECT 101.415 65.405 101.765 66.605 ;
        RECT 101.935 65.405 102.165 67.055 ;
        RECT 102.415 66.605 102.645 68.405 ;
        RECT 102.895 68.255 103.125 68.405 ;
        RECT 102.865 67.055 103.215 68.255 ;
        RECT 102.365 65.405 102.715 66.605 ;
        RECT 102.895 65.405 103.125 67.055 ;
        RECT 103.375 66.605 103.605 68.405 ;
        RECT 103.315 65.405 103.665 66.605 ;
        RECT 96.115 64.905 96.665 65.255 ;
        RECT 97.915 65.055 103.215 65.255 ;
        RECT 99.745 65.015 100.035 65.055 ;
        RECT 100.705 65.015 100.995 65.055 ;
        RECT 101.665 65.015 101.955 65.055 ;
        RECT 102.625 65.015 102.915 65.055 ;
        RECT 93.815 63.155 104.415 64.755 ;
        RECT 94.170 62.175 95.770 63.155 ;
        RECT 106.195 61.345 107.170 69.470 ;
        RECT 85.245 51.980 92.800 51.985 ;
        RECT 85.190 51.750 92.800 51.980 ;
        RECT 83.760 51.150 92.800 51.750 ;
        RECT 83.760 51.140 86.190 51.150 ;
        RECT 83.760 51.070 84.760 51.140 ;
        RECT 85.190 50.980 86.190 51.140 ;
        RECT 91.400 51.135 92.800 51.150 ;
        RECT 95.295 60.370 107.170 61.345 ;
        RECT 81.540 50.860 83.520 50.930 ;
        RECT 72.480 50.830 73.220 50.860 ;
        RECT 64.290 50.660 72.290 50.810 ;
        RECT 64.050 50.580 72.290 50.660 ;
        RECT 73.380 50.580 81.380 50.810 ;
        RECT 82.000 50.580 83.520 50.860 ;
        RECT 64.050 50.380 72.240 50.580 ;
        RECT 62.800 50.300 72.240 50.380 ;
        RECT 73.390 50.310 81.300 50.580 ;
        RECT 82.000 50.470 83.500 50.580 ;
        RECT 62.800 49.910 64.630 50.300 ;
        RECT 61.610 47.810 61.930 49.600 ;
        RECT 64.050 49.370 64.630 49.910 ;
        RECT 65.780 49.370 67.080 50.300 ;
        RECT 70.120 50.100 71.420 50.300 ;
        RECT 75.380 50.100 76.680 50.310 ;
        RECT 70.120 49.690 76.680 50.100 ;
        RECT 70.120 49.370 71.420 49.690 ;
        RECT 75.380 49.400 76.680 49.690 ;
        RECT 79.310 49.400 80.610 50.310 ;
        RECT 82.520 49.930 83.500 50.470 ;
        RECT 83.750 49.930 84.750 50.930 ;
        RECT 84.020 49.640 84.730 49.930 ;
        RECT 85.190 49.840 86.190 50.840 ;
        RECT 85.210 49.640 86.210 49.650 ;
        RECT 63.860 49.130 71.770 49.370 ;
        RECT 75.120 49.130 83.030 49.400 ;
        RECT 84.020 49.210 86.210 49.640 ;
        RECT 62.665 48.900 72.665 49.130 ;
        RECT 73.845 48.900 83.845 49.130 ;
        RECT 62.180 48.850 62.450 48.880 ;
        RECT 72.890 48.850 73.620 48.870 ;
        RECT 62.180 48.540 62.460 48.850 ;
        RECT 72.870 48.540 73.640 48.850 ;
        RECT 62.180 47.740 62.450 48.540 ;
        RECT 62.665 48.260 72.665 48.490 ;
        RECT 63.010 47.930 71.980 48.260 ;
        RECT 73.020 47.740 73.470 48.540 ;
        RECT 73.845 48.260 83.845 48.490 ;
        RECT 74.390 48.010 83.360 48.260 ;
        RECT 84.020 47.740 84.390 49.210 ;
        RECT 85.210 48.650 86.210 49.210 ;
        RECT 62.180 47.470 84.390 47.740 ;
        RECT 85.190 47.070 86.190 48.070 ;
        RECT 59.420 46.770 62.530 46.780 ;
        RECT 59.420 45.780 63.340 46.770 ;
        RECT 63.830 46.520 81.860 46.880 ;
        RECT 59.420 41.430 60.420 45.780 ;
        RECT 62.080 45.770 63.340 45.780 ;
        RECT 61.610 45.470 62.610 45.550 ;
        RECT 61.610 44.590 62.620 45.470 ;
        RECT 62.810 45.030 63.340 45.770 ;
        RECT 63.840 45.490 64.140 46.520 ;
        RECT 64.500 46.100 72.020 46.380 ;
        RECT 64.300 45.870 72.300 46.100 ;
        RECT 72.560 45.880 73.160 46.520 ;
        RECT 73.710 46.100 81.230 46.360 ;
        RECT 72.490 45.820 73.230 45.880 ;
        RECT 73.390 45.870 81.390 46.100 ;
        RECT 81.580 45.820 81.860 46.520 ;
        RECT 72.460 45.510 73.230 45.820 ;
        RECT 81.550 45.810 81.860 45.820 ;
        RECT 81.550 45.580 82.260 45.810 ;
        RECT 82.520 45.720 83.520 46.720 ;
        RECT 83.770 46.380 84.770 46.720 ;
        RECT 85.180 46.675 86.180 46.700 ;
        RECT 95.295 46.675 96.270 60.370 ;
        RECT 131.875 60.120 132.925 69.470 ;
        RECT 103.270 56.115 141.450 56.595 ;
        RECT 109.780 55.235 110.100 55.295 ;
        RECT 111.175 55.235 111.465 55.280 ;
        RECT 109.780 55.095 111.465 55.235 ;
        RECT 109.780 55.035 110.100 55.095 ;
        RECT 111.175 55.050 111.465 55.095 ;
        RECT 108.400 54.215 108.720 54.275 ;
        RECT 110.255 54.215 110.545 54.260 ;
        RECT 108.400 54.075 110.545 54.215 ;
        RECT 108.400 54.015 108.720 54.075 ;
        RECT 110.255 54.030 110.545 54.075 ;
        RECT 103.270 53.395 141.450 53.875 ;
        RECT 103.270 50.675 141.450 51.155 ;
        RECT 105.640 49.795 105.960 49.855 ;
        RECT 107.955 49.795 108.245 49.840 ;
        RECT 105.640 49.655 108.245 49.795 ;
        RECT 105.640 49.595 105.960 49.655 ;
        RECT 107.955 49.610 108.245 49.655 ;
        RECT 108.400 49.255 108.720 49.515 ;
        RECT 109.795 49.115 110.085 49.160 ;
        RECT 112.080 49.115 112.400 49.175 ;
        RECT 109.795 48.975 112.400 49.115 ;
        RECT 109.795 48.930 110.085 48.975 ;
        RECT 112.080 48.915 112.400 48.975 ;
        RECT 103.270 47.955 141.450 48.435 ;
        RECT 109.780 47.415 110.070 47.460 ;
        RECT 111.350 47.415 111.640 47.460 ;
        RECT 113.450 47.415 113.740 47.460 ;
        RECT 109.780 47.275 113.740 47.415 ;
        RECT 109.780 47.230 110.070 47.275 ;
        RECT 111.350 47.230 111.640 47.275 ;
        RECT 113.450 47.230 113.740 47.275 ;
        RECT 109.345 47.075 109.635 47.120 ;
        RECT 111.865 47.075 112.155 47.120 ;
        RECT 113.055 47.075 113.345 47.120 ;
        RECT 109.345 46.935 113.345 47.075 ;
        RECT 109.345 46.890 109.635 46.935 ;
        RECT 111.865 46.890 112.155 46.935 ;
        RECT 113.055 46.890 113.345 46.935 ;
        RECT 85.180 46.380 96.270 46.675 ;
        RECT 108.860 46.735 109.180 46.795 ;
        RECT 113.935 46.735 114.225 46.780 ;
        RECT 108.860 46.595 114.225 46.735 ;
        RECT 108.860 46.535 109.180 46.595 ;
        RECT 113.935 46.550 114.225 46.595 ;
        RECT 83.770 45.815 96.270 46.380 ;
        RECT 112.080 46.395 112.400 46.455 ;
        RECT 112.600 46.395 112.890 46.440 ;
        RECT 112.080 46.255 112.890 46.395 ;
        RECT 112.080 46.195 112.400 46.255 ;
        RECT 112.600 46.210 112.890 46.255 ;
        RECT 105.640 46.055 105.960 46.115 ;
        RECT 107.035 46.055 107.325 46.100 ;
        RECT 105.640 45.915 107.325 46.055 ;
        RECT 105.640 45.855 105.960 45.915 ;
        RECT 107.035 45.870 107.325 45.915 ;
        RECT 83.770 45.810 95.250 45.815 ;
        RECT 83.770 45.720 86.180 45.810 ;
        RECT 85.180 45.700 86.180 45.720 ;
        RECT 81.550 45.510 83.530 45.580 ;
        RECT 72.490 45.480 73.230 45.510 ;
        RECT 64.300 45.310 72.300 45.460 ;
        RECT 64.060 45.230 72.300 45.310 ;
        RECT 73.390 45.230 81.390 45.460 ;
        RECT 82.010 45.230 83.530 45.510 ;
        RECT 64.060 45.030 72.250 45.230 ;
        RECT 62.810 44.950 72.250 45.030 ;
        RECT 73.400 44.960 81.310 45.230 ;
        RECT 82.010 45.120 83.510 45.230 ;
        RECT 61.610 44.550 62.610 44.590 ;
        RECT 62.810 44.560 64.640 44.950 ;
        RECT 61.630 42.420 61.950 44.210 ;
        RECT 64.060 44.020 64.640 44.560 ;
        RECT 65.790 44.020 67.090 44.950 ;
        RECT 70.130 44.750 71.430 44.950 ;
        RECT 75.390 44.750 76.690 44.960 ;
        RECT 70.130 44.340 76.690 44.750 ;
        RECT 70.130 44.020 71.430 44.340 ;
        RECT 75.390 44.050 76.690 44.340 ;
        RECT 79.320 44.050 80.620 44.960 ;
        RECT 82.530 44.580 83.510 45.120 ;
        RECT 83.760 44.580 84.760 45.580 ;
        RECT 84.030 44.370 84.760 44.580 ;
        RECT 85.190 44.540 86.190 45.540 ;
        RECT 103.270 45.235 141.450 45.715 ;
        RECT 106.080 45.035 106.370 45.080 ;
        RECT 113.000 45.035 113.320 45.095 ;
        RECT 106.080 44.895 113.320 45.035 ;
        RECT 106.080 44.850 106.370 44.895 ;
        RECT 113.000 44.835 113.320 44.895 ;
        RECT 108.400 44.695 108.720 44.755 ;
        RECT 105.270 44.555 108.720 44.695 ;
        RECT 105.270 44.400 105.410 44.555 ;
        RECT 108.400 44.495 108.720 44.555 ;
        RECT 63.870 43.780 71.780 44.020 ;
        RECT 75.130 43.780 83.040 44.050 ;
        RECT 84.030 43.980 86.200 44.370 ;
        RECT 105.195 44.170 105.485 44.400 ;
        RECT 105.640 44.155 105.960 44.415 ;
        RECT 112.540 44.400 112.860 44.415 ;
        RECT 106.575 44.170 106.865 44.400 ;
        RECT 112.540 44.170 112.890 44.400 ;
        RECT 62.675 43.550 72.675 43.780 ;
        RECT 73.855 43.550 83.855 43.780 ;
        RECT 62.190 43.500 62.460 43.530 ;
        RECT 72.900 43.500 73.630 43.520 ;
        RECT 62.190 43.190 62.470 43.500 ;
        RECT 72.880 43.190 73.650 43.500 ;
        RECT 62.190 42.390 62.460 43.190 ;
        RECT 62.675 42.910 72.675 43.140 ;
        RECT 63.020 42.580 71.990 42.910 ;
        RECT 73.030 42.390 73.480 43.190 ;
        RECT 73.855 42.910 83.855 43.140 ;
        RECT 74.400 42.660 83.370 42.910 ;
        RECT 84.030 42.390 84.400 43.980 ;
        RECT 85.200 43.370 86.200 43.980 ;
        RECT 106.100 43.675 106.420 43.735 ;
        RECT 106.650 43.675 106.790 44.170 ;
        RECT 112.540 44.155 112.860 44.170 ;
        RECT 109.345 44.015 109.635 44.060 ;
        RECT 111.865 44.015 112.155 44.060 ;
        RECT 113.055 44.015 113.345 44.060 ;
        RECT 109.345 43.875 113.345 44.015 ;
        RECT 109.345 43.830 109.635 43.875 ;
        RECT 111.865 43.830 112.155 43.875 ;
        RECT 113.055 43.830 113.345 43.875 ;
        RECT 113.935 43.830 114.225 44.060 ;
        RECT 107.035 43.675 107.325 43.720 ;
        RECT 106.100 43.535 107.325 43.675 ;
        RECT 106.100 43.475 106.420 43.535 ;
        RECT 107.035 43.490 107.325 43.535 ;
        RECT 109.780 43.675 110.070 43.720 ;
        RECT 111.350 43.675 111.640 43.720 ;
        RECT 113.450 43.675 113.740 43.720 ;
        RECT 109.780 43.535 113.740 43.675 ;
        RECT 109.780 43.490 110.070 43.535 ;
        RECT 111.350 43.490 111.640 43.535 ;
        RECT 113.450 43.490 113.740 43.535 ;
        RECT 108.860 43.335 109.180 43.395 ;
        RECT 114.010 43.335 114.150 43.830 ;
        RECT 108.860 43.195 114.150 43.335 ;
        RECT 108.860 43.135 109.180 43.195 ;
        RECT 103.270 42.515 141.450 42.995 ;
        RECT 62.190 42.120 84.400 42.390 ;
        RECT 106.100 42.315 106.420 42.375 ;
        RECT 109.795 42.315 110.085 42.360 ;
        RECT 106.100 42.175 110.085 42.315 ;
        RECT 106.100 42.115 106.420 42.175 ;
        RECT 109.795 42.130 110.085 42.175 ;
        RECT 112.540 42.315 112.860 42.375 ;
        RECT 113.015 42.315 113.305 42.360 ;
        RECT 112.540 42.175 113.305 42.315 ;
        RECT 112.540 42.115 112.860 42.175 ;
        RECT 113.015 42.130 113.305 42.175 ;
        RECT 112.080 41.635 112.400 41.695 ;
        RECT 112.555 41.635 112.845 41.680 ;
        RECT 59.420 41.420 62.350 41.430 ;
        RECT 59.420 40.430 63.310 41.420 ;
        RECT 63.800 41.170 81.830 41.530 ;
        RECT 112.080 41.495 114.150 41.635 ;
        RECT 59.420 36.140 60.420 40.430 ;
        RECT 62.050 40.420 63.310 40.430 ;
        RECT 61.580 40.130 62.580 40.200 ;
        RECT 61.580 39.250 62.590 40.130 ;
        RECT 62.780 39.680 63.310 40.420 ;
        RECT 63.810 40.140 64.110 41.170 ;
        RECT 64.470 40.750 71.990 41.030 ;
        RECT 64.270 40.520 72.270 40.750 ;
        RECT 72.530 40.530 73.130 41.170 ;
        RECT 73.680 40.750 81.200 41.010 ;
        RECT 72.460 40.470 73.200 40.530 ;
        RECT 73.360 40.520 81.360 40.750 ;
        RECT 81.550 40.470 81.830 41.170 ;
        RECT 72.430 40.160 73.200 40.470 ;
        RECT 81.520 40.460 81.830 40.470 ;
        RECT 81.520 40.230 82.230 40.460 ;
        RECT 82.490 40.370 83.490 41.370 ;
        RECT 83.740 41.220 84.740 41.370 ;
        RECT 85.160 41.220 86.160 41.480 ;
        RECT 112.080 41.435 112.400 41.495 ;
        RECT 112.555 41.450 112.845 41.495 ;
        RECT 83.740 41.165 86.160 41.220 ;
        RECT 83.740 40.645 97.300 41.165 ;
        RECT 113.000 41.095 113.320 41.355 ;
        RECT 114.010 41.340 114.150 41.495 ;
        RECT 113.935 41.110 114.225 41.340 ;
        RECT 105.180 40.955 105.500 41.015 ;
        RECT 108.875 40.955 109.165 41.000 ;
        RECT 111.635 40.955 111.925 41.000 ;
        RECT 105.180 40.815 109.165 40.955 ;
        RECT 105.180 40.755 105.500 40.815 ;
        RECT 108.875 40.770 109.165 40.815 ;
        RECT 110.790 40.815 111.925 40.955 ;
        RECT 83.740 40.490 86.160 40.645 ;
        RECT 83.740 40.370 84.740 40.490 ;
        RECT 85.160 40.480 86.160 40.490 ;
        RECT 81.520 40.160 83.500 40.230 ;
        RECT 72.460 40.130 73.200 40.160 ;
        RECT 64.270 39.960 72.270 40.110 ;
        RECT 64.030 39.880 72.270 39.960 ;
        RECT 73.360 39.880 81.360 40.110 ;
        RECT 81.980 39.880 83.500 40.160 ;
        RECT 64.030 39.680 72.220 39.880 ;
        RECT 62.780 39.600 72.220 39.680 ;
        RECT 73.370 39.610 81.280 39.880 ;
        RECT 81.980 39.770 83.480 39.880 ;
        RECT 61.580 39.200 62.580 39.250 ;
        RECT 62.780 39.210 64.610 39.600 ;
        RECT 61.590 37.070 61.910 38.860 ;
        RECT 64.030 38.670 64.610 39.210 ;
        RECT 65.760 38.670 67.060 39.600 ;
        RECT 70.100 39.400 71.400 39.600 ;
        RECT 75.360 39.400 76.660 39.610 ;
        RECT 70.100 38.990 76.660 39.400 ;
        RECT 70.100 38.670 71.400 38.990 ;
        RECT 75.360 38.700 76.660 38.990 ;
        RECT 79.290 38.700 80.590 39.610 ;
        RECT 82.500 39.230 83.480 39.770 ;
        RECT 83.730 39.230 84.730 40.230 ;
        RECT 85.170 39.310 86.170 40.310 ;
        RECT 84.000 39.010 84.720 39.230 ;
        RECT 85.170 39.010 86.170 39.140 ;
        RECT 63.840 38.430 71.750 38.670 ;
        RECT 75.100 38.430 83.010 38.700 ;
        RECT 84.000 38.570 86.170 39.010 ;
        RECT 62.645 38.200 72.645 38.430 ;
        RECT 73.825 38.200 83.825 38.430 ;
        RECT 62.160 38.150 62.430 38.180 ;
        RECT 72.870 38.150 73.600 38.170 ;
        RECT 62.160 37.840 62.440 38.150 ;
        RECT 72.850 37.840 73.620 38.150 ;
        RECT 62.160 37.040 62.430 37.840 ;
        RECT 62.645 37.560 72.645 37.790 ;
        RECT 62.990 37.230 71.960 37.560 ;
        RECT 73.000 37.040 73.450 37.840 ;
        RECT 73.825 37.560 83.825 37.790 ;
        RECT 74.370 37.310 83.340 37.560 ;
        RECT 84.000 37.040 84.370 38.570 ;
        RECT 85.170 38.140 86.170 38.570 ;
        RECT 62.160 36.770 84.370 37.040 ;
        RECT 59.420 35.140 63.350 36.140 ;
        RECT 63.840 35.890 81.870 36.250 ;
        RECT 85.230 36.120 86.230 36.330 ;
        RECT 85.230 36.090 94.010 36.120 ;
        RECT 59.420 9.060 60.420 35.140 ;
        RECT 61.620 33.920 62.620 34.920 ;
        RECT 62.820 34.400 63.350 35.140 ;
        RECT 63.850 34.860 64.150 35.890 ;
        RECT 64.510 35.470 72.030 35.750 ;
        RECT 64.310 35.240 72.310 35.470 ;
        RECT 72.570 35.250 73.170 35.890 ;
        RECT 73.720 35.470 81.240 35.730 ;
        RECT 72.500 35.190 73.240 35.250 ;
        RECT 73.400 35.240 81.400 35.470 ;
        RECT 81.590 35.190 81.870 35.890 ;
        RECT 72.470 34.880 73.240 35.190 ;
        RECT 81.560 35.180 81.870 35.190 ;
        RECT 81.560 34.950 82.270 35.180 ;
        RECT 82.530 35.090 83.530 36.090 ;
        RECT 83.780 35.565 94.010 36.090 ;
        RECT 83.780 35.330 86.230 35.565 ;
        RECT 83.780 35.090 84.780 35.330 ;
        RECT 81.560 34.880 83.540 34.950 ;
        RECT 72.500 34.850 73.240 34.880 ;
        RECT 64.310 34.680 72.310 34.830 ;
        RECT 64.070 34.600 72.310 34.680 ;
        RECT 73.400 34.600 81.400 34.830 ;
        RECT 82.020 34.600 83.540 34.880 ;
        RECT 64.070 34.400 72.260 34.600 ;
        RECT 62.820 34.320 72.260 34.400 ;
        RECT 73.410 34.330 81.320 34.600 ;
        RECT 82.020 34.490 83.520 34.600 ;
        RECT 62.820 33.930 64.650 34.320 ;
        RECT 61.630 31.890 61.950 33.680 ;
        RECT 64.070 33.390 64.650 33.930 ;
        RECT 65.800 33.390 67.100 34.320 ;
        RECT 70.140 34.120 71.440 34.320 ;
        RECT 75.400 34.120 76.700 34.330 ;
        RECT 70.140 33.710 76.700 34.120 ;
        RECT 70.140 33.390 71.440 33.710 ;
        RECT 75.400 33.420 76.700 33.710 ;
        RECT 79.330 33.420 80.630 34.330 ;
        RECT 82.540 33.950 83.520 34.490 ;
        RECT 83.770 33.960 84.770 34.950 ;
        RECT 85.230 34.190 86.230 35.190 ;
        RECT 85.230 33.960 86.230 33.970 ;
        RECT 83.770 33.950 86.230 33.960 ;
        RECT 63.880 33.150 71.790 33.390 ;
        RECT 75.140 33.150 83.050 33.420 ;
        RECT 84.040 33.340 86.230 33.950 ;
        RECT 62.685 32.920 72.685 33.150 ;
        RECT 73.865 32.920 83.865 33.150 ;
        RECT 62.200 32.870 62.470 32.900 ;
        RECT 72.910 32.870 73.640 32.890 ;
        RECT 62.200 32.560 62.480 32.870 ;
        RECT 72.890 32.560 73.660 32.870 ;
        RECT 62.200 31.760 62.470 32.560 ;
        RECT 62.685 32.280 72.685 32.510 ;
        RECT 63.030 31.950 72.000 32.280 ;
        RECT 73.040 31.760 73.490 32.560 ;
        RECT 73.865 32.280 83.865 32.510 ;
        RECT 74.410 32.030 83.380 32.280 ;
        RECT 84.040 31.760 84.410 33.340 ;
        RECT 85.230 32.970 86.230 33.340 ;
        RECT 62.200 31.490 84.410 31.760 ;
        RECT 93.455 11.700 94.010 35.565 ;
        RECT 96.780 12.865 97.300 40.645 ;
        RECT 108.400 40.615 108.720 40.675 ;
        RECT 110.790 40.660 110.930 40.815 ;
        RECT 111.635 40.770 111.925 40.815 ;
        RECT 109.875 40.615 110.165 40.660 ;
        RECT 108.400 40.475 110.165 40.615 ;
        RECT 108.400 40.415 108.720 40.475 ;
        RECT 109.875 40.430 110.165 40.475 ;
        RECT 110.715 40.430 111.005 40.660 ;
        RECT 103.270 39.795 141.450 40.275 ;
        RECT 103.270 37.075 141.450 37.555 ;
        RECT 108.860 36.675 109.180 36.935 ;
        RECT 127.735 35.855 128.025 35.900 ;
        RECT 131.860 35.855 132.180 35.915 ;
        RECT 127.735 35.715 132.180 35.855 ;
        RECT 127.735 35.670 128.025 35.715 ;
        RECT 131.860 35.655 132.180 35.715 ;
        RECT 115.315 35.330 115.605 35.560 ;
        RECT 115.390 35.175 115.530 35.330 ;
        RECT 121.295 35.175 121.585 35.220 ;
        RECT 124.960 35.175 125.280 35.235 ;
        RECT 115.390 35.035 125.280 35.175 ;
        RECT 121.295 34.990 121.585 35.035 ;
        RECT 124.960 34.975 125.280 35.035 ;
        RECT 103.270 34.355 141.450 34.835 ;
        RECT 119.455 34.155 119.745 34.200 ;
        RECT 129.100 34.155 129.420 34.215 ;
        RECT 130.495 34.155 130.785 34.200 ;
        RECT 119.455 34.015 130.785 34.155 ;
        RECT 119.455 33.970 119.745 34.015 ;
        RECT 129.100 33.955 129.420 34.015 ;
        RECT 130.495 33.970 130.785 34.015 ;
        RECT 125.130 33.815 125.420 33.860 ;
        RECT 126.800 33.815 127.120 33.875 ;
        RECT 125.130 33.675 127.120 33.815 ;
        RECT 125.130 33.630 125.420 33.675 ;
        RECT 126.800 33.615 127.120 33.675 ;
        RECT 127.735 33.475 128.025 33.520 ;
        RECT 119.070 33.335 128.025 33.475 ;
        RECT 119.070 33.180 119.210 33.335 ;
        RECT 127.735 33.290 128.025 33.335 ;
        RECT 128.180 33.475 128.500 33.535 ;
        RECT 130.955 33.475 131.245 33.520 ;
        RECT 128.180 33.335 131.245 33.475 ;
        RECT 128.180 33.275 128.500 33.335 ;
        RECT 130.955 33.290 131.245 33.335 ;
        RECT 131.415 33.475 131.705 33.520 ;
        RECT 131.860 33.475 132.180 33.535 ;
        RECT 136.475 33.475 136.765 33.520 ;
        RECT 131.415 33.335 132.180 33.475 ;
        RECT 131.415 33.290 131.705 33.335 ;
        RECT 131.860 33.275 132.180 33.335 ;
        RECT 135.170 33.335 136.765 33.475 ;
        RECT 116.695 32.950 116.985 33.180 ;
        RECT 118.995 32.950 119.285 33.180 ;
        RECT 121.765 33.135 122.055 33.180 ;
        RECT 124.285 33.135 124.575 33.180 ;
        RECT 125.475 33.135 125.765 33.180 ;
        RECT 121.765 32.995 125.765 33.135 ;
        RECT 121.765 32.950 122.055 32.995 ;
        RECT 124.285 32.950 124.575 32.995 ;
        RECT 125.475 32.950 125.765 32.995 ;
        RECT 116.770 32.455 116.910 32.950 ;
        RECT 126.340 32.935 126.660 33.195 ;
        RECT 132.780 32.935 133.100 33.195 ;
        RECT 135.170 33.180 135.310 33.335 ;
        RECT 136.475 33.290 136.765 33.335 ;
        RECT 135.095 32.950 135.385 33.180 ;
        RECT 118.520 32.595 118.840 32.855 ;
        RECT 122.200 32.795 122.490 32.840 ;
        RECT 123.770 32.795 124.060 32.840 ;
        RECT 125.870 32.795 126.160 32.840 ;
        RECT 119.070 32.655 120.130 32.795 ;
        RECT 119.070 32.455 119.210 32.655 ;
        RECT 119.990 32.515 120.130 32.655 ;
        RECT 122.200 32.655 126.160 32.795 ;
        RECT 122.200 32.610 122.490 32.655 ;
        RECT 123.770 32.610 124.060 32.655 ;
        RECT 125.870 32.610 126.160 32.655 ;
        RECT 126.800 32.595 127.120 32.855 ;
        RECT 127.720 32.795 128.040 32.855 ;
        RECT 129.575 32.795 129.865 32.840 ;
        RECT 127.720 32.655 129.865 32.795 ;
        RECT 127.720 32.595 128.040 32.655 ;
        RECT 129.575 32.610 129.865 32.655 ;
        RECT 134.635 32.795 134.925 32.840 ;
        RECT 134.635 32.655 135.310 32.795 ;
        RECT 134.635 32.610 134.925 32.655 ;
        RECT 135.170 32.515 135.310 32.655 ;
        RECT 116.770 32.315 119.210 32.455 ;
        RECT 119.900 32.455 120.220 32.515 ;
        RECT 132.335 32.455 132.625 32.500 ;
        RECT 119.900 32.315 132.625 32.455 ;
        RECT 119.900 32.255 120.220 32.315 ;
        RECT 132.335 32.270 132.625 32.315 ;
        RECT 135.080 32.255 135.400 32.515 ;
        RECT 135.540 32.255 135.860 32.515 ;
        RECT 103.270 31.635 141.450 32.115 ;
        RECT 112.080 31.435 112.400 31.495 ;
        RECT 128.180 31.435 128.500 31.495 ;
        RECT 112.080 31.295 128.500 31.435 ;
        RECT 112.080 31.235 112.400 31.295 ;
        RECT 128.180 31.235 128.500 31.295 ;
        RECT 109.360 31.095 109.650 31.140 ;
        RECT 111.460 31.095 111.750 31.140 ;
        RECT 113.030 31.095 113.320 31.140 ;
        RECT 109.360 30.955 113.320 31.095 ;
        RECT 109.360 30.910 109.650 30.955 ;
        RECT 111.460 30.910 111.750 30.955 ;
        RECT 113.030 30.910 113.320 30.955 ;
        RECT 115.300 31.095 115.620 31.155 ;
        RECT 115.775 31.095 116.065 31.140 ;
        RECT 124.960 31.095 125.280 31.155 ;
        RECT 127.720 31.095 128.040 31.155 ;
        RECT 115.300 30.955 128.040 31.095 ;
        RECT 115.300 30.895 115.620 30.955 ;
        RECT 115.775 30.910 116.065 30.955 ;
        RECT 124.960 30.895 125.280 30.955 ;
        RECT 127.720 30.895 128.040 30.955 ;
        RECT 108.860 30.555 109.180 30.815 ;
        RECT 109.755 30.755 110.045 30.800 ;
        RECT 110.945 30.755 111.235 30.800 ;
        RECT 113.465 30.755 113.755 30.800 ;
        RECT 122.200 30.755 122.520 30.815 ;
        RECT 109.755 30.615 113.755 30.755 ;
        RECT 109.755 30.570 110.045 30.615 ;
        RECT 110.945 30.570 111.235 30.615 ;
        RECT 113.465 30.570 113.755 30.615 ;
        RECT 119.070 30.615 122.520 30.755 ;
        RECT 107.495 30.230 107.785 30.460 ;
        RECT 108.415 30.415 108.705 30.460 ;
        RECT 112.540 30.415 112.860 30.475 ;
        RECT 119.070 30.460 119.210 30.615 ;
        RECT 122.200 30.555 122.520 30.615 ;
        RECT 123.135 30.755 123.425 30.800 ;
        RECT 128.640 30.755 128.960 30.815 ;
        RECT 123.135 30.615 128.960 30.755 ;
        RECT 123.135 30.570 123.425 30.615 ;
        RECT 128.640 30.555 128.960 30.615 ;
        RECT 108.415 30.275 112.860 30.415 ;
        RECT 108.415 30.230 108.705 30.275 ;
        RECT 107.570 30.075 107.710 30.230 ;
        RECT 112.540 30.215 112.860 30.275 ;
        RECT 118.995 30.230 119.285 30.460 ;
        RECT 119.900 30.215 120.220 30.475 ;
        RECT 121.295 30.415 121.585 30.460 ;
        RECT 121.740 30.415 122.060 30.475 ;
        RECT 122.675 30.415 122.965 30.460 ;
        RECT 124.990 30.415 125.280 30.460 ;
        RECT 121.295 30.275 122.965 30.415 ;
        RECT 121.295 30.230 121.585 30.275 ;
        RECT 121.740 30.215 122.060 30.275 ;
        RECT 122.675 30.230 122.965 30.275 ;
        RECT 123.210 30.275 125.280 30.415 ;
        RECT 110.210 30.075 110.500 30.120 ;
        RECT 113.000 30.075 113.320 30.135 ;
        RECT 123.210 30.075 123.350 30.275 ;
        RECT 124.990 30.230 125.280 30.275 ;
        RECT 125.880 30.415 126.200 30.475 ;
        RECT 126.355 30.415 126.645 30.460 ;
        RECT 125.880 30.275 126.645 30.415 ;
        RECT 125.880 30.215 126.200 30.275 ;
        RECT 126.355 30.230 126.645 30.275 ;
        RECT 107.570 29.935 108.630 30.075 ;
        RECT 104.720 29.735 105.040 29.795 ;
        RECT 107.955 29.735 108.245 29.780 ;
        RECT 104.720 29.595 108.245 29.735 ;
        RECT 108.490 29.735 108.630 29.935 ;
        RECT 110.210 29.935 113.320 30.075 ;
        RECT 110.210 29.890 110.500 29.935 ;
        RECT 113.000 29.875 113.320 29.935 ;
        RECT 119.070 29.935 123.350 30.075 ;
        RECT 119.070 29.795 119.210 29.935 ;
        RECT 112.080 29.735 112.400 29.795 ;
        RECT 108.490 29.595 112.400 29.735 ;
        RECT 104.720 29.535 105.040 29.595 ;
        RECT 107.955 29.550 108.245 29.595 ;
        RECT 112.080 29.535 112.400 29.595 ;
        RECT 118.980 29.535 119.300 29.795 ;
        RECT 122.200 29.535 122.520 29.795 ;
        RECT 124.975 29.735 125.265 29.780 ;
        RECT 125.420 29.735 125.740 29.795 ;
        RECT 124.975 29.595 125.740 29.735 ;
        RECT 124.975 29.550 125.265 29.595 ;
        RECT 125.420 29.535 125.740 29.595 ;
        RECT 125.880 29.535 126.200 29.795 ;
        RECT 126.340 29.735 126.660 29.795 ;
        RECT 130.940 29.735 131.260 29.795 ;
        RECT 132.795 29.735 133.085 29.780 ;
        RECT 126.340 29.595 133.085 29.735 ;
        RECT 126.340 29.535 126.660 29.595 ;
        RECT 130.940 29.535 131.260 29.595 ;
        RECT 132.795 29.550 133.085 29.595 ;
        RECT 103.270 28.915 141.450 29.395 ;
        RECT 112.540 28.715 112.860 28.775 ;
        RECT 113.015 28.715 113.305 28.760 ;
        RECT 112.540 28.575 113.305 28.715 ;
        RECT 112.540 28.515 112.860 28.575 ;
        RECT 113.015 28.530 113.305 28.575 ;
        RECT 119.900 28.715 120.220 28.775 ;
        RECT 131.860 28.715 132.180 28.775 ;
        RECT 119.900 28.575 132.180 28.715 ;
        RECT 119.900 28.515 120.220 28.575 ;
        RECT 131.860 28.515 132.180 28.575 ;
        RECT 107.940 28.375 108.260 28.435 ;
        RECT 108.860 28.375 109.180 28.435 ;
        RECT 119.990 28.375 120.130 28.515 ;
        RECT 106.190 28.235 109.180 28.375 ;
        RECT 104.720 27.835 105.040 28.095 ;
        RECT 105.640 27.835 105.960 28.095 ;
        RECT 106.190 28.080 106.330 28.235 ;
        RECT 107.940 28.175 108.260 28.235 ;
        RECT 108.860 28.175 109.180 28.235 ;
        RECT 119.070 28.235 120.130 28.375 ;
        RECT 122.200 28.375 122.520 28.435 ;
        RECT 122.980 28.375 123.270 28.420 ;
        RECT 122.200 28.235 123.270 28.375 ;
        RECT 106.115 27.850 106.405 28.080 ;
        RECT 107.395 28.035 107.685 28.080 ;
        RECT 106.650 27.895 107.685 28.035 ;
        RECT 105.195 27.695 105.485 27.740 ;
        RECT 106.650 27.695 106.790 27.895 ;
        RECT 107.395 27.850 107.685 27.895 ;
        RECT 115.300 27.835 115.620 28.095 ;
        RECT 105.195 27.555 106.790 27.695 ;
        RECT 106.995 27.695 107.285 27.740 ;
        RECT 108.185 27.695 108.475 27.740 ;
        RECT 110.705 27.695 110.995 27.740 ;
        RECT 106.995 27.555 110.995 27.695 ;
        RECT 105.195 27.510 105.485 27.555 ;
        RECT 106.995 27.510 107.285 27.555 ;
        RECT 108.185 27.510 108.475 27.555 ;
        RECT 110.705 27.510 110.995 27.555 ;
        RECT 113.000 27.695 113.320 27.755 ;
        RECT 113.475 27.695 113.765 27.740 ;
        RECT 113.000 27.555 113.765 27.695 ;
        RECT 113.000 27.495 113.320 27.555 ;
        RECT 113.475 27.510 113.765 27.555 ;
        RECT 115.775 27.510 116.065 27.740 ;
        RECT 106.600 27.355 106.890 27.400 ;
        RECT 108.700 27.355 108.990 27.400 ;
        RECT 110.270 27.355 110.560 27.400 ;
        RECT 106.600 27.215 110.560 27.355 ;
        RECT 115.850 27.355 115.990 27.510 ;
        RECT 118.520 27.495 118.840 27.755 ;
        RECT 119.070 27.695 119.210 28.235 ;
        RECT 122.200 28.175 122.520 28.235 ;
        RECT 122.980 28.190 123.270 28.235 ;
        RECT 132.290 28.375 132.580 28.420 ;
        RECT 135.540 28.375 135.860 28.435 ;
        RECT 132.290 28.235 135.860 28.375 ;
        RECT 132.290 28.190 132.580 28.235 ;
        RECT 135.540 28.175 135.860 28.235 ;
        RECT 120.835 28.035 121.125 28.080 ;
        RECT 121.280 28.035 121.600 28.095 ;
        RECT 128.180 28.035 128.500 28.095 ;
        RECT 129.100 28.035 129.420 28.095 ;
        RECT 120.835 27.895 129.420 28.035 ;
        RECT 120.835 27.850 121.125 27.895 ;
        RECT 121.280 27.835 121.600 27.895 ;
        RECT 128.180 27.835 128.500 27.895 ;
        RECT 129.100 27.835 129.420 27.895 ;
        RECT 130.940 27.835 131.260 28.095 ;
        RECT 119.455 27.695 119.745 27.740 ;
        RECT 119.070 27.555 119.745 27.695 ;
        RECT 119.455 27.510 119.745 27.555 ;
        RECT 119.915 27.510 120.205 27.740 ;
        RECT 118.980 27.355 119.300 27.415 ;
        RECT 115.850 27.215 119.300 27.355 ;
        RECT 119.990 27.355 120.130 27.510 ;
        RECT 120.360 27.495 120.680 27.755 ;
        RECT 121.755 27.510 122.045 27.740 ;
        RECT 122.635 27.695 122.925 27.740 ;
        RECT 123.825 27.695 124.115 27.740 ;
        RECT 126.345 27.695 126.635 27.740 ;
        RECT 122.635 27.555 126.635 27.695 ;
        RECT 122.635 27.510 122.925 27.555 ;
        RECT 123.825 27.510 124.115 27.555 ;
        RECT 126.345 27.510 126.635 27.555 ;
        RECT 131.835 27.695 132.125 27.740 ;
        RECT 133.025 27.695 133.315 27.740 ;
        RECT 135.545 27.695 135.835 27.740 ;
        RECT 131.835 27.555 135.835 27.695 ;
        RECT 131.835 27.510 132.125 27.555 ;
        RECT 133.025 27.510 133.315 27.555 ;
        RECT 135.545 27.510 135.835 27.555 ;
        RECT 120.820 27.355 121.140 27.415 ;
        RECT 119.990 27.215 121.140 27.355 ;
        RECT 106.600 27.170 106.890 27.215 ;
        RECT 108.700 27.170 108.990 27.215 ;
        RECT 110.270 27.170 110.560 27.215 ;
        RECT 118.980 27.155 119.300 27.215 ;
        RECT 120.820 27.155 121.140 27.215 ;
        RECT 121.830 27.015 121.970 27.510 ;
        RECT 122.240 27.355 122.530 27.400 ;
        RECT 124.340 27.355 124.630 27.400 ;
        RECT 125.910 27.355 126.200 27.400 ;
        RECT 122.240 27.215 126.200 27.355 ;
        RECT 122.240 27.170 122.530 27.215 ;
        RECT 124.340 27.170 124.630 27.215 ;
        RECT 125.910 27.170 126.200 27.215 ;
        RECT 131.440 27.355 131.730 27.400 ;
        RECT 133.540 27.355 133.830 27.400 ;
        RECT 135.110 27.355 135.400 27.400 ;
        RECT 131.440 27.215 135.400 27.355 ;
        RECT 131.440 27.170 131.730 27.215 ;
        RECT 133.540 27.170 133.830 27.215 ;
        RECT 135.110 27.170 135.400 27.215 ;
        RECT 126.340 27.015 126.660 27.075 ;
        RECT 121.830 26.875 126.660 27.015 ;
        RECT 126.340 26.815 126.660 26.875 ;
        RECT 128.655 27.015 128.945 27.060 ;
        RECT 129.100 27.015 129.420 27.075 ;
        RECT 128.655 26.875 129.420 27.015 ;
        RECT 128.655 26.830 128.945 26.875 ;
        RECT 129.100 26.815 129.420 26.875 ;
        RECT 137.855 27.015 138.145 27.060 ;
        RECT 139.220 27.015 139.540 27.075 ;
        RECT 137.855 26.875 139.540 27.015 ;
        RECT 137.855 26.830 138.145 26.875 ;
        RECT 139.220 26.815 139.540 26.875 ;
        RECT 103.270 26.195 141.450 26.675 ;
        RECT 112.080 25.995 112.400 26.055 ;
        RECT 115.760 25.995 116.080 26.055 ;
        RECT 119.900 25.995 120.220 26.055 ;
        RECT 112.080 25.855 116.910 25.995 ;
        RECT 112.080 25.795 112.400 25.855 ;
        RECT 115.760 25.795 116.080 25.855 ;
        RECT 107.980 25.655 108.270 25.700 ;
        RECT 110.080 25.655 110.370 25.700 ;
        RECT 111.650 25.655 111.940 25.700 ;
        RECT 107.980 25.515 111.940 25.655 ;
        RECT 107.980 25.470 108.270 25.515 ;
        RECT 110.080 25.470 110.370 25.515 ;
        RECT 111.650 25.470 111.940 25.515 ;
        RECT 116.770 25.360 116.910 25.855 ;
        RECT 117.690 25.855 120.220 25.995 ;
        RECT 108.375 25.315 108.665 25.360 ;
        RECT 109.565 25.315 109.855 25.360 ;
        RECT 112.085 25.315 112.375 25.360 ;
        RECT 108.375 25.175 112.375 25.315 ;
        RECT 108.375 25.130 108.665 25.175 ;
        RECT 109.565 25.130 109.855 25.175 ;
        RECT 112.085 25.130 112.375 25.175 ;
        RECT 116.695 25.130 116.985 25.360 ;
        RECT 107.495 24.975 107.785 25.020 ;
        RECT 107.940 24.975 108.260 25.035 ;
        RECT 107.495 24.835 108.260 24.975 ;
        RECT 107.495 24.790 107.785 24.835 ;
        RECT 107.940 24.775 108.260 24.835 ;
        RECT 108.830 24.635 109.120 24.680 ;
        RECT 109.780 24.635 110.100 24.695 ;
        RECT 108.830 24.495 110.100 24.635 ;
        RECT 116.770 24.635 116.910 25.130 ;
        RECT 117.690 25.020 117.830 25.855 ;
        RECT 119.900 25.795 120.220 25.855 ;
        RECT 120.835 25.995 121.125 26.040 ;
        RECT 121.740 25.995 122.060 26.055 ;
        RECT 120.835 25.855 122.060 25.995 ;
        RECT 120.835 25.810 121.125 25.855 ;
        RECT 121.740 25.795 122.060 25.855 ;
        RECT 122.200 25.795 122.520 26.055 ;
        RECT 128.180 25.995 128.500 26.055 ;
        RECT 130.020 25.995 130.340 26.055 ;
        RECT 128.180 25.855 130.340 25.995 ;
        RECT 128.180 25.795 128.500 25.855 ;
        RECT 130.020 25.795 130.340 25.855 ;
        RECT 118.535 25.655 118.825 25.700 ;
        RECT 118.980 25.655 119.300 25.715 ;
        RECT 118.535 25.515 119.300 25.655 ;
        RECT 118.535 25.470 118.825 25.515 ;
        RECT 118.980 25.455 119.300 25.515 ;
        RECT 121.295 25.470 121.585 25.700 ;
        RECT 124.080 25.655 124.370 25.700 ;
        RECT 126.180 25.655 126.470 25.700 ;
        RECT 127.750 25.655 128.040 25.700 ;
        RECT 124.080 25.515 128.040 25.655 ;
        RECT 124.080 25.470 124.370 25.515 ;
        RECT 126.180 25.470 126.470 25.515 ;
        RECT 127.750 25.470 128.040 25.515 ;
        RECT 131.440 25.655 131.730 25.700 ;
        RECT 133.540 25.655 133.830 25.700 ;
        RECT 135.110 25.655 135.400 25.700 ;
        RECT 131.440 25.515 135.400 25.655 ;
        RECT 131.440 25.470 131.730 25.515 ;
        RECT 133.540 25.470 133.830 25.515 ;
        RECT 135.110 25.470 135.400 25.515 ;
        RECT 117.615 24.975 117.905 25.020 ;
        RECT 118.520 24.975 118.840 25.035 ;
        RECT 121.370 24.975 121.510 25.470 ;
        RECT 124.475 25.315 124.765 25.360 ;
        RECT 125.665 25.315 125.955 25.360 ;
        RECT 128.185 25.315 128.475 25.360 ;
        RECT 124.475 25.175 128.475 25.315 ;
        RECT 124.475 25.130 124.765 25.175 ;
        RECT 125.665 25.130 125.955 25.175 ;
        RECT 128.185 25.130 128.475 25.175 ;
        RECT 131.835 25.315 132.125 25.360 ;
        RECT 133.025 25.315 133.315 25.360 ;
        RECT 135.545 25.315 135.835 25.360 ;
        RECT 131.835 25.175 135.835 25.315 ;
        RECT 131.835 25.130 132.125 25.175 ;
        RECT 133.025 25.130 133.315 25.175 ;
        RECT 135.545 25.130 135.835 25.175 ;
        RECT 117.615 24.835 118.840 24.975 ;
        RECT 120.150 24.850 121.510 24.975 ;
        RECT 117.615 24.790 117.905 24.835 ;
        RECT 118.520 24.775 118.840 24.835 ;
        RECT 120.145 24.835 121.510 24.850 ;
        RECT 123.595 24.975 123.885 25.020 ;
        RECT 126.340 24.975 126.660 25.035 ;
        RECT 130.955 24.975 131.245 25.020 ;
        RECT 131.400 24.975 131.720 25.035 ;
        RECT 123.595 24.835 131.720 24.975 ;
        RECT 118.995 24.635 119.285 24.680 ;
        RECT 116.770 24.495 119.285 24.635 ;
        RECT 120.145 24.620 120.435 24.835 ;
        RECT 123.595 24.790 123.885 24.835 ;
        RECT 126.340 24.775 126.660 24.835 ;
        RECT 130.955 24.790 131.245 24.835 ;
        RECT 131.400 24.775 131.720 24.835 ;
        RECT 122.110 24.635 122.400 24.680 ;
        RECT 122.660 24.635 122.980 24.695 ;
        RECT 108.830 24.450 109.120 24.495 ;
        RECT 109.780 24.435 110.100 24.495 ;
        RECT 118.995 24.450 119.285 24.495 ;
        RECT 122.110 24.495 122.980 24.635 ;
        RECT 122.110 24.450 122.400 24.495 ;
        RECT 113.000 24.295 113.320 24.355 ;
        RECT 114.395 24.295 114.685 24.340 ;
        RECT 113.000 24.155 114.685 24.295 ;
        RECT 119.070 24.295 119.210 24.450 ;
        RECT 122.660 24.435 122.980 24.495 ;
        RECT 123.135 24.635 123.425 24.680 ;
        RECT 124.040 24.635 124.360 24.695 ;
        RECT 123.135 24.495 124.360 24.635 ;
        RECT 123.135 24.450 123.425 24.495 ;
        RECT 124.040 24.435 124.360 24.495 ;
        RECT 124.930 24.635 125.220 24.680 ;
        RECT 125.880 24.635 126.200 24.695 ;
        RECT 129.560 24.635 129.880 24.695 ;
        RECT 124.930 24.495 126.200 24.635 ;
        RECT 124.930 24.450 125.220 24.495 ;
        RECT 125.880 24.435 126.200 24.495 ;
        RECT 128.270 24.495 129.880 24.635 ;
        RECT 120.820 24.295 121.140 24.355 ;
        RECT 128.270 24.295 128.410 24.495 ;
        RECT 129.560 24.435 129.880 24.495 ;
        RECT 132.290 24.635 132.580 24.680 ;
        RECT 136.000 24.635 136.320 24.695 ;
        RECT 132.290 24.495 136.320 24.635 ;
        RECT 132.290 24.450 132.580 24.495 ;
        RECT 136.000 24.435 136.320 24.495 ;
        RECT 119.070 24.155 128.410 24.295 ;
        RECT 128.640 24.295 128.960 24.355 ;
        RECT 130.495 24.295 130.785 24.340 ;
        RECT 135.540 24.295 135.860 24.355 ;
        RECT 128.640 24.155 135.860 24.295 ;
        RECT 113.000 24.095 113.320 24.155 ;
        RECT 114.395 24.110 114.685 24.155 ;
        RECT 120.820 24.095 121.140 24.155 ;
        RECT 128.640 24.095 128.960 24.155 ;
        RECT 130.495 24.110 130.785 24.155 ;
        RECT 135.540 24.095 135.860 24.155 ;
        RECT 137.840 24.095 138.160 24.355 ;
        RECT 103.270 23.475 141.450 23.955 ;
        RECT 109.780 23.075 110.100 23.335 ;
        RECT 118.520 23.075 118.840 23.335 ;
        RECT 125.420 23.275 125.740 23.335 ;
        RECT 130.495 23.275 130.785 23.320 ;
        RECT 125.420 23.135 130.785 23.275 ;
        RECT 125.420 23.075 125.740 23.135 ;
        RECT 130.495 23.090 130.785 23.135 ;
        RECT 130.955 23.275 131.245 23.320 ;
        RECT 131.860 23.275 132.180 23.335 ;
        RECT 134.160 23.275 134.480 23.335 ;
        RECT 130.955 23.135 134.480 23.275 ;
        RECT 130.955 23.090 131.245 23.135 ;
        RECT 105.640 22.935 105.960 22.995 ;
        RECT 116.220 22.935 116.540 22.995 ;
        RECT 126.355 22.935 126.645 22.980 ;
        RECT 128.640 22.935 128.960 22.995 ;
        RECT 105.640 22.795 112.310 22.935 ;
        RECT 105.640 22.735 105.960 22.795 ;
        RECT 112.170 22.640 112.310 22.795 ;
        RECT 113.090 22.795 117.830 22.935 ;
        RECT 113.090 22.655 113.230 22.795 ;
        RECT 116.220 22.735 116.540 22.795 ;
        RECT 110.715 22.595 111.005 22.640 ;
        RECT 110.715 22.455 111.620 22.595 ;
        RECT 110.715 22.410 111.005 22.455 ;
        RECT 111.480 21.575 111.620 22.455 ;
        RECT 112.095 22.410 112.385 22.640 ;
        RECT 112.170 22.255 112.310 22.410 ;
        RECT 113.000 22.395 113.320 22.655 ;
        RECT 114.395 22.595 114.685 22.640 ;
        RECT 115.760 22.595 116.080 22.655 ;
        RECT 117.690 22.640 117.830 22.795 ;
        RECT 126.355 22.795 128.960 22.935 ;
        RECT 126.355 22.750 126.645 22.795 ;
        RECT 128.640 22.735 128.960 22.795 ;
        RECT 114.395 22.455 116.080 22.595 ;
        RECT 114.395 22.410 114.685 22.455 ;
        RECT 115.760 22.395 116.080 22.455 ;
        RECT 117.615 22.410 117.905 22.640 ;
        RECT 122.660 22.595 122.980 22.655 ;
        RECT 126.800 22.595 127.120 22.655 ;
        RECT 122.660 22.455 127.120 22.595 ;
        RECT 122.660 22.395 122.980 22.455 ;
        RECT 126.800 22.395 127.120 22.455 ;
        RECT 127.260 22.595 127.580 22.655 ;
        RECT 130.020 22.595 130.340 22.655 ;
        RECT 127.260 22.455 130.340 22.595 ;
        RECT 127.260 22.395 127.580 22.455 ;
        RECT 130.020 22.395 130.340 22.455 ;
        RECT 113.475 22.255 113.765 22.300 ;
        RECT 112.170 22.115 113.765 22.255 ;
        RECT 113.475 22.070 113.765 22.115 ;
        RECT 115.315 22.255 115.605 22.300 ;
        RECT 116.695 22.255 116.985 22.300 ;
        RECT 115.315 22.115 116.985 22.255 ;
        RECT 126.890 22.255 127.030 22.395 ;
        RECT 129.100 22.255 129.420 22.315 ;
        RECT 126.890 22.115 129.420 22.255 ;
        RECT 115.315 22.070 115.605 22.115 ;
        RECT 116.695 22.070 116.985 22.115 ;
        RECT 112.540 21.915 112.860 21.975 ;
        RECT 115.390 21.915 115.530 22.070 ;
        RECT 129.100 22.055 129.420 22.115 ;
        RECT 112.540 21.775 115.530 21.915 ;
        RECT 125.880 21.915 126.200 21.975 ;
        RECT 127.260 21.915 127.580 21.975 ;
        RECT 125.880 21.775 127.580 21.915 ;
        RECT 112.540 21.715 112.860 21.775 ;
        RECT 125.880 21.715 126.200 21.775 ;
        RECT 127.260 21.715 127.580 21.775 ;
        RECT 128.195 21.730 128.485 21.960 ;
        RECT 130.570 21.915 130.710 23.090 ;
        RECT 131.860 23.075 132.180 23.135 ;
        RECT 134.160 23.075 134.480 23.135 ;
        RECT 135.080 23.275 135.400 23.335 ;
        RECT 135.555 23.275 135.845 23.320 ;
        RECT 135.080 23.135 135.845 23.275 ;
        RECT 135.080 23.075 135.400 23.135 ;
        RECT 135.555 23.090 135.845 23.135 ;
        RECT 132.335 22.935 132.625 22.980 ;
        RECT 139.220 22.935 139.540 22.995 ;
        RECT 132.335 22.795 139.540 22.935 ;
        RECT 132.335 22.750 132.625 22.795 ;
        RECT 130.940 22.595 131.260 22.655 ;
        RECT 133.330 22.640 133.470 22.795 ;
        RECT 139.220 22.735 139.540 22.795 ;
        RECT 131.415 22.595 131.705 22.640 ;
        RECT 130.940 22.455 131.705 22.595 ;
        RECT 130.940 22.395 131.260 22.455 ;
        RECT 131.415 22.410 131.705 22.455 ;
        RECT 133.255 22.410 133.545 22.640 ;
        RECT 131.490 22.255 131.630 22.410 ;
        RECT 137.840 22.395 138.160 22.655 ;
        RECT 133.715 22.255 134.005 22.300 ;
        RECT 131.490 22.115 134.005 22.255 ;
        RECT 133.715 22.070 134.005 22.115 ;
        RECT 134.160 22.055 134.480 22.315 ;
        RECT 134.635 22.070 134.925 22.300 ;
        RECT 134.710 21.915 134.850 22.070 ;
        RECT 136.000 22.055 136.320 22.315 ;
        RECT 137.395 22.255 137.685 22.300 ;
        RECT 136.550 22.115 137.685 22.255 ;
        RECT 130.570 21.775 134.850 21.915 ;
        RECT 118.980 21.575 119.300 21.635 ;
        RECT 111.480 21.435 119.300 21.575 ;
        RECT 118.980 21.375 119.300 21.435 ;
        RECT 124.960 21.575 125.280 21.635 ;
        RECT 128.270 21.575 128.410 21.730 ;
        RECT 124.960 21.435 128.410 21.575 ;
        RECT 129.575 21.575 129.865 21.620 ;
        RECT 132.780 21.575 133.100 21.635 ;
        RECT 136.550 21.575 136.690 22.115 ;
        RECT 137.395 22.070 137.685 22.115 ;
        RECT 129.575 21.435 136.690 21.575 ;
        RECT 124.960 21.375 125.280 21.435 ;
        RECT 129.575 21.390 129.865 21.435 ;
        RECT 132.780 21.375 133.100 21.435 ;
        RECT 103.270 20.755 141.450 21.235 ;
        RECT 138.315 20.215 138.605 20.260 ;
        RECT 142.900 20.215 143.220 20.275 ;
        RECT 138.315 20.075 143.220 20.215 ;
        RECT 138.315 20.030 138.605 20.075 ;
        RECT 142.900 20.015 143.220 20.075 ;
        RECT 105.180 19.535 105.500 19.595 ;
        RECT 105.655 19.535 105.945 19.580 ;
        RECT 105.180 19.395 105.945 19.535 ;
        RECT 105.180 19.335 105.500 19.395 ;
        RECT 105.655 19.350 105.945 19.395 ;
        RECT 106.100 19.535 106.420 19.595 ;
        RECT 107.495 19.535 107.785 19.580 ;
        RECT 106.100 19.395 107.785 19.535 ;
        RECT 106.100 19.335 106.420 19.395 ;
        RECT 107.495 19.350 107.785 19.395 ;
        RECT 112.095 19.535 112.385 19.580 ;
        RECT 112.540 19.535 112.860 19.595 ;
        RECT 112.095 19.395 112.860 19.535 ;
        RECT 112.095 19.350 112.385 19.395 ;
        RECT 112.540 19.335 112.860 19.395 ;
        RECT 116.220 19.535 116.540 19.595 ;
        RECT 117.615 19.535 117.905 19.580 ;
        RECT 116.220 19.395 117.905 19.535 ;
        RECT 116.220 19.335 116.540 19.395 ;
        RECT 117.615 19.350 117.905 19.395 ;
        RECT 121.295 19.535 121.585 19.580 ;
        RECT 124.960 19.535 125.280 19.595 ;
        RECT 121.295 19.395 125.280 19.535 ;
        RECT 121.295 19.350 121.585 19.395 ;
        RECT 124.960 19.335 125.280 19.395 ;
        RECT 125.880 19.335 126.200 19.595 ;
        RECT 126.800 19.535 127.120 19.595 ;
        RECT 130.495 19.535 130.785 19.580 ;
        RECT 126.800 19.395 130.785 19.535 ;
        RECT 126.800 19.335 127.120 19.395 ;
        RECT 130.495 19.350 130.785 19.395 ;
        RECT 135.095 19.535 135.385 19.580 ;
        RECT 135.540 19.535 135.860 19.595 ;
        RECT 135.095 19.395 135.860 19.535 ;
        RECT 135.095 19.350 135.385 19.395 ;
        RECT 135.540 19.335 135.860 19.395 ;
        RECT 137.395 19.535 137.685 19.580 ;
        RECT 138.300 19.535 138.620 19.595 ;
        RECT 137.395 19.395 138.620 19.535 ;
        RECT 137.395 19.350 137.685 19.395 ;
        RECT 138.300 19.335 138.620 19.395 ;
        RECT 139.220 19.535 139.540 19.595 ;
        RECT 139.695 19.535 139.985 19.580 ;
        RECT 139.220 19.395 139.985 19.535 ;
        RECT 139.220 19.335 139.540 19.395 ;
        RECT 139.695 19.350 139.985 19.395 ;
        RECT 101.500 18.855 101.820 18.915 ;
        RECT 104.735 18.855 105.025 18.900 ;
        RECT 101.500 18.715 105.025 18.855 ;
        RECT 101.500 18.655 101.820 18.715 ;
        RECT 104.735 18.670 105.025 18.715 ;
        RECT 106.100 18.855 106.420 18.915 ;
        RECT 106.575 18.855 106.865 18.900 ;
        RECT 106.100 18.715 106.865 18.855 ;
        RECT 106.100 18.655 106.420 18.715 ;
        RECT 106.575 18.670 106.865 18.715 ;
        RECT 110.700 18.855 111.020 18.915 ;
        RECT 111.175 18.855 111.465 18.900 ;
        RECT 110.700 18.715 111.465 18.855 ;
        RECT 110.700 18.655 111.020 18.715 ;
        RECT 111.175 18.670 111.465 18.715 ;
        RECT 115.300 18.855 115.620 18.915 ;
        RECT 116.695 18.855 116.985 18.900 ;
        RECT 115.300 18.715 116.985 18.855 ;
        RECT 115.300 18.655 115.620 18.715 ;
        RECT 116.695 18.670 116.985 18.715 ;
        RECT 119.440 18.855 119.760 18.915 ;
        RECT 120.375 18.855 120.665 18.900 ;
        RECT 119.440 18.715 120.665 18.855 ;
        RECT 119.440 18.655 119.760 18.715 ;
        RECT 120.375 18.670 120.665 18.715 ;
        RECT 124.500 18.855 124.820 18.915 ;
        RECT 124.975 18.855 125.265 18.900 ;
        RECT 124.500 18.715 125.265 18.855 ;
        RECT 124.500 18.655 124.820 18.715 ;
        RECT 124.975 18.670 125.265 18.715 ;
        RECT 129.100 18.855 129.420 18.915 ;
        RECT 129.575 18.855 129.865 18.900 ;
        RECT 129.100 18.715 129.865 18.855 ;
        RECT 129.100 18.655 129.420 18.715 ;
        RECT 129.575 18.670 129.865 18.715 ;
        RECT 132.780 18.855 133.100 18.915 ;
        RECT 134.175 18.855 134.465 18.900 ;
        RECT 132.780 18.715 134.465 18.855 ;
        RECT 132.780 18.655 133.100 18.715 ;
        RECT 134.175 18.670 134.465 18.715 ;
        RECT 138.760 18.655 139.080 18.915 ;
        RECT 103.270 18.035 141.450 18.515 ;
        RECT 96.780 12.345 115.750 12.865 ;
        RECT 93.455 11.150 134.165 11.700 ;
        RECT 59.420 8.060 133.490 9.060 ;
        RECT 36.590 5.060 113.990 6.165 ;
        RECT 112.885 4.085 113.990 5.060 ;
        RECT 132.490 4.745 133.490 8.060 ;
        RECT 150.175 5.430 151.785 103.510 ;
        RECT 93.705 3.490 94.895 3.515 ;
        RECT 34.370 2.410 94.895 3.490 ;
        RECT 112.885 2.890 114.280 4.085 ;
        RECT 132.345 3.765 133.540 4.745 ;
        RECT 150.175 4.375 153.055 5.430 ;
        RECT 150.185 3.840 153.055 4.375 ;
        RECT 112.965 2.830 114.280 2.890 ;
        RECT 132.315 2.570 133.570 3.765 ;
        RECT 93.705 2.385 94.895 2.410 ;
      LAYER met2 ;
        RECT 127.070 223.020 128.050 224.290 ;
        RECT 129.770 223.520 130.590 224.220 ;
        RECT 51.970 132.845 52.850 209.350 ;
        RECT 54.610 133.180 55.610 211.660 ;
        RECT 127.070 211.630 128.070 223.020 ;
        RECT 127.040 210.630 128.100 211.630 ;
        RECT 129.740 208.410 130.620 223.520 ;
        RECT 132.610 223.110 133.275 224.215 ;
        RECT 135.385 223.215 136.020 224.410 ;
        RECT 138.175 223.245 138.745 224.375 ;
        RECT 89.610 174.380 133.305 175.045 ;
        RECT 135.355 172.535 136.050 172.550 ;
        RECT 90.895 171.925 136.050 172.535 ;
        RECT 135.355 171.915 136.050 171.925 ;
        RECT 92.220 169.760 138.795 170.425 ;
        RECT 90.015 165.530 90.345 165.560 ;
        RECT 90.940 165.530 91.270 165.545 ;
        RECT 90.015 165.200 91.270 165.530 ;
        RECT 91.440 165.245 91.770 165.555 ;
        RECT 90.015 165.170 90.345 165.200 ;
        RECT 87.900 162.715 89.460 162.815 ;
        RECT 87.870 161.675 89.490 162.715 ;
        RECT 87.900 161.570 89.460 161.675 ;
        RECT 57.725 155.540 58.395 155.555 ;
        RECT 57.715 154.620 58.545 155.540 ;
        RECT 54.610 130.545 55.610 130.570 ;
        RECT 51.970 130.365 52.850 130.390 ;
        RECT 51.950 129.535 52.870 130.365 ;
        RECT 54.590 129.595 55.630 130.545 ;
        RECT 39.430 123.425 40.430 124.485 ;
        RECT 37.220 86.650 38.220 122.515 ;
        RECT 39.435 87.965 40.430 123.425 ;
        RECT 51.970 122.515 52.855 129.535 ;
        RECT 54.610 123.425 55.610 129.595 ;
        RECT 51.950 121.455 52.950 122.515 ;
        RECT 57.725 117.810 58.395 154.620 ;
        RECT 62.995 152.790 63.375 153.230 ;
        RECT 67.165 152.550 71.710 152.560 ;
        RECT 61.875 152.360 66.420 152.370 ;
        RECT 61.855 152.040 66.420 152.360 ;
        RECT 67.145 152.230 71.710 152.550 ;
        RECT 67.145 152.040 67.755 152.230 ;
        RECT 61.855 151.850 62.465 152.040 ;
        RECT 61.285 151.300 62.485 151.850 ;
        RECT 61.295 151.150 62.485 151.300 ;
        RECT 61.305 147.410 61.635 151.150 ;
        RECT 61.795 149.770 62.605 150.700 ;
        RECT 62.835 149.860 63.525 150.590 ;
        RECT 61.835 149.760 62.575 149.770 ;
        RECT 65.225 148.670 65.685 150.530 ;
        RECT 66.090 148.670 66.420 152.040 ;
        RECT 66.575 151.490 67.775 152.040 ;
        RECT 66.585 151.340 67.775 151.490 ;
        RECT 61.885 147.410 62.365 148.390 ;
        RECT 61.305 141.630 62.365 147.410 ;
        RECT 65.225 144.160 66.420 148.670 ;
        RECT 65.225 141.660 65.685 144.160 ;
        RECT 61.305 138.670 61.635 141.630 ;
        RECT 61.885 140.970 62.365 141.630 ;
        RECT 61.865 138.670 62.345 139.180 ;
        RECT 61.305 132.890 62.345 138.670 ;
        RECT 61.305 132.170 61.635 132.890 ;
        RECT 61.865 131.760 62.345 132.890 ;
        RECT 65.305 138.310 65.765 139.150 ;
        RECT 66.090 138.310 66.420 144.160 ;
        RECT 65.305 133.800 66.420 138.310 ;
        RECT 65.305 130.280 65.765 133.800 ;
        RECT 66.090 133.785 66.420 133.800 ;
        RECT 66.595 147.600 66.925 151.340 ;
        RECT 68.075 151.280 68.945 152.050 ;
        RECT 67.075 150.870 67.805 150.910 ;
        RECT 67.075 149.970 67.875 150.870 ;
        RECT 68.135 150.070 68.795 150.750 ;
        RECT 67.075 149.940 67.805 149.970 ;
        RECT 70.515 148.860 70.975 150.720 ;
        RECT 71.380 148.860 71.710 152.230 ;
        RECT 73.515 150.810 74.395 155.565 ;
        RECT 90.940 154.580 91.270 165.200 ;
        RECT 91.410 164.915 91.800 165.245 ;
        RECT 91.950 163.390 92.280 166.050 ;
        RECT 93.125 164.880 99.345 165.310 ;
        RECT 99.835 164.890 100.185 165.370 ;
        RECT 93.050 164.080 93.310 164.400 ;
        RECT 96.745 164.300 96.925 164.520 ;
        RECT 91.635 162.235 92.015 162.260 ;
        RECT 91.615 161.905 92.035 162.235 ;
        RECT 90.865 153.735 91.345 154.580 ;
        RECT 91.635 152.775 92.015 161.905 ;
        RECT 92.675 160.610 92.945 161.800 ;
        RECT 92.715 158.220 92.865 160.610 ;
        RECT 93.085 160.430 93.280 164.080 ;
        RECT 96.745 163.950 97.075 164.300 ;
        RECT 93.745 163.330 94.145 163.770 ;
        RECT 95.385 163.750 95.725 163.810 ;
        RECT 93.055 160.060 93.335 160.430 ;
        RECT 93.495 159.010 93.665 161.630 ;
        RECT 93.905 160.790 94.145 163.330 ;
        RECT 95.315 163.370 95.725 163.750 ;
        RECT 96.775 163.390 97.075 163.950 ;
        RECT 93.825 160.350 94.145 160.790 ;
        RECT 94.795 162.170 95.105 162.620 ;
        RECT 92.660 157.900 92.920 158.220 ;
        RECT 92.715 156.225 92.865 157.900 ;
        RECT 93.055 156.730 94.625 157.160 ;
        RECT 94.795 156.710 95.095 162.170 ;
        RECT 95.315 161.330 95.565 163.370 ;
        RECT 96.105 161.720 96.365 162.040 ;
        RECT 96.805 161.910 97.055 163.390 ;
        RECT 97.215 162.180 99.655 162.610 ;
        RECT 95.310 161.010 95.570 161.330 ;
        RECT 95.735 158.460 96.015 159.260 ;
        RECT 95.775 156.575 95.925 158.460 ;
        RECT 96.170 158.300 96.320 161.720 ;
        RECT 96.765 161.530 97.085 161.910 ;
        RECT 97.525 161.400 97.785 161.720 ;
        RECT 98.465 161.550 98.725 161.870 ;
        RECT 97.570 160.345 97.740 161.400 ;
        RECT 98.005 161.080 98.265 161.400 ;
        RECT 98.030 160.710 98.240 161.080 ;
        RECT 97.975 160.450 98.295 160.710 ;
        RECT 97.525 160.025 97.785 160.345 ;
        RECT 96.605 159.440 98.235 159.870 ;
        RECT 97.105 158.460 97.365 159.250 ;
        RECT 96.115 157.980 96.375 158.300 ;
        RECT 92.685 152.815 92.895 156.225 ;
        RECT 95.735 153.340 95.970 156.575 ;
        RECT 96.170 156.530 96.320 157.980 ;
        RECT 97.165 156.540 97.315 158.460 ;
        RECT 98.485 158.320 98.705 161.550 ;
        RECT 99.865 159.460 100.165 164.890 ;
        RECT 101.745 164.830 102.095 165.330 ;
        RECT 101.175 164.525 101.495 164.695 ;
        RECT 101.125 164.385 101.545 164.525 ;
        RECT 100.705 163.815 101.620 164.385 ;
        RECT 100.395 162.170 101.565 162.600 ;
        RECT 101.255 160.950 101.595 161.930 ;
        RECT 98.955 158.440 99.245 159.150 ;
        RECT 99.915 158.840 100.175 159.160 ;
        RECT 101.255 158.840 101.515 160.950 ;
        RECT 101.795 160.240 102.095 164.830 ;
        RECT 102.635 162.540 102.925 162.590 ;
        RECT 101.755 159.400 102.155 160.240 ;
        RECT 98.485 157.920 98.815 158.320 ;
        RECT 98.510 156.540 98.680 157.920 ;
        RECT 96.145 153.755 96.350 156.530 ;
        RECT 97.130 154.190 97.350 156.540 ;
        RECT 98.475 154.805 98.720 156.540 ;
        RECT 99.015 156.470 99.165 158.440 ;
        RECT 99.940 158.300 100.150 158.840 ;
        RECT 99.915 157.980 100.175 158.300 ;
        RECT 99.965 156.600 100.130 157.980 ;
        RECT 100.405 157.420 100.715 158.280 ;
        RECT 98.970 155.260 99.210 156.470 ;
        RECT 99.905 155.840 100.185 156.600 ;
        RECT 100.425 156.545 100.590 157.420 ;
        RECT 100.825 156.730 102.395 157.160 ;
        RECT 102.625 156.730 102.925 162.540 ;
        RECT 100.340 156.210 102.930 156.545 ;
        RECT 100.425 156.190 100.590 156.210 ;
        RECT 99.905 155.560 102.335 155.840 ;
        RECT 98.970 155.020 101.715 155.260 ;
        RECT 98.475 154.560 101.195 154.805 ;
        RECT 97.130 153.970 100.535 154.190 ;
        RECT 96.145 153.550 99.915 153.755 ;
        RECT 98.955 153.340 99.205 153.350 ;
        RECT 95.735 153.105 99.205 153.340 ;
        RECT 92.685 152.605 98.590 152.815 ;
        RECT 95.665 152.410 96.215 152.420 ;
        RECT 95.515 152.400 96.215 152.410 ;
        RECT 76.535 152.070 96.215 152.400 ;
        RECT 77.255 151.840 83.035 152.070 ;
        RECT 76.125 151.360 83.545 151.840 ;
        RECT 85.995 151.820 91.775 152.070 ;
        RECT 85.335 151.340 92.755 151.820 ;
        RECT 94.375 151.450 94.925 151.920 ;
        RECT 95.515 151.850 96.215 152.070 ;
        RECT 95.515 151.830 96.725 151.850 ;
        RECT 95.515 151.240 96.735 151.830 ;
        RECT 95.515 151.220 96.215 151.240 ;
        RECT 73.395 150.030 74.395 150.810 ;
        RECT 94.255 150.220 94.805 150.780 ;
        RECT 73.515 149.730 74.395 150.030 ;
        RECT 73.175 149.610 74.395 149.730 ;
        RECT 67.175 147.600 67.655 148.580 ;
        RECT 66.595 141.820 67.655 147.600 ;
        RECT 70.515 144.350 71.710 148.860 ;
        RECT 73.145 147.920 74.395 149.610 ;
        RECT 74.645 147.940 83.515 148.400 ;
        RECT 86.025 148.020 94.895 148.480 ;
        RECT 73.175 147.790 74.395 147.920 ;
        RECT 73.615 145.480 74.395 147.790 ;
        RECT 78.165 147.615 82.675 147.940 ;
        RECT 88.525 147.615 93.035 148.020 ;
        RECT 96.405 147.615 96.735 151.240 ;
        RECT 96.955 150.495 97.505 150.740 ;
        RECT 98.380 150.495 98.590 152.605 ;
        RECT 98.955 152.620 99.205 153.105 ;
        RECT 99.710 152.620 99.915 153.550 ;
        RECT 100.315 152.620 100.535 153.970 ;
        RECT 98.955 152.265 99.220 152.620 ;
        RECT 96.955 150.285 98.590 150.495 ;
        RECT 96.955 150.180 97.505 150.285 ;
        RECT 78.150 147.285 96.735 147.615 ;
        RECT 96.935 147.310 97.485 148.010 ;
        RECT 95.675 147.060 96.225 147.070 ;
        RECT 95.525 147.050 96.225 147.060 ;
        RECT 76.545 146.720 96.225 147.050 ;
        RECT 77.265 146.490 83.045 146.720 ;
        RECT 76.135 146.010 83.555 146.490 ;
        RECT 86.005 146.470 91.785 146.720 ;
        RECT 85.345 145.990 92.765 146.470 ;
        RECT 94.355 146.070 94.905 146.540 ;
        RECT 95.525 146.500 96.225 146.720 ;
        RECT 95.525 146.480 96.735 146.500 ;
        RECT 95.525 145.890 96.745 146.480 ;
        RECT 95.525 145.870 96.225 145.890 ;
        RECT 73.435 144.700 74.395 145.480 ;
        RECT 94.355 144.920 94.945 145.390 ;
        RECT 73.615 144.390 74.395 144.700 ;
        RECT 70.515 141.850 70.975 144.350 ;
        RECT 66.595 138.860 66.925 141.820 ;
        RECT 67.175 141.160 67.655 141.820 ;
        RECT 67.155 138.860 67.635 139.370 ;
        RECT 66.595 133.080 67.635 138.860 ;
        RECT 66.595 132.360 66.925 133.080 ;
        RECT 67.155 131.950 67.635 133.080 ;
        RECT 70.595 138.500 71.055 139.340 ;
        RECT 71.380 138.500 71.710 144.350 ;
        RECT 73.175 144.220 74.395 144.390 ;
        RECT 73.165 142.530 74.395 144.220 ;
        RECT 74.655 142.590 83.525 143.050 ;
        RECT 86.035 142.670 94.905 143.130 ;
        RECT 73.175 142.450 74.395 142.530 ;
        RECT 73.615 140.140 74.395 142.450 ;
        RECT 78.175 142.265 82.685 142.590 ;
        RECT 88.535 142.265 93.045 142.670 ;
        RECT 96.415 142.265 96.745 145.890 ;
        RECT 96.945 144.910 97.535 145.380 ;
        RECT 78.160 141.935 96.745 142.265 ;
        RECT 95.645 141.710 96.195 141.720 ;
        RECT 95.495 141.700 96.195 141.710 ;
        RECT 76.515 141.370 96.195 141.700 ;
        RECT 77.235 141.140 83.015 141.370 ;
        RECT 76.105 140.660 83.525 141.140 ;
        RECT 85.975 141.120 91.755 141.370 ;
        RECT 85.315 140.640 92.735 141.120 ;
        RECT 94.325 140.710 94.875 141.180 ;
        RECT 95.495 141.150 96.195 141.370 ;
        RECT 95.495 141.130 96.705 141.150 ;
        RECT 95.495 140.540 96.715 141.130 ;
        RECT 95.495 140.520 96.195 140.540 ;
        RECT 73.405 139.360 74.395 140.140 ;
        RECT 94.315 139.550 94.905 140.070 ;
        RECT 73.615 139.020 74.395 139.360 ;
        RECT 73.155 138.870 74.395 139.020 ;
        RECT 70.595 133.990 71.710 138.500 ;
        RECT 73.125 137.180 74.395 138.870 ;
        RECT 74.625 137.240 83.495 137.700 ;
        RECT 86.005 137.320 94.875 137.780 ;
        RECT 73.155 137.080 74.395 137.180 ;
        RECT 73.615 134.890 74.395 137.080 ;
        RECT 78.145 136.915 82.655 137.240 ;
        RECT 88.505 136.915 93.015 137.320 ;
        RECT 96.385 136.915 96.715 140.540 ;
        RECT 96.935 139.550 97.525 140.070 ;
        RECT 78.130 136.585 96.715 136.915 ;
        RECT 95.685 136.430 96.235 136.440 ;
        RECT 95.535 136.420 96.235 136.430 ;
        RECT 76.555 136.090 96.235 136.420 ;
        RECT 77.275 135.860 83.055 136.090 ;
        RECT 76.145 135.380 83.565 135.860 ;
        RECT 86.015 135.840 91.795 136.090 ;
        RECT 95.535 135.870 96.235 136.090 ;
        RECT 95.535 135.850 96.745 135.870 ;
        RECT 85.355 135.360 92.775 135.840 ;
        RECT 94.355 135.350 94.905 135.820 ;
        RECT 95.535 135.260 96.755 135.850 ;
        RECT 95.535 135.240 96.235 135.260 ;
        RECT 73.395 134.880 74.395 134.890 ;
        RECT 70.595 130.470 71.055 133.990 ;
        RECT 71.380 133.975 71.710 133.990 ;
        RECT 73.155 133.970 74.395 134.880 ;
        RECT 94.115 134.190 95.045 134.880 ;
        RECT 73.155 133.960 74.365 133.970 ;
        RECT 62.845 128.690 63.595 129.795 ;
        RECT 68.180 128.690 68.930 129.985 ;
        RECT 73.155 129.390 74.085 133.960 ;
        RECT 74.665 131.960 83.535 132.420 ;
        RECT 86.045 132.040 94.915 132.500 ;
        RECT 78.185 131.635 82.695 131.960 ;
        RECT 88.545 131.635 93.055 132.040 ;
        RECT 96.425 131.635 96.755 135.260 ;
        RECT 97.015 134.360 97.665 134.830 ;
        RECT 78.170 131.305 96.755 131.635 ;
        RECT 95.675 130.840 96.225 130.850 ;
        RECT 95.525 130.830 96.225 130.840 ;
        RECT 76.545 130.500 96.225 130.830 ;
        RECT 77.265 130.270 83.045 130.500 ;
        RECT 76.135 129.790 83.555 130.270 ;
        RECT 86.005 130.250 91.785 130.500 ;
        RECT 85.345 129.770 92.765 130.250 ;
        RECT 94.385 129.880 94.935 130.350 ;
        RECT 95.525 130.280 96.225 130.500 ;
        RECT 95.525 130.260 96.735 130.280 ;
        RECT 95.525 129.670 96.745 130.260 ;
        RECT 95.525 129.650 96.225 129.670 ;
        RECT 73.155 128.690 74.405 129.390 ;
        RECT 62.845 127.940 74.405 128.690 ;
        RECT 94.265 128.650 94.815 129.210 ;
        RECT 71.180 127.545 71.930 127.575 ;
        RECT 60.290 126.795 71.930 127.545 ;
        RECT 71.180 126.765 71.930 126.795 ;
        RECT 66.840 126.300 67.840 126.330 ;
        RECT 69.400 126.300 70.400 126.345 ;
        RECT 73.155 126.340 74.405 127.940 ;
        RECT 74.655 126.370 83.525 126.830 ;
        RECT 86.035 126.450 94.905 126.910 ;
        RECT 66.840 125.300 70.400 126.300 ;
        RECT 73.185 126.220 74.405 126.340 ;
        RECT 66.840 125.270 67.840 125.300 ;
        RECT 69.400 125.255 70.400 125.300 ;
        RECT 73.625 123.910 74.405 126.220 ;
        RECT 78.175 126.045 82.685 126.370 ;
        RECT 88.535 126.045 93.045 126.450 ;
        RECT 96.415 126.045 96.745 129.670 ;
        RECT 96.965 128.935 97.515 129.170 ;
        RECT 98.380 128.935 98.590 150.285 ;
        RECT 98.985 149.360 99.220 152.265 ;
        RECT 99.700 152.030 99.915 152.620 ;
        RECT 100.295 152.240 100.535 152.620 ;
        RECT 98.975 149.040 99.235 149.360 ;
        RECT 96.965 128.725 98.590 128.935 ;
        RECT 96.965 128.610 97.515 128.725 ;
        RECT 96.995 127.850 97.755 128.010 ;
        RECT 98.985 127.850 99.220 149.040 ;
        RECT 99.700 145.290 99.905 152.030 ;
        RECT 99.675 144.970 99.935 145.290 ;
        RECT 96.995 127.615 99.220 127.850 ;
        RECT 96.995 127.310 97.755 127.615 ;
        RECT 78.160 125.715 96.745 126.045 ;
        RECT 96.945 125.740 97.495 126.440 ;
        RECT 95.685 125.490 96.235 125.500 ;
        RECT 95.535 125.480 96.235 125.490 ;
        RECT 76.555 125.150 96.235 125.480 ;
        RECT 77.275 124.920 83.055 125.150 ;
        RECT 76.145 124.440 83.565 124.920 ;
        RECT 86.015 124.900 91.795 125.150 ;
        RECT 85.355 124.420 92.775 124.900 ;
        RECT 94.365 124.500 94.915 124.970 ;
        RECT 95.535 124.930 96.235 125.150 ;
        RECT 95.535 124.910 96.745 124.930 ;
        RECT 95.535 124.320 96.755 124.910 ;
        RECT 95.535 124.300 96.235 124.320 ;
        RECT 59.040 123.345 65.260 123.775 ;
        RECT 65.750 123.355 66.100 123.835 ;
        RECT 58.965 122.545 59.225 122.865 ;
        RECT 62.660 122.765 62.840 122.985 ;
        RECT 58.590 119.075 58.860 120.265 ;
        RECT 43.975 112.805 44.405 112.825 ;
        RECT 43.950 110.345 44.430 112.805 ;
        RECT 57.820 112.280 58.300 117.810 ;
        RECT 58.630 116.685 58.780 119.075 ;
        RECT 59.000 118.895 59.195 122.545 ;
        RECT 62.660 122.415 62.990 122.765 ;
        RECT 59.660 121.795 60.060 122.235 ;
        RECT 61.300 122.215 61.640 122.275 ;
        RECT 58.970 118.525 59.250 118.895 ;
        RECT 59.410 117.475 59.580 120.095 ;
        RECT 59.820 119.255 60.060 121.795 ;
        RECT 61.230 121.835 61.640 122.215 ;
        RECT 62.690 121.855 62.990 122.415 ;
        RECT 59.740 118.815 60.060 119.255 ;
        RECT 60.710 120.635 61.020 121.085 ;
        RECT 58.575 116.365 58.835 116.685 ;
        RECT 58.630 112.200 58.780 116.365 ;
        RECT 58.970 115.195 60.540 115.625 ;
        RECT 60.710 115.175 61.010 120.635 ;
        RECT 61.230 119.795 61.480 121.835 ;
        RECT 62.020 120.185 62.280 120.505 ;
        RECT 62.720 120.375 62.970 121.855 ;
        RECT 63.130 120.645 65.570 121.075 ;
        RECT 61.225 119.475 61.485 119.795 ;
        RECT 61.650 116.925 61.930 117.725 ;
        RECT 61.690 112.570 61.840 116.925 ;
        RECT 62.085 116.765 62.235 120.185 ;
        RECT 62.680 119.995 63.000 120.375 ;
        RECT 63.440 119.865 63.700 120.185 ;
        RECT 64.380 120.015 64.640 120.335 ;
        RECT 63.485 118.810 63.655 119.865 ;
        RECT 63.920 119.545 64.180 119.865 ;
        RECT 63.945 119.175 64.155 119.545 ;
        RECT 63.890 118.915 64.210 119.175 ;
        RECT 63.440 118.490 63.700 118.810 ;
        RECT 62.520 117.905 64.150 118.335 ;
        RECT 63.020 116.925 63.280 117.715 ;
        RECT 62.030 116.445 62.290 116.765 ;
        RECT 62.085 114.815 62.235 116.445 ;
        RECT 63.080 114.860 63.230 116.925 ;
        RECT 64.400 116.785 64.620 120.015 ;
        RECT 65.780 117.925 66.080 123.355 ;
        RECT 67.660 123.295 68.010 123.795 ;
        RECT 66.310 120.635 67.480 121.065 ;
        RECT 67.170 119.415 67.510 120.395 ;
        RECT 64.870 116.905 65.160 117.615 ;
        RECT 65.830 117.305 66.090 117.625 ;
        RECT 67.170 117.305 67.430 119.415 ;
        RECT 67.710 118.705 68.010 123.295 ;
        RECT 73.445 123.130 74.405 123.910 ;
        RECT 94.365 123.350 94.955 123.820 ;
        RECT 73.625 122.820 74.405 123.130 ;
        RECT 73.185 122.650 74.405 122.820 ;
        RECT 68.550 121.005 68.840 121.055 ;
        RECT 67.670 117.865 68.070 118.705 ;
        RECT 64.400 116.385 64.730 116.785 ;
        RECT 62.080 112.935 62.245 114.815 ;
        RECT 63.060 113.335 63.255 114.860 ;
        RECT 64.425 114.835 64.595 116.385 ;
        RECT 64.930 114.855 65.080 116.905 ;
        RECT 65.855 116.765 66.065 117.305 ;
        RECT 65.830 116.445 66.090 116.765 ;
        RECT 65.880 114.970 66.045 116.445 ;
        RECT 66.320 115.885 66.630 116.745 ;
        RECT 66.340 114.975 66.505 115.885 ;
        RECT 66.740 115.195 68.310 115.625 ;
        RECT 68.540 115.195 68.840 121.005 ;
        RECT 73.175 120.960 74.405 122.650 ;
        RECT 74.665 121.020 83.535 121.480 ;
        RECT 86.045 121.100 94.915 121.560 ;
        RECT 73.185 120.880 74.405 120.960 ;
        RECT 73.625 118.570 74.405 120.880 ;
        RECT 78.185 120.695 82.695 121.020 ;
        RECT 88.545 120.695 93.055 121.100 ;
        RECT 96.425 120.695 96.755 124.320 ;
        RECT 96.955 123.665 97.545 123.810 ;
        RECT 99.700 123.665 99.905 144.970 ;
        RECT 100.295 144.070 100.515 152.240 ;
        RECT 100.275 143.750 100.535 144.070 ;
        RECT 96.955 123.460 99.905 123.665 ;
        RECT 96.955 123.340 97.545 123.460 ;
        RECT 96.995 123.290 97.200 123.340 ;
        RECT 96.965 122.450 97.725 122.710 ;
        RECT 100.295 122.450 100.515 143.750 ;
        RECT 100.950 140.050 101.195 154.560 ;
        RECT 100.945 139.730 101.205 140.050 ;
        RECT 96.965 122.230 100.515 122.450 ;
        RECT 96.965 122.010 97.725 122.230 ;
        RECT 78.170 120.365 96.755 120.695 ;
        RECT 95.655 120.140 96.205 120.150 ;
        RECT 95.505 120.130 96.205 120.140 ;
        RECT 76.525 119.800 96.205 120.130 ;
        RECT 77.245 119.570 83.025 119.800 ;
        RECT 76.115 119.090 83.535 119.570 ;
        RECT 85.985 119.550 91.765 119.800 ;
        RECT 85.325 119.070 92.745 119.550 ;
        RECT 94.335 119.140 94.885 119.610 ;
        RECT 95.505 119.580 96.205 119.800 ;
        RECT 95.505 119.560 96.715 119.580 ;
        RECT 95.505 118.970 96.725 119.560 ;
        RECT 95.505 118.950 96.205 118.970 ;
        RECT 73.415 117.790 74.405 118.570 ;
        RECT 94.325 117.980 94.915 118.500 ;
        RECT 73.625 117.450 74.405 117.790 ;
        RECT 73.165 117.300 74.405 117.450 ;
        RECT 73.135 115.610 74.405 117.300 ;
        RECT 74.635 115.670 83.505 116.130 ;
        RECT 86.015 115.750 94.885 116.210 ;
        RECT 73.165 115.510 74.405 115.610 ;
        RECT 64.410 113.730 64.615 114.835 ;
        RECT 64.905 114.115 65.105 114.855 ;
        RECT 65.865 114.495 66.065 114.970 ;
        RECT 66.310 114.740 70.635 114.975 ;
        RECT 66.340 114.655 66.505 114.740 ;
        RECT 65.865 114.295 70.250 114.495 ;
        RECT 64.905 113.915 69.880 114.115 ;
        RECT 64.410 113.525 69.470 113.730 ;
        RECT 63.060 113.140 69.065 113.335 ;
        RECT 62.070 112.745 68.655 112.935 ;
        RECT 61.670 112.380 68.265 112.570 ;
        RECT 58.620 112.025 67.915 112.200 ;
        RECT 65.430 111.795 65.980 111.805 ;
        RECT 65.280 111.785 65.980 111.795 ;
        RECT 46.300 111.455 65.980 111.785 ;
        RECT 47.020 111.225 52.800 111.455 ;
        RECT 45.890 110.745 53.310 111.225 ;
        RECT 55.760 111.205 61.540 111.455 ;
        RECT 55.100 110.725 62.520 111.205 ;
        RECT 64.140 110.835 64.690 111.305 ;
        RECT 65.280 111.235 65.980 111.455 ;
        RECT 65.280 111.215 66.490 111.235 ;
        RECT 65.280 110.625 66.500 111.215 ;
        RECT 65.280 110.605 65.980 110.625 ;
        RECT 43.380 110.195 44.430 110.345 ;
        RECT 43.160 109.415 44.430 110.195 ;
        RECT 64.020 109.605 64.570 110.165 ;
        RECT 43.380 109.345 44.430 109.415 ;
        RECT 43.380 109.115 44.160 109.345 ;
        RECT 42.940 108.995 44.160 109.115 ;
        RECT 42.910 107.305 44.160 108.995 ;
        RECT 44.410 107.325 53.280 107.785 ;
        RECT 55.790 107.405 64.660 107.865 ;
        RECT 42.940 107.175 44.160 107.305 ;
        RECT 43.380 104.865 44.160 107.175 ;
        RECT 47.930 107.000 52.440 107.325 ;
        RECT 58.290 107.000 62.800 107.405 ;
        RECT 66.170 107.000 66.500 110.625 ;
        RECT 66.720 109.885 67.270 110.125 ;
        RECT 67.740 109.885 67.915 112.025 ;
        RECT 66.720 109.710 67.915 109.885 ;
        RECT 66.720 109.565 67.270 109.710 ;
        RECT 66.680 108.770 67.220 108.925 ;
        RECT 68.075 108.770 68.265 112.380 ;
        RECT 66.680 108.555 68.280 108.770 ;
        RECT 66.680 108.335 67.220 108.555 ;
        RECT 47.915 106.670 66.500 107.000 ;
        RECT 66.700 106.695 67.250 107.395 ;
        RECT 65.440 106.445 65.990 106.455 ;
        RECT 65.290 106.435 65.990 106.445 ;
        RECT 46.310 106.105 65.990 106.435 ;
        RECT 47.030 105.875 52.810 106.105 ;
        RECT 45.900 105.395 53.320 105.875 ;
        RECT 55.770 105.855 61.550 106.105 ;
        RECT 55.110 105.375 62.530 105.855 ;
        RECT 64.120 105.455 64.670 105.925 ;
        RECT 65.290 105.885 65.990 106.105 ;
        RECT 65.290 105.865 66.500 105.885 ;
        RECT 65.290 105.275 66.510 105.865 ;
        RECT 66.750 105.295 67.450 106.055 ;
        RECT 65.290 105.255 65.990 105.275 ;
        RECT 43.200 104.085 44.160 104.865 ;
        RECT 64.120 104.305 64.710 104.775 ;
        RECT 43.380 103.775 44.160 104.085 ;
        RECT 42.940 103.605 44.160 103.775 ;
        RECT 42.930 101.915 44.160 103.605 ;
        RECT 44.420 101.975 53.290 102.435 ;
        RECT 55.800 102.055 64.670 102.515 ;
        RECT 42.940 101.835 44.160 101.915 ;
        RECT 43.380 99.525 44.160 101.835 ;
        RECT 47.940 101.650 52.450 101.975 ;
        RECT 58.300 101.650 62.810 102.055 ;
        RECT 66.180 101.650 66.510 105.275 ;
        RECT 66.710 104.640 67.300 104.765 ;
        RECT 68.465 104.640 68.655 112.745 ;
        RECT 66.710 104.450 68.655 104.640 ;
        RECT 66.710 104.295 67.300 104.450 ;
        RECT 66.815 104.290 67.005 104.295 ;
        RECT 66.720 103.385 67.560 103.625 ;
        RECT 68.870 103.385 69.065 113.140 ;
        RECT 66.720 103.190 69.065 103.385 ;
        RECT 66.720 102.915 67.560 103.190 ;
        RECT 47.925 101.320 66.510 101.650 ;
        RECT 65.410 101.095 65.960 101.105 ;
        RECT 65.260 101.085 65.960 101.095 ;
        RECT 46.280 100.755 65.960 101.085 ;
        RECT 47.000 100.525 52.780 100.755 ;
        RECT 45.870 100.045 53.290 100.525 ;
        RECT 55.740 100.505 61.520 100.755 ;
        RECT 55.080 100.025 62.500 100.505 ;
        RECT 64.090 100.095 64.640 100.565 ;
        RECT 65.260 100.535 65.960 100.755 ;
        RECT 65.260 100.515 66.470 100.535 ;
        RECT 65.260 99.925 66.480 100.515 ;
        RECT 65.260 99.905 65.960 99.925 ;
        RECT 43.170 98.745 44.160 99.525 ;
        RECT 64.080 98.935 64.670 99.455 ;
        RECT 43.380 98.405 44.160 98.745 ;
        RECT 42.920 98.255 44.160 98.405 ;
        RECT 42.890 96.565 44.160 98.255 ;
        RECT 44.390 96.625 53.260 97.085 ;
        RECT 55.770 96.705 64.640 97.165 ;
        RECT 42.920 96.465 44.160 96.565 ;
        RECT 43.380 94.275 44.160 96.465 ;
        RECT 47.910 96.300 52.420 96.625 ;
        RECT 58.270 96.300 62.780 96.705 ;
        RECT 66.150 96.300 66.480 99.925 ;
        RECT 66.700 99.400 67.290 99.455 ;
        RECT 69.265 99.400 69.470 113.525 ;
        RECT 66.700 99.195 69.470 99.400 ;
        RECT 66.700 98.935 67.290 99.195 ;
        RECT 66.800 98.245 67.430 98.475 ;
        RECT 69.680 98.245 69.880 113.915 ;
        RECT 66.750 98.045 69.880 98.245 ;
        RECT 66.800 97.705 67.430 98.045 ;
        RECT 47.895 95.970 66.480 96.300 ;
        RECT 65.450 95.815 66.000 95.825 ;
        RECT 65.300 95.805 66.000 95.815 ;
        RECT 46.320 95.475 66.000 95.805 ;
        RECT 47.040 95.245 52.820 95.475 ;
        RECT 45.910 94.765 53.330 95.245 ;
        RECT 55.780 95.225 61.560 95.475 ;
        RECT 65.300 95.255 66.000 95.475 ;
        RECT 65.300 95.235 66.510 95.255 ;
        RECT 55.120 94.745 62.540 95.225 ;
        RECT 64.120 94.735 64.670 95.205 ;
        RECT 65.300 94.645 66.520 95.235 ;
        RECT 65.300 94.625 66.000 94.645 ;
        RECT 43.160 93.505 44.160 94.275 ;
        RECT 63.880 93.575 64.810 94.265 ;
        RECT 42.940 93.355 44.160 93.505 ;
        RECT 42.940 93.345 44.130 93.355 ;
        RECT 42.940 93.075 43.390 93.345 ;
        RECT 42.930 91.385 43.390 93.075 ;
        RECT 42.940 91.185 43.390 91.385 ;
        RECT 44.430 91.345 53.300 91.805 ;
        RECT 55.810 91.425 64.680 91.885 ;
        RECT 47.950 91.020 52.460 91.345 ;
        RECT 58.310 91.020 62.820 91.425 ;
        RECT 66.190 91.020 66.520 94.645 ;
        RECT 66.780 94.185 67.430 94.215 ;
        RECT 70.050 94.185 70.250 114.295 ;
        RECT 66.780 93.985 70.250 94.185 ;
        RECT 66.780 93.745 67.430 93.985 ;
        RECT 66.750 93.055 67.520 93.245 ;
        RECT 70.400 93.055 70.635 114.740 ;
        RECT 73.625 113.320 74.405 115.510 ;
        RECT 78.155 115.345 82.665 115.670 ;
        RECT 88.515 115.345 93.025 115.750 ;
        RECT 96.395 115.345 96.725 118.970 ;
        RECT 96.945 118.445 97.535 118.500 ;
        RECT 100.950 118.445 101.195 139.730 ;
        RECT 101.475 138.890 101.715 155.020 ;
        RECT 101.465 138.570 101.725 138.890 ;
        RECT 96.945 118.200 101.195 118.445 ;
        RECT 96.945 117.980 97.535 118.200 ;
        RECT 96.965 117.390 97.725 117.500 ;
        RECT 101.475 117.390 101.715 138.570 ;
        RECT 96.935 117.150 101.715 117.390 ;
        RECT 96.935 117.000 97.725 117.150 ;
        RECT 96.965 116.800 97.725 117.000 ;
        RECT 78.140 115.015 96.725 115.345 ;
        RECT 95.695 114.860 96.245 114.870 ;
        RECT 95.545 114.850 96.245 114.860 ;
        RECT 76.565 114.520 96.245 114.850 ;
        RECT 77.285 114.290 83.065 114.520 ;
        RECT 76.155 113.810 83.575 114.290 ;
        RECT 86.025 114.270 91.805 114.520 ;
        RECT 95.545 114.300 96.245 114.520 ;
        RECT 95.545 114.280 96.755 114.300 ;
        RECT 85.365 113.790 92.785 114.270 ;
        RECT 94.365 113.780 94.915 114.250 ;
        RECT 95.545 113.690 96.765 114.280 ;
        RECT 95.545 113.670 96.245 113.690 ;
        RECT 73.405 112.550 74.405 113.320 ;
        RECT 94.125 112.620 95.055 113.310 ;
        RECT 73.185 112.400 74.405 112.550 ;
        RECT 73.185 112.390 74.375 112.400 ;
        RECT 73.185 112.120 73.635 112.390 ;
        RECT 71.565 111.565 72.515 111.585 ;
        RECT 70.950 110.565 72.540 111.565 ;
        RECT 71.565 110.545 72.515 110.565 ;
        RECT 73.175 110.430 73.635 112.120 ;
        RECT 73.185 110.230 73.635 110.430 ;
        RECT 74.675 110.390 83.545 110.850 ;
        RECT 86.055 110.470 94.925 110.930 ;
        RECT 78.195 110.065 82.705 110.390 ;
        RECT 88.555 110.065 93.065 110.470 ;
        RECT 96.435 110.065 96.765 113.690 ;
        RECT 97.025 113.240 97.675 113.260 ;
        RECT 102.055 113.240 102.335 155.560 ;
        RECT 96.945 112.960 102.335 113.240 ;
        RECT 97.025 112.790 97.675 112.960 ;
        RECT 97.035 112.150 97.795 112.340 ;
        RECT 102.595 112.150 102.930 156.210 ;
        RECT 103.395 153.615 104.285 153.625 ;
        RECT 104.915 153.615 105.865 153.645 ;
        RECT 103.335 152.665 105.865 153.615 ;
        RECT 103.395 152.645 104.285 152.665 ;
        RECT 104.915 152.635 105.865 152.665 ;
        RECT 111.470 151.240 117.830 154.460 ;
        RECT 105.560 146.905 106.780 148.625 ;
        RECT 105.565 145.935 106.720 146.905 ;
        RECT 104.010 124.715 105.200 126.965 ;
        RECT 104.010 123.750 105.190 124.715 ;
        RECT 96.990 111.815 102.930 112.150 ;
        RECT 97.035 111.640 97.795 111.815 ;
        RECT 78.180 109.735 96.765 110.065 ;
        RECT 71.950 108.850 105.190 108.875 ;
        RECT 71.950 108.795 105.210 108.850 ;
        RECT 71.840 107.720 105.210 108.795 ;
        RECT 71.840 107.695 105.190 107.720 ;
        RECT 71.840 106.785 73.400 107.695 ;
        RECT 74.305 106.750 106.730 106.775 ;
        RECT 74.305 105.645 106.745 106.750 ;
        RECT 74.305 105.625 106.730 105.645 ;
        RECT 74.305 105.620 103.750 105.625 ;
        RECT 105.550 105.620 106.730 105.625 ;
        RECT 74.305 104.910 75.990 105.620 ;
        RECT 105.550 105.615 105.830 105.620 ;
        RECT 74.310 104.575 75.990 104.910 ;
        RECT 102.295 104.605 103.280 104.625 ;
        RECT 105.755 104.605 106.885 104.620 ;
        RECT 102.275 103.570 106.885 104.605 ;
        RECT 102.295 103.550 103.280 103.570 ;
        RECT 105.755 103.550 106.885 103.570 ;
        RECT 66.750 92.820 70.635 93.055 ;
        RECT 66.750 92.575 67.520 92.820 ;
        RECT 47.935 90.690 66.520 91.020 ;
        RECT 64.485 89.000 65.475 89.015 ;
        RECT 64.485 87.965 65.485 89.000 ;
        RECT 37.220 85.650 39.680 86.650 ;
        RECT 63.190 85.620 64.190 86.680 ;
        RECT 60.105 82.140 63.060 83.650 ;
        RECT 60.255 74.535 61.465 82.140 ;
        RECT 63.575 79.525 64.165 85.620 ;
        RECT 60.130 73.075 62.640 74.535 ;
        RECT 60.255 66.615 61.465 73.075 ;
        RECT 60.145 66.530 62.765 66.615 ;
        RECT 59.795 65.250 62.770 66.530 ;
        RECT 60.145 65.180 62.765 65.250 ;
        RECT 60.255 50.915 61.470 65.180 ;
        RECT 63.605 62.340 64.135 79.525 ;
        RECT 64.800 79.375 65.485 87.965 ;
        RECT 95.250 87.430 96.650 87.460 ;
        RECT 90.920 86.030 96.650 87.430 ;
        RECT 95.250 86.000 96.650 86.030 ;
        RECT 119.190 86.000 120.590 167.405 ;
        RECT 94.170 82.055 95.810 83.695 ;
        RECT 113.295 83.240 114.205 83.260 ;
        RECT 121.530 83.240 122.490 166.765 ;
        RECT 96.115 81.055 96.615 81.455 ;
        RECT 64.835 62.950 65.450 79.375 ;
        RECT 68.445 60.760 69.835 70.690 ;
        RECT 71.475 68.900 71.825 71.735 ;
        RECT 72.500 65.255 85.400 74.655 ;
        RECT 96.215 71.805 96.515 81.055 ;
        RECT 99.415 78.155 103.815 83.055 ;
        RECT 109.460 82.280 114.230 83.240 ;
        RECT 119.660 82.280 122.490 83.240 ;
        RECT 89.450 71.405 89.850 71.805 ;
        RECT 96.115 71.405 96.615 71.805 ;
        RECT 89.500 69.305 89.800 71.405 ;
        RECT 99.415 70.805 103.815 74.755 ;
        RECT 99.415 69.355 104.815 70.805 ;
        RECT 89.470 69.005 89.830 69.305 ;
        RECT 96.115 68.505 96.665 68.905 ;
        RECT 96.215 65.305 96.515 68.505 ;
        RECT 99.415 67.005 103.815 69.355 ;
        RECT 96.115 64.905 96.665 65.305 ;
        RECT 77.690 63.900 83.910 64.330 ;
        RECT 84.400 63.910 84.750 64.390 ;
        RECT 77.615 63.100 77.875 63.420 ;
        RECT 81.310 63.320 81.490 63.540 ;
        RECT 77.240 59.630 77.510 60.820 ;
        RECT 76.385 58.930 76.925 58.950 ;
        RECT 76.385 58.720 76.950 58.930 ;
        RECT 76.355 58.390 76.950 58.720 ;
        RECT 62.625 53.360 63.055 53.380 ;
        RECT 60.255 50.900 62.160 50.915 ;
        RECT 62.600 50.900 63.080 53.360 ;
        RECT 76.470 52.835 76.950 58.390 ;
        RECT 77.280 57.240 77.430 59.630 ;
        RECT 77.650 59.450 77.845 63.100 ;
        RECT 81.310 62.970 81.640 63.320 ;
        RECT 78.310 62.350 78.710 62.790 ;
        RECT 79.950 62.770 80.290 62.830 ;
        RECT 77.620 59.080 77.900 59.450 ;
        RECT 78.060 58.030 78.230 60.650 ;
        RECT 78.470 59.810 78.710 62.350 ;
        RECT 79.880 62.390 80.290 62.770 ;
        RECT 81.340 62.410 81.640 62.970 ;
        RECT 78.390 59.370 78.710 59.810 ;
        RECT 79.360 61.190 79.670 61.640 ;
        RECT 77.225 56.920 77.485 57.240 ;
        RECT 77.280 52.755 77.430 56.920 ;
        RECT 77.620 55.750 79.190 56.180 ;
        RECT 79.360 55.730 79.660 61.190 ;
        RECT 79.880 60.350 80.130 62.390 ;
        RECT 80.670 60.740 80.930 61.060 ;
        RECT 81.370 60.930 81.620 62.410 ;
        RECT 81.780 61.200 84.220 61.630 ;
        RECT 79.875 60.030 80.135 60.350 ;
        RECT 80.300 57.480 80.580 58.280 ;
        RECT 80.340 53.125 80.490 57.480 ;
        RECT 80.735 57.320 80.885 60.740 ;
        RECT 81.330 60.550 81.650 60.930 ;
        RECT 82.090 60.420 82.350 60.740 ;
        RECT 83.030 60.570 83.290 60.890 ;
        RECT 82.135 59.365 82.305 60.420 ;
        RECT 82.570 60.100 82.830 60.420 ;
        RECT 82.595 59.730 82.805 60.100 ;
        RECT 82.540 59.470 82.860 59.730 ;
        RECT 82.090 59.045 82.350 59.365 ;
        RECT 81.170 58.460 82.800 58.890 ;
        RECT 81.670 57.480 81.930 58.270 ;
        RECT 80.680 57.000 80.940 57.320 ;
        RECT 80.735 55.370 80.885 57.000 ;
        RECT 81.730 55.415 81.880 57.480 ;
        RECT 83.050 57.340 83.270 60.570 ;
        RECT 84.430 58.480 84.730 63.910 ;
        RECT 86.310 63.850 86.660 64.350 ;
        RECT 84.960 61.190 86.130 61.620 ;
        RECT 85.820 59.970 86.160 60.950 ;
        RECT 83.520 57.460 83.810 58.170 ;
        RECT 84.480 57.860 84.740 58.180 ;
        RECT 85.820 57.860 86.080 59.970 ;
        RECT 86.360 59.260 86.660 63.850 ;
        RECT 94.140 62.205 95.800 63.805 ;
        RECT 99.415 63.605 103.815 66.655 ;
        RECT 87.200 61.560 87.490 61.610 ;
        RECT 86.320 58.420 86.720 59.260 ;
        RECT 83.050 56.940 83.380 57.340 ;
        RECT 80.730 53.490 80.895 55.370 ;
        RECT 81.710 53.890 81.905 55.415 ;
        RECT 83.075 55.390 83.245 56.940 ;
        RECT 83.580 55.410 83.730 57.460 ;
        RECT 84.505 57.320 84.715 57.860 ;
        RECT 84.480 57.000 84.740 57.320 ;
        RECT 84.530 55.525 84.695 57.000 ;
        RECT 84.970 56.440 85.280 57.300 ;
        RECT 84.990 55.530 85.155 56.440 ;
        RECT 85.390 55.750 86.960 56.180 ;
        RECT 87.190 55.750 87.490 61.560 ;
        RECT 94.170 56.530 95.770 62.205 ;
        RECT 101.200 58.280 102.400 63.605 ;
        RECT 109.600 59.975 110.285 82.280 ;
        RECT 113.295 82.260 114.205 82.280 ;
        RECT 132.340 61.200 132.620 61.345 ;
        RECT 131.845 60.150 132.955 61.200 ;
        RECT 101.180 57.130 102.420 58.280 ;
        RECT 109.800 57.825 110.080 59.975 ;
        RECT 101.200 57.105 102.400 57.130 ;
        RECT 106.800 56.170 108.340 56.540 ;
        RECT 83.060 54.285 83.265 55.390 ;
        RECT 83.555 54.670 83.755 55.410 ;
        RECT 84.515 55.050 84.715 55.525 ;
        RECT 84.960 55.295 89.285 55.530 ;
        RECT 109.870 55.325 110.010 57.825 ;
        RECT 132.340 57.345 132.620 60.150 ;
        RECT 132.340 57.275 132.550 57.345 ;
        RECT 113.400 56.170 114.940 56.540 ;
        RECT 120.000 56.170 121.540 56.540 ;
        RECT 126.600 56.170 128.140 56.540 ;
        RECT 84.990 55.210 85.155 55.295 ;
        RECT 84.515 54.850 88.900 55.050 ;
        RECT 83.555 54.470 88.530 54.670 ;
        RECT 83.060 54.080 88.120 54.285 ;
        RECT 81.710 53.695 87.715 53.890 ;
        RECT 80.720 53.300 87.305 53.490 ;
        RECT 80.320 52.935 86.915 53.125 ;
        RECT 77.270 52.580 86.565 52.755 ;
        RECT 84.080 52.350 84.630 52.360 ;
        RECT 83.930 52.340 84.630 52.350 ;
        RECT 64.950 52.010 84.630 52.340 ;
        RECT 65.670 51.780 71.450 52.010 ;
        RECT 64.540 51.300 71.960 51.780 ;
        RECT 74.410 51.760 80.190 52.010 ;
        RECT 73.750 51.280 81.170 51.760 ;
        RECT 82.790 51.390 83.340 51.860 ;
        RECT 83.930 51.790 84.630 52.010 ;
        RECT 83.930 51.770 85.140 51.790 ;
        RECT 83.930 51.180 85.150 51.770 ;
        RECT 83.930 51.160 84.630 51.180 ;
        RECT 60.255 49.900 63.080 50.900 ;
        RECT 82.670 50.160 83.220 50.720 ;
        RECT 60.255 47.595 62.810 49.900 ;
        RECT 63.060 47.880 71.930 48.340 ;
        RECT 74.440 47.960 83.310 48.420 ;
        RECT 60.255 45.495 61.470 47.595 ;
        RECT 62.030 45.495 62.810 47.595 ;
        RECT 66.580 47.555 71.090 47.880 ;
        RECT 76.940 47.555 81.450 47.960 ;
        RECT 84.820 47.555 85.150 51.180 ;
        RECT 85.370 50.440 85.920 50.680 ;
        RECT 86.390 50.440 86.565 52.580 ;
        RECT 85.370 50.265 86.565 50.440 ;
        RECT 85.370 50.120 85.920 50.265 ;
        RECT 85.330 49.325 85.870 49.480 ;
        RECT 86.725 49.325 86.915 52.935 ;
        RECT 85.330 49.110 86.930 49.325 ;
        RECT 85.330 48.890 85.870 49.110 ;
        RECT 66.565 47.225 85.150 47.555 ;
        RECT 85.350 47.250 85.900 47.950 ;
        RECT 84.090 47.000 84.640 47.010 ;
        RECT 83.940 46.990 84.640 47.000 ;
        RECT 64.960 46.660 84.640 46.990 ;
        RECT 65.680 46.430 71.460 46.660 ;
        RECT 64.550 45.950 71.970 46.430 ;
        RECT 74.420 46.410 80.200 46.660 ;
        RECT 73.760 45.930 81.180 46.410 ;
        RECT 82.770 46.010 83.320 46.480 ;
        RECT 83.940 46.440 84.640 46.660 ;
        RECT 83.940 46.420 85.150 46.440 ;
        RECT 83.940 45.830 85.160 46.420 ;
        RECT 83.940 45.810 84.640 45.830 ;
        RECT 60.255 42.175 62.810 45.495 ;
        RECT 82.770 44.860 83.360 45.330 ;
        RECT 63.070 42.530 71.940 42.990 ;
        RECT 74.450 42.610 83.320 43.070 ;
        RECT 66.590 42.205 71.100 42.530 ;
        RECT 76.950 42.205 81.460 42.610 ;
        RECT 84.830 42.205 85.160 45.830 ;
        RECT 85.360 45.195 85.950 45.320 ;
        RECT 87.115 45.195 87.305 53.300 ;
        RECT 85.360 45.005 87.305 45.195 ;
        RECT 85.360 44.850 85.950 45.005 ;
        RECT 85.465 44.845 85.655 44.850 ;
        RECT 85.370 43.940 86.210 44.180 ;
        RECT 87.520 43.940 87.715 53.695 ;
        RECT 85.370 43.745 87.715 43.940 ;
        RECT 85.370 43.470 86.210 43.745 ;
        RECT 60.255 40.105 61.470 42.175 ;
        RECT 62.030 40.105 62.810 42.175 ;
        RECT 66.575 41.875 85.160 42.205 ;
        RECT 84.060 41.650 84.610 41.660 ;
        RECT 83.910 41.640 84.610 41.650 ;
        RECT 64.930 41.310 84.610 41.640 ;
        RECT 65.650 41.080 71.430 41.310 ;
        RECT 64.520 40.600 71.940 41.080 ;
        RECT 74.390 41.060 80.170 41.310 ;
        RECT 73.730 40.580 81.150 41.060 ;
        RECT 82.740 40.650 83.290 41.120 ;
        RECT 83.910 41.090 84.610 41.310 ;
        RECT 83.910 41.070 85.120 41.090 ;
        RECT 83.910 40.480 85.130 41.070 ;
        RECT 83.910 40.460 84.610 40.480 ;
        RECT 60.255 36.785 62.810 40.105 ;
        RECT 82.730 39.490 83.320 40.010 ;
        RECT 63.040 37.180 71.910 37.640 ;
        RECT 74.420 37.260 83.290 37.720 ;
        RECT 66.560 36.855 71.070 37.180 ;
        RECT 76.920 36.855 81.430 37.260 ;
        RECT 84.800 36.855 85.130 40.480 ;
        RECT 85.350 39.955 85.940 40.010 ;
        RECT 87.915 39.955 88.120 54.080 ;
        RECT 85.350 39.750 88.120 39.955 ;
        RECT 85.350 39.490 85.940 39.750 ;
        RECT 85.450 38.800 86.080 39.030 ;
        RECT 88.330 38.800 88.530 54.470 ;
        RECT 85.400 38.600 88.530 38.800 ;
        RECT 85.450 38.260 86.080 38.600 ;
        RECT 60.255 35.425 61.470 36.785 ;
        RECT 62.030 35.425 62.810 36.785 ;
        RECT 66.545 36.525 85.130 36.855 ;
        RECT 84.100 36.370 84.650 36.380 ;
        RECT 83.950 36.360 84.650 36.370 ;
        RECT 64.970 36.030 84.650 36.360 ;
        RECT 65.690 35.800 71.470 36.030 ;
        RECT 60.255 33.910 62.810 35.425 ;
        RECT 64.560 35.320 71.980 35.800 ;
        RECT 74.430 35.780 80.210 36.030 ;
        RECT 83.950 35.810 84.650 36.030 ;
        RECT 83.950 35.790 85.160 35.810 ;
        RECT 73.770 35.300 81.190 35.780 ;
        RECT 82.770 35.290 83.320 35.760 ;
        RECT 83.950 35.200 85.170 35.790 ;
        RECT 83.950 35.180 84.650 35.200 ;
        RECT 82.530 34.130 83.460 34.820 ;
        RECT 60.255 33.900 62.780 33.910 ;
        RECT 60.255 31.740 62.040 33.900 ;
        RECT 63.080 31.900 71.950 32.360 ;
        RECT 74.460 31.980 83.330 32.440 ;
        RECT 60.255 31.525 62.020 31.740 ;
        RECT 66.600 31.575 71.110 31.900 ;
        RECT 76.960 31.575 81.470 31.980 ;
        RECT 84.840 31.575 85.170 35.200 ;
        RECT 85.430 34.740 86.080 34.770 ;
        RECT 88.700 34.740 88.900 54.850 ;
        RECT 85.430 34.540 88.900 34.740 ;
        RECT 85.430 34.300 86.080 34.540 ;
        RECT 85.400 33.610 86.170 33.800 ;
        RECT 89.050 33.610 89.285 55.295 ;
        RECT 109.810 55.005 110.070 55.325 ;
        RECT 108.430 53.985 108.690 54.305 ;
        RECT 103.500 53.450 105.040 53.820 ;
        RECT 106.800 50.730 108.340 51.100 ;
        RECT 105.670 49.565 105.930 49.885 ;
        RECT 103.500 48.010 105.040 48.380 ;
        RECT 105.730 46.145 105.870 49.565 ;
        RECT 108.490 49.545 108.630 53.985 ;
        RECT 110.100 53.450 111.640 53.820 ;
        RECT 116.700 53.450 118.240 53.820 ;
        RECT 123.300 53.450 124.840 53.820 ;
        RECT 129.900 53.450 131.440 53.820 ;
        RECT 113.400 50.730 114.940 51.100 ;
        RECT 120.000 50.730 121.540 51.100 ;
        RECT 126.600 50.730 128.140 51.100 ;
        RECT 108.430 49.225 108.690 49.545 ;
        RECT 105.670 45.825 105.930 46.145 ;
        RECT 105.730 44.445 105.870 45.825 ;
        RECT 106.800 45.290 108.340 45.660 ;
        RECT 108.490 44.785 108.630 49.225 ;
        RECT 112.110 48.885 112.370 49.205 ;
        RECT 110.100 48.010 111.640 48.380 ;
        RECT 108.890 46.505 109.150 46.825 ;
        RECT 108.430 44.465 108.690 44.785 ;
        RECT 105.670 44.125 105.930 44.445 ;
        RECT 103.500 42.570 105.040 42.940 ;
        RECT 105.730 41.965 105.870 44.125 ;
        RECT 106.130 43.445 106.390 43.765 ;
        RECT 106.190 42.405 106.330 43.445 ;
        RECT 106.130 42.085 106.390 42.405 ;
        RECT 105.270 41.825 105.870 41.965 ;
        RECT 105.270 41.045 105.410 41.825 ;
        RECT 105.210 40.725 105.470 41.045 ;
        RECT 103.500 37.130 105.040 37.500 ;
        RECT 85.400 33.375 89.285 33.610 ;
        RECT 85.400 33.130 86.170 33.375 ;
        RECT 103.500 31.690 105.040 32.060 ;
        RECT 60.255 17.535 61.470 31.525 ;
        RECT 66.585 31.245 85.170 31.575 ;
        RECT 104.750 29.505 105.010 29.825 ;
        RECT 104.810 28.125 104.950 29.505 ;
        RECT 104.750 27.805 105.010 28.125 ;
        RECT 103.500 26.250 105.040 26.620 ;
        RECT 103.500 20.810 105.040 21.180 ;
        RECT 105.270 19.625 105.410 40.725 ;
        RECT 105.670 27.805 105.930 28.125 ;
        RECT 105.730 23.025 105.870 27.805 ;
        RECT 105.670 22.705 105.930 23.025 ;
        RECT 106.190 19.625 106.330 42.085 ;
        RECT 108.490 40.705 108.630 44.465 ;
        RECT 108.950 43.425 109.090 46.505 ;
        RECT 112.170 46.485 112.310 48.885 ;
        RECT 116.700 48.010 118.240 48.380 ;
        RECT 123.300 48.010 124.840 48.380 ;
        RECT 129.900 48.010 131.440 48.380 ;
        RECT 112.110 46.165 112.370 46.485 ;
        RECT 113.400 45.290 114.940 45.660 ;
        RECT 120.000 45.290 121.540 45.660 ;
        RECT 126.600 45.290 128.140 45.660 ;
        RECT 113.030 44.805 113.290 45.125 ;
        RECT 112.570 44.125 112.830 44.445 ;
        RECT 108.890 43.105 109.150 43.425 ;
        RECT 108.430 40.385 108.690 40.705 ;
        RECT 106.800 39.850 108.340 40.220 ;
        RECT 108.950 36.965 109.090 43.105 ;
        RECT 110.100 42.570 111.640 42.940 ;
        RECT 112.630 42.405 112.770 44.125 ;
        RECT 112.570 42.085 112.830 42.405 ;
        RECT 112.110 41.405 112.370 41.725 ;
        RECT 110.100 37.130 111.640 37.500 ;
        RECT 108.890 36.645 109.150 36.965 ;
        RECT 106.800 34.410 108.340 34.780 ;
        RECT 108.950 30.845 109.090 36.645 ;
        RECT 110.100 31.690 111.640 32.060 ;
        RECT 112.170 31.525 112.310 41.405 ;
        RECT 113.090 41.385 113.230 44.805 ;
        RECT 116.700 42.570 118.240 42.940 ;
        RECT 123.300 42.570 124.840 42.940 ;
        RECT 129.900 42.570 131.440 42.940 ;
        RECT 132.410 41.805 132.550 57.275 ;
        RECT 133.200 56.170 134.740 56.540 ;
        RECT 139.800 56.170 141.340 56.540 ;
        RECT 136.500 53.450 138.040 53.820 ;
        RECT 133.200 50.730 134.740 51.100 ;
        RECT 139.800 50.730 141.340 51.100 ;
        RECT 136.500 48.010 138.040 48.380 ;
        RECT 133.200 45.290 134.740 45.660 ;
        RECT 139.800 45.290 141.340 45.660 ;
        RECT 136.500 42.570 138.040 42.940 ;
        RECT 131.950 41.665 132.550 41.805 ;
        RECT 113.030 41.065 113.290 41.385 ;
        RECT 113.400 39.850 114.940 40.220 ;
        RECT 120.000 39.850 121.540 40.220 ;
        RECT 126.600 39.850 128.140 40.220 ;
        RECT 116.700 37.130 118.240 37.500 ;
        RECT 123.300 37.130 124.840 37.500 ;
        RECT 129.900 37.130 131.440 37.500 ;
        RECT 131.950 35.945 132.090 41.665 ;
        RECT 133.200 39.850 134.740 40.220 ;
        RECT 139.800 39.850 141.340 40.220 ;
        RECT 136.500 37.130 138.040 37.500 ;
        RECT 131.890 35.625 132.150 35.945 ;
        RECT 124.990 35.005 125.250 35.265 ;
        RECT 124.990 34.945 125.650 35.005 ;
        RECT 125.050 34.865 125.650 34.945 ;
        RECT 113.400 34.410 114.940 34.780 ;
        RECT 120.000 34.410 121.540 34.780 ;
        RECT 125.510 34.325 125.650 34.865 ;
        RECT 126.600 34.410 128.140 34.780 ;
        RECT 133.200 34.410 134.740 34.780 ;
        RECT 139.800 34.410 141.340 34.780 ;
        RECT 125.510 34.185 126.110 34.325 ;
        RECT 118.550 32.565 118.810 32.885 ;
        RECT 116.700 31.690 118.240 32.060 ;
        RECT 112.110 31.205 112.370 31.525 ;
        RECT 108.890 30.525 109.150 30.845 ;
        RECT 106.800 28.970 108.340 29.340 ;
        RECT 108.950 28.465 109.090 30.525 ;
        RECT 112.170 29.825 112.310 31.205 ;
        RECT 115.330 30.865 115.590 31.185 ;
        RECT 112.570 30.185 112.830 30.505 ;
        RECT 112.110 29.505 112.370 29.825 ;
        RECT 107.970 28.145 108.230 28.465 ;
        RECT 108.890 28.145 109.150 28.465 ;
        RECT 108.030 25.065 108.170 28.145 ;
        RECT 110.100 26.250 111.640 26.620 ;
        RECT 112.170 26.085 112.310 29.505 ;
        RECT 112.630 28.805 112.770 30.185 ;
        RECT 113.030 29.845 113.290 30.165 ;
        RECT 112.570 28.485 112.830 28.805 ;
        RECT 112.110 25.765 112.370 26.085 ;
        RECT 107.970 24.745 108.230 25.065 ;
        RECT 109.810 24.405 110.070 24.725 ;
        RECT 106.800 23.530 108.340 23.900 ;
        RECT 109.870 23.365 110.010 24.405 ;
        RECT 109.810 23.045 110.070 23.365 ;
        RECT 112.630 22.005 112.770 28.485 ;
        RECT 113.090 27.785 113.230 29.845 ;
        RECT 113.400 28.970 114.940 29.340 ;
        RECT 115.390 28.125 115.530 30.865 ;
        RECT 115.330 27.805 115.590 28.125 ;
        RECT 118.610 27.785 118.750 32.565 ;
        RECT 119.930 32.225 120.190 32.545 ;
        RECT 119.990 30.505 120.130 32.225 ;
        RECT 123.300 31.690 124.840 32.060 ;
        RECT 124.990 30.865 125.250 31.185 ;
        RECT 122.230 30.525 122.490 30.845 ;
        RECT 119.930 30.185 120.190 30.505 ;
        RECT 121.770 30.185 122.030 30.505 ;
        RECT 122.290 30.245 122.430 30.525 ;
        RECT 119.010 29.505 119.270 29.825 ;
        RECT 113.030 27.465 113.290 27.785 ;
        RECT 118.550 27.465 118.810 27.785 ;
        RECT 119.070 27.445 119.210 29.505 ;
        RECT 120.000 28.970 121.540 29.340 ;
        RECT 119.930 28.485 120.190 28.805 ;
        RECT 119.010 27.125 119.270 27.445 ;
        RECT 116.700 26.250 118.240 26.620 ;
        RECT 115.790 25.765 116.050 26.085 ;
        RECT 113.030 24.065 113.290 24.385 ;
        RECT 113.090 22.685 113.230 24.065 ;
        RECT 113.400 23.530 114.940 23.900 ;
        RECT 115.850 22.685 115.990 25.765 ;
        RECT 119.070 25.745 119.210 27.125 ;
        RECT 119.990 26.085 120.130 28.485 ;
        RECT 121.310 27.805 121.570 28.125 ;
        RECT 120.390 27.640 120.650 27.785 ;
        RECT 120.380 27.270 120.660 27.640 ;
        RECT 120.850 27.125 121.110 27.445 ;
        RECT 119.930 25.765 120.190 26.085 ;
        RECT 119.010 25.425 119.270 25.745 ;
        RECT 118.550 24.745 118.810 25.065 ;
        RECT 118.610 23.365 118.750 24.745 ;
        RECT 118.550 23.045 118.810 23.365 ;
        RECT 116.250 22.705 116.510 23.025 ;
        RECT 113.030 22.365 113.290 22.685 ;
        RECT 115.790 22.365 116.050 22.685 ;
        RECT 112.570 21.685 112.830 22.005 ;
        RECT 110.100 20.810 111.640 21.180 ;
        RECT 112.630 19.625 112.770 21.685 ;
        RECT 116.310 19.625 116.450 22.705 ;
        RECT 119.070 21.665 119.210 25.425 ;
        RECT 120.910 24.385 121.050 27.125 ;
        RECT 121.370 25.485 121.510 27.805 ;
        RECT 121.830 26.085 121.970 30.185 ;
        RECT 122.290 30.105 122.890 30.245 ;
        RECT 122.230 29.505 122.490 29.825 ;
        RECT 122.290 28.465 122.430 29.505 ;
        RECT 122.230 28.145 122.490 28.465 ;
        RECT 121.770 25.765 122.030 26.085 ;
        RECT 122.230 25.765 122.490 26.085 ;
        RECT 122.290 25.485 122.430 25.765 ;
        RECT 121.370 25.345 122.430 25.485 ;
        RECT 122.750 24.725 122.890 30.105 ;
        RECT 125.050 27.640 125.190 30.865 ;
        RECT 125.970 30.505 126.110 34.185 ;
        RECT 129.130 33.925 129.390 34.245 ;
        RECT 126.830 33.585 127.090 33.905 ;
        RECT 126.370 32.905 126.630 33.225 ;
        RECT 125.910 30.185 126.170 30.505 ;
        RECT 126.430 29.825 126.570 32.905 ;
        RECT 126.890 32.885 127.030 33.585 ;
        RECT 128.210 33.245 128.470 33.565 ;
        RECT 126.830 32.565 127.090 32.885 ;
        RECT 127.750 32.565 128.010 32.885 ;
        RECT 127.810 31.185 127.950 32.565 ;
        RECT 128.270 31.525 128.410 33.245 ;
        RECT 128.210 31.205 128.470 31.525 ;
        RECT 127.750 30.865 128.010 31.185 ;
        RECT 128.670 30.525 128.930 30.845 ;
        RECT 125.450 29.505 125.710 29.825 ;
        RECT 125.910 29.505 126.170 29.825 ;
        RECT 126.370 29.505 126.630 29.825 ;
        RECT 124.980 27.270 125.260 27.640 ;
        RECT 123.300 26.250 124.840 26.620 ;
        RECT 122.690 24.405 122.950 24.725 ;
        RECT 124.070 24.635 124.330 24.725 ;
        RECT 125.050 24.635 125.190 27.270 ;
        RECT 124.070 24.495 125.190 24.635 ;
        RECT 124.070 24.405 124.330 24.495 ;
        RECT 120.850 24.065 121.110 24.385 ;
        RECT 120.000 23.530 121.540 23.900 ;
        RECT 122.750 22.685 122.890 24.405 ;
        RECT 122.690 22.365 122.950 22.685 ;
        RECT 125.050 21.665 125.190 24.495 ;
        RECT 125.510 23.365 125.650 29.505 ;
        RECT 125.970 24.725 126.110 29.505 ;
        RECT 126.600 28.970 128.140 29.340 ;
        RECT 128.210 27.805 128.470 28.125 ;
        RECT 126.370 26.785 126.630 27.105 ;
        RECT 126.430 25.065 126.570 26.785 ;
        RECT 128.270 26.085 128.410 27.805 ;
        RECT 128.210 25.765 128.470 26.085 ;
        RECT 126.370 24.745 126.630 25.065 ;
        RECT 125.910 24.405 126.170 24.725 ;
        RECT 128.730 24.385 128.870 30.525 ;
        RECT 129.190 28.125 129.330 33.925 ;
        RECT 131.890 33.245 132.150 33.565 ;
        RECT 129.900 31.690 131.440 32.060 ;
        RECT 130.970 29.505 131.230 29.825 ;
        RECT 131.030 28.125 131.170 29.505 ;
        RECT 131.950 28.805 132.090 33.245 ;
        RECT 132.810 32.905 133.070 33.225 ;
        RECT 131.890 28.485 132.150 28.805 ;
        RECT 131.950 28.205 132.090 28.485 ;
        RECT 129.130 27.805 129.390 28.125 ;
        RECT 130.970 27.805 131.230 28.125 ;
        RECT 131.950 28.065 132.550 28.205 ;
        RECT 131.030 27.525 131.170 27.805 ;
        RECT 131.030 27.385 132.090 27.525 ;
        RECT 129.130 26.785 129.390 27.105 ;
        RECT 128.670 24.065 128.930 24.385 ;
        RECT 126.600 23.530 128.140 23.900 ;
        RECT 125.450 23.045 125.710 23.365 ;
        RECT 128.730 23.025 128.870 24.065 ;
        RECT 128.670 22.705 128.930 23.025 ;
        RECT 126.830 22.365 127.090 22.685 ;
        RECT 127.290 22.365 127.550 22.685 ;
        RECT 125.910 21.685 126.170 22.005 ;
        RECT 119.010 21.345 119.270 21.665 ;
        RECT 124.990 21.345 125.250 21.665 ;
        RECT 116.700 20.810 118.240 21.180 ;
        RECT 123.300 20.810 124.840 21.180 ;
        RECT 125.050 19.625 125.190 21.345 ;
        RECT 125.970 19.625 126.110 21.685 ;
        RECT 126.890 19.625 127.030 22.365 ;
        RECT 127.350 22.005 127.490 22.365 ;
        RECT 129.190 22.345 129.330 26.785 ;
        RECT 129.900 26.250 131.440 26.620 ;
        RECT 130.050 25.765 130.310 26.085 ;
        RECT 129.590 24.405 129.850 24.725 ;
        RECT 129.130 22.025 129.390 22.345 ;
        RECT 129.650 22.085 129.790 24.405 ;
        RECT 130.110 22.685 130.250 25.765 ;
        RECT 131.950 25.485 132.090 27.385 ;
        RECT 131.490 25.345 132.090 25.485 ;
        RECT 131.490 25.065 131.630 25.345 ;
        RECT 131.430 24.745 131.690 25.065 ;
        RECT 132.410 24.805 132.550 28.065 ;
        RECT 131.950 24.665 132.550 24.805 ;
        RECT 131.950 23.365 132.090 24.665 ;
        RECT 131.890 23.045 132.150 23.365 ;
        RECT 130.050 22.365 130.310 22.685 ;
        RECT 130.970 22.365 131.230 22.685 ;
        RECT 131.030 22.085 131.170 22.365 ;
        RECT 127.290 21.685 127.550 22.005 ;
        RECT 129.650 21.945 131.170 22.085 ;
        RECT 132.870 21.665 133.010 32.905 ;
        RECT 135.110 32.225 135.370 32.545 ;
        RECT 135.570 32.225 135.830 32.545 ;
        RECT 133.200 28.970 134.740 29.340 ;
        RECT 133.200 23.530 134.740 23.900 ;
        RECT 135.170 23.365 135.310 32.225 ;
        RECT 135.630 28.465 135.770 32.225 ;
        RECT 136.500 31.690 138.040 32.060 ;
        RECT 139.800 28.970 141.340 29.340 ;
        RECT 135.570 28.145 135.830 28.465 ;
        RECT 139.250 26.785 139.510 27.105 ;
        RECT 136.500 26.250 138.040 26.620 ;
        RECT 136.030 24.405 136.290 24.725 ;
        RECT 135.570 24.065 135.830 24.385 ;
        RECT 134.190 23.045 134.450 23.365 ;
        RECT 135.110 23.045 135.370 23.365 ;
        RECT 134.250 22.345 134.390 23.045 ;
        RECT 134.190 22.025 134.450 22.345 ;
        RECT 132.810 21.345 133.070 21.665 ;
        RECT 129.900 20.810 131.440 21.180 ;
        RECT 135.630 19.625 135.770 24.065 ;
        RECT 136.090 22.345 136.230 24.405 ;
        RECT 137.870 24.065 138.130 24.385 ;
        RECT 137.930 22.685 138.070 24.065 ;
        RECT 139.310 23.025 139.450 26.785 ;
        RECT 139.800 23.530 141.340 23.900 ;
        RECT 139.250 22.705 139.510 23.025 ;
        RECT 137.870 22.365 138.130 22.685 ;
        RECT 136.030 22.025 136.290 22.345 ;
        RECT 137.930 22.085 138.070 22.365 ;
        RECT 137.930 21.945 138.530 22.085 ;
        RECT 136.500 20.810 138.040 21.180 ;
        RECT 138.390 19.625 138.530 21.945 ;
        RECT 139.310 19.625 139.450 22.705 ;
        RECT 142.930 19.985 143.190 20.305 ;
        RECT 105.210 19.305 105.470 19.625 ;
        RECT 106.130 19.305 106.390 19.625 ;
        RECT 112.570 19.305 112.830 19.625 ;
        RECT 116.250 19.305 116.510 19.625 ;
        RECT 124.990 19.305 125.250 19.625 ;
        RECT 125.910 19.305 126.170 19.625 ;
        RECT 126.830 19.305 127.090 19.625 ;
        RECT 135.570 19.305 135.830 19.625 ;
        RECT 138.330 19.305 138.590 19.625 ;
        RECT 139.250 19.305 139.510 19.625 ;
        RECT 101.530 18.625 101.790 18.945 ;
        RECT 106.130 18.625 106.390 18.945 ;
        RECT 110.730 18.625 110.990 18.945 ;
        RECT 115.330 18.625 115.590 18.945 ;
        RECT 119.470 18.625 119.730 18.945 ;
        RECT 124.530 18.625 124.790 18.945 ;
        RECT 129.130 18.625 129.390 18.945 ;
        RECT 132.810 18.625 133.070 18.945 ;
        RECT 138.790 18.855 139.050 18.945 ;
        RECT 138.390 18.715 139.050 18.855 ;
        RECT 60.255 17.520 62.525 17.535 ;
        RECT 60.255 16.305 62.550 17.520 ;
        RECT 101.590 16.305 101.730 18.625 ;
        RECT 106.190 16.305 106.330 18.625 ;
        RECT 106.800 18.090 108.340 18.460 ;
        RECT 110.790 16.305 110.930 18.625 ;
        RECT 113.400 18.090 114.940 18.460 ;
        RECT 115.390 16.305 115.530 18.625 ;
        RECT 119.530 17.355 119.670 18.625 ;
        RECT 120.000 18.090 121.540 18.460 ;
        RECT 119.530 17.215 120.130 17.355 ;
        RECT 119.530 17.205 119.670 17.215 ;
        RECT 119.990 16.305 120.130 17.215 ;
        RECT 124.590 16.305 124.730 18.625 ;
        RECT 126.600 18.090 128.140 18.460 ;
        RECT 129.190 16.305 129.330 18.625 ;
        RECT 132.870 17.155 133.010 18.625 ;
        RECT 133.200 18.090 134.740 18.460 ;
        RECT 132.870 17.015 133.930 17.155 ;
        RECT 133.790 16.305 133.930 17.015 ;
        RECT 138.390 16.305 138.530 18.715 ;
        RECT 138.790 18.625 139.050 18.715 ;
        RECT 139.800 18.090 141.340 18.460 ;
        RECT 142.990 16.305 143.130 19.985 ;
        RECT 61.360 16.280 62.525 16.305 ;
        RECT 101.520 12.305 101.800 16.305 ;
        RECT 106.120 12.305 106.400 16.305 ;
        RECT 110.720 12.305 111.000 16.305 ;
        RECT 115.320 15.175 115.600 16.305 ;
        RECT 115.200 12.315 115.720 15.175 ;
        RECT 115.320 12.305 115.600 12.315 ;
        RECT 119.920 12.305 120.200 16.305 ;
        RECT 124.520 12.305 124.800 16.305 ;
        RECT 129.120 12.305 129.400 16.305 ;
        RECT 133.720 15.150 134.000 16.305 ;
        RECT 133.585 11.120 134.135 15.150 ;
        RECT 138.320 12.305 138.600 16.305 ;
        RECT 142.920 12.305 143.200 16.305 ;
        RECT 93.735 1.425 94.865 3.545 ;
        RECT 112.995 1.695 114.250 4.115 ;
        RECT 132.345 1.570 133.540 3.795 ;
        RECT 151.575 2.225 152.950 5.355 ;
      LAYER met3 ;
        RECT 124.450 224.455 124.880 224.460 ;
        RECT 119.190 219.415 120.590 219.420 ;
        RECT 121.285 219.415 122.375 224.345 ;
        RECT 119.190 218.325 122.375 219.415 ;
        RECT 119.190 207.820 120.590 218.325 ;
        RECT 124.180 217.465 125.155 224.455 ;
        RECT 127.170 223.690 127.675 224.615 ;
        RECT 129.885 223.515 130.480 224.720 ;
        RECT 132.710 223.650 133.175 224.655 ;
        RECT 135.445 223.835 135.955 224.685 ;
        RECT 138.230 223.860 138.690 224.660 ;
        RECT 121.525 216.490 125.155 217.465 ;
        RECT 121.525 215.835 122.500 216.490 ;
        RECT 121.525 214.065 122.500 214.070 ;
        RECT 121.500 213.100 122.525 214.065 ;
        RECT 119.190 205.145 120.590 205.150 ;
        RECT 119.165 203.755 120.615 205.145 ;
        RECT 119.190 167.385 120.590 203.755 ;
        RECT 119.165 165.935 120.615 167.385 ;
        RECT 121.525 166.745 122.500 213.100 ;
        RECT 121.505 165.735 122.515 166.745 ;
        RECT 92.865 164.870 102.985 165.350 ;
        RECT 100.725 164.290 101.345 164.410 ;
        RECT 94.385 163.910 101.345 164.290 ;
        RECT 94.385 163.350 94.765 163.910 ;
        RECT 100.725 163.790 101.345 163.910 ;
        RECT 27.270 163.300 30.890 163.320 ;
        RECT 26.795 160.770 89.510 163.300 ;
        RECT 91.635 162.970 94.765 163.350 ;
        RECT 91.635 161.880 92.015 162.970 ;
        RECT 149.580 162.815 153.650 163.230 ;
        RECT 102.260 162.630 154.260 162.815 ;
        RECT 92.865 162.150 154.260 162.630 ;
        RECT 102.260 161.970 154.260 162.150 ;
        RECT 149.580 161.690 153.650 161.970 ;
        RECT 27.270 160.630 30.890 160.770 ;
        RECT 88.105 160.225 89.260 160.770 ;
        RECT 88.105 159.910 89.880 160.225 ;
        RECT 88.105 159.430 102.995 159.910 ;
        RECT 88.105 159.355 89.880 159.430 ;
        RECT 26.920 155.520 60.725 155.665 ;
        RECT 73.490 155.520 74.420 155.545 ;
        RECT 88.105 155.520 89.260 159.355 ;
        RECT 102.160 157.190 103.150 157.235 ;
        RECT 92.875 156.710 103.150 157.190 ;
        RECT 102.160 156.305 103.150 156.710 ;
        RECT 26.920 154.640 89.995 155.520 ;
        RECT 26.920 154.500 60.725 154.640 ;
        RECT 73.490 154.615 74.420 154.640 ;
        RECT 27.270 154.480 30.450 154.500 ;
        RECT 90.840 154.240 91.370 154.285 ;
        RECT 64.035 153.795 91.370 154.240 ;
        RECT 69.585 153.730 70.145 153.795 ;
        RECT 90.840 153.755 91.370 153.795 ;
        RECT 102.190 153.605 103.120 153.630 ;
        RECT 91.610 153.200 92.040 153.225 ;
        RECT 62.995 152.820 92.040 153.200 ;
        RECT 91.610 152.795 92.040 152.820 ;
        RECT 102.185 152.665 104.310 153.605 ;
        RECT 102.190 152.640 103.120 152.665 ;
        RECT 68.100 151.980 68.920 152.100 ;
        RECT 68.100 151.940 69.895 151.980 ;
        RECT 68.100 151.430 70.150 151.940 ;
        RECT 93.355 151.930 93.895 152.110 ;
        RECT 94.400 151.930 94.900 151.970 ;
        RECT 93.355 151.440 94.900 151.930 ;
        RECT 68.100 151.390 69.895 151.430 ;
        RECT 68.100 151.230 68.920 151.390 ;
        RECT 67.120 150.860 67.850 150.920 ;
        RECT 64.015 150.785 64.575 150.790 ;
        RECT 61.890 150.750 62.620 150.775 ;
        RECT 61.820 149.720 62.620 150.750 ;
        RECT 63.990 150.440 64.600 150.785 ;
        RECT 62.945 150.235 64.600 150.440 ;
        RECT 62.945 149.880 64.575 150.235 ;
        RECT 67.120 149.920 67.860 150.860 ;
        RECT 68.160 150.020 68.770 150.800 ;
        RECT 61.890 148.030 62.620 149.720 ;
        RECT 67.215 148.030 67.860 149.920 ;
        RECT 93.355 148.030 93.895 151.440 ;
        RECT 94.400 151.400 94.900 151.440 ;
        RECT 114.580 151.060 154.090 154.520 ;
        RECT 94.280 150.750 94.780 150.830 ;
        RECT 96.980 150.750 97.480 150.790 ;
        RECT 94.195 150.300 97.480 150.750 ;
        RECT 94.280 150.170 94.780 150.300 ;
        RECT 96.980 150.130 97.480 150.300 ;
        RECT 96.960 148.030 97.460 148.060 ;
        RECT 61.830 148.025 97.460 148.030 ;
        RECT 97.965 148.025 103.155 148.050 ;
        RECT 61.830 147.180 103.155 148.025 ;
        RECT 93.355 146.550 93.895 147.180 ;
        RECT 95.860 147.135 103.155 147.180 ;
        RECT 97.965 147.110 103.155 147.135 ;
        RECT 94.380 146.550 94.880 146.590 ;
        RECT 93.355 146.060 94.880 146.550 ;
        RECT 93.355 141.190 93.895 146.060 ;
        RECT 94.380 146.020 94.880 146.060 ;
        RECT 94.380 145.390 94.920 145.440 ;
        RECT 96.970 145.390 97.510 145.430 ;
        RECT 94.255 144.890 97.510 145.390 ;
        RECT 94.380 144.870 94.920 144.890 ;
        RECT 96.970 144.860 97.510 144.890 ;
        RECT 94.350 141.190 94.850 141.230 ;
        RECT 93.355 140.700 94.855 141.190 ;
        RECT 93.355 135.840 93.895 140.700 ;
        RECT 94.350 140.660 94.850 140.700 ;
        RECT 94.340 140.080 94.880 140.120 ;
        RECT 96.960 140.080 97.500 140.120 ;
        RECT 94.275 139.540 97.515 140.080 ;
        RECT 94.340 139.500 94.880 139.540 ;
        RECT 96.960 139.500 97.500 139.540 ;
        RECT 94.380 135.840 94.880 135.870 ;
        RECT 93.355 135.350 94.880 135.840 ;
        RECT 93.355 135.280 93.895 135.350 ;
        RECT 94.380 135.300 94.880 135.350 ;
        RECT 54.585 133.945 55.635 134.995 ;
        RECT 94.300 134.900 94.950 134.920 ;
        RECT 94.175 134.880 97.625 134.900 ;
        RECT 94.175 134.310 97.640 134.880 ;
        RECT 94.175 134.300 97.625 134.310 ;
        RECT 51.945 132.865 52.875 133.795 ;
        RECT 51.970 129.510 52.850 132.865 ;
        RECT 54.610 129.570 55.610 133.945 ;
        RECT 93.365 130.360 93.905 130.540 ;
        RECT 94.410 130.360 94.910 130.400 ;
        RECT 93.365 129.870 94.910 130.360 ;
        RECT 93.365 126.460 93.905 129.870 ;
        RECT 94.410 129.830 94.910 129.870 ;
        RECT 94.290 129.180 94.790 129.260 ;
        RECT 96.990 129.180 97.490 129.220 ;
        RECT 94.205 128.730 97.490 129.180 ;
        RECT 94.290 128.600 94.790 128.730 ;
        RECT 96.990 128.560 97.490 128.730 ;
        RECT 96.970 126.460 97.470 126.490 ;
        RECT 97.965 126.460 98.905 147.110 ;
        RECT 105.540 145.955 106.745 147.160 ;
        RECT 69.375 126.300 70.425 126.325 ;
        RECT 69.375 125.300 73.110 126.300 ;
        RECT 69.375 125.275 70.425 125.300 ;
        RECT 58.780 123.335 68.900 123.815 ;
        RECT 58.780 120.615 68.900 121.095 ;
        RECT 57.760 118.375 58.310 118.415 ;
        RECT 57.760 117.895 68.910 118.375 ;
        RECT 57.760 117.805 58.310 117.895 ;
        RECT 67.805 115.655 70.025 115.720 ;
        RECT 58.790 115.175 70.025 115.655 ;
        RECT 67.805 114.870 70.025 115.175 ;
        RECT 26.590 112.940 31.340 113.080 ;
        RECT 26.590 112.805 44.525 112.940 ;
        RECT 57.795 112.805 58.325 112.830 ;
        RECT 26.590 112.325 58.325 112.805 ;
        RECT 26.590 112.190 44.525 112.325 ;
        RECT 57.795 112.300 58.325 112.325 ;
        RECT 26.590 112.050 31.340 112.190 ;
        RECT 63.120 111.315 63.660 111.495 ;
        RECT 64.165 111.315 64.665 111.355 ;
        RECT 63.120 110.825 64.665 111.315 ;
        RECT 63.120 107.415 63.660 110.825 ;
        RECT 64.165 110.785 64.665 110.825 ;
        RECT 64.045 110.135 64.545 110.215 ;
        RECT 66.745 110.135 67.245 110.175 ;
        RECT 63.960 109.685 67.245 110.135 ;
        RECT 64.045 109.555 64.545 109.685 ;
        RECT 66.745 109.515 67.245 109.685 ;
        RECT 67.815 107.645 68.665 114.870 ;
        RECT 72.110 111.565 73.110 125.300 ;
        RECT 93.365 125.610 98.905 126.460 ;
        RECT 93.365 124.980 93.905 125.610 ;
        RECT 94.390 124.980 94.890 125.020 ;
        RECT 93.365 124.490 94.890 124.980 ;
        RECT 93.365 119.620 93.905 124.490 ;
        RECT 94.390 124.450 94.890 124.490 ;
        RECT 94.390 123.820 94.930 123.870 ;
        RECT 96.980 123.820 97.520 123.860 ;
        RECT 94.265 123.320 97.520 123.820 ;
        RECT 94.390 123.300 94.930 123.320 ;
        RECT 96.980 123.290 97.520 123.320 ;
        RECT 94.360 119.620 94.860 119.660 ;
        RECT 93.365 119.130 94.865 119.620 ;
        RECT 93.365 114.270 93.905 119.130 ;
        RECT 94.360 119.090 94.860 119.130 ;
        RECT 94.350 118.510 94.890 118.550 ;
        RECT 96.970 118.510 97.510 118.550 ;
        RECT 94.285 117.970 97.525 118.510 ;
        RECT 94.350 117.930 94.890 117.970 ;
        RECT 96.970 117.930 97.510 117.970 ;
        RECT 94.390 114.270 94.890 114.300 ;
        RECT 93.365 113.780 94.890 114.270 ;
        RECT 93.365 113.710 93.905 113.780 ;
        RECT 94.390 113.730 94.890 113.780 ;
        RECT 94.310 113.330 94.960 113.350 ;
        RECT 94.185 113.310 97.635 113.330 ;
        RECT 94.185 112.740 97.650 113.310 ;
        RECT 94.185 112.730 97.635 112.740 ;
        RECT 71.540 110.565 73.110 111.565 ;
        RECT 97.965 107.645 98.905 125.610 ;
        RECT 103.985 123.770 105.215 125.000 ;
        RECT 104.010 107.695 105.190 123.770 ;
        RECT 66.725 107.415 67.225 107.445 ;
        RECT 67.815 107.415 98.905 107.645 ;
        RECT 63.120 106.715 98.905 107.415 ;
        RECT 63.120 106.565 68.665 106.715 ;
        RECT 94.915 106.710 98.905 106.715 ;
        RECT 63.120 105.935 63.660 106.565 ;
        RECT 66.530 106.055 67.530 106.145 ;
        RECT 64.145 105.935 64.645 105.975 ;
        RECT 63.120 105.445 64.645 105.935 ;
        RECT 63.120 100.575 63.660 105.445 ;
        RECT 64.145 105.405 64.645 105.445 ;
        RECT 66.530 105.375 73.260 106.055 ;
        RECT 105.570 105.620 106.725 145.955 ;
        RECT 66.530 105.295 100.430 105.375 ;
        RECT 66.530 105.145 67.530 105.295 ;
        RECT 64.145 104.775 64.685 104.825 ;
        RECT 66.735 104.775 67.275 104.815 ;
        RECT 64.020 104.275 67.275 104.775 ;
        RECT 72.390 104.605 100.430 105.295 ;
        RECT 72.390 104.390 103.305 104.605 ;
        RECT 64.145 104.255 64.685 104.275 ;
        RECT 66.735 104.245 67.275 104.275 ;
        RECT 99.425 103.570 103.305 104.390 ;
        RECT 64.115 100.575 64.615 100.615 ;
        RECT 63.120 100.085 64.620 100.575 ;
        RECT 63.120 95.225 63.660 100.085 ;
        RECT 64.115 100.045 64.615 100.085 ;
        RECT 66.510 99.925 67.510 100.925 ;
        RECT 64.105 99.465 64.645 99.505 ;
        RECT 66.725 99.465 67.265 99.505 ;
        RECT 64.040 98.925 67.280 99.465 ;
        RECT 64.105 98.885 64.645 98.925 ;
        RECT 66.725 98.885 67.265 98.925 ;
        RECT 89.760 97.680 153.710 100.940 ;
        RECT 64.145 95.225 64.645 95.255 ;
        RECT 63.120 94.735 64.645 95.225 ;
        RECT 66.580 94.775 67.580 95.775 ;
        RECT 63.120 94.665 63.660 94.735 ;
        RECT 64.145 94.685 64.645 94.735 ;
        RECT 64.065 94.285 64.715 94.305 ;
        RECT 63.940 94.265 67.390 94.285 ;
        RECT 63.940 93.695 67.405 94.265 ;
        RECT 63.940 93.685 67.390 93.695 ;
        RECT 26.890 83.825 31.040 84.120 ;
        RECT 26.650 83.650 65.690 83.825 ;
        RECT 26.650 82.140 95.755 83.650 ;
        RECT 119.945 83.240 120.955 83.265 ;
        RECT 113.270 82.280 120.955 83.240 ;
        RECT 119.945 82.255 120.955 82.280 ;
        RECT 26.650 81.965 65.690 82.140 ;
        RECT 26.890 81.550 31.040 81.965 ;
        RECT 27.090 66.710 31.400 67.120 ;
        RECT 26.610 65.070 61.300 66.710 ;
        RECT 27.090 64.630 31.400 65.070 ;
        RECT 77.430 63.890 87.550 64.370 ;
        RECT 68.420 61.855 69.940 61.885 ;
        RECT 68.420 60.875 90.220 61.855 ;
        RECT 68.420 59.705 69.940 60.875 ;
        RECT 76.410 58.930 76.960 58.970 ;
        RECT 76.410 58.450 87.560 58.930 ;
        RECT 76.410 58.360 76.960 58.450 ;
        RECT 89.240 57.585 90.220 60.875 ;
        RECT 139.680 58.920 141.370 61.850 ;
        RECT 139.680 58.695 154.180 58.920 ;
        RECT 94.145 57.585 95.795 58.200 ;
        RECT 101.200 57.585 102.400 58.305 ;
        RECT 106.750 57.585 154.180 58.695 ;
        RECT 89.240 57.115 154.180 57.585 ;
        RECT 89.240 56.605 108.170 57.115 ;
        RECT 89.240 56.275 90.220 56.605 ;
        RECT 94.145 56.550 95.795 56.605 ;
        RECT 101.200 56.495 102.400 56.605 ;
        RECT 106.750 56.520 108.170 56.605 ;
        RECT 86.455 56.210 90.220 56.275 ;
        RECT 77.440 55.730 90.220 56.210 ;
        RECT 106.750 56.190 108.360 56.520 ;
        RECT 106.750 55.945 108.170 56.190 ;
        RECT 86.455 55.425 90.220 55.730 ;
        RECT 26.900 53.635 31.250 53.840 ;
        RECT 26.575 53.360 63.810 53.635 ;
        RECT 76.445 53.360 76.975 53.385 ;
        RECT 26.575 52.880 76.975 53.360 ;
        RECT 26.575 52.605 63.810 52.880 ;
        RECT 76.445 52.855 76.975 52.880 ;
        RECT 26.900 52.310 31.250 52.605 ;
        RECT 81.770 51.870 82.310 52.050 ;
        RECT 82.815 51.870 83.315 51.910 ;
        RECT 81.770 51.380 83.315 51.870 ;
        RECT 81.770 47.970 82.310 51.380 ;
        RECT 82.815 51.340 83.315 51.380 ;
        RECT 82.695 50.690 83.195 50.770 ;
        RECT 85.395 50.690 85.895 50.730 ;
        RECT 82.610 50.240 85.895 50.690 ;
        RECT 82.695 50.110 83.195 50.240 ;
        RECT 85.395 50.070 85.895 50.240 ;
        RECT 85.375 47.970 85.875 48.000 ;
        RECT 86.465 47.970 87.315 55.425 ;
        RECT 89.240 55.405 90.220 55.425 ;
        RECT 113.360 55.145 115.040 57.115 ;
        RECT 120.010 56.520 121.590 57.115 ;
        RECT 126.610 56.520 128.190 57.115 ;
        RECT 133.200 56.520 134.780 57.115 ;
        RECT 139.680 56.900 154.180 57.115 ;
        RECT 139.680 56.665 141.370 56.900 ;
        RECT 119.980 56.190 121.590 56.520 ;
        RECT 126.580 56.190 128.190 56.520 ;
        RECT 133.180 56.190 134.780 56.520 ;
        RECT 120.010 55.255 121.590 56.190 ;
        RECT 126.610 55.325 128.190 56.190 ;
        RECT 133.200 55.365 134.780 56.190 ;
        RECT 139.780 55.395 141.360 56.665 ;
        RECT 103.480 53.470 105.060 53.800 ;
        RECT 110.080 53.470 111.660 53.800 ;
        RECT 116.680 53.470 118.260 53.800 ;
        RECT 123.280 53.470 124.860 53.800 ;
        RECT 129.880 53.470 131.460 53.800 ;
        RECT 136.480 53.470 138.060 53.800 ;
        RECT 106.780 50.750 108.360 51.080 ;
        RECT 113.380 50.750 114.960 51.080 ;
        RECT 119.980 50.750 121.560 51.080 ;
        RECT 126.580 50.750 128.160 51.080 ;
        RECT 133.180 50.750 134.760 51.080 ;
        RECT 139.780 49.620 153.990 51.890 ;
        RECT 103.480 48.030 105.060 48.360 ;
        RECT 110.080 48.030 111.660 48.360 ;
        RECT 116.680 48.030 118.260 48.360 ;
        RECT 123.280 48.030 124.860 48.360 ;
        RECT 129.880 48.030 131.460 48.360 ;
        RECT 136.480 48.030 138.060 48.360 ;
        RECT 81.770 47.120 87.315 47.970 ;
        RECT 81.770 46.490 82.310 47.120 ;
        RECT 82.795 46.490 83.295 46.530 ;
        RECT 81.770 46.000 83.295 46.490 ;
        RECT 81.770 41.130 82.310 46.000 ;
        RECT 82.795 45.960 83.295 46.000 ;
        RECT 85.180 45.700 86.180 46.700 ;
        RECT 82.795 45.330 83.335 45.380 ;
        RECT 85.385 45.330 85.925 45.370 ;
        RECT 82.670 44.830 85.925 45.330 ;
        RECT 106.780 45.310 108.360 45.640 ;
        RECT 113.380 45.310 114.960 45.640 ;
        RECT 119.980 45.310 121.560 45.640 ;
        RECT 126.580 45.310 128.160 45.640 ;
        RECT 133.180 45.310 134.760 45.640 ;
        RECT 139.780 45.310 141.360 45.640 ;
        RECT 82.795 44.810 83.335 44.830 ;
        RECT 85.385 44.800 85.925 44.830 ;
        RECT 103.480 42.590 105.060 42.920 ;
        RECT 110.080 42.590 111.660 42.920 ;
        RECT 116.680 42.590 118.260 42.920 ;
        RECT 123.280 42.590 124.860 42.920 ;
        RECT 129.880 42.590 131.460 42.920 ;
        RECT 136.480 42.590 138.060 42.920 ;
        RECT 82.765 41.130 83.265 41.170 ;
        RECT 81.770 40.640 83.270 41.130 ;
        RECT 81.770 35.780 82.310 40.640 ;
        RECT 82.765 40.600 83.265 40.640 ;
        RECT 85.160 40.480 86.160 41.480 ;
        RECT 82.755 40.020 83.295 40.060 ;
        RECT 85.375 40.020 85.915 40.060 ;
        RECT 82.690 39.480 85.930 40.020 ;
        RECT 106.780 39.870 108.360 40.200 ;
        RECT 113.380 39.870 114.960 40.200 ;
        RECT 119.980 39.870 121.560 40.200 ;
        RECT 126.580 39.870 128.160 40.200 ;
        RECT 133.180 39.870 134.760 40.200 ;
        RECT 139.780 39.870 141.360 40.200 ;
        RECT 82.755 39.440 83.295 39.480 ;
        RECT 85.375 39.440 85.915 39.480 ;
        RECT 103.480 37.150 105.060 37.480 ;
        RECT 110.080 37.150 111.660 37.480 ;
        RECT 116.680 37.150 118.260 37.480 ;
        RECT 123.280 37.150 124.860 37.480 ;
        RECT 129.880 37.150 131.460 37.480 ;
        RECT 136.480 37.150 138.060 37.480 ;
        RECT 82.795 35.780 83.295 35.810 ;
        RECT 81.770 35.290 83.295 35.780 ;
        RECT 85.230 35.330 86.230 36.330 ;
        RECT 81.770 35.220 82.310 35.290 ;
        RECT 82.795 35.240 83.295 35.290 ;
        RECT 82.715 34.840 83.365 34.860 ;
        RECT 82.590 34.820 86.040 34.840 ;
        RECT 82.590 34.250 86.055 34.820 ;
        RECT 106.780 34.430 108.360 34.760 ;
        RECT 113.380 34.430 114.960 34.760 ;
        RECT 119.980 34.430 121.560 34.760 ;
        RECT 126.580 34.430 128.160 34.760 ;
        RECT 133.180 34.430 134.760 34.760 ;
        RECT 82.590 34.240 86.040 34.250 ;
        RECT 139.730 33.600 153.940 35.870 ;
        RECT 103.480 31.710 105.060 32.040 ;
        RECT 110.080 31.710 111.660 32.040 ;
        RECT 116.680 31.710 118.260 32.040 ;
        RECT 123.280 31.710 124.860 32.040 ;
        RECT 129.880 31.710 131.460 32.040 ;
        RECT 136.480 31.710 138.060 32.040 ;
        RECT 106.780 28.990 108.360 29.320 ;
        RECT 113.380 28.990 114.960 29.320 ;
        RECT 119.980 28.990 121.560 29.320 ;
        RECT 126.580 28.990 128.160 29.320 ;
        RECT 133.180 28.990 134.760 29.320 ;
        RECT 139.780 28.990 141.360 29.320 ;
        RECT 120.355 27.605 120.685 27.620 ;
        RECT 124.955 27.605 125.285 27.620 ;
        RECT 120.355 27.305 125.285 27.605 ;
        RECT 120.355 27.290 120.685 27.305 ;
        RECT 124.955 27.290 125.285 27.305 ;
        RECT 103.480 26.270 105.060 26.600 ;
        RECT 110.080 26.270 111.660 26.600 ;
        RECT 116.680 26.270 118.260 26.600 ;
        RECT 123.280 26.270 124.860 26.600 ;
        RECT 129.880 26.270 131.460 26.600 ;
        RECT 136.480 26.270 138.060 26.600 ;
        RECT 106.780 23.550 108.360 23.880 ;
        RECT 113.380 23.550 114.960 23.880 ;
        RECT 119.980 23.550 121.560 23.880 ;
        RECT 126.580 23.550 128.160 23.880 ;
        RECT 133.180 23.550 134.760 23.880 ;
        RECT 139.750 22.470 153.960 24.740 ;
        RECT 103.460 21.160 105.040 21.245 ;
        RECT 110.060 21.160 111.640 21.235 ;
        RECT 116.660 21.160 118.240 21.225 ;
        RECT 123.270 21.160 124.850 21.235 ;
        RECT 129.810 21.160 131.390 21.305 ;
        RECT 136.520 21.160 138.100 21.305 ;
        RECT 103.460 20.830 105.060 21.160 ;
        RECT 110.060 20.830 111.660 21.160 ;
        RECT 116.660 20.830 118.260 21.160 ;
        RECT 123.270 20.830 124.860 21.160 ;
        RECT 129.810 20.830 131.460 21.160 ;
        RECT 136.480 20.830 138.100 21.160 ;
        RECT 26.740 18.100 31.370 18.280 ;
        RECT 103.460 18.100 105.040 20.830 ;
        RECT 106.780 18.110 108.360 18.440 ;
        RECT 26.640 17.725 105.040 18.100 ;
        RECT 110.060 17.725 111.640 20.830 ;
        RECT 113.380 18.110 114.960 18.440 ;
        RECT 116.660 17.725 118.240 20.830 ;
        RECT 119.980 18.110 121.560 18.440 ;
        RECT 123.270 17.725 124.850 20.830 ;
        RECT 126.580 18.110 128.160 18.440 ;
        RECT 129.810 17.725 131.390 20.830 ;
        RECT 133.180 18.110 134.760 18.440 ;
        RECT 136.520 17.725 138.100 20.830 ;
        RECT 139.780 18.110 141.360 18.440 ;
        RECT 26.640 16.145 138.100 17.725 ;
        RECT 26.640 15.590 104.505 16.145 ;
        RECT 26.740 15.270 31.370 15.590 ;
        RECT 93.780 0.790 94.820 2.510 ;
        RECT 113.065 0.985 114.175 2.875 ;
        RECT 132.390 0.790 133.495 2.720 ;
        RECT 151.645 1.235 152.875 3.525 ;
      LAYER met4 ;
        RECT 124.810 224.760 124.815 225.235 ;
        RECT 30.670 222.660 30.970 224.760 ;
        RECT 33.430 222.660 33.730 224.760 ;
        RECT 36.190 222.660 36.490 224.760 ;
        RECT 38.950 222.660 39.250 224.760 ;
        RECT 41.710 222.660 42.010 224.760 ;
        RECT 44.470 222.660 44.770 224.760 ;
        RECT 47.230 222.660 47.530 224.760 ;
        RECT 49.990 222.660 50.290 224.760 ;
        RECT 52.750 222.660 53.050 224.760 ;
        RECT 55.510 222.660 55.810 224.760 ;
        RECT 58.270 222.660 58.570 224.760 ;
        RECT 61.030 222.660 61.330 224.760 ;
        RECT 63.790 222.660 64.090 224.760 ;
        RECT 66.550 222.660 66.850 224.760 ;
        RECT 69.310 222.660 69.610 224.760 ;
        RECT 72.070 222.660 72.370 224.760 ;
        RECT 74.830 222.660 75.130 224.760 ;
        RECT 77.590 222.660 77.890 224.760 ;
        RECT 80.350 222.660 80.650 224.760 ;
        RECT 83.110 222.660 83.410 224.760 ;
        RECT 85.870 222.660 86.170 224.760 ;
        RECT 88.630 222.660 88.930 224.760 ;
        RECT 91.390 222.660 91.690 224.760 ;
        RECT 94.150 222.660 94.450 224.760 ;
        RECT 113.470 224.680 113.770 224.760 ;
        RECT 116.230 224.680 116.530 224.760 ;
        RECT 121.750 224.755 122.050 224.760 ;
        RECT 121.670 223.710 122.135 224.755 ;
        RECT 124.510 224.460 124.815 224.760 ;
        RECT 127.270 224.525 127.570 224.760 ;
        RECT 130.030 224.585 130.330 224.760 ;
        RECT 132.790 224.585 133.090 224.760 ;
        RECT 135.550 224.595 135.850 224.760 ;
        RECT 138.310 224.595 138.610 224.760 ;
        RECT 124.450 224.030 124.880 224.460 ;
        RECT 127.255 224.195 127.585 224.525 ;
        RECT 130.015 224.255 130.345 224.585 ;
        RECT 132.775 224.255 133.105 224.585 ;
        RECT 135.535 224.265 135.865 224.595 ;
        RECT 138.295 224.265 138.625 224.595 ;
        RECT 30.530 222.340 154.130 222.660 ;
        RECT 30.530 219.560 148.900 222.340 ;
        RECT 153.990 220.880 154.130 222.340 ;
        RECT 26.400 216.500 31.730 216.690 ;
        RECT 31.500 3.740 31.730 216.500 ;
        RECT 121.520 215.860 122.505 216.845 ;
        RECT 121.525 213.095 122.500 215.860 ;
        RECT 119.185 207.845 120.595 209.255 ;
        RECT 119.190 203.750 120.590 207.845 ;
        RECT 88.075 160.230 89.230 162.360 ;
        RECT 88.075 158.020 89.855 160.230 ;
        RECT 88.075 156.865 89.885 158.020 ;
        RECT 88.100 156.860 89.855 156.865 ;
        RECT 88.975 155.525 89.855 156.860 ;
        RECT 88.970 154.635 89.860 155.525 ;
        RECT 64.060 153.790 64.515 154.245 ;
        RECT 64.070 150.790 64.515 153.790 ;
        RECT 68.210 152.815 68.600 153.205 ;
        RECT 64.015 149.915 64.575 150.790 ;
        RECT 68.215 150.755 68.595 152.815 ;
        RECT 69.610 151.945 70.120 154.235 ;
        RECT 69.605 151.425 70.125 151.945 ;
        RECT 68.180 150.065 68.750 150.755 ;
        RECT 102.185 148.055 103.125 157.240 ;
        RECT 102.180 147.105 103.130 148.055 ;
        RECT 89.940 100.395 91.320 107.870 ;
        RECT 89.925 97.845 91.355 100.395 ;
        RECT 89.940 97.710 91.320 97.845 ;
        RECT 106.750 57.115 141.360 58.695 ;
        RECT 106.750 56.795 108.690 57.115 ;
        RECT 103.450 18.155 105.070 56.595 ;
        RECT 106.750 56.515 108.390 56.795 ;
        RECT 103.460 18.035 105.070 18.155 ;
        RECT 106.770 18.485 108.390 56.515 ;
        RECT 110.070 20.835 111.670 56.595 ;
        RECT 113.360 56.515 115.040 57.115 ;
        RECT 116.770 56.595 118.170 56.735 ;
        RECT 120.100 56.595 121.500 57.115 ;
        RECT 123.390 56.595 124.790 56.775 ;
        RECT 126.610 56.595 128.190 57.115 ;
        RECT 133.200 56.595 134.780 57.115 ;
        RECT 136.550 56.595 137.950 56.715 ;
        RECT 139.780 56.595 141.360 57.115 ;
        RECT 106.770 18.035 108.370 18.485 ;
        RECT 110.060 18.035 111.670 20.835 ;
        RECT 113.370 18.035 114.970 56.515 ;
        RECT 116.670 20.835 118.270 56.595 ;
        RECT 116.660 18.035 118.270 20.835 ;
        RECT 119.970 18.035 121.570 56.595 ;
        RECT 123.270 18.035 124.870 56.595 ;
        RECT 126.570 56.515 128.190 56.595 ;
        RECT 126.570 18.035 128.170 56.515 ;
        RECT 129.870 20.835 131.470 56.595 ;
        RECT 129.810 18.035 131.470 20.835 ;
        RECT 133.170 56.515 134.780 56.595 ;
        RECT 133.170 18.035 134.770 56.515 ;
        RECT 136.470 20.835 138.070 56.595 ;
        RECT 136.470 18.035 138.100 20.835 ;
        RECT 139.770 18.035 141.370 56.595 ;
        RECT 103.460 17.725 105.040 18.035 ;
        RECT 110.060 17.725 111.640 18.035 ;
        RECT 116.660 17.725 118.240 18.035 ;
        RECT 123.270 17.725 124.850 18.035 ;
        RECT 129.810 17.725 131.390 18.035 ;
        RECT 136.520 17.725 138.100 18.035 ;
        RECT 103.420 16.145 138.100 17.725 ;
        RECT 153.990 7.040 154.230 220.880 ;
        RECT 93.850 1.000 94.750 1.760 ;
        RECT 113.170 1.000 114.070 1.990 ;
        RECT 132.490 1.000 133.390 1.790 ;
        RECT 151.810 1.000 152.710 2.300 ;
  END
END tt_um_patdeegan_anamux
END LIBRARY

