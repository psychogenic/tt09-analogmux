* NGSPICE file created from muxtest_parax.ext - technology: sky130A

.subckt muxtest_parax SELECT0 RSEL2 VRES LADDEROUT RSEL1 RSEL0 SELECT1 OUT VDD VSS
X0 R7R8.t3 R6R7.t1 VSS.t50 sky130_fd_pr__res_high_po_1p41 l=1.75
X1 R4R5.t3 x1.x3.GP4.t4 x1.x5.A.t4 VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X2 R1R2.t0 VRES.t0 VSS.t11 sky130_fd_pr__res_high_po_1p41 l=1.75
X3 x1.x4.A x1.x3.GN1.t2 R3R4.t1 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X4 VSS.t106 VDD.t152 VSS.t105 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X5 a_13269_n10181# SELECT0.t0 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X6 x1.x5.A.t11 RSEL2.t0 LADDEROUT.t9 VDD.t74 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X7 a_13269_n10869# a_13269_n10693# a_13295_n10741# VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X8 a_4962_n3364# RSEL1.t0 a_5016_n3226# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X9 x1.x5.A.t1 x1.x3.GN4.t2 R4R5.t0 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X10 R7R8.t7 x2.x2.GP4.t4 OUT.t13 VDD.t84 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X11 VSS.t97 x1.x3.GN3 x1.x3.GP3 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X12 VSS.t85 x2.x2.GN1.t2 x2.x2.GP1.t1 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X13 VSS.t3 RSEL1.t1 x1.x1.nSEL1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X14 a_13295_n11293# SELECT0.t1 VSS.t103 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X15 VSS.t113 a_13269_n11421# x2.x2.GN2 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X16 VDD.t129 x2.x2.GN4.t2 x2.x2.GP4.t1 VDD.t128 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X17 x1.x5.A.t2 x1.x3.GN4.t3 R4R5.t1 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X18 VSS.t137 RSEL0.t0 x1.x1.nSEL0 VSS.t136 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X19 x1.x3.GP1.t1 x1.x3.GN1.t3 VSS.t123 VSS.t122 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X20 VSS.t63 x1.x3.GN2 x1.x3.GP2.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X21 VRES.t6 x2.x2.GP2.t4 OUT.t6 VDD.t101 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X22 VSS.t70 RSEL0.t1 a_4962_n3876# VSS.t69 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X23 R1R2.t5 x1.x3.GP3 x1.x4.A VDD.t134 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X24 a_4962_n4052# a_4962_n3876# a_4988_n3924# VSS.t144 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X25 VSS.t24 x1.x3.GN1.t4 x1.x3.GP1.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X26 x1.x5.A.t15 x1.x3.GN3 R5R6.t1 VSS.t92 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X27 a_4962_n5020# x1.x1.nSEL1 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X28 LADDEROUT.t11 RSEL2.t1 x1.x4.A VSS.t79 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X29 VRES.t2 x1.x3.GP4.t5 x1.x4.A VDD.t33 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X30 a_4962_n4604# RSEL0.t2 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X31 a_4988_n4476# RSEL0.t3 VSS.t72 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X32 VSS.t27 a_4962_n4604# x1.x3.GN2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X33 VDD.t149 x1.x1.nSEL0 a_4962_n5020# VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X34 VSS.t14 a_13269_n10181# x2.x2.GN4.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X35 VDD.t23 VSS.t153 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X36 x1.x5.A.t9 x1.x3.GN2 R6R7.t3 VSS.t61 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X37 R2R3.t4 x1.x3.GP2.t4 x1.x4.A VDD.t35 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X38 R5R6.t4 x1.x3.GP3 x1.x5.A.t18 VDD.t135 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X39 OUT.t15 x2.x2.GN3 R3R4.t8 VSS.t151 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X40 x2.nselect2 VDD.t80 VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X41 R7R8.t8 x1.x3.GP1.t4 x1.x5.A.t16 VDD.t32 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X42 VSS.t75 VDD.t153 VSS.t74 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X43 x2.x1.nSEL0 SELECT0.t2 VSS.t130 VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X44 VSS.t140 SELECT1.t0 x2.x1.nSEL1 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X45 x1.x1.nSEL0 RSEL0.t4 VSS.t134 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X46 x1.x5.A.t5 x1.x3.GN1.t5 R7R8.t2 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X47 VSS.t78 VDD.t154 VSS.t77 VSS.t76 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X48 x1.x3.GP4.t3 x1.x3.GN4.t4 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X49 VDD.t20 VSS.t154 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X50 a_13269_n11837# x2.x1.nSEL0 a_13323_n11699# VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X51 x2.x2.GP4.t0 x2.x2.GN4.t3 VSS.t115 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X52 x1.x4.A x1.x3.GN4.t5 VRES.t5 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X53 VSS.t47 a_4962_n3364# x1.x3.GN4.t0 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X54 x1.x5.GN RSEL2.t2 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X55 VSS.t132 SELECT0.t3 x2.x1.nSEL0 VSS.t131 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X56 x2.x2.GP3 x2.x2.GN3 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X57 VDD.t116 a_13269_n11421# x2.x2.GN2 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X58 x1.x3.GP3 x1.x3.GN3 VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X59 VDD.t61 x1.x3.GN4.t6 x1.x3.GP4.t0 VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X60 x1.x1.nSEL1 RSEL1.t2 VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X61 LADDEROUT.t1 x2.x2.GP1.t4 OUT.t2 VDD.t83 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X62 VDD.t73 RSEL2.t3 x1.x5.GN VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X63 VSS.t32 VDD.t155 VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X64 x1.x4.A x1.x3.GN3 R1R2.t3 VSS.t95 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X65 x1.x5.A.t7 RSEL2.t4 LADDEROUT.t8 VDD.t55 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X66 VSS.t99 a_13269_n10869# x2.x2.GN3 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X67 a_13269_n10869# SELECT1.t1 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X68 a_5016_n4882# x1.x1.nSEL1 VSS.t111 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X69 VDD.t17 VSS.t155 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X70 x2.x2.GP2.t3 x2.x2.GN2 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X71 x1.x3.GP2.t3 x1.x3.GN2 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X72 VDD.t14 VSS.t156 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X73 a_13269_n11837# x2.x1.nSEL1 VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X74 VSS.t146 x2.x2.GN4.t4 x2.x2.GP4.t2 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X75 x2.x2.GP1.t3 x2.x2.GN1.t3 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X76 VDD.t11 VSS.t157 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X77 a_4962_n5020# x1.x1.nSEL0 a_5016_n4882# VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X78 R3R4.t9 x1.x3.GP1.t5 x1.x4.A VDD.t142 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X79 VDD.t124 x2.x2.GN2 x2.x2.GP2.t2 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X80 R4R5.t4 R3R4.t5 VSS.t141 sky130_fd_pr__res_high_po_1p41 l=1.75
X81 VDD.t139 a_4962_n5020# x1.x3.GN1.t1 VDD.t138 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X82 VSS.t9 SELECT1.t2 a_13269_n11245# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X83 a_4962_n3876# RSEL0.t5 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X84 VSS.t35 VDD.t156 VSS.t34 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X85 a_13269_n11421# a_13269_n11245# a_13295_n11293# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X86 a_13269_n11245# SELECT1.t3 VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X87 VSS.t108 R7R8.t6 VSS.t107 sky130_fd_pr__res_high_po_1p41 l=1.75
X88 VDD.t141 a_4962_n3876# a_4962_n4052# VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X89 OUT.t9 x2.x2.GN2 VRES.t8 VSS.t126 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X90 VDD.t37 a_13269_n10181# x2.x2.GN4.t1 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X91 VDD.t88 a_13269_n11245# a_13269_n11421# VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X92 a_4962_n3364# RSEL0.t6 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X93 x1.x5.A.t8 x1.x3.GN2 R6R7.t2 VSS.t61 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X94 OUT.t14 x2.x2.GN3 R3R4.t7 VSS.t151 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X95 R2R3.t3 x1.x3.GP2.t5 x1.x4.A VDD.t35 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X96 LADDEROUT.t10 RSEL2.t5 x1.x4.A VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X97 VDD.t43 a_4962_n4052# x1.x3.GN3 VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X98 R5R6.t3 x1.x3.GP3 x1.x5.A.t17 VDD.t135 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X99 R7R8.t4 x2.x2.GP4.t5 OUT.t12 VDD.t84 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X100 OUT.t4 x2.x2.GN4.t5 R7R8.t5 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X101 VSS.t19 VDD.t157 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X102 LADDEROUT.t3 x1.x5.GN x1.x5.A.t13 VSS.t89 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X103 VSS.t40 RSEL1.t3 a_4962_n4428# VSS.t39 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X104 R3R4.t2 x2.x2.GP3 OUT.t11 VDD.t127 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X105 VSS.t22 VDD.t158 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X106 R1R2.t4 x1.x3.GP3 x1.x4.A VDD.t134 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X107 a_4962_n4604# a_4962_n4428# a_4988_n4476# VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X108 x1.x5.A.t19 x1.x3.GN1.t6 R7R8.t9 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X109 x1.x4.A x1.x3.GN4.t7 VRES.t3 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X110 x2.nselect2 VDD.t159 VSS.t65 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X111 VSS.t91 a_13269_n11837# x2.x2.GN1.t0 VSS.t90 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X112 VDD.t79 VDD.t77 x2.nselect2 VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X113 a_13323_n10043# SELECT0.t4 VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X114 x1.x4.A x1.x3.GN3 R1R2.t2 VSS.t95 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X115 VDD.t98 a_13269_n10869# x2.x2.GN3 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X116 R6R7.t0 x1.x3.GP2.t6 x1.x5.A.t6 VDD.t44 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X117 VRES.t4 x2.x2.GP2.t5 OUT.t3 VDD.t101 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X118 x2.x1.nSEL1 SELECT1.t4 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X119 x2.x2.GP3 x2.x2.GN3 VSS.t150 VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X120 VDD.t8 VSS.t158 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X121 VDD.t145 x2.x2.GN3 x2.x2.GP3 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X122 x1.x4.A x1.x3.GN2 R2R3.t2 VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X123 a_13295_n10741# SELECT1.t5 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X124 R6R7.t5 R5R6.t2 VSS.t109 sky130_fd_pr__res_high_po_1p41 l=1.75
X125 VDD.t94 x1.x3.GN3 x1.x3.GP3 VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X126 VDD.t144 RSEL1.t4 x1.x1.nSEL1 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X127 x1.x3.GP4.t1 x1.x3.GN4.t8 VSS.t81 VSS.t80 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X128 x1.x5.GN RSEL2.t6 VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X129 R3R4.t6 x1.x3.GP1.t6 x1.x4.A VDD.t142 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X130 x2.x2.GP2.t1 x2.x2.GN2 VSS.t128 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X131 R7R8.t1 x1.x3.GP1.t7 x1.x5.A.t0 VDD.t32 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X132 a_5016_n3226# RSEL0.t7 VSS.t49 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X133 x1.x4.A x1.x3.GN2 R2R3.t1 VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X134 R5R6.t5 R4R5.t5 VSS.t50 sky130_fd_pr__res_high_po_1p41 l=1.75
X135 VDD.t133 RSEL0.t8 x1.x1.nSEL0 VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X136 OUT.t8 x2.x2.GN2 VRES.t7 VSS.t126 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X137 x1.x3.GP3 x1.x3.GN3 VSS.t94 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X138 x2.x2.GP1.t0 x2.x2.GN1.t4 VSS.t117 VSS.t116 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X139 VSS.t83 x1.x3.GN4.t9 x1.x3.GP4.t2 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X140 VSS.t57 RSEL2.t7 x1.x5.GN VSS.t56 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X141 VDD.t65 x1.x3.GN2 x1.x3.GP2.t2 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X142 x1.x1.nSEL1 RSEL1.t5 VSS.t38 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X143 x1.x3.GP1.t3 x1.x3.GN1.t7 VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X144 R3R4.t3 x2.x2.GP3 OUT.t10 VDD.t127 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X145 VSS.t125 x2.x2.GN2 x2.x2.GP2.t0 VSS.t124 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X146 VSS.t143 a_4962_n5020# x1.x3.GN1.t0 VSS.t142 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X147 R4R5.t2 x1.x3.GP4.t6 x1.x5.A.t3 VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X148 VDD.t29 x2.x1.nSEL0 a_13269_n11837# VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X149 VDD.t52 x2.x2.GN1.t5 x2.x2.GP1.t2 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X150 a_4988_n3924# RSEL1.t6 VSS.t101 VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X151 VDD.t27 x1.x3.GN1.t8 x1.x3.GP1.t2 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X152 x1.x4.A x1.x3.GN1.t9 R3R4.t0 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X153 a_4962_n4052# RSEL1.t7 VDD.t102 VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X154 x1.x3.GP2.t0 x1.x3.GN2 VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X155 OUT.t0 x2.x2.GN4.t6 R7R8.t0 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X156 a_13269_n11421# SELECT0.t5 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X157 VSS.t42 SELECT0.t6 a_13269_n10693# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X158 a_13269_n10693# SELECT0.t7 VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X159 VDD.t131 a_13269_n10693# a_13269_n10869# VDD.t130 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X160 VDD.t112 RSEL1.t8 a_4962_n3364# VDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X161 a_13269_n10181# SELECT1.t6 a_13323_n10043# VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X162 VSS.t68 VDD.t160 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X163 VSS.t29 a_4962_n4052# x1.x3.GN3 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X164 VDD.t92 a_13269_n11837# x2.x2.GN1.t1 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X165 a_4962_n4428# RSEL1.t9 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X166 LADDEROUT.t6 x2.x2.GP1.t5 OUT.t5 VDD.t83 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X167 VDD.t114 SELECT1.t7 a_13269_n10181# VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X168 VDD.t86 a_4962_n4428# a_4962_n4604# VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X169 VDD.t41 a_4962_n4604# x1.x3.GN2 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X170 x1.x5.A.t14 x1.x3.GN3 R5R6.t0 VSS.t92 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X171 VDD.t5 VSS.t159 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X172 VRES.t1 x1.x3.GP4.t7 x1.x4.A VDD.t33 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X173 R3R4.t4 R2R3.t5 VSS.t138 sky130_fd_pr__res_high_po_1p41 l=1.75
X174 R6R7.t4 x1.x3.GP2.t7 x1.x5.A.t10 VDD.t44 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X175 VSS.t53 VDD.t161 x2.nselect2 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X176 x1.x1.nSEL0 RSEL0.t9 VDD.t76 VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X177 VDD.t2 VSS.t160 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X178 OUT.t7 x2.x2.GN1.t6 LADDEROUT.t7 VSS.t119 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X179 LADDEROUT.t2 x1.x5.GN x1.x5.A.t12 VSS.t88 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X180 x2.x1.nSEL1 SELECT1.t8 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X181 x1.x4.A x1.x5.GN LADDEROUT.t5 VDD.t90 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X182 x2.x1.nSEL0 SELECT0.t8 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X183 a_13323_n11699# x2.x1.nSEL1 VSS.t121 VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X184 VDD.t120 SELECT1.t9 x2.x1.nSEL1 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X185 VSS.t148 x2.x2.GN3 x2.x2.GP3 VSS.t147 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X186 x1.x4.A x1.x5.GN LADDEROUT.t4 VDD.t89 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X187 OUT.t1 x2.x2.GN1.t7 LADDEROUT.t0 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X188 R2R3.t0 R1R2.t1 VSS.t43 sky130_fd_pr__res_high_po_1p41 l=1.75
X189 x2.x2.GP4.t3 x2.x2.GN4.t7 VDD.t151 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X190 VDD.t57 a_4962_n3364# x1.x3.GN4.t1 VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X191 VDD.t48 SELECT0.t9 x2.x1.nSEL0 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
R0 R7R8.n6 R7R8.t4 26.3998
R1 R7R8.n1 R7R8.t1 26.3998
R2 R7R8.n6 R7R8.t7 23.5483
R3 R7R8.n1 R7R8.t8 23.5483
R4 R7R8.n5 R7R8.t0 12.7127
R5 R7R8.n0 R7R8.t9 12.7127
R6 R7R8.n5 R7R8.t5 10.8578
R7 R7R8.n0 R7R8.t2 10.8578
R8 R7R8.n4 R7R8.t6 10.7774
R9 R7R8.n4 R7R8.t3 10.6159
R10 R7R8.n9 R7R8 8.70294
R11 R7R8.n7 R7R8.n6 3.12177
R12 R7R8.n2 R7R8.n1 3.12177
R13 R7R8.n7 R7R8.n5 1.81453
R14 R7R8.n2 R7R8.n0 1.81453
R15 R7R8.n8 R7R8.n7 1.1255
R16 R7R8.n3 R7R8.n2 1.1255
R17 R7R8.n10 R7R8 1.11113
R18 R7R8.n10 R7R8.n9 0.427375
R19 R7R8.n9 R7R8.n4 0.230945
R20 R7R8 R7R8.n3 0.148615
R21 R7R8 R7R8.n8 0.134513
R22 R7R8.n8 R7R8 0.0655
R23 R7R8.n3 R7R8 0.0655
R24 R7R8 R7R8.n10 0.008625
R25 R6R7.n2 R6R7.t0 26.3998
R26 R6R7.n2 R6R7.t4 23.5483
R27 R6R7.n0 R6R7.t5 17.5523
R28 R6R7.n1 R6R7.t2 12.7127
R29 R6R7.n1 R6R7.t3 10.8578
R30 R6R7.n0 R6R7.t1 10.5295
R31 R6R7.n3 R6R7.n2 3.12177
R32 R6R7.n3 R6R7.n1 1.81453
R33 R6R7.n4 R6R7.n3 1.1255
R34 R6R7 R6R7.n0 0.411443
R35 R6R7 R6R7.n4 0.138152
R36 R6R7.n4 R6R7 0.0655
R37 VSS.n173 VSS.n171 3.3198e+06
R38 VSS.n442 VSS.n441 2.3452e+06
R39 VSS.n173 VSS.n172 2.3386e+06
R40 VSS.n172 VSS.n47 2.1428e+06
R41 VSS.n398 VSS.n154 1.2298e+06
R42 VSS.n381 VSS.n367 1.19185e+06
R43 VSS.n441 VSS.t23 1.17724e+06
R44 VSS.n172 VSS.t114 1.17707e+06
R45 VSS.n397 VSS.n396 1.177e+06
R46 VSS.n398 VSS.n397 1.177e+06
R47 VSS.n465 VSS.n154 1.177e+06
R48 VSS.n171 VSS.n33 392333
R49 VSS.n382 VSS.n381 392333
R50 VSS.n441 VSS.n422 392333
R51 VSS.n171 VSS.n40 387200
R52 VSS.n396 VSS.n382 387200
R53 VSS.n441 VSS.n433 387200
R54 VSS.n173 VSS.n170 331554
R55 VSS.n367 VSS.n366 297447
R56 VSS.n304 VSS.n14 28658
R57 VSS.n466 VSS.n465 16580.8
R58 VSS.n462 VSS.n417 11744.7
R59 VSS.n458 VSS.n417 11744.7
R60 VSS.n462 VSS.n418 11744.7
R61 VSS.n458 VSS.n418 11744.7
R62 VSS.n416 VSS.n155 11744.7
R63 VSS.n412 VSS.n156 11744.7
R64 VSS.n416 VSS.n156 11744.7
R65 VSS.n400 VSS.n399 11744.7
R66 VSS.n163 VSS.n162 11744.7
R67 VSS.n399 VSS.n163 11744.7
R68 VSS.n169 VSS.n31 11744.7
R69 VSS.n536 VSS.n31 11744.7
R70 VSS.n169 VSS.n32 11744.7
R71 VSS.n536 VSS.n32 11744.7
R72 VSS.n533 VSS.n34 11744.7
R73 VSS.n529 VSS.n34 11744.7
R74 VSS.n533 VSS.n35 11744.7
R75 VSS.n529 VSS.n35 11744.7
R76 VSS.n526 VSS.n41 11744.7
R77 VSS.n522 VSS.n41 11744.7
R78 VSS.n526 VSS.n42 11744.7
R79 VSS.n522 VSS.n42 11744.7
R80 VSS.n512 VSS.n48 11744.7
R81 VSS.n512 VSS.n49 11744.7
R82 VSS.n519 VSS.n48 11744.7
R83 VSS.n519 VSS.n49 11744.7
R84 VSS.n473 VSS.n16 11744.7
R85 VSS.n556 VSS.n16 11744.7
R86 VSS.n473 VSS.n17 11744.7
R87 VSS.n556 VSS.n17 11744.7
R88 VSS.n567 VSS.n9 11744.7
R89 VSS.n562 VSS.n9 11744.7
R90 VSS.n562 VSS.n8 11744.7
R91 VSS.n567 VSS.n8 11744.7
R92 VSS.n455 VSS.n423 11744.7
R93 VSS.n451 VSS.n423 11744.7
R94 VSS.n455 VSS.n424 11744.7
R95 VSS.n451 VSS.n424 11744.7
R96 VSS.n444 VSS.n434 11744.7
R97 VSS.n444 VSS.n435 11744.7
R98 VSS.n448 VSS.n435 11744.7
R99 VSS.n448 VSS.n434 11744.7
R100 VSS.n151 VSS.n140 11744.7
R101 VSS.n146 VSS.n140 11744.7
R102 VSS.n151 VSS.n142 11744.7
R103 VSS.n146 VSS.n142 11744.7
R104 VSS.n380 VSS.n368 11744.7
R105 VSS.n376 VSS.n369 11744.7
R106 VSS.n380 VSS.n369 11744.7
R107 VSS.n395 VSS.n383 11744.7
R108 VSS.n395 VSS.n384 11744.7
R109 VSS.n391 VSS.n383 11744.7
R110 VSS.n558 VSS.n15 9851.18
R111 VSS.n174 VSS.n153 7320.68
R112 VSS.n152 VSS.t88 7065.1
R113 VSS.t89 VSS.n15 7065.1
R114 VSS.n141 VSS.t88 6710.74
R115 VSS.n141 VSS.t89 6710.74
R116 VSS.n457 VSS.n456 6049.9
R117 VSS.n443 VSS.n13 6004.3
R118 VSS.n464 VSS.n463 5972.7
R119 VSS.n450 VSS.n449 5963.12
R120 VSS.n521 VSS.n520 5875.08
R121 VSS.n329 VSS.n315 5452.26
R122 VSS.n335 VSS.n315 5452.26
R123 VSS.n335 VSS.n314 5452.26
R124 VSS.n329 VSS.n314 5452.26
R125 VSS.n197 VSS.n190 5452.26
R126 VSS.n197 VSS.n191 5452.26
R127 VSS.n196 VSS.n191 5452.26
R128 VSS.n196 VSS.n190 5452.26
R129 VSS.n327 VSS.n318 5452.26
R130 VSS.n319 VSS.n318 5452.26
R131 VSS.n327 VSS.n320 5452.26
R132 VSS.n320 VSS.n319 5452.26
R133 VSS.n354 VSS.n186 5452.26
R134 VSS.n350 VSS.n186 5452.26
R135 VSS.n354 VSS.n187 5452.26
R136 VSS.n350 VSS.n187 5452.26
R137 VSS.n347 VSS.n308 5452.26
R138 VSS.n307 VSS.n306 5452.26
R139 VSS.n308 VSS.n306 5452.26
R140 VSS.n358 VSS.n182 5452.26
R141 VSS.n358 VSS.n183 5452.26
R142 VSS.n359 VSS.n182 5452.26
R143 VSS.n359 VSS.n183 5452.26
R144 VSS.n365 VSS.n175 5452.26
R145 VSS.n178 VSS.n175 5452.26
R146 VSS.n365 VSS.n176 5452.26
R147 VSS.n178 VSS.n176 5452.26
R148 VSS.n338 VSS.n204 5452.26
R149 VSS.n338 VSS.n205 5452.26
R150 VSS.n341 VSS.n205 5452.26
R151 VSS.n341 VSS.n204 5452.26
R152 VSS.n535 VSS.n534 5045.58
R153 VSS.n528 VSS.n527 4989.46
R154 VSS.n305 VSS 3384.3
R155 VSS.n467 VSS.n152 2857.05
R156 VSS VSS.n466 2525.55
R157 VSS.n475 VSS.n469 2384.59
R158 VSS.n558 VSS.n557 1919.2
R159 VSS.n466 VSS.n153 1685.21
R160 VSS.n397 VSS.n153 1610.68
R161 VSS.n520 VSS.t119 1455.01
R162 VSS.n477 VSS.n476 1363.79
R163 VSS.n478 VSS.n477 1342.5
R164 VSS VSS.t41 1289.66
R165 VSS VSS.t69 1289.66
R166 VSS.n584 VSS.n583 1198.25
R167 VSS.n98 VSS.n51 1198.25
R168 VSS.n480 VSS.n479 1198.25
R169 VSS.n293 VSS.n259 1198.25
R170 VSS.n489 VSS.n75 1194.5
R171 VSS.n303 VSS.n302 1194.5
R172 VSS.n510 VSS.n509 1171.32
R173 VSS.n570 VSS.n569 1171.32
R174 VSS.n560 VSS.n559 1121.18
R175 VSS.n366 VSS.t11 938.872
R176 VSS VSS.n75 918.774
R177 VSS.t90 VSS 918.774
R178 VSS.n303 VSS 918.774
R179 VSS.t142 VSS 918.774
R180 VSS.n474 VSS.t79 915.591
R181 VSS.n557 VSS.t45 915.591
R182 VSS.t79 VSS.n470 869.668
R183 VSS.n470 VSS.t45 869.668
R184 VSS.n475 VSS.n474 850.534
R185 VSS.t0 VSS.t98 826.054
R186 VSS.t102 VSS.t112 826.054
R187 VSS.t100 VSS.t28 826.054
R188 VSS.t71 VSS.t26 826.054
R189 VSS.t8 VSS.t139 792.337
R190 VSS.t39 VSS.t2 792.337
R191 VSS.n559 VSS.n558 789.042
R192 VSS.n414 VSS.n413 767.294
R193 VSS.n454 VSS.n453 767.294
R194 VSS.n532 VSS.n531 767.294
R195 VSS.n518 VSS.n50 767.294
R196 VSS.n563 VSS.n12 767.294
R197 VSS.n393 VSS.n392 767.294
R198 VSS.n461 VSS.n460 763.106
R199 VSS.n447 VSS.n446 763.106
R200 VSS.n168 VSS.n30 763.106
R201 VSS.n525 VSS.n524 763.106
R202 VSS.n378 VSS.n377 763.106
R203 VSS.n164 VSS.n160 763.106
R204 VSS.n472 VSS.n471 763.09
R205 VSS.n150 VSS.n143 763.09
R206 VSS.n413 VSS.n410 732.236
R207 VSS.n461 VSS.n419 732.236
R208 VSS.n454 VSS.n425 732.236
R209 VSS.n447 VSS.n436 732.236
R210 VSS.n471 VSS.n18 732.236
R211 VSS.n145 VSS.n143 732.236
R212 VSS.n168 VSS.n28 732.236
R213 VSS.n532 VSS.n36 732.236
R214 VSS.n525 VSS.n43 732.236
R215 VSS.n514 VSS.n50 732.236
R216 VSS.n12 VSS.n10 732.236
R217 VSS.n377 VSS.n374 732.236
R218 VSS.n392 VSS.n389 732.236
R219 VSS.n402 VSS.n160 732.236
R220 VSS.n469 VSS.n75 708.047
R221 VSS.t52 VSS.t64 708.047
R222 VSS.t139 VSS.t6 708.047
R223 VSS.t131 VSS.t129 708.047
R224 VSS.t10 VSS.t120 708.047
R225 VSS.n304 VSS.n303 708.047
R226 VSS.t56 VSS.t54 708.047
R227 VSS.t2 VSS.t37 708.047
R228 VSS.t136 VSS.t133 708.047
R229 VSS.t152 VSS.t110 708.047
R230 VSS.n510 VSS.t33 681.482
R231 VSS.n366 VSS.n365 631.774
R232 VSS.n569 VSS.t73 606.351
R233 VSS.n355 VSS.n185 601.636
R234 VSS.n559 VSS.n14 595.21
R235 VSS.t64 VSS 564.751
R236 VSS.t129 VSS 564.751
R237 VSS VSS.t10 564.751
R238 VSS VSS.n478 564.751
R239 VSS.t54 VSS 564.751
R240 VSS.t133 VSS 564.751
R241 VSS VSS.t152 564.751
R242 VSS VSS.n14 564.751
R243 VSS.n382 VSS.n166 558.457
R244 VSS.t43 VSS.n192 538.306
R245 VSS.t138 VSS.n184 538.306
R246 VSS.n203 VSS.t141 538.306
R247 VSS.n349 VSS.t50 538.306
R248 VSS.n174 VSS.t17 529.082
R249 VSS.t120 VSS.t104 522.606
R250 VSS.t110 VSS.t20 522.606
R251 VSS.n476 VSS.n475 481.236
R252 VSS.t87 VSS 480.461
R253 VSS.t86 VSS 480.461
R254 VSS.n192 VSS.n184 474.976
R255 VSS.n349 VSS.n203 474.976
R256 VSS VSS.t33 459.26
R257 VSS.t48 VSS.t46 425.807
R258 VSS.t138 VSS.n355 411.646
R259 VSS.t46 VSS.n304 394.265
R260 VSS.n206 VSS.t76 393.586
R261 VSS.t104 VSS.t90 387.74
R262 VSS.t20 VSS.t142 387.74
R263 VSS.n568 VSS 384.901
R264 VSS VSS.t147 370.37
R265 VSS VSS.t84 370.37
R266 VSS.t11 VSS.n166 365.587
R267 VSS.t43 VSS.n167 365.587
R268 VSS.n326 VSS.n325 354.26
R269 VSS.n325 VSS.n324 354.26
R270 VSS.n353 VSS.n352 354.26
R271 VSS.n352 VSS.n351 354.26
R272 VSS.n346 VSS.n345 354.26
R273 VSS.n346 VSS.n309 354.26
R274 VSS.n357 VSS.n180 354.26
R275 VSS.n357 VSS.n356 354.26
R276 VSS.n339 VSS.n312 354.26
R277 VSS.n340 VSS.n339 354.26
R278 VSS.n195 VSS.n188 354.26
R279 VSS.n334 VSS.n316 354.26
R280 VSS.n334 VSS.n333 354.26
R281 VSS.n367 VSS.n174 342.298
R282 VSS.n479 VSS.t135 337.166
R283 VSS.n259 VSS.t144 337.166
R284 VSS.n511 VSS.n51 334.815
R285 VSS.n561 VSS.n560 332.642
R286 VSS.t44 VSS.t48 331.183
R287 VSS.t141 VSS.n154 326.726
R288 VSS.n415 VSS.n414 325.502
R289 VSS.n453 VSS.n452 325.502
R290 VSS.n531 VSS.n530 325.502
R291 VSS.n518 VSS.n517 325.502
R292 VSS.n564 VSS.n563 325.502
R293 VSS.n394 VSS.n393 325.502
R294 VSS.n479 VSS.t0 320.307
R295 VSS.n259 VSS.t100 320.307
R296 VSS.n472 VSS.n19 304.553
R297 VSS.n150 VSS.n149 304.553
R298 VSS.n460 VSS.n459 304.204
R299 VSS.n446 VSS.n445 304.204
R300 VSS.n537 VSS.n30 304.204
R301 VSS.n524 VSS.n523 304.204
R302 VSS.n379 VSS.n378 304.204
R303 VSS.n165 VSS.n164 304.204
R304 VSS.t135 VSS 295.019
R305 VSS.t144 VSS 295.019
R306 VSS.n554 VSS.n19 266.349
R307 VSS.n149 VSS.n148 266.349
R308 VSS VSS.t44 264.159
R309 VSS VSS.t8 261.303
R310 VSS VSS.t39 261.303
R311 VSS.n194 VSS.n179 255.839
R312 VSS.n195 VSS.n194 253.365
R313 VSS.t147 VSS.t149 248.889
R314 VSS.t124 VSS.t127 248.889
R315 VSS.t84 VSS.t116 248.889
R316 VSS.t30 VSS 244.445
R317 VSS.t66 VSS 244.445
R318 VSS.n415 VSS.n157 242.448
R319 VSS.n459 VSS.n421 242.448
R320 VSS.n452 VSS.n432 242.448
R321 VSS.n445 VSS.n440 242.448
R322 VSS.n538 VSS.n537 242.448
R323 VSS.n530 VSS.n39 242.448
R324 VSS.n523 VSS.n46 242.448
R325 VSS.n517 VSS.n516 242.448
R326 VSS.n565 VSS.n564 242.448
R327 VSS.n379 VSS.n370 242.448
R328 VSS.n394 VSS.n385 242.448
R329 VSS.n165 VSS.n159 242.448
R330 VSS.n496 VSS.t9 240.575
R331 VSS.n286 VSS.t40 240.575
R332 VSS.n137 VSS.t42 237.327
R333 VSS.n298 VSS.t70 237.327
R334 VSS.n469 VSS.n468 223.726
R335 VSS VSS.n51 222.222
R336 VSS VSS.n510 222.222
R337 VSS.t23 VSS.t122 221.451
R338 VSS.n233 VSS.t155 218.308
R339 VSS.n211 VSS.t157 218.308
R340 VSS.n116 VSS.t154 218.308
R341 VSS.n79 VSS.t156 218.308
R342 VSS.n483 VSS.t153 218.308
R343 VSS.n60 VSS.t159 218.308
R344 VSS.n268 VSS.t158 218.308
R345 VSS.n255 VSS.t160 218.308
R346 VSS.n230 VSS.t74 214.456
R347 VSS.n232 VSS.t75 214.456
R348 VSS.n243 VSS.t77 214.456
R349 VSS.n212 VSS.t78 214.456
R350 VSS.n113 VSS.t34 214.456
R351 VSS.n115 VSS.t35 214.456
R352 VSS.n126 VSS.t18 214.456
R353 VSS.n80 VSS.t19 214.456
R354 VSS.n488 VSS.t31 214.456
R355 VSS.n482 VSS.t32 214.456
R356 VSS.n55 VSS.t105 214.456
R357 VSS.n59 VSS.t106 214.456
R358 VSS.n264 VSS.t21 214.456
R359 VSS.n267 VSS.t22 214.456
R360 VSS.n208 VSS.t67 214.456
R361 VSS.n256 VSS.t68 214.456
R362 VSS.n328 VSS.t109 208.017
R363 VSS.t107 VSS.n313 208.017
R364 VSS.n131 VSS.n130 204.457
R365 VSS.n250 VSS.n249 204.457
R366 VSS.n68 VSS.n67 200.231
R367 VSS.n73 VSS.n72 200.231
R368 VSS.n280 VSS.n277 200.231
R369 VSS.n258 VSS.n257 200.231
R370 VSS.n62 VSS.n57 200.105
R371 VSS.n270 VSS.n265 200.105
R372 VSS.t114 VSS 198.519
R373 VSS.t149 VSS 198.519
R374 VSS.t127 VSS 198.519
R375 VSS.t116 VSS 198.519
R376 VSS.n569 VSS 197.724
R377 VSS.t15 VSS.t118 195.97
R378 VSS.n453 VSS.n424 195
R379 VSS.n424 VSS.t92 195
R380 VSS.n431 VSS.n423 195
R381 VSS.n423 VSS.t92 195
R382 VSS.n437 VSS.n434 195
R383 VSS.n434 VSS.t61 195
R384 VSS.n446 VSS.n435 195
R385 VSS.n435 VSS.t61 195
R386 VSS.n147 VSS.n146 195
R387 VSS.n146 VSS.n15 195
R388 VSS.n151 VSS.n150 195
R389 VSS.n152 VSS.n151 195
R390 VSS.n567 VSS.n566 195
R391 VSS.n568 VSS.n567 195
R392 VSS.n563 VSS.n562 195
R393 VSS.n562 VSS.t25 195
R394 VSS.n556 VSS.n555 195
R395 VSS.n557 VSS.n556 195
R396 VSS.n473 VSS.n472 195
R397 VSS.n474 VSS.n473 195
R398 VSS.n519 VSS.n518 195
R399 VSS.n520 VSS.n519 195
R400 VSS.n513 VSS.n512 195
R401 VSS.n512 VSS.n511 195
R402 VSS.n524 VSS.n42 195
R403 VSS.n42 VSS.t126 195
R404 VSS.n44 VSS.n41 195
R405 VSS.n41 VSS.t126 195
R406 VSS.n531 VSS.n35 195
R407 VSS.n35 VSS.t151 195
R408 VSS.n37 VSS.n34 195
R409 VSS.n34 VSS.t151 195
R410 VSS.n32 VSS.n30 195
R411 VSS.t4 VSS.n32 195
R412 VSS.n31 VSS.n29 195
R413 VSS.t4 VSS.n31 195
R414 VSS.n378 VSS.n369 195
R415 VSS.n369 VSS.t51 195
R416 VSS.n373 VSS.n368 195
R417 VSS.n388 VSS.n383 195
R418 VSS.n383 VSS.t95 195
R419 VSS.n393 VSS.n384 195
R420 VSS.n164 VSS.n163 195
R421 VSS.t60 VSS.n163 195
R422 VSS.n401 VSS.n400 195
R423 VSS.n414 VSS.n156 195
R424 VSS.n156 VSS.t5 195
R425 VSS.n409 VSS.n155 195
R426 VSS.n460 VSS.n418 195
R427 VSS.n418 VSS.t12 195
R428 VSS.n420 VSS.n417 195
R429 VSS.n417 VSS.t12 195
R430 VSS.n411 VSS.n155 188.989
R431 VSS.n400 VSS.n161 188.988
R432 VSS.n390 VSS.n384 188.986
R433 VSS.n375 VSS.n368 188.984
R434 VSS.t50 VSS.n305 188.119
R435 VSS.t25 VSS.n13 183.936
R436 VSS.n468 VSS.n467 183.457
R437 VSS VSS.t102 177.012
R438 VSS VSS.t71 177.012
R439 VSS.t122 VSS 176.633
R440 VSS.n560 VSS 176.633
R441 VSS.n376 VSS.n375 173.373
R442 VSS.n391 VSS.n390 173.304
R443 VSS.n162 VSS.n161 173.167
R444 VSS.n412 VSS.n411 173.097
R445 VSS.n223 VSS.t83 162.471
R446 VSS.n218 VSS.t97 162.471
R447 VSS.n582 VSS.t63 162.471
R448 VSS.n577 VSS.t24 162.471
R449 VSS.n106 VSS.t146 162.471
R450 VSS.n101 VSS.t148 162.471
R451 VSS.n97 VSS.t125 162.471
R452 VSS.n92 VSS.t85 162.471
R453 VSS.n497 VSS.t140 162.471
R454 VSS.n260 VSS.t3 162.471
R455 VSS.n68 VSS.t132 160.046
R456 VSS.n73 VSS.t53 160.046
R457 VSS.n280 VSS.t137 160.046
R458 VSS.n258 VSS.t57 160.046
R459 VSS.n214 VSS.t81 160.017
R460 VSS.n0 VSS.t94 160.017
R461 VSS.n3 VSS.t59 160.017
R462 VSS.n575 VSS.t123 160.017
R463 VSS.n82 VSS.t115 160.017
R464 VSS.n99 VSS.t150 160.017
R465 VSS.n87 VSS.t128 160.017
R466 VSS.n90 VSS.t117 160.017
R467 VSS.n504 VSS.t130 160.017
R468 VSS.n499 VSS.t7 160.017
R469 VSS.n275 VSS.t134 160.017
R470 VSS.n281 VSS.t38 160.017
R471 VSS.n496 VSS.t65 158.534
R472 VSS.n286 VSS.t55 158.534
R473 VSS.t118 VSS 156.31
R474 VSS.n456 VSS.t92 155.954
R475 VSS.n463 VSS.t12 155.954
R476 VSS.n449 VSS.t61 155.831
R477 VSS.n534 VSS.t151 153.75
R478 VSS.n170 VSS.t4 153.75
R479 VSS.n527 VSS.t126 153.63
R480 VSS VSS.t76 140.185
R481 VSS.n332 VSS.n330 139.727
R482 VSS.t25 VSS.n561 139.648
R483 VSS.t17 VSS 131.004
R484 VSS.n584 VSS.t62 128.429
R485 VSS.n341 VSS.n206 127.624
R486 VSS.n342 VSS.n340 123.882
R487 VSS.t36 VSS 121.481
R488 VSS.n381 VSS.n380 118.54
R489 VSS.n365 VSS.n364 117.121
R490 VSS.n179 VSS.n178 117.001
R491 VSS.n178 VSS.n167 117.001
R492 VSS.n356 VSS.n183 117.001
R493 VSS.n185 VSS.n183 117.001
R494 VSS.n182 VSS.n180 117.001
R495 VSS.n192 VSS.n182 117.001
R496 VSS.n309 VSS.n308 117.001
R497 VSS.n308 VSS.n203 117.001
R498 VSS.n351 VSS.n350 117.001
R499 VSS.n350 VSS.n349 117.001
R500 VSS.n354 VSS.n353 117.001
R501 VSS.n355 VSS.n354 117.001
R502 VSS.n345 VSS.n307 117.001
R503 VSS.n324 VSS.n319 117.001
R504 VSS.t109 VSS.n319 117.001
R505 VSS.n327 VSS.n326 117.001
R506 VSS.t109 VSS.n327 117.001
R507 VSS.n312 VSS.n204 117.001
R508 VSS.t50 VSS.n204 117.001
R509 VSS.n340 VSS.n205 117.001
R510 VSS.t50 VSS.n205 117.001
R511 VSS.n193 VSS.n190 117.001
R512 VSS.n190 VSS.n166 117.001
R513 VSS.n191 VSS.n188 117.001
R514 VSS.n191 VSS.n184 117.001
R515 VSS.n316 VSS.n314 117.001
R516 VSS.t107 VSS.n314 117.001
R517 VSS.n333 VSS.n315 117.001
R518 VSS.t107 VSS.n315 117.001
R519 VSS.n348 VSS.n307 113.879
R520 VSS VSS.t82 113.052
R521 VSS VSS.t96 113.052
R522 VSS.n396 VSS.n395 111.895
R523 VSS.n399 VSS.n398 111.808
R524 VSS VSS.t145 105.647
R525 VSS.n457 VSS.n422 99.881
R526 VSS.n535 VSS.n33 98.4693
R527 VSS.n450 VSS.n433 93.748
R528 VSS.n443 VSS.n442 93.6734
R529 VSS.n528 VSS.n40 92.423
R530 VSS.n521 VSS.n47 92.3504
R531 VSS.n465 VSS.t5 89.4314
R532 VSS.n382 VSS.n167 89.2383
R533 VSS.n345 VSS.n344 89.224
R534 VSS.n310 VSS.n309 89.224
R535 VSS.n361 VSS.n180 89.224
R536 VSS.n356 VSS.n181 89.224
R537 VSS.n343 VSS.n312 89.224
R538 VSS.n317 VSS.n316 89.224
R539 VSS.n362 VSS.n179 88.4711
R540 VSS.n511 VSS.t124 85.9264
R541 VSS.n185 VSS.n154 84.9204
R542 VSS.n199 VSS.n188 84.7064
R543 VSS.t6 VSS.t87 84.2917
R544 VSS.t37 VSS.t86 84.2917
R545 VSS.n337 VSS.n336 81.3982
R546 VSS.n326 VSS.n321 80.1887
R547 VSS.n324 VSS.n323 80.1887
R548 VSS.n353 VSS.n200 80.1887
R549 VSS.n351 VSS.n202 80.1887
R550 VSS.t82 VSS.t80 75.9717
R551 VSS.t96 VSS.t93 75.9717
R552 VSS.t58 VSS.t62 75.9717
R553 VSS.n130 VSS.t16 72.8576
R554 VSS.n57 VSS.t121 72.8576
R555 VSS.n265 VSS.t111 72.8576
R556 VSS.n249 VSS.t49 72.8576
R557 VSS.n465 VSS.n464 72.6343
R558 VSS VSS.n584 67.8319
R559 VSS.n396 VSS.t95 66.9242
R560 VSS.n398 VSS.t60 66.8669
R561 VSS.n198 VSS.n189 64.8307
R562 VSS.n433 VSS.t92 62.2068
R563 VSS.n442 VSS.t61 62.1573
R564 VSS.n40 VSS.t151 61.3275
R565 VSS.n47 VSS.t126 61.2794
R566 VSS.n467 VSS.t15 60.658
R567 VSS.t80 VSS 60.5966
R568 VSS.t93 VSS 60.5966
R569 VSS VSS.t58 60.5966
R570 VSS.n381 VSS.t51 60.352
R571 VSS.n177 VSS.n175 58.7133
R572 VSS.n67 VSS.t103 58.5719
R573 VSS.n72 VSS.t1 58.5719
R574 VSS.n277 VSS.t72 58.5719
R575 VSS.n257 VSS.t101 58.5719
R576 VSS.n422 VSS.t12 56.0738
R577 VSS.t4 VSS.n33 55.2812
R578 VSS.n555 VSS.n554 54.2123
R579 VSS.n148 VSS.n147 54.2123
R580 VSS.n328 VSS.n318 54.2066
R581 VSS.n364 VSS.n363 52.1725
R582 VSS.t98 VSS.t52 50.5752
R583 VSS.t112 VSS.t131 50.5752
R584 VSS.t28 VSS.t56 50.5752
R585 VSS.t26 VSS.t136 50.5752
R586 VSS.t145 VSS.n173 47.3305
R587 VSS.n129 VSS 43.9579
R588 VSS.n247 VSS 43.9579
R589 VSS.n561 VSS.n9 42.2329
R590 VSS.n199 VSS.n198 42.1089
R591 VSS.n201 VSS.n200 42.1089
R592 VSS.n202 VSS.n201 42.1089
R593 VSS.n322 VSS.n321 42.1089
R594 VSS.n323 VSS.n322 42.1089
R595 VSS.n330 VSS.n317 42.1089
R596 VSS.n337 VSS.n305 41.6038
R597 VSS.n200 VSS.n199 39.4771
R598 VSS.n321 VSS.n202 35.2902
R599 VSS.n363 VSS.n362 34.659
R600 VSS.n361 VSS.n360 34.659
R601 VSS.n360 VSS.n181 34.659
R602 VSS.n311 VSS.n310 34.659
R603 VSS.n344 VSS.n311 34.659
R604 VSS.n343 VSS.n342 34.659
R605 VSS.n132 VSS.n129 34.6358
R606 VSS.n136 VSS.n76 34.6358
R607 VSS.n248 VSS.n247 34.6358
R608 VSS.n251 VSS.n207 34.6358
R609 VSS.n358 VSS.n357 32.5005
R610 VSS.t138 VSS.n358 32.5005
R611 VSS.n347 VSS.n346 32.5005
R612 VSS.n352 VSS.n187 32.5005
R613 VSS.t141 VSS.n187 32.5005
R614 VSS.n325 VSS.n320 32.5005
R615 VSS.n320 VSS.n313 32.5005
R616 VSS.n339 VSS.n338 32.5005
R617 VSS.n338 VSS.n337 32.5005
R618 VSS.n363 VSS.n176 32.5005
R619 VSS.n176 VSS.t11 32.5005
R620 VSS.n360 VSS.n359 32.5005
R621 VSS.n359 VSS.t138 32.5005
R622 VSS.n311 VSS.n306 32.5005
R623 VSS.t50 VSS.n306 32.5005
R624 VSS.n342 VSS.n341 32.5005
R625 VSS.n175 VSS.t11 32.5005
R626 VSS.n196 VSS.n195 32.5005
R627 VSS.t43 VSS.n196 32.5005
R628 VSS.n198 VSS.n197 32.5005
R629 VSS.n197 VSS.t43 32.5005
R630 VSS.n201 VSS.n186 32.5005
R631 VSS.t141 VSS.n186 32.5005
R632 VSS.n322 VSS.n318 32.5005
R633 VSS.n330 VSS.n329 32.5005
R634 VSS.n329 VSS.n328 32.5005
R635 VSS.n335 VSS.n334 32.5005
R636 VSS.n336 VSS.n335 32.5005
R637 VSS.n310 VSS.n181 32.4928
R638 VSS.n348 VSS.n347 31.6336
R639 VSS.n362 VSS.n361 30.9174
R640 VSS.n410 VSS.n409 30.8711
R641 VSS.n420 VSS.n419 30.8711
R642 VSS.n431 VSS.n425 30.8711
R643 VSS.n437 VSS.n436 30.8711
R644 VSS.n555 VSS.n18 30.8711
R645 VSS.n147 VSS.n145 30.8711
R646 VSS.n29 VSS.n28 30.8711
R647 VSS.n37 VSS.n36 30.8711
R648 VSS.n44 VSS.n43 30.8711
R649 VSS.n514 VSS.n513 30.8711
R650 VSS.n566 VSS.n10 30.8711
R651 VSS.n374 VSS.n373 30.8711
R652 VSS.n389 VSS.n388 30.8711
R653 VSS.n402 VSS.n401 30.8711
R654 VSS.n333 VSS.n332 30.8711
R655 VSS.n323 VSS.n317 30.7444
R656 VSS.n441 VSS 29.8463
R657 VSS.n344 VSS.n343 28.259
R658 VSS.n509 VSS.n52 26.9246
R659 VSS.n570 VSS.n5 26.9246
R660 VSS.n478 VSS.t36 26.1252
R661 VSS.n489 VSS.n136 25.6926
R662 VSS.n302 VSS.n207 25.6926
R663 VSS.n67 VSS.t113 25.4291
R664 VSS.n72 VSS.t99 25.4291
R665 VSS.n277 VSS.t27 25.4291
R666 VSS.n257 VSS.t29 25.4291
R667 VSS.n223 VSS.n222 25.224
R668 VSS.n222 VSS.n214 25.224
R669 VSS.n218 VSS.n217 25.224
R670 VSS.n217 VSS.n0 25.224
R671 VSS.n582 VSS.n581 25.224
R672 VSS.n581 VSS.n3 25.224
R673 VSS.n577 VSS.n576 25.224
R674 VSS.n576 VSS.n575 25.224
R675 VSS.n106 VSS.n105 25.224
R676 VSS.n105 VSS.n82 25.224
R677 VSS.n101 VSS.n100 25.224
R678 VSS.n100 VSS.n99 25.224
R679 VSS.n97 VSS.n96 25.224
R680 VSS.n96 VSS.n87 25.224
R681 VSS.n92 VSS.n91 25.224
R682 VSS.n91 VSS.n90 25.224
R683 VSS.n504 VSS.n503 25.224
R684 VSS.n498 VSS.n497 25.224
R685 VSS.n499 VSS.n498 25.224
R686 VSS.n276 VSS.n275 25.224
R687 VSS.n282 VSS.n260 25.224
R688 VSS.n282 VSS.n281 25.224
R689 VSS.n496 VSS.n495 24.0946
R690 VSS.n287 VSS.n286 24.0946
R691 VSS.t73 VSS.n568 23.7273
R692 VSS.n364 VSS.n177 23.3238
R693 VSS.n130 VSS.t14 22.3257
R694 VSS.n57 VSS.t91 22.3257
R695 VSS.n265 VSS.t143 22.3257
R696 VSS.n249 VSS.t47 22.3257
R697 VSS.t109 VSS.t107 21.7066
R698 VSS.n336 VSS.n313 21.7066
R699 VSS.n194 VSS.n193 21.6752
R700 VSS.n503 VSS.n68 21.4593
R701 VSS.n495 VSS.n73 21.4593
R702 VSS.n280 VSS.n276 21.4593
R703 VSS.n287 VSS.n258 21.4593
R704 VSS.n218 VSS.n214 20.3299
R705 VSS.n577 VSS.n3 20.3299
R706 VSS.n101 VSS.n82 20.3299
R707 VSS.n92 VSS.n87 20.3299
R708 VSS.n224 VSS.n223 19.2926
R709 VSS.n107 VSS.n106 19.2926
R710 VSS.n476 VSS.t119 18.2451
R711 VSS.n504 VSS.n66 17.7867
R712 VSS.n275 VSS.n262 17.7867
R713 VSS.n583 VSS.n582 17.3181
R714 VSS.n98 VSS.n97 17.3181
R715 VSS.t41 VSS.t30 16.8587
R716 VSS.t69 VSS.t66 16.8587
R717 VSS.n583 VSS.n0 15.8123
R718 VSS.n575 VSS.n5 15.8123
R719 VSS.n99 VSS.n98 15.8123
R720 VSS.n90 VSS.n52 15.8123
R721 VSS.n464 VSS.n416 15.1478
R722 VSS.t50 VSS.n206 14.9893
R723 VSS.n229 VSS.n5 14.775
R724 VSS.n112 VSS.n52 14.775
R725 VSS.n481 VSS.n480 14.775
R726 VSS.n294 VSS.n293 14.775
R727 VSS.n497 VSS.n496 13.5534
R728 VSS.n286 VSS.n260 13.5534
R729 VSS.n128 VSS.n127 11.2844
R730 VSS.n245 VSS.n244 11.2844
R731 VSS.n452 VSS.n451 11.0382
R732 VSS.n451 VSS.n450 11.0382
R733 VSS.n455 VSS.n454 11.0382
R734 VSS.n456 VSS.n455 11.0382
R735 VSS.n448 VSS.n447 11.0382
R736 VSS.n449 VSS.n448 11.0382
R737 VSS.n445 VSS.n444 11.0382
R738 VSS.n444 VSS.n443 11.0382
R739 VSS.n149 VSS.n142 11.0382
R740 VSS.n142 VSS.n141 11.0382
R741 VSS.n143 VSS.n140 11.0382
R742 VSS.n141 VSS.n140 11.0382
R743 VSS.n564 VSS.n9 11.0382
R744 VSS.n12 VSS.n8 11.0382
R745 VSS.n13 VSS.n8 11.0382
R746 VSS.n19 VSS.n17 11.0382
R747 VSS.n470 VSS.n17 11.0382
R748 VSS.n471 VSS.n16 11.0382
R749 VSS.n470 VSS.n16 11.0382
R750 VSS.n517 VSS.n49 11.0382
R751 VSS.n477 VSS.n49 11.0382
R752 VSS.n50 VSS.n48 11.0382
R753 VSS.n477 VSS.n48 11.0382
R754 VSS.n523 VSS.n522 11.0382
R755 VSS.n522 VSS.n521 11.0382
R756 VSS.n526 VSS.n525 11.0382
R757 VSS.n527 VSS.n526 11.0382
R758 VSS.n530 VSS.n529 11.0382
R759 VSS.n529 VSS.n528 11.0382
R760 VSS.n533 VSS.n532 11.0382
R761 VSS.n534 VSS.n533 11.0382
R762 VSS.n537 VSS.n536 11.0382
R763 VSS.n536 VSS.n535 11.0382
R764 VSS.n169 VSS.n168 11.0382
R765 VSS.n170 VSS.n169 11.0382
R766 VSS.n380 VSS.n379 11.0382
R767 VSS.n377 VSS.n376 11.0382
R768 VSS.n392 VSS.n391 11.0382
R769 VSS.n395 VSS.n394 11.0382
R770 VSS.n399 VSS.n165 11.0382
R771 VSS.n162 VSS.n160 11.0382
R772 VSS.n416 VSS.n415 11.0382
R773 VSS.n413 VSS.n412 11.0382
R774 VSS.n459 VSS.n458 11.0382
R775 VSS.n458 VSS.n457 11.0382
R776 VSS.n462 VSS.n461 11.0382
R777 VSS.n463 VSS.n462 11.0382
R778 VSS.n409 VSS.n157 10.9181
R779 VSS.n421 VSS.n420 10.9181
R780 VSS.n432 VSS.n431 10.9181
R781 VSS.n440 VSS.n437 10.9181
R782 VSS.n538 VSS.n29 10.9181
R783 VSS.n39 VSS.n37 10.9181
R784 VSS.n46 VSS.n44 10.9181
R785 VSS.n516 VSS.n513 10.9181
R786 VSS.n566 VSS.n565 10.9181
R787 VSS.n373 VSS.n370 10.9181
R788 VSS.n388 VSS.n385 10.9181
R789 VSS.n401 VSS.n159 10.9181
R790 VSS.n331 VSS.t108 10.7858
R791 VSS.n410 VSS.n408 10.4476
R792 VSS.n426 VSS.n419 10.4476
R793 VSS.n430 VSS.n425 10.4476
R794 VSS.n439 VSS.n436 10.4476
R795 VSS.n553 VSS.n18 10.4476
R796 VSS.n145 VSS.n144 10.4476
R797 VSS.n539 VSS.n28 10.4476
R798 VSS.n38 VSS.n36 10.4476
R799 VSS.n45 VSS.n43 10.4476
R800 VSS.n515 VSS.n514 10.4476
R801 VSS.n11 VSS.n10 10.4476
R802 VSS.n374 VSS.n372 10.4476
R803 VSS.n389 VSS.n387 10.4476
R804 VSS.n403 VSS.n402 10.4476
R805 VSS.n499 VSS.n68 10.1652
R806 VSS.n281 VSS.n280 10.1652
R807 VSS.n232 VSS.n227 9.70901
R808 VSS.n244 VSS.n243 9.70901
R809 VSS.n115 VSS.n110 9.70901
R810 VSS.n127 VSS.n126 9.70901
R811 VSS.n59 VSS.n58 9.70901
R812 VSS.n267 VSS.n266 9.70901
R813 VSS.n131 VSS.n76 9.41227
R814 VSS.n251 VSS.n250 9.41227
R815 VSS.n490 VSS.n489 9.3005
R816 VSS.n487 VSS.n486 9.3005
R817 VSS.n74 VSS.n73 9.3005
R818 VSS.n496 VSS.n71 9.3005
R819 VSS.n501 VSS.n68 9.3005
R820 VSS.n61 VSS.n56 9.3005
R821 VSS.n64 VSS.n63 9.3005
R822 VSS.n66 VSS.n65 9.3005
R823 VSS.n505 VSS.n504 9.3005
R824 VSS.n503 VSS.n502 9.3005
R825 VSS.n500 VSS.n499 9.3005
R826 VSS.n498 VSS.n69 9.3005
R827 VSS.n497 VSS.n70 9.3005
R828 VSS.n495 VSS.n494 9.3005
R829 VSS.n480 VSS.n139 9.3005
R830 VSS.n481 VSS.n138 9.3005
R831 VSS.n485 VSS.n484 9.3005
R832 VSS.n136 VSS.n135 9.3005
R833 VSS.n134 VSS.n76 9.3005
R834 VSS.n133 VSS.n132 9.3005
R835 VSS.n129 VSS.n77 9.3005
R836 VSS.n509 VSS.n508 9.3005
R837 VSS.n90 VSS.n89 9.3005
R838 VSS.n94 VSS.n87 9.3005
R839 VSS.n98 VSS.n85 9.3005
R840 VSS.n99 VSS.n84 9.3005
R841 VSS.n103 VSS.n82 9.3005
R842 VSS.n108 VSS.n107 9.3005
R843 VSS.n124 VSS.n123 9.3005
R844 VSS.n125 VSS.n78 9.3005
R845 VSS.n106 VSS.n81 9.3005
R846 VSS.n105 VSS.n104 9.3005
R847 VSS.n102 VSS.n101 9.3005
R848 VSS.n100 VSS.n83 9.3005
R849 VSS.n97 VSS.n86 9.3005
R850 VSS.n96 VSS.n95 9.3005
R851 VSS.n93 VSS.n92 9.3005
R852 VSS.n91 VSS.n88 9.3005
R853 VSS.n118 VSS.n117 9.3005
R854 VSS.n114 VSS.n109 9.3005
R855 VSS.n112 VSS.n111 9.3005
R856 VSS.n54 VSS.n52 9.3005
R857 VSS.n571 VSS.n570 9.3005
R858 VSS.n575 VSS.n574 9.3005
R859 VSS.n579 VSS.n3 9.3005
R860 VSS.n583 VSS.n1 9.3005
R861 VSS.n215 VSS.n0 9.3005
R862 VSS.n220 VSS.n214 9.3005
R863 VSS.n225 VSS.n224 9.3005
R864 VSS.n241 VSS.n240 9.3005
R865 VSS.n242 VSS.n210 9.3005
R866 VSS.n223 VSS.n213 9.3005
R867 VSS.n222 VSS.n221 9.3005
R868 VSS.n219 VSS.n218 9.3005
R869 VSS.n217 VSS.n216 9.3005
R870 VSS.n582 VSS.n2 9.3005
R871 VSS.n581 VSS.n580 9.3005
R872 VSS.n578 VSS.n577 9.3005
R873 VSS.n576 VSS.n4 9.3005
R874 VSS.n235 VSS.n234 9.3005
R875 VSS.n231 VSS.n226 9.3005
R876 VSS.n229 VSS.n228 9.3005
R877 VSS.n573 VSS.n5 9.3005
R878 VSS.n302 VSS.n301 9.3005
R879 VSS.n300 VSS.n299 9.3005
R880 VSS.n291 VSS.n258 9.3005
R881 VSS.n286 VSS.n285 9.3005
R882 VSS.n280 VSS.n279 9.3005
R883 VSS.n269 VSS.n263 9.3005
R884 VSS.n272 VSS.n271 9.3005
R885 VSS.n273 VSS.n262 9.3005
R886 VSS.n275 VSS.n274 9.3005
R887 VSS.n278 VSS.n276 9.3005
R888 VSS.n281 VSS.n261 9.3005
R889 VSS.n283 VSS.n282 9.3005
R890 VSS.n284 VSS.n260 9.3005
R891 VSS.n288 VSS.n287 9.3005
R892 VSS.n295 VSS.n294 9.3005
R893 VSS.n297 VSS.n296 9.3005
R894 VSS.n253 VSS.n207 9.3005
R895 VSS.n252 VSS.n251 9.3005
R896 VSS.n248 VSS.n209 9.3005
R897 VSS.n247 VSS.n246 9.3005
R898 VSS.n293 VSS.n292 9.3005
R899 VSS.n428 VSS.n427 8.45078
R900 VSS.n541 VSS.n540 8.45078
R901 VSS.n371 VSS.n158 8.45078
R902 VSS.n407 VSS.n406 8.30267
R903 VSS.n543 VSS.n25 8.30267
R904 VSS.n550 VSS.n549 8.30267
R905 VSS.n438 VSS.n21 7.97888
R906 VSS.n542 VSS.n26 7.97888
R907 VSS.n405 VSS.n404 7.97888
R908 VSS.n429 VSS.n428 7.97601
R909 VSS.n541 VSS.n27 7.97601
R910 VSS.n386 VSS.n158 7.97601
R911 VSS.n408 VSS.n407 7.16724
R912 VSS.n427 VSS.n426 7.16724
R913 VSS.n430 VSS.n429 7.16724
R914 VSS.n439 VSS.n438 7.16724
R915 VSS.n553 VSS.n552 7.16724
R916 VSS.n144 VSS.n20 7.16724
R917 VSS.n540 VSS.n539 7.16724
R918 VSS.n38 VSS.n27 7.16724
R919 VSS.n45 VSS.n26 7.16724
R920 VSS.n515 VSS.n25 7.16724
R921 VSS.n549 VSS.n11 7.16724
R922 VSS.n372 VSS.n371 7.16724
R923 VSS.n387 VSS.n386 7.16724
R924 VSS.n404 VSS.n403 7.16724
R925 VSS.n480 VSS.n73 7.15344
R926 VSS.n293 VSS.n258 7.15344
R927 VSS.n507 VSS.n506 6.50373
R928 VSS.n572 VSS.n7 6.50373
R929 VSS.n132 VSS.n131 6.4005
R930 VSS.n250 VSS.n248 6.4005
R931 VSS.n234 VSS.n231 6.26433
R932 VSS.n242 VSS.n241 6.26433
R933 VSS.n117 VSS.n114 6.26433
R934 VSS.n125 VSS.n124 6.26433
R935 VSS.n231 VSS.n230 5.85582
R936 VSS.n243 VSS.n242 5.85582
R937 VSS.n114 VSS.n113 5.85582
R938 VSS.n126 VSS.n125 5.85582
R939 VSS.n63 VSS.n55 5.85582
R940 VSS.n488 VSS.n487 5.85582
R941 VSS.n484 VSS.n137 5.85582
R942 VSS.n271 VSS.n264 5.85582
R943 VSS.n299 VSS.n208 5.85582
R944 VSS.n298 VSS.n297 5.85582
R945 VSS.n507 VSS.n54 4.788
R946 VSS.n573 VSS.n572 4.788
R947 VSS.n408 VSS.n157 4.73093
R948 VSS.n426 VSS.n421 4.73093
R949 VSS.n432 VSS.n430 4.73093
R950 VSS.n440 VSS.n439 4.73093
R951 VSS.n539 VSS.n538 4.73093
R952 VSS.n39 VSS.n38 4.73093
R953 VSS.n46 VSS.n45 4.73093
R954 VSS.n516 VSS.n515 4.73093
R955 VSS.n565 VSS.n11 4.73093
R956 VSS.n372 VSS.n370 4.73093
R957 VSS.n387 VSS.n385 4.73093
R958 VSS.n403 VSS.n159 4.73093
R959 VSS.n332 VSS.n331 4.5578
R960 VSS.n508 VSS.n507 4.50726
R961 VSS.n572 VSS.n571 4.50726
R962 VSS.n468 VSS.t13 4.31383
R963 VSS.n548 VSS 4.01425
R964 VSS.n23 VSS 4.01425
R965 VSS.n544 VSS 4.01425
R966 VSS.n554 VSS.n553 3.78485
R967 VSS.n148 VSS.n144 3.78485
R968 VSS.n193 VSS.n189 3.75517
R969 VSS.n62 VSS.n61 3.40476
R970 VSS.n270 VSS.n269 3.40476
R971 VSS.n234 VSS.n233 3.13241
R972 VSS.n241 VSS.n211 3.13241
R973 VSS.n117 VSS.n116 3.13241
R974 VSS.n124 VSS.n79 3.13241
R975 VSS.n61 VSS.n60 3.13241
R976 VSS.n484 VSS.n483 3.13241
R977 VSS.n269 VSS.n268 3.13241
R978 VSS.n297 VSS.n255 3.13241
R979 VSS.n492 VSS.n491 2.88636
R980 VSS.n289 VSS.n254 2.88636
R981 VSS.n375 VSS.t51 2.87953
R982 VSS.n390 VSS.t95 2.87839
R983 VSS.t60 VSS.n161 2.87611
R984 VSS.n411 VSS.t5 2.87497
R985 VSS.n63 VSS.n62 2.86007
R986 VSS.n271 VSS.n270 2.86007
R987 VSS.n233 VSS.n232 2.7239
R988 VSS.n212 VSS.n211 2.7239
R989 VSS.n116 VSS.n115 2.7239
R990 VSS.n80 VSS.n79 2.7239
R991 VSS.n60 VSS.n59 2.7239
R992 VSS.n483 VSS.n482 2.7239
R993 VSS.n268 VSS.n267 2.7239
R994 VSS.n256 VSS.n255 2.7239
R995 VSS VSS.n22 2.56367
R996 VSS.n546 VSS.n545 2.44167
R997 VSS.n552 VSS.n551 2.03666
R998 VSS.n551 VSS.n20 1.77451
R999 VSS.n122 VSS.n121 1.753
R1000 VSS.n120 VSS.n119 1.753
R1001 VSS.n239 VSS.n238 1.753
R1002 VSS.n237 VSS.n236 1.753
R1003 VSS.n551 VSS.n550 1.44312
R1004 VSS.n547 VSS.n22 1.318
R1005 VSS.n493 VSS.n492 1.21169
R1006 VSS.n290 VSS.n289 1.21169
R1007 VSS.n189 VSS.n177 1.15795
R1008 VSS.n547 VSS.n546 1.07775
R1009 VSS.n238 VSS 0.95037
R1010 VSS.n238 VSS.n237 0.761313
R1011 VSS.n121 VSS.n120 0.761313
R1012 VSS.t50 VSS.n348 0.679804
R1013 VSS.n121 VSS.n24 0.591917
R1014 VSS.n492 VSS 0.531208
R1015 VSS.n289 VSS 0.531208
R1016 VSS.n428 VSS.n21 0.467019
R1017 VSS.n542 VSS.n541 0.467019
R1018 VSS.n405 VSS.n158 0.467019
R1019 VSS.n545 VSS.n24 0.4235
R1020 VSS.n230 VSS.n229 0.409011
R1021 VSS.n224 VSS.n212 0.409011
R1022 VSS.n113 VSS.n112 0.409011
R1023 VSS.n107 VSS.n80 0.409011
R1024 VSS.n66 VSS.n55 0.409011
R1025 VSS.n489 VSS.n488 0.409011
R1026 VSS.n487 VSS.n137 0.409011
R1027 VSS.n482 VSS.n481 0.409011
R1028 VSS.n264 VSS.n262 0.409011
R1029 VSS.n302 VSS.n208 0.409011
R1030 VSS.n299 VSS.n298 0.409011
R1031 VSS.n294 VSS.n256 0.409011
R1032 VSS.n331 VSS 0.26347
R1033 VSS.n406 VSS.n23 0.198729
R1034 VSS.n544 VSS.n543 0.198729
R1035 VSS.n550 VSS.n548 0.194976
R1036 VSS VSS.n22 0.16375
R1037 VSS.n508 VSS.n53 0.1255
R1038 VSS.n571 VSS.n6 0.1255
R1039 VSS.n133 VSS.n77 0.120292
R1040 VSS.n134 VSS.n133 0.120292
R1041 VSS.n135 VSS.n134 0.120292
R1042 VSS.n485 VSS.n138 0.120292
R1043 VSS.n70 VSS.n69 0.120292
R1044 VSS.n500 VSS.n69 0.120292
R1045 VSS.n502 VSS.n501 0.120292
R1046 VSS.n65 VSS.n64 0.120292
R1047 VSS.n64 VSS.n56 0.120292
R1048 VSS.n58 VSS.n56 0.120292
R1049 VSS.n127 VSS.n78 0.120292
R1050 VSS.n123 VSS.n78 0.120292
R1051 VSS.n104 VSS.n81 0.120292
R1052 VSS.n104 VSS.n103 0.120292
R1053 VSS.n102 VSS.n83 0.120292
R1054 VSS.n84 VSS.n83 0.120292
R1055 VSS.n95 VSS.n86 0.120292
R1056 VSS.n95 VSS.n94 0.120292
R1057 VSS.n93 VSS.n88 0.120292
R1058 VSS.n89 VSS.n88 0.120292
R1059 VSS.n111 VSS.n109 0.120292
R1060 VSS.n118 VSS.n110 0.120292
R1061 VSS.n244 VSS.n210 0.120292
R1062 VSS.n240 VSS.n210 0.120292
R1063 VSS.n221 VSS.n213 0.120292
R1064 VSS.n221 VSS.n220 0.120292
R1065 VSS.n219 VSS.n216 0.120292
R1066 VSS.n216 VSS.n215 0.120292
R1067 VSS.n580 VSS.n2 0.120292
R1068 VSS.n580 VSS.n579 0.120292
R1069 VSS.n578 VSS.n4 0.120292
R1070 VSS.n574 VSS.n4 0.120292
R1071 VSS.n228 VSS.n226 0.120292
R1072 VSS.n235 VSS.n227 0.120292
R1073 VSS.n246 VSS.n209 0.120292
R1074 VSS.n252 VSS.n209 0.120292
R1075 VSS.n253 VSS.n252 0.120292
R1076 VSS.n296 VSS.n295 0.120292
R1077 VSS.n284 VSS.n283 0.120292
R1078 VSS.n283 VSS.n261 0.120292
R1079 VSS.n279 VSS.n278 0.120292
R1080 VSS.n273 VSS.n272 0.120292
R1081 VSS.n272 VSS.n263 0.120292
R1082 VSS.n266 VSS.n263 0.120292
R1083 VSS VSS.n485 0.0981562
R1084 VSS.n296 VSS 0.0981562
R1085 VSS VSS.n128 0.09425
R1086 VSS.n245 VSS 0.09425
R1087 VSS.n237 VSS 0.0881354
R1088 VSS.n120 VSS 0.0881354
R1089 VSS.n550 VSS.n21 0.0766574
R1090 VSS.n543 VSS.n542 0.0766574
R1091 VSS.n406 VSS.n405 0.0766574
R1092 VSS.n119 VSS.n118 0.0721146
R1093 VSS.n236 VSS.n235 0.0721146
R1094 VSS.n494 VSS.n493 0.0708125
R1095 VSS.n290 VSS.n288 0.0708125
R1096 VSS.n545 VSS.n544 0.0654424
R1097 VSS.n407 VSS 0.064875
R1098 VSS.n429 VSS 0.064875
R1099 VSS.n438 VSS 0.064875
R1100 VSS.n27 VSS 0.064875
R1101 VSS.n26 VSS 0.064875
R1102 VSS.n25 VSS 0.064875
R1103 VSS.n549 VSS 0.064875
R1104 VSS.n386 VSS 0.064875
R1105 VSS.n404 VSS 0.064875
R1106 VSS.n427 VSS 0.063625
R1107 VSS.n540 VSS 0.063625
R1108 VSS.n371 VSS 0.063625
R1109 VSS.n123 VSS.n122 0.0616979
R1110 VSS.n240 VSS.n239 0.0616979
R1111 VSS.n552 VSS 0.061125
R1112 VSS.n20 VSS 0.061125
R1113 VSS.n135 VSS 0.0603958
R1114 VSS.n486 VSS 0.0603958
R1115 VSS.n139 VSS 0.0603958
R1116 VSS VSS.n74 0.0603958
R1117 VSS.n494 VSS 0.0603958
R1118 VSS VSS.n71 0.0603958
R1119 VSS VSS.n70 0.0603958
R1120 VSS.n501 VSS 0.0603958
R1121 VSS.n502 VSS 0.0603958
R1122 VSS.n65 VSS 0.0603958
R1123 VSS.n81 VSS 0.0603958
R1124 VSS VSS.n102 0.0603958
R1125 VSS.n85 VSS 0.0603958
R1126 VSS.n86 VSS 0.0603958
R1127 VSS VSS.n93 0.0603958
R1128 VSS VSS.n54 0.0603958
R1129 VSS.n111 VSS 0.0603958
R1130 VSS.n213 VSS 0.0603958
R1131 VSS VSS.n219 0.0603958
R1132 VSS VSS.n1 0.0603958
R1133 VSS.n2 VSS 0.0603958
R1134 VSS VSS.n578 0.0603958
R1135 VSS VSS.n573 0.0603958
R1136 VSS.n228 VSS 0.0603958
R1137 VSS VSS.n253 0.0603958
R1138 VSS VSS.n300 0.0603958
R1139 VSS.n292 VSS 0.0603958
R1140 VSS VSS.n291 0.0603958
R1141 VSS.n288 VSS 0.0603958
R1142 VSS.n285 VSS 0.0603958
R1143 VSS VSS.n284 0.0603958
R1144 VSS.n279 VSS 0.0603958
R1145 VSS.n278 VSS 0.0603958
R1146 VSS VSS.n273 0.0603958
R1147 VSS.n506 VSS 0.0590938
R1148 VSS.n122 VSS.n108 0.0590938
R1149 VSS.n239 VSS.n225 0.0590938
R1150 VSS VSS.n7 0.0590938
R1151 VSS.n493 VSS.n74 0.0499792
R1152 VSS.n291 VSS.n290 0.0499792
R1153 VSS.n119 VSS.n109 0.0486771
R1154 VSS.n236 VSS.n226 0.0486771
R1155 VSS.n491 VSS 0.0460729
R1156 VSS.n254 VSS 0.0460729
R1157 VSS.n546 VSS.n23 0.0416941
R1158 VSS.n548 VSS.n547 0.040297
R1159 VSS.n490 VSS 0.0343542
R1160 VSS.n301 VSS 0.0343542
R1161 VSS.n139 VSS 0.0330521
R1162 VSS VSS.n85 0.0330521
R1163 VSS VSS.n1 0.0330521
R1164 VSS.n292 VSS 0.0330521
R1165 VSS VSS.n53 0.03175
R1166 VSS VSS.n6 0.03175
R1167 VSS.n24 VSS 0.0292529
R1168 VSS.n486 VSS 0.0226354
R1169 VSS VSS.n138 0.0226354
R1170 VSS.n71 VSS 0.0226354
R1171 VSS VSS.n500 0.0226354
R1172 VSS.n505 VSS 0.0226354
R1173 VSS.n58 VSS 0.0226354
R1174 VSS.n108 VSS 0.0226354
R1175 VSS.n103 VSS 0.0226354
R1176 VSS VSS.n84 0.0226354
R1177 VSS.n94 VSS 0.0226354
R1178 VSS.n89 VSS 0.0226354
R1179 VSS.n110 VSS 0.0226354
R1180 VSS.n225 VSS 0.0226354
R1181 VSS.n220 VSS 0.0226354
R1182 VSS.n215 VSS 0.0226354
R1183 VSS.n579 VSS 0.0226354
R1184 VSS.n574 VSS 0.0226354
R1185 VSS.n227 VSS 0.0226354
R1186 VSS.n300 VSS 0.0226354
R1187 VSS.n295 VSS 0.0226354
R1188 VSS.n285 VSS 0.0226354
R1189 VSS VSS.n261 0.0226354
R1190 VSS.n274 VSS 0.0226354
R1191 VSS.n266 VSS 0.0226354
R1192 VSS.n491 VSS.n490 0.0148229
R1193 VSS.n301 VSS.n254 0.0148229
R1194 VSS.n128 VSS.n77 0.00440625
R1195 VSS.n246 VSS.n245 0.00440625
R1196 VSS.n506 VSS.n505 0.00180208
R1197 VSS.n54 VSS.n53 0.00180208
R1198 VSS.n573 VSS.n6 0.00180208
R1199 VSS.n274 VSS.n7 0.00180208
R1200 x1.x3.GP4.n3 x1.x3.GP4.t6 450.938
R1201 x1.x3.GP4.n2 x1.x3.GP4.t7 450.938
R1202 x1.x3.GP4.n3 x1.x3.GP4.t4 445.666
R1203 x1.x3.GP4.n2 x1.x3.GP4.t5 445.666
R1204 x1.x1.x14.Y x1.x3.GP4.n6 203.923
R1205 x1.x3.GP4.n0 x1.x3.GP4.n1 101.49
R1206 x1.x3.GP4.n6 x1.x3.GP4.t0 26.5955
R1207 x1.x3.GP4.n6 x1.x3.GP4.t3 26.5955
R1208 x1.x3.GP4.n1 x1.x3.GP4.t2 24.9236
R1209 x1.x3.GP4.n1 x1.x3.GP4.t1 24.9236
R1210 x1.x3.GP4.n4 x1.x3.x4.GP 11.0619
R1211 x1.x3.GP4.n5 x1.x1.x14.Y 10.7525
R1212 x1.x1.gpo3 x1.x3.GP4.n4 9.34192
R1213 x1.x3.GP4.n0 x1.x1.gpo3 7.73829
R1214 x1.x3.GP4.n5 x1.x1.x14.Y 6.6565
R1215 x1.x3.GP4.n4 x1.x2.x4.GP 5.84951
R1216 x1.x1.x14.Y x1.x3.GP4.n5 5.04292
R1217 x1.x2.x4.GP x1.x3.GP4.n3 2.95993
R1218 x1.x3.x4.GP x1.x3.GP4.n2 2.95993
R1219 x1.x1.x14.Y x1.x3.GP4.n0 2.5605
R1220 x1.x3.GP4.n0 x1.x1.x14.Y 1.93989
R1221 x1.x5.A.n15 x1.x5.A.t7 26.3998
R1222 x1.x5.A.n18 x1.x5.A.t10 23.6581
R1223 x1.x5.A.n11 x1.x5.A.t4 23.6581
R1224 x1.x5.A.n9 x1.x5.A.t17 23.6581
R1225 x1.x5.A.n13 x1.x5.A.t16 23.6581
R1226 x1.x5.A.n15 x1.x5.A.t11 23.5483
R1227 x1.x5.A.n0 x1.x5.A.t3 23.3739
R1228 x1.x5.A.n2 x1.x5.A.t18 23.3739
R1229 x1.x5.A.n4 x1.x5.A.t0 23.3739
R1230 x1.x5.A.n6 x1.x5.A.t6 23.3739
R1231 x1.x5.A.n16 x1.x5.A.t12 12.7127
R1232 x1.x5.A.n16 x1.x5.A.t13 10.8578
R1233 x1.x5.A.n11 x1.x5.A.t2 10.7528
R1234 x1.x5.A.n9 x1.x5.A.t14 10.7528
R1235 x1.x5.A.n13 x1.x5.A.t5 10.7528
R1236 x1.x5.A.n18 x1.x5.A.t9 10.7528
R1237 x1.x5.A.n17 x1.x5.A.n15 3.06895
R1238 x1.x5.A.n12 x1.x5.A 1.85764
R1239 x1.x5.A.n17 x1.x5.A.n16 1.84731
R1240 x1.x5.A.n1 x1.x5.A.n11 1.5062
R1241 x1.x5.A.n3 x1.x5.A.n9 1.5062
R1242 x1.x5.A.n5 x1.x5.A.n13 1.5062
R1243 x1.x5.A.n14 x1.x5.A 1.28884
R1244 x1.x5.A.n8 x1.x5.A.n14 1.26452
R1245 x1.x5.A x1.x5.A.n0 1.26165
R1246 x1.x5.A.n8 x1.x5.A.n10 1.254
R1247 x1.x5.A.n10 x1.x5.A.n12 1.25206
R1248 x1.x5.A x1.x5.A.n17 1.12636
R1249 x1.x5.A x1.x5.A.n4 0.983856
R1250 x1.x5.A x1.x5.A.n6 0.936641
R1251 x1.x5.A x1.x5.A.n2 0.924585
R1252 x1.x5.A.n0 x1.x5.A.n1 0.231183
R1253 x1.x5.A.n2 x1.x5.A.n3 0.231183
R1254 x1.x5.A.n4 x1.x5.A.n5 0.231183
R1255 x1.x5.A.n7 x1.x5.A.n6 0.231183
R1256 x1.x5.A.n7 x1.x5.A.t8 10.8045
R1257 x1.x5.A.n7 x1.x5.A.n18 1.5062
R1258 x1.x5.A.n5 x1.x5.A.t19 10.8045
R1259 x1.x5.A.n3 x1.x5.A.t15 10.8045
R1260 x1.x5.A.n1 x1.x5.A.t1 10.8045
R1261 x1.x5.A.n12 x1.x5.A 0.416271
R1262 x1.x5.A x1.x5.A.n8 0.260839
R1263 x1.x5.A.n14 x1.x5.A 0.257416
R1264 x1.x5.A.n10 x1.x5.A 0.237533
R1265 R4R5.n1 R4R5.t2 26.3998
R1266 R4R5.n1 R4R5.t3 23.5483
R1267 R4R5.n0 R4R5.t0 12.7127
R1268 R4R5.n4 R4R5.t4 10.8674
R1269 R4R5.n0 R4R5.t1 10.8578
R1270 R4R5.n4 R4R5.t5 10.5285
R1271 R4R5.n2 R4R5.n1 3.12177
R1272 R4R5.n2 R4R5.n0 1.81453
R1273 R4R5.n3 R4R5.n2 1.1255
R1274 R4R5.n5 R4R5.n4 0.785021
R1275 R4R5 R4R5.n3 0.134513
R1276 R4R5.n3 R4R5 0.0655
R1277 R4R5 R4R5.n5 0.053625
R1278 R4R5.n5 R4R5 0.0055
R1279 VDD.n344 VDD.n342 8629.41
R1280 VDD.n347 VDD.n341 8629.41
R1281 VDD.n329 VDD.n328 8629.41
R1282 VDD.n331 VDD.n326 8629.41
R1283 VDD.n312 VDD.n311 8629.41
R1284 VDD.n314 VDD.n309 8629.41
R1285 VDD.n295 VDD.n293 8629.41
R1286 VDD.n298 VDD.n292 8629.41
R1287 VDD.n230 VDD.n223 8629.41
R1288 VDD.n227 VDD.n224 8629.41
R1289 VDD.n272 VDD.n271 8629.41
R1290 VDD.n274 VDD.n269 8629.41
R1291 VDD.n255 VDD.n254 8629.41
R1292 VDD.n257 VDD.n252 8629.41
R1293 VDD.n238 VDD.n236 8629.41
R1294 VDD.n241 VDD.n235 8629.41
R1295 VDD.n201 VDD.n195 8629.41
R1296 VDD.n201 VDD.n196 8629.41
R1297 VDD.n199 VDD.n195 8629.41
R1298 VDD.n199 VDD.n196 8629.41
R1299 VDD.n214 VDD.n208 8629.41
R1300 VDD.n214 VDD.n209 8629.41
R1301 VDD.n212 VDD.n208 8629.41
R1302 VDD.n212 VDD.n209 8629.41
R1303 VDD.n57 VDD.n55 8629.41
R1304 VDD.n60 VDD.n54 8629.41
R1305 VDD.n40 VDD.n39 8629.41
R1306 VDD.n42 VDD.n37 8629.41
R1307 VDD.n23 VDD.n22 8629.41
R1308 VDD.n25 VDD.n20 8629.41
R1309 VDD.n6 VDD.n4 8629.41
R1310 VDD.n9 VDD.n3 8629.41
R1311 VDD.n201 VDD.t90 2459.29
R1312 VDD.t89 VDD.n199 2459.29
R1313 VDD.n214 VDD.t55 2459.29
R1314 VDD.t74 VDD.n212 2459.29
R1315 VDD.t90 VDD.n200 2298.92
R1316 VDD.n200 VDD.t89 2298.92
R1317 VDD.t55 VDD.n213 2298.92
R1318 VDD.n213 VDD.t74 2298.92
R1319 VDD.n343 VDD.n340 920.471
R1320 VDD.n332 VDD.n325 920.471
R1321 VDD.n315 VDD.n308 920.471
R1322 VDD.n294 VDD.n291 920.471
R1323 VDD.n226 VDD.n225 920.471
R1324 VDD.n275 VDD.n268 920.471
R1325 VDD.n258 VDD.n251 920.471
R1326 VDD.n237 VDD.n234 920.471
R1327 VDD.n198 VDD.n197 920.471
R1328 VDD.n211 VDD.n210 920.471
R1329 VDD.n56 VDD.n53 920.471
R1330 VDD.n43 VDD.n36 920.471
R1331 VDD.n26 VDD.n19 920.471
R1332 VDD.n5 VDD.n2 920.471
R1333 VDD.n349 VDD.n340 914.447
R1334 VDD.n334 VDD.n332 914.447
R1335 VDD.n317 VDD.n315 914.447
R1336 VDD.n300 VDD.n291 914.447
R1337 VDD.n225 VDD.n222 914.447
R1338 VDD.n277 VDD.n275 914.447
R1339 VDD.n260 VDD.n258 914.447
R1340 VDD.n243 VDD.n234 914.447
R1341 VDD.n197 VDD.n193 914.447
R1342 VDD.n210 VDD.n206 914.447
R1343 VDD.n62 VDD.n53 914.447
R1344 VDD.n45 VDD.n43 914.447
R1345 VDD.n28 VDD.n26 914.447
R1346 VDD.n11 VDD.n2 914.447
R1347 VDD.t4 VDD.n126 804.731
R1348 VDD.t7 VDD.n417 804.731
R1349 VDD.n128 VDD.t4 751.692
R1350 VDD.n419 VDD.t7 751.692
R1351 VDD.n100 VDD.t114 671.408
R1352 VDD.n89 VDD.t29 671.408
R1353 VDD.n391 VDD.t112 671.408
R1354 VDD.n380 VDD.t149 671.408
R1355 VDD VDD.t3 630.375
R1356 VDD VDD.t6 630.375
R1357 VDD.n159 VDD.n158 602.456
R1358 VDD.n181 VDD.n69 602.456
R1359 VDD.n450 VDD.n449 602.456
R1360 VDD.n472 VDD.n360 602.456
R1361 VDD.n73 VDD.n72 585
R1362 VDD.n75 VDD.n74 585
R1363 VDD.n364 VDD.n363 585
R1364 VDD.n366 VDD.n365 585
R1365 VDD.n198 VDD.n194 480.764
R1366 VDD.n211 VDD.n207 480.764
R1367 VDD.n343 VDD.n339 480.764
R1368 VDD.n325 VDD.n323 480.764
R1369 VDD.n308 VDD.n306 480.764
R1370 VDD.n294 VDD.n289 480.764
R1371 VDD.n226 VDD.n221 480.764
R1372 VDD.n268 VDD.n266 480.764
R1373 VDD.n251 VDD.n249 480.764
R1374 VDD.n237 VDD.n233 480.764
R1375 VDD.n56 VDD.n51 480.764
R1376 VDD.n36 VDD.n34 480.764
R1377 VDD.n19 VDD.n17 480.764
R1378 VDD.n5 VDD.n1 480.764
R1379 VDD VDD.t21 458.724
R1380 VDD.t3 VDD 458.724
R1381 VDD VDD.t0 458.724
R1382 VDD.t6 VDD 458.724
R1383 VDD.n121 VDD.t78 420.25
R1384 VDD.n412 VDD.t72 420.25
R1385 VDD.n117 VDD.t22 388.656
R1386 VDD.n152 VDD.t23 388.656
R1387 VDD.n130 VDD.t5 388.656
R1388 VDD.n103 VDD.t13 388.656
R1389 VDD.n112 VDD.t14 388.656
R1390 VDD.n77 VDD.t19 388.656
R1391 VDD.n82 VDD.t20 388.656
R1392 VDD.n408 VDD.t1 388.656
R1393 VDD.n443 VDD.t2 388.656
R1394 VDD.n421 VDD.t8 388.656
R1395 VDD.n394 VDD.t10 388.656
R1396 VDD.n403 VDD.t11 388.656
R1397 VDD.n368 VDD.t16 388.656
R1398 VDD.n373 VDD.t17 388.656
R1399 VDD.n351 VDD.n339 379.2
R1400 VDD.n336 VDD.n323 379.2
R1401 VDD.n319 VDD.n306 379.2
R1402 VDD.n302 VDD.n289 379.2
R1403 VDD.n285 VDD.n221 379.2
R1404 VDD.n279 VDD.n266 379.2
R1405 VDD.n262 VDD.n249 379.2
R1406 VDD.n245 VDD.n233 379.2
R1407 VDD.n203 VDD.n194 379.2
R1408 VDD.n216 VDD.n207 379.2
R1409 VDD.n64 VDD.n51 379.2
R1410 VDD.n47 VDD.n34 379.2
R1411 VDD.n30 VDD.n17 379.2
R1412 VDD.n13 VDD.n1 379.2
R1413 VDD VDD.t119 369.938
R1414 VDD VDD.t47 369.938
R1415 VDD VDD.t143 369.938
R1416 VDD VDD.t132 369.938
R1417 VDD.n106 VDD.n99 322.329
R1418 VDD.n84 VDD.n80 322.329
R1419 VDD.n397 VDD.n390 322.329
R1420 VDD.n375 VDD.n371 322.329
R1421 VDD.n163 VDD.n161 259.697
R1422 VDD.n454 VDD.n452 259.697
R1423 VDD.n139 VDD.t48 255.905
R1424 VDD.n144 VDD.t120 255.905
R1425 VDD.n120 VDD.t79 255.905
R1426 VDD.n160 VDD.t145 255.905
R1427 VDD.n430 VDD.t133 255.905
R1428 VDD.n435 VDD.t144 255.905
R1429 VDD.n411 VDD.t73 255.905
R1430 VDD.n451 VDD.t94 255.905
R1431 VDD.n110 VDD.t129 254.475
R1432 VDD.n401 VDD.t61 254.475
R1433 VDD.n135 VDD.t46 252.95
R1434 VDD.n140 VDD.t106 252.95
R1435 VDD.n145 VDD.t82 252.95
R1436 VDD.n180 VDD.t126 252.95
R1437 VDD.n426 VDD.t76 252.95
R1438 VDD.n431 VDD.t118 252.95
R1439 VDD.n436 VDD.t71 252.95
R1440 VDD.n471 VDD.t67 252.95
R1441 VDD.n159 VDD.t151 251.516
R1442 VDD.n450 VDD.t108 251.516
R1443 VDD.n70 VDD.t52 250.724
R1444 VDD.n68 VDD.t124 250.724
R1445 VDD.n361 VDD.t27 250.724
R1446 VDD.n359 VDD.t65 250.724
R1447 VDD.t78 VDD.t81 248.599
R1448 VDD.t119 VDD.t105 248.599
R1449 VDD.t47 VDD.t45 248.599
R1450 VDD.t72 VDD.t70 248.599
R1451 VDD.t143 VDD.t117 248.599
R1452 VDD.t132 VDD.t75 248.599
R1453 VDD.n175 VDD.t63 248.219
R1454 VDD.n162 VDD.t147 248.219
R1455 VDD.n466 VDD.t137 248.219
R1456 VDD.n453 VDD.t96 248.219
R1457 VDD.n121 VDD 221.964
R1458 VDD.n412 VDD 221.964
R1459 VDD.n128 VDD.t152 215.827
R1460 VDD.n419 VDD.t158 215.827
R1461 VDD.n110 VDD.n109 213.119
R1462 VDD.n401 VDD.n400 213.119
R1463 VDD.n150 VDD.n121 213.119
R1464 VDD.n441 VDD.n412 213.119
R1465 VDD.n188 VDD.t80 212.081
R1466 VDD.n187 VDD.t77 212.081
R1467 VDD.n118 VDD.t155 210.964
R1468 VDD.n104 VDD.t157 210.964
R1469 VDD.n79 VDD.t156 210.964
R1470 VDD.n409 VDD.t160 210.964
R1471 VDD.n395 VDD.t154 210.964
R1472 VDD.n370 VDD.t153 210.964
R1473 VDD.n170 VDD.n169 209.368
R1474 VDD.n461 VDD.n460 209.368
R1475 VDD.t81 VDD 198.287
R1476 VDD.t105 VDD 198.287
R1477 VDD.t45 VDD 198.287
R1478 VDD.t70 VDD 198.287
R1479 VDD.t117 VDD 198.287
R1480 VDD.t75 VDD 198.287
R1481 VDD.n172 VDD.n171 183.673
R1482 VDD.n463 VDD.n462 183.673
R1483 VDD.n189 VDD.n188 183.441
R1484 VDD VDD.t36 182.952
R1485 VDD VDD.n170 182.952
R1486 VDD.t91 VDD 182.952
R1487 VDD VDD.t56 182.952
R1488 VDD VDD.n461 182.952
R1489 VDD.t138 VDD 182.952
R1490 VDD.n74 VDD.n73 159.476
R1491 VDD.n365 VDD.n364 159.476
R1492 VDD.n161 VDD.t25 157.014
R1493 VDD.n452 VDD.t102 157.014
R1494 VDD.t51 VDD.t38 154.417
R1495 VDD.t26 VDD.t68 154.417
R1496 VDD.t130 VDD.t24 147.703
R1497 VDD.t140 VDD.t93 147.703
R1498 VDD.t103 VDD.t113 140.989
R1499 VDD.t24 VDD.t146 140.989
R1500 VDD.t125 VDD.t123 140.989
R1501 VDD.t62 VDD.t51 140.989
R1502 VDD.t28 VDD.t121 140.989
R1503 VDD.t30 VDD.t111 140.989
R1504 VDD.t93 VDD.t95 140.989
R1505 VDD.t66 VDD.t64 140.989
R1506 VDD.t136 VDD.t26 140.989
R1507 VDD.t148 VDD.t109 140.989
R1508 VDD.n188 VDD.t159 139.78
R1509 VDD.n187 VDD.t161 139.78
R1510 VDD.n161 VDD.t98 137.079
R1511 VDD.n452 VDD.t43 137.079
R1512 VDD.n109 VDD 125.883
R1513 VDD.n171 VDD 125.883
R1514 VDD.n400 VDD 125.883
R1515 VDD.n462 VDD 125.883
R1516 VDD.n99 VDD.t104 116.341
R1517 VDD.n80 VDD.t122 116.341
R1518 VDD.n390 VDD.t31 116.341
R1519 VDD.n371 VDD.t110 116.341
R1520 VDD.t113 VDD 112.457
R1521 VDD.t146 VDD 112.457
R1522 VDD VDD.t28 112.457
R1523 VDD.t111 VDD 112.457
R1524 VDD.t95 VDD 112.457
R1525 VDD VDD.t148 112.457
R1526 VDD VDD.t115 109.1
R1527 VDD VDD.t40 109.1
R1528 VDD.n204 VDD.n193 105.788
R1529 VDD.n217 VDD.n206 105.788
R1530 VDD.t12 VDD.t103 104.064
R1531 VDD.t121 VDD.t18 104.064
R1532 VDD.t9 VDD.t30 104.064
R1533 VDD.t109 VDD.t15 104.064
R1534 VDD.t53 VDD 102.385
R1535 VDD.t99 VDD 102.385
R1536 VDD.t128 VDD 99.0288
R1537 VDD.t60 VDD 99.0288
R1538 VDD.n158 VDD.t131 96.1553
R1539 VDD.n69 VDD.t88 96.1553
R1540 VDD.n449 VDD.t141 96.1553
R1541 VDD.n360 VDD.t86 96.1553
R1542 VDD VDD.t87 92.315
R1543 VDD VDD.t85 92.315
R1544 VDD.n73 VDD.t39 86.7743
R1545 VDD.n364 VDD.t69 86.7743
R1546 VDD.n109 VDD.t128 83.9228
R1547 VDD.n400 VDD.t60 83.9228
R1548 VDD.n170 VDD.t97 80.5659
R1549 VDD.n461 VDD.t42 80.5659
R1550 VDD.t36 VDD.t12 77.209
R1551 VDD.t18 VDD.t91 77.209
R1552 VDD.t56 VDD.t9 77.209
R1553 VDD.t15 VDD.t138 77.209
R1554 VDD.n74 VDD.t116 66.8398
R1555 VDD.n365 VDD.t41 66.8398
R1556 VDD.n350 VDD.n349 66.6358
R1557 VDD.n335 VDD.n334 66.6358
R1558 VDD.n318 VDD.n317 66.6358
R1559 VDD.n301 VDD.n300 66.6358
R1560 VDD.n284 VDD.n222 66.6358
R1561 VDD.n278 VDD.n277 66.6358
R1562 VDD.n261 VDD.n260 66.6358
R1563 VDD.n244 VDD.n243 66.6358
R1564 VDD.n63 VDD.n62 66.6358
R1565 VDD.n46 VDD.n45 66.6358
R1566 VDD.n29 VDD.n28 66.6358
R1567 VDD.n12 VDD.n11 66.6358
R1568 VDD.n203 VDD.n202 63.3551
R1569 VDD.n216 VDD.n215 63.3551
R1570 VDD.n158 VDD.t54 63.3219
R1571 VDD.n69 VDD.t50 63.3219
R1572 VDD.n449 VDD.t100 63.3219
R1573 VDD.n360 VDD.t59 63.3219
R1574 VDD VDD.t130 62.103
R1575 VDD VDD.t140 62.103
R1576 VDD.n344 VDD.n343 61.6672
R1577 VDD.n348 VDD.n347 61.6672
R1578 VDD.n329 VDD.n325 61.6672
R1579 VDD.n326 VDD.n324 61.6672
R1580 VDD.n312 VDD.n308 61.6672
R1581 VDD.n309 VDD.n307 61.6672
R1582 VDD.n295 VDD.n294 61.6672
R1583 VDD.n299 VDD.n298 61.6672
R1584 VDD.n231 VDD.n230 61.6672
R1585 VDD.n227 VDD.n226 61.6672
R1586 VDD.n272 VDD.n268 61.6672
R1587 VDD.n269 VDD.n267 61.6672
R1588 VDD.n255 VDD.n251 61.6672
R1589 VDD.n252 VDD.n250 61.6672
R1590 VDD.n238 VDD.n237 61.6672
R1591 VDD.n242 VDD.n241 61.6672
R1592 VDD.n199 VDD.n198 61.6672
R1593 VDD.n202 VDD.n201 61.6672
R1594 VDD.n212 VDD.n211 61.6672
R1595 VDD.n215 VDD.n214 61.6672
R1596 VDD.n57 VDD.n56 61.6672
R1597 VDD.n61 VDD.n60 61.6672
R1598 VDD.n40 VDD.n36 61.6672
R1599 VDD.n37 VDD.n35 61.6672
R1600 VDD.n23 VDD.n19 61.6672
R1601 VDD.n20 VDD.n18 61.6672
R1602 VDD.n6 VDD.n5 61.6672
R1603 VDD.n10 VDD.n9 61.6672
R1604 VDD.n188 VDD.n187 61.346
R1605 VDD.n345 VDD.n344 60.9564
R1606 VDD.n347 VDD.n346 60.9564
R1607 VDD.n330 VDD.n329 60.9564
R1608 VDD.n327 VDD.n326 60.9564
R1609 VDD.n313 VDD.n312 60.9564
R1610 VDD.n310 VDD.n309 60.9564
R1611 VDD.n296 VDD.n295 60.9564
R1612 VDD.n298 VDD.n297 60.9564
R1613 VDD.n230 VDD.n229 60.9564
R1614 VDD.n228 VDD.n227 60.9564
R1615 VDD.n273 VDD.n272 60.9564
R1616 VDD.n270 VDD.n269 60.9564
R1617 VDD.n256 VDD.n255 60.9564
R1618 VDD.n253 VDD.n252 60.9564
R1619 VDD.n239 VDD.n238 60.9564
R1620 VDD.n241 VDD.n240 60.9564
R1621 VDD.n58 VDD.n57 60.9564
R1622 VDD.n60 VDD.n59 60.9564
R1623 VDD.n41 VDD.n40 60.9564
R1624 VDD.n38 VDD.n37 60.9564
R1625 VDD.n24 VDD.n23 60.9564
R1626 VDD.n21 VDD.n20 60.9564
R1627 VDD.n7 VDD.n6 60.9564
R1628 VDD.n9 VDD.n8 60.9564
R1629 VDD.n335 VDD.n324 60.6123
R1630 VDD.n318 VDD.n307 60.6123
R1631 VDD.n278 VDD.n267 60.6123
R1632 VDD.n261 VDD.n250 60.6123
R1633 VDD.n46 VDD.n35 60.6123
R1634 VDD.n29 VDD.n18 60.6123
R1635 VDD.n350 VDD.n192 59.4829
R1636 VDD.n284 VDD.n283 59.4829
R1637 VDD.n63 VDD.n52 59.4829
R1638 VDD.n301 VDD.n290 58.7299
R1639 VDD.n244 VDD.n232 58.7299
R1640 VDD.n12 VDD.n0 58.7299
R1641 VDD.t38 VDD 55.3892
R1642 VDD.t68 VDD 55.3892
R1643 VDD.t49 VDD 52.0323
R1644 VDD.t58 VDD 52.0323
R1645 VDD VDD.t97 45.3185
R1646 VDD VDD.t42 45.3185
R1647 VDD VDD.t150 41.9616
R1648 VDD VDD.t107 41.9616
R1649 VDD.n345 VDD.n341 38.5759
R1650 VDD.n346 VDD.n342 38.5759
R1651 VDD.n331 VDD.n330 38.5759
R1652 VDD.n328 VDD.n327 38.5759
R1653 VDD.n314 VDD.n313 38.5759
R1654 VDD.n311 VDD.n310 38.5759
R1655 VDD.n296 VDD.n292 38.5759
R1656 VDD.n297 VDD.n293 38.5759
R1657 VDD.n228 VDD.n223 38.5759
R1658 VDD.n229 VDD.n224 38.5759
R1659 VDD.n274 VDD.n273 38.5759
R1660 VDD.n271 VDD.n270 38.5759
R1661 VDD.n257 VDD.n256 38.5759
R1662 VDD.n254 VDD.n253 38.5759
R1663 VDD.n239 VDD.n235 38.5759
R1664 VDD.n240 VDD.n236 38.5759
R1665 VDD.n58 VDD.n54 38.5759
R1666 VDD.n59 VDD.n55 38.5759
R1667 VDD.n42 VDD.n41 38.5759
R1668 VDD.n39 VDD.n38 38.5759
R1669 VDD.n25 VDD.n24 38.5759
R1670 VDD.n22 VDD.n21 38.5759
R1671 VDD.n7 VDD.n3 38.5759
R1672 VDD.n8 VDD.n4 38.5759
R1673 VDD.n169 VDD.n91 34.6358
R1674 VDD.n169 VDD.n92 34.6358
R1675 VDD.n174 VDD.n173 34.6358
R1676 VDD.n460 VDD.n382 34.6358
R1677 VDD.n460 VDD.n383 34.6358
R1678 VDD.n465 VDD.n464 34.6358
R1679 VDD.n171 VDD 28.5341
R1680 VDD.n462 VDD 28.5341
R1681 VDD.n99 VDD.t37 28.4453
R1682 VDD.n80 VDD.t92 28.4453
R1683 VDD.n390 VDD.t57 28.4453
R1684 VDD.n371 VDD.t139 28.4453
R1685 VDD.n176 VDD.n175 28.3534
R1686 VDD.n467 VDD.n466 28.3534
R1687 VDD.n173 VDD.n172 25.6953
R1688 VDD.n464 VDD.n463 25.6953
R1689 VDD.n139 VDD.n124 25.224
R1690 VDD.n135 VDD.n124 25.224
R1691 VDD.n144 VDD.n123 25.224
R1692 VDD.n140 VDD.n123 25.224
R1693 VDD.n146 VDD.n120 25.224
R1694 VDD.n146 VDD.n145 25.224
R1695 VDD.n164 VDD.n160 25.224
R1696 VDD.n430 VDD.n415 25.224
R1697 VDD.n426 VDD.n415 25.224
R1698 VDD.n435 VDD.n414 25.224
R1699 VDD.n431 VDD.n414 25.224
R1700 VDD.n437 VDD.n411 25.224
R1701 VDD.n437 VDD.n436 25.224
R1702 VDD.n455 VDD.n451 25.224
R1703 VDD.n110 VDD.n94 23.7181
R1704 VDD.n401 VDD.n385 23.7181
R1705 VDD VDD.n100 23.252
R1706 VDD VDD.n391 23.252
R1707 VDD.n159 VDD.n94 21.4593
R1708 VDD.n450 VDD.n385 21.4593
R1709 VDD.n140 VDD.n139 20.3299
R1710 VDD.n145 VDD.n144 20.3299
R1711 VDD.n431 VDD.n430 20.3299
R1712 VDD.n436 VDD.n435 20.3299
R1713 VDD.t87 VDD.t125 20.1418
R1714 VDD.t85 VDD.t66 20.1418
R1715 VDD.n181 VDD.n68 19.9534
R1716 VDD.n472 VDD.n359 19.9534
R1717 VDD.n180 VDD.n179 19.8181
R1718 VDD.n471 VDD.n470 19.8181
R1719 VDD.n150 VDD.n120 17.3181
R1720 VDD.n163 VDD.n162 17.3181
R1721 VDD.n441 VDD.n411 17.3181
R1722 VDD.n454 VDD.n453 17.3181
R1723 VDD.n160 VDD.n159 16.5652
R1724 VDD.n164 VDD.n163 16.5652
R1725 VDD.n451 VDD.n450 16.5652
R1726 VDD.n455 VDD.n454 16.5652
R1727 VDD.n135 VDD.n134 15.8123
R1728 VDD.n426 VDD.n425 15.8123
R1729 VDD.n151 VDD.n150 14.2735
R1730 VDD.n111 VDD.n110 14.2735
R1731 VDD.n442 VDD.n441 14.2735
R1732 VDD.n402 VDD.n401 14.2735
R1733 VDD.n173 VDD.n89 13.9299
R1734 VDD.n464 VDD.n380 13.9299
R1735 VDD.n181 VDD.n180 13.5534
R1736 VDD.n472 VDD.n471 13.5534
R1737 VDD.n116 VDD.n115 11.4366
R1738 VDD.n407 VDD.n406 11.4366
R1739 VDD VDD.n189 11.4331
R1740 VDD.n352 VDD.n351 11.3235
R1741 VDD.n337 VDD.n336 11.3235
R1742 VDD.n320 VDD.n319 11.3235
R1743 VDD.n303 VDD.n302 11.3235
R1744 VDD.n286 VDD.n285 11.3235
R1745 VDD.n280 VDD.n279 11.3235
R1746 VDD.n263 VDD.n262 11.3235
R1747 VDD.n246 VDD.n245 11.3235
R1748 VDD.n65 VDD.n64 11.3235
R1749 VDD.n48 VDD.n47 11.3235
R1750 VDD.n31 VDD.n30 11.3235
R1751 VDD.n14 VDD.n13 11.3235
R1752 VDD.n172 VDD.n90 11.2937
R1753 VDD.n463 VDD.n381 11.2937
R1754 VDD.n156 VDD.n155 11.2737
R1755 VDD.n447 VDD.n446 11.2737
R1756 VDD.n186 VDD.n66 10.2451
R1757 VDD.t150 VDD.t53 10.0712
R1758 VDD.t107 VDD.t99 10.0712
R1759 VDD.n130 VDD.n127 9.60526
R1760 VDD.n117 VDD.n116 9.60526
R1761 VDD.n82 VDD.n81 9.60526
R1762 VDD.n421 VDD.n418 9.60526
R1763 VDD.n408 VDD.n407 9.60526
R1764 VDD.n373 VDD.n372 9.60526
R1765 VDD.n119 VDD.n95 9.3005
R1766 VDD.n154 VDD.n153 9.3005
R1767 VDD.n151 VDD.n96 9.3005
R1768 VDD.n150 VDD.n149 9.3005
R1769 VDD.n145 VDD.n122 9.3005
R1770 VDD.n141 VDD.n140 9.3005
R1771 VDD.n136 VDD.n135 9.3005
R1772 VDD.n132 VDD.n131 9.3005
R1773 VDD.n137 VDD.n124 9.3005
R1774 VDD.n139 VDD.n138 9.3005
R1775 VDD.n142 VDD.n123 9.3005
R1776 VDD.n144 VDD.n143 9.3005
R1777 VDD.n147 VDD.n146 9.3005
R1778 VDD.n148 VDD.n120 9.3005
R1779 VDD.n177 VDD.n176 9.3005
R1780 VDD.n182 VDD.n181 9.3005
R1781 VDD.n166 VDD.n91 9.3005
R1782 VDD.n159 VDD.n157 9.3005
R1783 VDD.n110 VDD.n108 9.3005
R1784 VDD.n102 VDD.n101 9.3005
R1785 VDD.n105 VDD.n97 9.3005
R1786 VDD.n114 VDD.n113 9.3005
R1787 VDD.n111 VDD.n98 9.3005
R1788 VDD.n107 VDD.n94 9.3005
R1789 VDD.n160 VDD.n93 9.3005
R1790 VDD.n165 VDD.n164 9.3005
R1791 VDD.n169 VDD.n168 9.3005
R1792 VDD.n167 VDD.n92 9.3005
R1793 VDD.n180 VDD.n67 9.3005
R1794 VDD.n179 VDD.n178 9.3005
R1795 VDD.n174 VDD.n71 9.3005
R1796 VDD.n173 VDD.n76 9.3005
R1797 VDD.n88 VDD.n87 9.3005
R1798 VDD.n86 VDD.n85 9.3005
R1799 VDD.n83 VDD.n78 9.3005
R1800 VDD.n410 VDD.n386 9.3005
R1801 VDD.n445 VDD.n444 9.3005
R1802 VDD.n442 VDD.n387 9.3005
R1803 VDD.n441 VDD.n440 9.3005
R1804 VDD.n436 VDD.n413 9.3005
R1805 VDD.n432 VDD.n431 9.3005
R1806 VDD.n427 VDD.n426 9.3005
R1807 VDD.n423 VDD.n422 9.3005
R1808 VDD.n428 VDD.n415 9.3005
R1809 VDD.n430 VDD.n429 9.3005
R1810 VDD.n433 VDD.n414 9.3005
R1811 VDD.n435 VDD.n434 9.3005
R1812 VDD.n438 VDD.n437 9.3005
R1813 VDD.n439 VDD.n411 9.3005
R1814 VDD.n468 VDD.n467 9.3005
R1815 VDD.n473 VDD.n472 9.3005
R1816 VDD.n457 VDD.n382 9.3005
R1817 VDD.n450 VDD.n448 9.3005
R1818 VDD.n401 VDD.n399 9.3005
R1819 VDD.n393 VDD.n392 9.3005
R1820 VDD.n396 VDD.n388 9.3005
R1821 VDD.n405 VDD.n404 9.3005
R1822 VDD.n402 VDD.n389 9.3005
R1823 VDD.n398 VDD.n385 9.3005
R1824 VDD.n451 VDD.n384 9.3005
R1825 VDD.n456 VDD.n455 9.3005
R1826 VDD.n460 VDD.n459 9.3005
R1827 VDD.n458 VDD.n383 9.3005
R1828 VDD.n471 VDD.n358 9.3005
R1829 VDD.n470 VDD.n469 9.3005
R1830 VDD.n465 VDD.n362 9.3005
R1831 VDD.n464 VDD.n367 9.3005
R1832 VDD.n379 VDD.n378 9.3005
R1833 VDD.n377 VDD.n376 9.3005
R1834 VDD.n374 VDD.n369 9.3005
R1835 VDD.n247 VDD.n232 8.23557
R1836 VDD.n15 VDD.n0 8.23557
R1837 VDD.n355 VDD.n191 7.94898
R1838 VDD.n205 VDD.n204 7.54844
R1839 VDD.n218 VDD.n217 7.54407
R1840 VDD.n354 VDD.n192 6.88686
R1841 VDD.n75 VDD.n72 6.8005
R1842 VDD.n366 VDD.n363 6.8005
R1843 VDD.n134 VDD.n126 6.48583
R1844 VDD.n425 VDD.n417 6.48583
R1845 VDD.n349 VDD.n348 6.02403
R1846 VDD.n300 VDD.n299 6.02403
R1847 VDD.n231 VDD.n222 6.02403
R1848 VDD.n243 VDD.n242 6.02403
R1849 VDD.n202 VDD.n193 6.02403
R1850 VDD.n215 VDD.n206 6.02403
R1851 VDD.n62 VDD.n61 6.02403
R1852 VDD.n11 VDD.n10 6.02403
R1853 VDD.n129 VDD.n128 5.8885
R1854 VDD.n420 VDD.n419 5.8885
R1855 VDD.n189 VDD 5.6325
R1856 VDD.n204 VDD.n203 5.18145
R1857 VDD.n217 VDD.n216 5.18145
R1858 VDD.n333 VDD.n324 4.89462
R1859 VDD.n317 VDD.n316 4.89462
R1860 VDD.n276 VDD.n267 4.89462
R1861 VDD.n260 VDD.n259 4.89462
R1862 VDD.n44 VDD.n35 4.89462
R1863 VDD.n28 VDD.n27 4.89462
R1864 VDD.n153 VDD.n119 4.67352
R1865 VDD.n444 VDD.n410 4.67352
R1866 VDD.n134 VDD.n133 4.62124
R1867 VDD.n425 VDD.n424 4.62124
R1868 VDD.n191 VDD.n190 4.5005
R1869 VDD.n131 VDD.n130 4.36875
R1870 VDD.n153 VDD.n152 4.36875
R1871 VDD.n113 VDD.n112 4.36875
R1872 VDD.n83 VDD.n82 4.36875
R1873 VDD.n422 VDD.n421 4.36875
R1874 VDD.n444 VDD.n443 4.36875
R1875 VDD.n404 VDD.n403 4.36875
R1876 VDD.n374 VDD.n373 4.36875
R1877 VDD.n186 VDD.n185 3.4105
R1878 VDD.t123 VDD.t49 3.35739
R1879 VDD.t115 VDD.t62 3.35739
R1880 VDD.t64 VDD.t58 3.35739
R1881 VDD.t40 VDD.t136 3.35739
R1882 VDD.n333 VDD.n322 3.25464
R1883 VDD.n290 VDD.n288 3.24308
R1884 VDD.n276 VDD.n265 3.23917
R1885 VDD.n44 VDD.n33 3.23917
R1886 VDD.n316 VDD.n305 3.23136
R1887 VDD.n259 VDD.n248 3.23136
R1888 VDD.n27 VDD.n16 3.23136
R1889 VDD.n283 VDD.n282 3.22655
R1890 VDD.n52 VDD.n50 3.22655
R1891 VDD.n131 VDD.n129 3.2005
R1892 VDD.n422 VDD.n420 3.2005
R1893 VDD.n341 VDD.n340 2.84665
R1894 VDD.n342 VDD.n339 2.84665
R1895 VDD.n332 VDD.n331 2.84665
R1896 VDD.n328 VDD.n323 2.84665
R1897 VDD.n315 VDD.n314 2.84665
R1898 VDD.n311 VDD.n306 2.84665
R1899 VDD.n292 VDD.n291 2.84665
R1900 VDD.n293 VDD.n289 2.84665
R1901 VDD.n225 VDD.n223 2.84665
R1902 VDD.n224 VDD.n221 2.84665
R1903 VDD.n275 VDD.n274 2.84665
R1904 VDD.n271 VDD.n266 2.84665
R1905 VDD.n258 VDD.n257 2.84665
R1906 VDD.n254 VDD.n249 2.84665
R1907 VDD.n235 VDD.n234 2.84665
R1908 VDD.n236 VDD.n233 2.84665
R1909 VDD.n196 VDD.n194 2.84665
R1910 VDD.n200 VDD.n196 2.84665
R1911 VDD.n197 VDD.n195 2.84665
R1912 VDD.n200 VDD.n195 2.84665
R1913 VDD.n209 VDD.n207 2.84665
R1914 VDD.n213 VDD.n209 2.84665
R1915 VDD.n210 VDD.n208 2.84665
R1916 VDD.n213 VDD.n208 2.84665
R1917 VDD.n54 VDD.n53 2.84665
R1918 VDD.n55 VDD.n51 2.84665
R1919 VDD.n43 VDD.n42 2.84665
R1920 VDD.n39 VDD.n34 2.84665
R1921 VDD.n26 VDD.n25 2.84665
R1922 VDD.n22 VDD.n17 2.84665
R1923 VDD.n3 VDD.n2 2.84665
R1924 VDD.n4 VDD.n1 2.84665
R1925 VDD.n129 VDD.n126 2.8165
R1926 VDD.n420 VDD.n417 2.8165
R1927 VDD.n106 VDD.n105 2.54018
R1928 VDD.n85 VDD.n84 2.54018
R1929 VDD.n397 VDD.n396 2.54018
R1930 VDD.n376 VDD.n375 2.54018
R1931 VDD.n119 VDD.n118 2.33701
R1932 VDD.n105 VDD.n104 2.33701
R1933 VDD.n85 VDD.n79 2.33701
R1934 VDD.n410 VDD.n409 2.33701
R1935 VDD.n396 VDD.n395 2.33701
R1936 VDD.n376 VDD.n370 2.33701
R1937 VDD.n351 VDD.n350 2.28169
R1938 VDD.n336 VDD.n335 2.28169
R1939 VDD.n319 VDD.n318 2.28169
R1940 VDD.n302 VDD.n301 2.28169
R1941 VDD.n285 VDD.n284 2.28169
R1942 VDD.n279 VDD.n278 2.28169
R1943 VDD.n262 VDD.n261 2.28169
R1944 VDD.n245 VDD.n244 2.28169
R1945 VDD.n64 VDD.n63 2.28169
R1946 VDD.n47 VDD.n46 2.28169
R1947 VDD.n30 VDD.n29 2.28169
R1948 VDD.n13 VDD.n12 2.28169
R1949 VDD.n305 VDD.n304 2.13544
R1950 VDD.n113 VDD.n106 2.13383
R1951 VDD.n84 VDD.n83 2.13383
R1952 VDD.n404 VDD.n397 2.13383
R1953 VDD.n375 VDD.n374 2.13383
R1954 VDD.n219 VDD.n205 2.06883
R1955 VDD.n118 VDD.n117 2.03225
R1956 VDD.n104 VDD.n103 2.03225
R1957 VDD.n79 VDD.n77 2.03225
R1958 VDD.n409 VDD.n408 2.03225
R1959 VDD.n395 VDD.n394 2.03225
R1960 VDD.n370 VDD.n368 2.03225
R1961 VDD.n304 VDD.n288 1.95379
R1962 VDD.n299 VDD.n290 1.88285
R1963 VDD.n242 VDD.n232 1.88285
R1964 VDD.n10 VDD.n0 1.88285
R1965 VDD.n184 VDD.n183 1.753
R1966 VDD.n475 VDD.n474 1.753
R1967 VDD.n92 VDD.n68 1.50638
R1968 VDD.n383 VDD.n359 1.50638
R1969 VDD.n176 VDD.n75 1.4005
R1970 VDD.n467 VDD.n366 1.4005
R1971 VDD.n355 VDD.n354 1.39787
R1972 VDD.n102 VDD.n100 1.37193
R1973 VDD.n89 VDD.n88 1.37193
R1974 VDD.n393 VDD.n391 1.37193
R1975 VDD.n380 VDD.n379 1.37193
R1976 VDD.n219 VDD.n218 1.33758
R1977 VDD.n338 VDD.n337 1.143
R1978 VDD.n321 VDD.n320 1.143
R1979 VDD.n281 VDD.n280 1.143
R1980 VDD.n264 VDD.n263 1.143
R1981 VDD.n49 VDD.n48 1.143
R1982 VDD.n32 VDD.n31 1.143
R1983 VDD.n353 VDD.n352 1.13925
R1984 VDD.n287 VDD.n286 1.13925
R1985 VDD.n66 VDD.n65 1.13925
R1986 VDD.n304 VDD.n303 1.13675
R1987 VDD.n247 VDD.n246 1.13675
R1988 VDD.n15 VDD.n14 1.13675
R1989 VDD.n348 VDD.n192 1.12991
R1990 VDD.n334 VDD.n333 1.12991
R1991 VDD.n316 VDD.n307 1.12991
R1992 VDD.n283 VDD.n231 1.12991
R1993 VDD.n277 VDD.n276 1.12991
R1994 VDD.n259 VDD.n250 1.12991
R1995 VDD.n61 VDD.n52 1.12991
R1996 VDD.n45 VDD.n44 1.12991
R1997 VDD.n27 VDD.n18 1.12991
R1998 VDD.n125 VDD 1.06099
R1999 VDD.n416 VDD 1.06099
R2000 VDD.n265 VDD.n264 0.862816
R2001 VDD.n33 VDD.n32 0.862816
R2002 VDD.n353 VDD.n338 0.854667
R2003 VDD.n478 VDD.n477 0.853
R2004 VDD.n356 VDD.n355 0.84345
R2005 VDD.n248 VDD.n247 0.770881
R2006 VDD.n16 VDD.n15 0.770881
R2007 VDD.n477 VDD.n475 0.763912
R2008 VDD.n162 VDD.n91 0.753441
R2009 VDD.n175 VDD.n174 0.753441
R2010 VDD.n453 VDD.n382 0.753441
R2011 VDD.n466 VDD.n465 0.753441
R2012 VDD.n282 VDD.n281 0.747859
R2013 VDD.n50 VDD.n49 0.729231
R2014 VDD.n220 VDD.n219 0.704667
R2015 VDD.n191 VDD.n186 0.624567
R2016 VDD.n357 VDD 0.614909
R2017 VDD.n72 VDD.n70 0.6005
R2018 VDD.n363 VDD.n361 0.6005
R2019 VDD.n322 VDD.n321 0.588641
R2020 VDD.n288 VDD.n287 0.518882
R2021 VDD.n185 VDD.n184 0.511794
R2022 VDD.n184 VDD 0.460219
R2023 VDD.n475 VDD 0.460219
R2024 VDD.n478 VDD.n357 0.455174
R2025 VDD.n66 VDD.n50 0.405788
R2026 VDD.n179 VDD.n70 0.4005
R2027 VDD.n470 VDD.n361 0.4005
R2028 VDD VDD.n356 0.396619
R2029 VDD.n264 VDD.n248 0.392323
R2030 VDD.n32 VDD.n16 0.392323
R2031 VDD.n281 VDD.n265 0.360318
R2032 VDD.n49 VDD.n33 0.360318
R2033 VDD.n152 VDD.n151 0.305262
R2034 VDD.n103 VDD.n102 0.305262
R2035 VDD.n112 VDD.n111 0.305262
R2036 VDD.n88 VDD.n77 0.305262
R2037 VDD.n443 VDD.n442 0.305262
R2038 VDD.n394 VDD.n393 0.305262
R2039 VDD.n403 VDD.n402 0.305262
R2040 VDD.n379 VDD.n368 0.305262
R2041 VDD.t32 VDD.n345 0.27666
R2042 VDD.n346 VDD.t32 0.27666
R2043 VDD.n330 VDD.t44 0.27666
R2044 VDD.n327 VDD.t44 0.27666
R2045 VDD.n313 VDD.t135 0.27666
R2046 VDD.n310 VDD.t135 0.27666
R2047 VDD.t34 VDD.n296 0.27666
R2048 VDD.n297 VDD.t34 0.27666
R2049 VDD.t142 VDD.n228 0.27666
R2050 VDD.n229 VDD.t142 0.27666
R2051 VDD.n273 VDD.t35 0.27666
R2052 VDD.n270 VDD.t35 0.27666
R2053 VDD.n256 VDD.t134 0.27666
R2054 VDD.n253 VDD.t134 0.27666
R2055 VDD.t33 VDD.n239 0.27666
R2056 VDD.n240 VDD.t33 0.27666
R2057 VDD.t83 VDD.n58 0.27666
R2058 VDD.n59 VDD.t83 0.27666
R2059 VDD.n41 VDD.t101 0.27666
R2060 VDD.n38 VDD.t101 0.27666
R2061 VDD.n24 VDD.t127 0.27666
R2062 VDD.n21 VDD.t127 0.27666
R2063 VDD.t84 VDD.n7 0.27666
R2064 VDD.n8 VDD.t84 0.27666
R2065 VDD.n338 VDD.n322 0.268128
R2066 VDD.n321 VDD.n305 0.223986
R2067 VDD.n354 VDD.n353 0.202423
R2068 VDD.n133 VDD.n132 0.180304
R2069 VDD.n424 VDD.n423 0.180304
R2070 VDD.n190 VDD 0.163379
R2071 VDD.n133 VDD 0.120408
R2072 VDD.n424 VDD 0.120408
R2073 VDD.n116 VDD.n95 0.120292
R2074 VDD.n154 VDD.n96 0.120292
R2075 VDD.n148 VDD.n147 0.120292
R2076 VDD.n147 VDD.n122 0.120292
R2077 VDD.n143 VDD.n142 0.120292
R2078 VDD.n142 VDD.n141 0.120292
R2079 VDD.n138 VDD.n137 0.120292
R2080 VDD.n137 VDD.n136 0.120292
R2081 VDD.n132 VDD.n127 0.120292
R2082 VDD.n101 VDD.n97 0.120292
R2083 VDD.n114 VDD.n98 0.120292
R2084 VDD.n165 VDD.n93 0.120292
R2085 VDD.n166 VDD.n165 0.120292
R2086 VDD.n182 VDD.n67 0.120292
R2087 VDD.n178 VDD.n177 0.120292
R2088 VDD.n177 VDD.n71 0.120292
R2089 VDD.n87 VDD.n86 0.120292
R2090 VDD.n86 VDD.n78 0.120292
R2091 VDD.n81 VDD.n78 0.120292
R2092 VDD.n407 VDD.n386 0.120292
R2093 VDD.n445 VDD.n387 0.120292
R2094 VDD.n439 VDD.n438 0.120292
R2095 VDD.n438 VDD.n413 0.120292
R2096 VDD.n434 VDD.n433 0.120292
R2097 VDD.n433 VDD.n432 0.120292
R2098 VDD.n429 VDD.n428 0.120292
R2099 VDD.n428 VDD.n427 0.120292
R2100 VDD.n423 VDD.n418 0.120292
R2101 VDD.n392 VDD.n388 0.120292
R2102 VDD.n405 VDD.n389 0.120292
R2103 VDD.n456 VDD.n384 0.120292
R2104 VDD.n457 VDD.n456 0.120292
R2105 VDD.n473 VDD.n358 0.120292
R2106 VDD.n469 VDD.n468 0.120292
R2107 VDD.n468 VDD.n362 0.120292
R2108 VDD.n378 VDD.n377 0.120292
R2109 VDD.n377 VDD.n369 0.120292
R2110 VDD.n372 VDD.n369 0.120292
R2111 VDD.n155 VDD.n95 0.11899
R2112 VDD.n446 VDD.n386 0.11899
R2113 VDD.n282 VDD.n220 0.1125
R2114 VDD.n476 VDD.n356 0.102957
R2115 VDD.n101 VDD 0.0981562
R2116 VDD.n392 VDD 0.0981562
R2117 VDD.n156 VDD 0.0955521
R2118 VDD.n447 VDD 0.0955521
R2119 VDD.n115 VDD.n97 0.0916458
R2120 VDD.n406 VDD.n388 0.0916458
R2121 VDD.n190 VDD 0.0800455
R2122 VDD.n352 VDD 0.06425
R2123 VDD.n337 VDD 0.06425
R2124 VDD.n320 VDD 0.06425
R2125 VDD.n303 VDD 0.06425
R2126 VDD.n286 VDD 0.06425
R2127 VDD.n280 VDD 0.06425
R2128 VDD.n263 VDD 0.06425
R2129 VDD.n246 VDD 0.06425
R2130 VDD.n218 VDD 0.06425
R2131 VDD.n65 VDD 0.06425
R2132 VDD.n48 VDD 0.06425
R2133 VDD.n31 VDD 0.06425
R2134 VDD.n14 VDD 0.06425
R2135 VDD.n149 VDD 0.0603958
R2136 VDD VDD.n148 0.0603958
R2137 VDD.n143 VDD 0.0603958
R2138 VDD.n138 VDD 0.0603958
R2139 VDD.n108 VDD 0.0603958
R2140 VDD VDD.n107 0.0603958
R2141 VDD VDD.n93 0.0603958
R2142 VDD.n168 VDD 0.0603958
R2143 VDD VDD.n167 0.0603958
R2144 VDD.n178 VDD 0.0603958
R2145 VDD.n87 VDD 0.0603958
R2146 VDD.n440 VDD 0.0603958
R2147 VDD VDD.n439 0.0603958
R2148 VDD.n434 VDD 0.0603958
R2149 VDD.n429 VDD 0.0603958
R2150 VDD.n399 VDD 0.0603958
R2151 VDD VDD.n398 0.0603958
R2152 VDD VDD.n384 0.0603958
R2153 VDD.n459 VDD 0.0603958
R2154 VDD VDD.n458 0.0603958
R2155 VDD.n469 VDD 0.0603958
R2156 VDD.n378 VDD 0.0603958
R2157 VDD.n205 VDD 0.059875
R2158 VDD.n90 VDD 0.0590938
R2159 VDD.n381 VDD 0.0590938
R2160 VDD.n476 VDD.n357 0.0582836
R2161 VDD.n287 VDD.n220 0.054
R2162 VDD.n183 VDD 0.0525833
R2163 VDD.n474 VDD 0.0525833
R2164 VDD.n183 VDD.n182 0.0460729
R2165 VDD.n474 VDD.n473 0.0460729
R2166 VDD.n108 VDD 0.0382604
R2167 VDD.n399 VDD 0.0382604
R2168 VDD VDD.n125 0.0369583
R2169 VDD VDD.n416 0.0369583
R2170 VDD.n149 VDD 0.03175
R2171 VDD.n168 VDD 0.03175
R2172 VDD.n440 VDD 0.03175
R2173 VDD.n459 VDD 0.03175
R2174 VDD.n115 VDD.n114 0.0291458
R2175 VDD.n406 VDD.n405 0.0291458
R2176 VDD.n185 VDD 0.0236148
R2177 VDD VDD.n96 0.0226354
R2178 VDD VDD.n122 0.0226354
R2179 VDD.n141 VDD 0.0226354
R2180 VDD.n136 VDD 0.0226354
R2181 VDD.n127 VDD 0.0226354
R2182 VDD VDD.n98 0.0226354
R2183 VDD.n107 VDD 0.0226354
R2184 VDD.n157 VDD 0.0226354
R2185 VDD VDD.n166 0.0226354
R2186 VDD.n167 VDD 0.0226354
R2187 VDD VDD.n67 0.0226354
R2188 VDD VDD.n71 0.0226354
R2189 VDD VDD.n76 0.0226354
R2190 VDD.n81 VDD 0.0226354
R2191 VDD VDD.n387 0.0226354
R2192 VDD VDD.n413 0.0226354
R2193 VDD.n432 VDD 0.0226354
R2194 VDD.n427 VDD 0.0226354
R2195 VDD.n418 VDD 0.0226354
R2196 VDD VDD.n389 0.0226354
R2197 VDD.n398 VDD 0.0226354
R2198 VDD.n448 VDD 0.0226354
R2199 VDD VDD.n457 0.0226354
R2200 VDD.n458 VDD 0.0226354
R2201 VDD VDD.n358 0.0226354
R2202 VDD VDD.n362 0.0226354
R2203 VDD VDD.n367 0.0226354
R2204 VDD.n372 VDD 0.0226354
R2205 VDD VDD.n478 0.0134382
R2206 VDD.n477 VDD.n476 0.00887356
R2207 VDD.n157 VDD.n156 0.00310417
R2208 VDD.n448 VDD.n447 0.00310417
R2209 VDD.n155 VDD.n154 0.00180208
R2210 VDD.n125 VDD 0.00180208
R2211 VDD.n90 VDD.n76 0.00180208
R2212 VDD.n446 VDD.n445 0.00180208
R2213 VDD.n416 VDD 0.00180208
R2214 VDD.n381 VDD.n367 0.00180208
R2215 R1R2.n2 R1R2.t4 26.3998
R2216 R1R2.n2 R1R2.t5 23.5483
R2217 R1R2.n1 R1R2.t2 12.7127
R2218 R1R2.n1 R1R2.t3 10.8578
R2219 R1R2.n0 R1R2.t1 10.8194
R2220 R1R2.n0 R1R2.t0 10.5739
R2221 R1R2.n3 R1R2.n2 3.12177
R2222 R1R2.n3 R1R2.n1 1.81453
R2223 R1R2.n4 R1R2.n3 1.1255
R2224 R1R2 R1R2.n0 0.539965
R2225 R1R2 R1R2.n4 0.132418
R2226 R1R2.n4 R1R2 0.0655
R2227 VRES.n5 VRES.t1 26.3998
R2228 VRES.n1 VRES.t6 26.3998
R2229 VRES.n5 VRES.t2 23.5483
R2230 VRES.n1 VRES.t4 23.5483
R2231 VRES.n4 VRES.t3 12.7127
R2232 VRES.n0 VRES.t7 12.7127
R2233 VRES.n4 VRES.t5 10.8578
R2234 VRES.n0 VRES.t8 10.8578
R2235 VRES.n8 VRES.t0 10.5285
R2236 VRES.n9 VRES 6.58743
R2237 VRES.n6 VRES.n5 3.12177
R2238 VRES.n2 VRES.n1 3.12177
R2239 VRES.n6 VRES.n4 1.81453
R2240 VRES.n2 VRES.n0 1.81453
R2241 VRES.n8 VRES 1.39577
R2242 VRES.n7 VRES.n6 1.1255
R2243 VRES.n3 VRES.n2 1.1255
R2244 VRES VRES.n8 0.472894
R2245 VRES.n9 VRES.n3 0.160652
R2246 VRES VRES.n7 0.134513
R2247 VRES.n7 VRES 0.0655
R2248 VRES.n3 VRES 0.0655
R2249 VRES VRES.n9 0.05925
R2250 x1.x3.GN1.n2 x1.x3.GN1.t6 377.486
R2251 x1.x3.GN1.n3 x1.x3.GN1.t2 377.486
R2252 x1.x3.GN1.n2 x1.x3.GN1.t5 374.202
R2253 x1.x3.GN1.n3 x1.x3.GN1.t9 374.202
R2254 x1.x3.GN1.n10 x1.x3.GN1.t1 339.418
R2255 x1.x3.GN1.n1 x1.x3.GN1.t0 274.06
R2256 x1.x3.GN1.n7 x1.x3.GN1.t7 212.081
R2257 x1.x3.GN1.n6 x1.x3.GN1.t8 212.081
R2258 x1.x3.GN1.n8 x1.x3.GN1.n7 182.673
R2259 x1.x3.GN1.n7 x1.x3.GN1.t3 139.78
R2260 x1.x3.GN1.n6 x1.x3.GN1.t4 139.78
R2261 x1.x3.GN1.n7 x1.x3.GN1.n6 61.346
R2262 x1.x3.GN1.n5 x1.x3.GN1.n8 15.8606
R2263 x1.x3.GN1 x1.x3.GN1.n9 13.8044
R2264 x1.x3.GN1.n0 x1.x3.GN1.n4 13.4101
R2265 x1.x3.GN1.n0 x1.x3.GN1 11.5859
R2266 x1.x3.GN1.n4 x1.x3.GN1 11.5859
R2267 x1.x3.GN1 x1.x3.GN1.n1 11.0989
R2268 x1.x3.GN1.n9 x1.x3.GN1.n5 6.94768
R2269 x1.x3.GN1 x1.x3.GN1.n0 6.73859
R2270 x1.x3.GN1.n11 x1.x3.GN1 6.6565
R2271 x1.x3.GN1.n8 x1.x3.GN1 6.4005
R2272 x1.x3.GN1.n1 x1.x3.GN1 6.1445
R2273 x1.x3.GN1.n0 x1.x3.GN1 5.13959
R2274 x1.x3.GN1.n4 x1.x3.GN1 4.55738
R2275 x1.x3.GN1.n11 x1.x3.GN1.n10 4.0914
R2276 x1.x3.GN1 x1.x3.GN1.n11 3.61789
R2277 x1.x3.GN1.n9 x1.x3.GN1 3.26325
R2278 x1.x3.GN1.n1 x1.x3.GN1 2.86947
R2279 x1.x3.GN1 x1.x3.GN1.n2 2.04102
R2280 x1.x3.GN1 x1.x3.GN1.n3 2.04102
R2281 x1.x3.GN1.n10 x1.x3.GN1 1.74382
R2282 x1.x3.GN1.n5 x1.x3.GN1 1.47326
R2283 R3R4.n2 R3R4.t3 26.3998
R2284 R3R4.n8 R3R4.t9 26.3998
R2285 R3R4.n2 R3R4.t2 23.5483
R2286 R3R4.n8 R3R4.t6 23.5483
R2287 R3R4.n1 R3R4.t7 12.7127
R2288 R3R4.n7 R3R4.t1 12.7127
R2289 R3R4.n1 R3R4.t8 10.8578
R2290 R3R4.n7 R3R4.t0 10.8578
R2291 R3R4.n0 R3R4.t5 10.8241
R2292 R3R4.n0 R3R4.t4 10.5739
R2293 R3R4.n6 R3R4.n5 7.08509
R2294 R3R4.n3 R3R4.n2 3.12177
R2295 R3R4.n9 R3R4.n8 3.12177
R2296 R3R4.n3 R3R4.n1 1.81453
R2297 R3R4.n9 R3R4.n7 1.81453
R2298 R3R4.n4 R3R4.n3 1.1255
R2299 R3R4.n10 R3R4.n9 1.1255
R2300 R3R4.n5 R3R4 0.893357
R2301 R3R4 R3R4.n6 0.43675
R2302 R3R4.n5 R3R4.n4 0.355632
R2303 R3R4.n6 R3R4.n0 0.183423
R2304 R3R4 R3R4.n10 0.148615
R2305 R3R4.n4 R3R4 0.0655
R2306 R3R4.n10 R3R4 0.0655
R2307 R3R4.n5 R3R4 0.00907843
R2308 SELECT0.n5 SELECT0.t7 327.99
R2309 SELECT0.n9 SELECT0.t1 293.969
R2310 SELECT0.n3 SELECT0.t0 261.887
R2311 SELECT0.n1 SELECT0.t8 212.081
R2312 SELECT0.n0 SELECT0.t9 212.081
R2313 SELECT0.n5 SELECT0.t6 199.457
R2314 SELECT0.n2 SELECT0.n1 183.185
R2315 SELECT0.n3 SELECT0.t4 155.847
R2316 SELECT0 SELECT0.n9 154.065
R2317 SELECT0.n6 SELECT0.n5 152
R2318 SELECT0.n4 SELECT0.n3 152
R2319 SELECT0.n1 SELECT0.t2 139.78
R2320 SELECT0.n0 SELECT0.t3 139.78
R2321 SELECT0.n9 SELECT0.t5 138.338
R2322 SELECT0.n1 SELECT0.n0 61.346
R2323 SELECT0.n10 SELECT0 13.4199
R2324 SELECT0.n8 SELECT0.n4 11.9062
R2325 SELECT0.n11 SELECT0.n8 11.7395
R2326 SELECT0.n12 SELECT0.n11 11.5949
R2327 SELECT0.n12 SELECT0.n2 9.68118
R2328 SELECT0.n7 SELECT0 9.17383
R2329 SELECT0.n2 SELECT0 5.8885
R2330 SELECT0.n10 SELECT0 5.57469
R2331 SELECT0.n8 SELECT0.n7 4.6505
R2332 SELECT0.n11 SELECT0.n10 4.6505
R2333 SELECT0.n7 SELECT0.n6 2.98717
R2334 SELECT0.n6 SELECT0 2.34717
R2335 SELECT0.n4 SELECT0 2.07109
R2336 SELECT0 SELECT0.n12 0.559212
R2337 RSEL2.n3 RSEL2.t4 450.938
R2338 RSEL2.n3 RSEL2.t0 445.666
R2339 RSEL2.n0 RSEL2.t1 377.486
R2340 RSEL2.n0 RSEL2.t5 374.202
R2341 RSEL2.n7 RSEL2.t2 212.081
R2342 RSEL2.n6 RSEL2.t3 212.081
R2343 RSEL2.n8 RSEL2.n7 183.441
R2344 RSEL2.n7 RSEL2.t6 139.78
R2345 RSEL2.n6 RSEL2.t7 139.78
R2346 RSEL2.n7 RSEL2.n6 61.346
R2347 RSEL2.n5 RSEL2.n2 12.4093
R2348 RSEL2 RSEL2.n8 11.4331
R2349 RSEL2.n5 RSEL2.n4 9.10647
R2350 RSEL2.n9 RSEL2.n5 8.98648
R2351 RSEL2.n8 RSEL2 5.6325
R2352 RSEL2.n9 RSEL2 5.02323
R2353 RSEL2.n10 RSEL2 4.97651
R2354 RSEL2.n4 RSEL2.n3 3.1748
R2355 RSEL2.n2 RSEL2.n0 2.10165
R2356 RSEL2.n1 RSEL2 1.09425
R2357 RSEL2.n10 RSEL2.n9 0.890652
R2358 RSEL2.n4 RSEL2 0.063625
R2359 RSEL2.n2 RSEL2.n1 0.062375
R2360 RSEL2 RSEL2.n10 0.0516364
R2361 RSEL2.n1 RSEL2 0.003
R2362 LADDEROUT.n1 LADDEROUT.t1 26.3998
R2363 LADDEROUT.n5 LADDEROUT.t9 23.6581
R2364 LADDEROUT.n12 LADDEROUT.t4 23.6581
R2365 LADDEROUT.n1 LADDEROUT.t6 23.5483
R2366 LADDEROUT.n4 LADDEROUT.t8 23.3739
R2367 LADDEROUT.n11 LADDEROUT.t5 23.3739
R2368 LADDEROUT.n0 LADDEROUT.t7 12.7127
R2369 LADDEROUT.n0 LADDEROUT.t0 10.8578
R2370 LADDEROUT.n5 LADDEROUT.t3 10.7528
R2371 LADDEROUT.n12 LADDEROUT.t10 10.7528
R2372 LADDEROUT.n7 LADDEROUT.t2 10.6417
R2373 LADDEROUT.n14 LADDEROUT.t11 10.6417
R2374 LADDEROUT.n10 LADDEROUT 4.4752
R2375 LADDEROUT.n2 LADDEROUT.n1 3.12177
R2376 LADDEROUT.n2 LADDEROUT.n0 1.81453
R2377 LADDEROUT.n6 LADDEROUT.n5 1.30064
R2378 LADDEROUT.n13 LADDEROUT.n12 1.30064
R2379 LADDEROUT.n3 LADDEROUT.n2 1.1255
R2380 LADDEROUT.n16 LADDEROUT.n15 1.04212
R2381 LADDEROUT.n9 LADDEROUT.n8 0.859481
R2382 LADDEROUT.n6 LADDEROUT.n4 0.726502
R2383 LADDEROUT.n13 LADDEROUT.n11 0.726502
R2384 LADDEROUT.n18 LADDEROUT.n17 0.659371
R2385 LADDEROUT.n10 LADDEROUT.n9 0.584875
R2386 LADDEROUT.n17 LADDEROUT.n16 0.547124
R2387 LADDEROUT.n7 LADDEROUT.n6 0.512491
R2388 LADDEROUT.n14 LADDEROUT.n13 0.512491
R2389 LADDEROUT.n8 LADDEROUT.n7 0.359663
R2390 LADDEROUT.n15 LADDEROUT.n14 0.359663
R2391 LADDEROUT LADDEROUT.n10 0.3355
R2392 LADDEROUT.n18 LADDEROUT 0.329447
R2393 LADDEROUT LADDEROUT.n3 0.294448
R2394 LADDEROUT.n8 LADDEROUT.n4 0.216071
R2395 LADDEROUT.n15 LADDEROUT.n11 0.216071
R2396 LADDEROUT.n17 LADDEROUT 0.208
R2397 LADDEROUT.n3 LADDEROUT 0.0655
R2398 LADDEROUT LADDEROUT.n18 0.0241318
R2399 LADDEROUT.n16 LADDEROUT 0.0100278
R2400 LADDEROUT.n9 LADDEROUT 0.001125
R2401 RSEL1.n10 RSEL1.t9 327.99
R2402 RSEL1.n3 RSEL1.t6 293.969
R2403 RSEL1.n6 RSEL1.t8 256.07
R2404 RSEL1.n1 RSEL1.t2 212.081
R2405 RSEL1.n0 RSEL1.t4 212.081
R2406 RSEL1.n10 RSEL1.t3 199.457
R2407 RSEL1.n2 RSEL1.n1 182.929
R2408 RSEL1 RSEL1.n3 154.065
R2409 RSEL1.n11 RSEL1.n10 152
R2410 RSEL1.n7 RSEL1.n6 152
R2411 RSEL1.n6 RSEL1.t0 150.03
R2412 RSEL1.n1 RSEL1.t5 139.78
R2413 RSEL1.n0 RSEL1.t1 139.78
R2414 RSEL1.n3 RSEL1.t7 138.338
R2415 RSEL1.n1 RSEL1.n0 61.346
R2416 RSEL1.n5 RSEL1 22.1096
R2417 RSEL1.n14 RSEL1.n13 14.6836
R2418 RSEL1.n13 RSEL1.n12 14.6704
R2419 RSEL1.n12 RSEL1 13.8672
R2420 RSEL1.n4 RSEL1 13.8328
R2421 RSEL1.n11 RSEL1 12.1605
R2422 RSEL1.n14 RSEL1.n2 10.6811
R2423 RSEL1.n7 RSEL1.n5 10.4374
R2424 RSEL1.n9 RSEL1.n8 8.15359
R2425 RSEL1.n2 RSEL1 6.1445
R2426 RSEL1.n4 RSEL1 5.16179
R2427 RSEL1.n15 RSEL1 4.66338
R2428 RSEL1.n9 RSEL1.n4 4.65206
R2429 RSEL1.n8 RSEL1 3.93896
R2430 RSEL1.n16 RSEL1 2.5005
R2431 RSEL1 RSEL1.n11 2.34717
R2432 RSEL1.n5 RSEL1 2.16665
R2433 RSEL1.n8 RSEL1.n7 1.57588
R2434 RSEL1.n13 RSEL1.n9 0.79438
R2435 RSEL1.n12 RSEL1 0.6405
R2436 RSEL1.n15 RSEL1 0.606561
R2437 RSEL1.n16 RSEL1.n15 0.342759
R2438 RSEL1 RSEL1.n14 0.248606
R2439 RSEL1 RSEL1.n16 0.00359406
R2440 x1.x3.GN4.n3 x1.x3.GN4.t2 377.486
R2441 x1.x3.GN4.n1 x1.x3.GN4.t7 377.486
R2442 x1.x3.GN4.n3 x1.x3.GN4.t3 374.202
R2443 x1.x3.GN4.n1 x1.x3.GN4.t5 374.202
R2444 x1.x3.GN4.n9 x1.x3.GN4.t1 339.418
R2445 x1.x3.GN4.n0 x1.x3.GN4.t0 274.06
R2446 x1.x3.GN4.n6 x1.x3.GN4.t4 212.081
R2447 x1.x3.GN4.n5 x1.x3.GN4.t6 212.081
R2448 x1.x3.GN4.n7 x1.x3.GN4.n6 184.977
R2449 x1.x3.GN4.n6 x1.x3.GN4.t8 139.78
R2450 x1.x3.GN4.n5 x1.x3.GN4.t9 139.78
R2451 x1.x3.GN4.n6 x1.x3.GN4.n5 61.346
R2452 x1.x3.GN4.n8 x1.x3.GN4 18.2601
R2453 x1.x3.GN4 x1.x3.GN4.n7 13.8193
R2454 x1.x3.GN4 x1.x3.GN4.n4 11.7568
R2455 x1.x3.GN4.n4 x1.x3.GN4.n2 11.6628
R2456 x1.x3.GN4 x1.x3.GN4.n0 11.2645
R2457 x1.x3.GN4 x1.x3.GN4.n8 8.9605
R2458 x1.x3.GN4.n8 x1.x3.GN4 8.4485
R2459 x1.x3.GN4.n2 x1.x3.GN4 8.16743
R2460 x1.x3.GN4.n10 x1.x3.GN4 6.6565
R2461 x1.x3.GN4.n0 x1.x3.GN4 6.1445
R2462 x1.x3.GN4.n4 x1.x3.GN4 5.8185
R2463 x1.x3.GN4.n2 x1.x3.GN4 4.58237
R2464 x1.x3.GN4.n7 x1.x3.GN4 4.0965
R2465 x1.x3.GN4.n10 x1.x3.GN4.n9 4.0914
R2466 x1.x3.GN4 x1.x3.GN4.n10 3.61789
R2467 x1.x3.GN4.n0 x1.x3.GN4 2.86947
R2468 x1.x3.GN4 x1.x3.GN4.n3 2.04102
R2469 x1.x3.GN4 x1.x3.GN4.n1 2.04102
R2470 x1.x3.GN4.n9 x1.x3.GN4 1.74382
R2471 x2.x2.GP4.n2 x2.x2.GP4.t5 450.938
R2472 x2.x2.GP4.n2 x2.x2.GP4.t4 445.666
R2473 x2.x1.x14.Y x2.x2.GP4.n4 203.923
R2474 x2.x2.GP4.n0 x2.x2.GP4.n1 101.49
R2475 x2.x2.GP4.n4 x2.x2.GP4.t1 26.5955
R2476 x2.x2.GP4.n4 x2.x2.GP4.t3 26.5955
R2477 x2.x2.GP4.n1 x2.x2.GP4.t2 24.9236
R2478 x2.x2.GP4.n1 x2.x2.GP4.t0 24.9236
R2479 x2.x1.gpo3 x2.x2.x4.GP 16.5752
R2480 x2.x2.GP4.n3 x2.x1.x14.Y 10.7525
R2481 x2.x2.GP4.n0 x2.x1.gpo3 7.7042
R2482 x2.x2.GP4.n3 x2.x1.x14.Y 6.6565
R2483 x2.x1.x14.Y x2.x2.GP4.n3 5.04292
R2484 x2.x2.x4.GP x2.x2.GP4.n2 2.95993
R2485 x2.x1.x14.Y x2.x2.GP4.n0 2.5605
R2486 x2.x2.GP4.n0 x2.x1.x14.Y 1.93989
R2487 OUT.n19 OUT.t13 23.6581
R2488 OUT.n13 OUT.t11 23.6581
R2489 OUT.n7 OUT.t3 23.6581
R2490 OUT.n1 OUT.t5 23.6581
R2491 OUT.n21 OUT.t12 23.3739
R2492 OUT.n15 OUT.t10 23.3739
R2493 OUT.n9 OUT.t6 23.3739
R2494 OUT.n3 OUT.t2 23.3739
R2495 OUT.n19 OUT.t4 10.7528
R2496 OUT.n13 OUT.t15 10.7528
R2497 OUT.n7 OUT.t9 10.7528
R2498 OUT.n1 OUT.t1 10.7528
R2499 OUT.n18 OUT.t0 10.6417
R2500 OUT.n12 OUT.t14 10.6417
R2501 OUT.n6 OUT.t8 10.6417
R2502 OUT.n0 OUT.t7 10.6417
R2503 OUT.n20 OUT.n19 1.30064
R2504 OUT.n14 OUT.n13 1.30064
R2505 OUT.n8 OUT.n7 1.30064
R2506 OUT.n2 OUT.n1 1.30064
R2507 OUT OUT.n22 0.983856
R2508 OUT.n5 OUT.n4 0.956356
R2509 OUT.n11 OUT.n10 0.936641
R2510 OUT.n17 OUT.n16 0.924585
R2511 OUT.n23 OUT 0.76175
R2512 OUT.n21 OUT.n20 0.726502
R2513 OUT.n15 OUT.n14 0.726502
R2514 OUT.n9 OUT.n8 0.726502
R2515 OUT.n3 OUT.n2 0.726502
R2516 OUT.n25 OUT.n24 0.67425
R2517 OUT.n24 OUT.n23 0.66925
R2518 OUT.n27 OUT.n26 0.550998
R2519 OUT.n20 OUT.n18 0.512491
R2520 OUT.n14 OUT.n12 0.512491
R2521 OUT.n8 OUT.n6 0.512491
R2522 OUT.n2 OUT.n0 0.512491
R2523 OUT.n22 OUT.n18 0.359663
R2524 OUT.n16 OUT.n12 0.359663
R2525 OUT.n10 OUT.n6 0.359663
R2526 OUT.n4 OUT.n0 0.359663
R2527 OUT.n27 OUT 0.28175
R2528 OUT.n22 OUT.n21 0.216071
R2529 OUT.n16 OUT.n15 0.216071
R2530 OUT.n10 OUT.n9 0.216071
R2531 OUT.n4 OUT.n3 0.216071
R2532 OUT.n24 OUT 0.12425
R2533 OUT.n25 OUT 0.12175
R2534 OUT.n23 OUT 0.10175
R2535 OUT.n11 OUT 0.0776605
R2536 OUT.n17 OUT 0.0656042
R2537 OUT OUT.n11 0.0561931
R2538 OUT.n26 OUT 0.0529998
R2539 OUT OUT.n17 0.0376287
R2540 OUT OUT.n27 0.0282778
R2541 OUT.n5 OUT 0.028
R2542 OUT OUT.n5 0.0266905
R2543 OUT.n26 OUT.n25 0.01303
R2544 x2.x2.GN1.n1 x2.x2.GN1.t6 377.486
R2545 x2.x2.GN1.n1 x2.x2.GN1.t7 374.202
R2546 x2.x2.GN1.n7 x2.x2.GN1.t1 339.418
R2547 x2.x2.GN1.n0 x2.x2.GN1.t0 274.06
R2548 x2.x2.GN1.n4 x2.x2.GN1.t3 212.081
R2549 x2.x2.GN1.n3 x2.x2.GN1.t5 212.081
R2550 x2.x2.GN1.n5 x2.x2.GN1.n4 182.673
R2551 x2.x2.GN1.n4 x2.x2.GN1.t4 139.78
R2552 x2.x2.GN1.n3 x2.x2.GN1.t2 139.78
R2553 x2.x2.GN1.n4 x2.x2.GN1.n3 61.346
R2554 x2.x2.GN1 x2.x2.GN1.n5 15.8606
R2555 x2.x2.GN1 x2.x2.GN1.n6 13.8044
R2556 x2.x2.GN1.n2 x2.x2.GN1 11.5859
R2557 x2.x2.GN1 x2.x2.GN1.n0 11.0989
R2558 x2.x2.GN1 x2.x2.GN1.n2 10.8756
R2559 x2.x2.GN1.n6 x2.x2.GN1 8.1246
R2560 x2.x2.GN1.n8 x2.x2.GN1 6.6565
R2561 x2.x2.GN1.n5 x2.x2.GN1 6.4005
R2562 x2.x2.GN1.n0 x2.x2.GN1 6.1445
R2563 x2.x2.GN1.n2 x2.x2.GN1 4.55738
R2564 x2.x2.GN1.n8 x2.x2.GN1.n7 4.0914
R2565 x2.x2.GN1 x2.x2.GN1.n8 3.61789
R2566 x2.x2.GN1.n6 x2.x2.GN1 3.26325
R2567 x2.x2.GN1.n0 x2.x2.GN1 2.86947
R2568 x2.x2.GN1 x2.x2.GN1.n1 2.04102
R2569 x2.x2.GN1.n7 x2.x2.GN1 1.74382
R2570 x2.x2.GP1.n4 x2.x2.GP1.t4 450.938
R2571 x2.x2.GP1.n4 x2.x2.GP1.t5 445.666
R2572 x2.x2.GP1.n5 x2.x2.GP1.n3 195.832
R2573 x2.x2.GP1.n1 x2.x2.GP1.n0 101.49
R2574 x2.x2.GP1.n3 x2.x2.GP1.t2 26.5955
R2575 x2.x2.GP1.n3 x2.x2.GP1.t3 26.5955
R2576 x2.x2.GP1.n0 x2.x2.GP1.t1 24.9236
R2577 x2.x2.GP1.n0 x2.x2.GP1.t0 24.9236
R2578 x2.x2.GP1.n5 x2.x1.gpo0 11.8923
R2579 x2.x1.gpo0 x2.x2.x1.GP 11.5413
R2580 x2.x2.GP1.n2 x2.x1.x11.Y 10.7525
R2581 x2.x1.x11.Y x2.x2.GP1.n5 8.09215
R2582 x2.x2.GP1.n2 x2.x1.x11.Y 6.6565
R2583 x2.x1.x11.Y x2.x2.GP1.n2 5.04292
R2584 x2.x2.x1.GP x2.x2.GP1.n4 2.90754
R2585 x2.x1.x11.Y x2.x2.GP1.n1 2.5605
R2586 x2.x2.GP1.n1 x2.x1.x11.Y 1.93989
R2587 x2.x2.GN4.n1 x2.x2.GN4.t6 377.486
R2588 x2.x2.GN4.n1 x2.x2.GN4.t5 374.202
R2589 x2.x2.GN4.n7 x2.x2.GN4.t1 339.418
R2590 x2.x2.GN4.n0 x2.x2.GN4.t0 274.06
R2591 x2.x2.GN4.n4 x2.x2.GN4.t7 212.081
R2592 x2.x2.GN4.n3 x2.x2.GN4.t2 212.081
R2593 x2.x2.GN4.n5 x2.x2.GN4.n4 184.977
R2594 x2.x2.GN4.n4 x2.x2.GN4.t3 139.78
R2595 x2.x2.GN4.n3 x2.x2.GN4.t4 139.78
R2596 x2.x2.GN4.n4 x2.x2.GN4.n3 61.346
R2597 x2.x2.GN4.n6 x2.x2.GN4 18.2601
R2598 x2.x2.GN4 x2.x2.GN4.n2 17.2682
R2599 x2.x2.GN4 x2.x2.GN4.n5 15.0136
R2600 x2.x2.GN4 x2.x2.GN4.n0 11.2645
R2601 x2.x2.GN4 x2.x2.GN4.n6 8.9605
R2602 x2.x2.GN4.n6 x2.x2.GN4 8.4485
R2603 x2.x2.GN4.n2 x2.x2.GN4 8.16743
R2604 x2.x2.GN4.n8 x2.x2.GN4 6.6565
R2605 x2.x2.GN4.n0 x2.x2.GN4 6.1445
R2606 x2.x2.GN4.n2 x2.x2.GN4 4.58237
R2607 x2.x2.GN4.n5 x2.x2.GN4 4.0965
R2608 x2.x2.GN4.n8 x2.x2.GN4.n7 4.0914
R2609 x2.x2.GN4 x2.x2.GN4.n8 3.61789
R2610 x2.x2.GN4.n0 x2.x2.GN4 2.86947
R2611 x2.x2.GN4 x2.x2.GN4.n1 2.04102
R2612 x2.x2.GN4.n7 x2.x2.GN4 1.74382
R2613 RSEL0.n5 RSEL0.t5 327.99
R2614 RSEL0.n9 RSEL0.t3 293.969
R2615 RSEL0.n3 RSEL0.t6 261.887
R2616 RSEL0.n1 RSEL0.t9 212.081
R2617 RSEL0.n0 RSEL0.t8 212.081
R2618 RSEL0.n5 RSEL0.t1 199.457
R2619 RSEL0.n2 RSEL0.n1 183.185
R2620 RSEL0.n3 RSEL0.t7 155.847
R2621 RSEL0 RSEL0.n9 154.065
R2622 RSEL0.n6 RSEL0.n5 152
R2623 RSEL0.n4 RSEL0.n3 152
R2624 RSEL0.n1 RSEL0.t4 139.78
R2625 RSEL0.n0 RSEL0.t0 139.78
R2626 RSEL0.n9 RSEL0.t2 138.338
R2627 RSEL0.n1 RSEL0.n0 61.346
R2628 RSEL0.n10 RSEL0 13.4199
R2629 RSEL0.n8 RSEL0.n4 11.9062
R2630 RSEL0.n11 RSEL0.n8 11.7395
R2631 RSEL0.n12 RSEL0.n11 11.5949
R2632 RSEL0.n12 RSEL0.n2 9.68118
R2633 RSEL0.n7 RSEL0 9.17383
R2634 RSEL0.n2 RSEL0 5.8885
R2635 RSEL0.n10 RSEL0 5.57469
R2636 RSEL0.n8 RSEL0.n7 4.6505
R2637 RSEL0.n11 RSEL0.n10 4.6505
R2638 RSEL0.n7 RSEL0.n6 2.98717
R2639 RSEL0.n6 RSEL0 2.34717
R2640 RSEL0.n4 RSEL0 2.07109
R2641 RSEL0 RSEL0.n12 0.559212
R2642 x1.x3.GP1.n4 x1.x3.GP1.t7 450.938
R2643 x1.x3.GP1.n3 x1.x3.GP1.t5 450.938
R2644 x1.x3.GP1.n4 x1.x3.GP1.t4 445.666
R2645 x1.x3.GP1.n3 x1.x3.GP1.t6 445.666
R2646 x1.x3.GP1.n7 x1.x3.GP1.n6 195.832
R2647 x1.x3.GP1.n1 x1.x3.GP1.n0 101.49
R2648 x1.x3.GP1.n6 x1.x3.GP1.t2 26.5955
R2649 x1.x3.GP1.n6 x1.x3.GP1.t3 26.5955
R2650 x1.x3.GP1.n0 x1.x3.GP1.t0 24.9236
R2651 x1.x3.GP1.n0 x1.x3.GP1.t1 24.9236
R2652 x1.x3.GP1.n5 x1.x3.x1.GP 13.3282
R2653 x1.x3.GP1.n7 x1.x1.gpo0 11.8923
R2654 x1.x3.GP1.n2 x1.x1.x11.Y 10.7525
R2655 x1.x1.x11.Y x1.x3.GP1.n7 8.09215
R2656 x1.x3.GP1.n2 x1.x1.x11.Y 6.6565
R2657 x1.x1.gpo0 x1.x3.GP1.n5 5.46644
R2658 x1.x3.GP1.n5 x1.x2.GP1 5.31412
R2659 x1.x1.x11.Y x1.x3.GP1.n2 5.04292
R2660 x1.x2.GP1 x1.x3.GP1.n4 3.18415
R2661 x1.x3.x1.GP x1.x3.GP1.n3 2.90754
R2662 x1.x1.x11.Y x1.x3.GP1.n1 2.5605
R2663 x1.x3.GP1.n1 x1.x1.x11.Y 1.93989
R2664 x1.x3.GP2.n4 x1.x3.GP2.t6 450.938
R2665 x1.x3.GP2.n3 x1.x3.GP2.t4 450.938
R2666 x1.x3.GP2.n4 x1.x3.GP2.t7 445.666
R2667 x1.x3.GP2.n3 x1.x3.GP2.t5 445.666
R2668 x1.x3.GP2.n7 x1.x3.GP2.n6 195.958
R2669 x1.x3.GP2.n1 x1.x3.GP2.n0 101.49
R2670 x1.x3.GP2.n6 x1.x3.GP2.t2 26.5955
R2671 x1.x3.GP2.n6 x1.x3.GP2.t3 26.5955
R2672 x1.x3.GP2.n0 x1.x3.GP2.t1 24.9236
R2673 x1.x3.GP2.n0 x1.x3.GP2.t0 24.9236
R2674 x1.x3.GP2.n5 x1.x3.x2.GP 14.964
R2675 x1.x3.GP2.n7 x1.x1.gpo1 11.8408
R2676 x1.x3.GP2.n2 x1.x1.x12.Y 10.7525
R2677 x1.x1.gpo1 x1.x3.GP2.n5 8.86265
R2678 x1.x1.x12.Y x1.x3.GP2.n7 7.96524
R2679 x1.x3.GP2.n2 x1.x1.x12.Y 6.6565
R2680 x1.x3.GP2.n5 x1.x2.x2.GP 5.75481
R2681 x1.x1.x12.Y x1.x3.GP2.n2 5.04292
R2682 x1.x2.x2.GP x1.x3.GP2.n4 2.94361
R2683 x1.x3.x2.GP x1.x3.GP2.n3 2.94361
R2684 x1.x1.x12.Y x1.x3.GP2.n1 2.5605
R2685 x1.x3.GP2.n1 x1.x1.x12.Y 1.93989
R2686 x2.x2.GP2.n4 x2.x2.GP2.t4 450.938
R2687 x2.x2.GP2.n4 x2.x2.GP2.t5 445.666
R2688 x2.x2.GP2.n5 x2.x2.GP2.n3 195.958
R2689 x2.x2.GP2.n1 x2.x2.GP2.n0 101.49
R2690 x2.x2.GP2.n3 x2.x2.GP2.t2 26.5955
R2691 x2.x2.GP2.n3 x2.x2.GP2.t3 26.5955
R2692 x2.x2.GP2.n0 x2.x2.GP2.t0 24.9236
R2693 x2.x2.GP2.n0 x2.x2.GP2.t1 24.9236
R2694 x2.x1.gpo1 x2.x2.x2.GP 13.129
R2695 x2.x2.GP2.n5 x2.x1.gpo1 11.995
R2696 x2.x2.GP2.n2 x2.x1.x12.Y 10.7525
R2697 x2.x1.x12.Y x2.x2.GP2.n5 7.96524
R2698 x2.x2.GP2.n2 x2.x1.x12.Y 6.6565
R2699 x2.x1.x12.Y x2.x2.GP2.n2 5.04292
R2700 x2.x2.x2.GP x2.x2.GP2.n4 2.94361
R2701 x2.x1.x12.Y x2.x2.GP2.n1 2.5605
R2702 x2.x2.GP2.n1 x2.x1.x12.Y 1.93989
R2703 R5R6.n1 R5R6.t4 26.3998
R2704 R5R6.n1 R5R6.t3 23.5483
R2705 R5R6.n0 R5R6.t1 12.7127
R2706 R5R6.n4 R5R6.t2 10.885
R2707 R5R6.n0 R5R6.t0 10.8578
R2708 R5R6.n4 R5R6.t5 10.5949
R2709 R5R6.n2 R5R6.n1 3.12177
R2710 R5R6.n2 R5R6.n0 1.81453
R2711 R5R6.n3 R5R6.n2 1.1255
R2712 R5R6.n5 R5R6.n4 0.78425
R2713 R5R6.n5 R5R6 0.758625
R2714 R5R6 R5R6.n3 0.132418
R2715 R5R6.n3 R5R6 0.0655
R2716 R5R6 R5R6.n5 0.024875
R2717 R2R3.n1 R2R3.t4 26.3998
R2718 R2R3.n1 R2R3.t3 23.5483
R2719 R2R3.n0 R2R3.t2 12.7127
R2720 R2R3.n4 R2R3.t0 10.861
R2721 R2R3.n0 R2R3.t1 10.8578
R2722 R2R3.n4 R2R3.t5 10.5285
R2723 R2R3.n2 R2R3.n1 3.12177
R2724 R2R3.n2 R2R3.n0 1.81453
R2725 R2R3.n3 R2R3.n2 1.1255
R2726 R2R3.n5 R2R3.n4 0.69002
R2727 R2R3 R2R3.n3 0.138152
R2728 R2R3.n3 R2R3 0.0655
R2729 R2R3 R2R3.n5 0.053625
R2730 R2R3.n5 R2R3 0.02675
R2731 SELECT1.n10 SELECT1.t3 327.99
R2732 SELECT1.n3 SELECT1.t5 293.969
R2733 SELECT1.n6 SELECT1.t7 256.07
R2734 SELECT1.n1 SELECT1.t4 212.081
R2735 SELECT1.n0 SELECT1.t9 212.081
R2736 SELECT1.n10 SELECT1.t2 199.457
R2737 SELECT1.n2 SELECT1.n1 182.929
R2738 SELECT1 SELECT1.n3 154.065
R2739 SELECT1.n11 SELECT1.n10 152
R2740 SELECT1.n7 SELECT1.n6 152
R2741 SELECT1.n6 SELECT1.t6 150.03
R2742 SELECT1.n1 SELECT1.t8 139.78
R2743 SELECT1.n0 SELECT1.t0 139.78
R2744 SELECT1.n3 SELECT1.t1 138.338
R2745 SELECT1.n1 SELECT1.n0 61.346
R2746 SELECT1.n5 SELECT1 22.1096
R2747 SELECT1.n14 SELECT1.n13 14.6836
R2748 SELECT1.n13 SELECT1.n12 14.6704
R2749 SELECT1.n12 SELECT1 13.8672
R2750 SELECT1.n4 SELECT1 13.8328
R2751 SELECT1.n11 SELECT1 12.1605
R2752 SELECT1.n14 SELECT1.n2 10.6811
R2753 SELECT1.n7 SELECT1.n5 10.4374
R2754 SELECT1.n9 SELECT1.n8 8.15359
R2755 SELECT1.n2 SELECT1 6.1445
R2756 SELECT1.n4 SELECT1 5.16179
R2757 SELECT1.n9 SELECT1.n4 4.65206
R2758 SELECT1.n8 SELECT1 3.93896
R2759 SELECT1 SELECT1.n11 2.34717
R2760 SELECT1.n5 SELECT1 2.16665
R2761 SELECT1.n8 SELECT1.n7 1.57588
R2762 SELECT1.n13 SELECT1.n9 0.79438
R2763 SELECT1.n12 SELECT1 0.6405
R2764 SELECT1 SELECT1.n14 0.248606
C0 a_13269_n10693# x2.x2.GN1 3.78e-20
C1 VDD x1.x4.A 15.0138f
C2 x1.x3.GP3 LADDEROUT 0.023203f
C3 x1.x3.GN3 a_4962_n3364# 1.07e-20
C4 RSEL0 a_4962_n4604# 0.246189f
C5 x1.x4.A x1.x3.GN2 0.429208f
C6 R4R5 R7R8 0.286971f
C7 SELECT0 m2_13400_n11836# 0.130999f
C8 x2.x2.GN3 a_13269_n10181# 1.07e-20
C9 x2.x2.GN2 R3R4 0.015379f
C10 x1.x3.GN3 a_4988_n3924# 0.001073f
C11 a_13269_n10869# a_13295_n10741# 0.004764f
C12 SELECT1 x2.x1.nSEL0 0.137679f
C13 a_4988_n4476# x1.x3.GN1 1.22e-20
C14 x2.x1.nSEL1 a_13323_n11699# 0.00175f
C15 VDD x1.x3.GN4 1.35534f
C16 R7R8 x1.x3.GN1 4.45992f
C17 x1.x3.GN4 x1.x3.GN2 0.057602f
C18 VDD m2_13400_n11836# 0.139985f
C19 x2.x1.nSEL1 x2.x2.GN2 0.209956f
C20 R6R7 R7R8 2.27687f
C21 a_13269_n11837# a_13323_n11699# 0.006584f
C22 VDD R1R2 1.61319f
C23 R1R2 x1.x3.GN2 0.006941f
C24 x2.x1.nSEL1 x2.x2.GN1 0.034891f
C25 a_4962_n4052# x1.x3.GN1 7.37e-20
C26 x1.x3.GP3 x1.x4.A 0.358391f
C27 x2.x2.GN2 a_13269_n11837# 0.039612f
C28 x2.x2.GN3 m3_18264_n10402# 0.016026f
C29 x2.x2.GN3 SELECT0 0.254198f
C30 a_13269_n10869# x2.x1.nSEL0 1.91e-20
C31 x2.x2.GN1 a_13269_n11837# 0.12869f
C32 VDD a_5016_n4882# 0.001272f
C33 a_13269_n11245# x2.x2.GN2 0.017018f
C34 a_5016_n4882# x1.x3.GN2 8.86e-19
C35 a_4962_n3876# x1.x1.nSEL0 1.21e-20
C36 x1.x3.GN4 x1.x3.GP3 5.60371f
C37 a_4962_n4604# x1.x5.GN 3.56e-19
C38 x2.x2.GN2 a_13295_n11293# 0.002418f
C39 a_13269_n11245# x2.x2.GN1 1.46e-19
C40 VDD x2.x2.GN3 0.651371f
C41 a_13295_n11293# x2.x2.GN1 1.22e-20
C42 R1R2 x1.x3.GP3 4.25867f
C43 x2.x2.GN4 VRES 0.046938f
C44 RSEL0 x1.x3.GN1 0.020521f
C45 R7R8 VRES 2.33155f
C46 x2.x2.GP3 x2.x2.GN4 3.44338f
C47 a_13269_n11421# LADDEROUT 1.21e-19
C48 OUT SELECT0 4.1e-22
C49 x2.x2.GP3 R7R8 0.17349f
C50 VDD RSEL1 2.66244f
C51 x1.x1.nSEL1 a_4988_n4476# 9.57e-19
C52 RSEL1 x1.x3.GN2 0.108644f
C53 x2.x2.GN4 LADDEROUT 0.085877f
C54 a_13269_n10693# SELECT1 0.127717f
C55 x1.x3.GN3 a_4962_n4604# 6.68e-19
C56 x2.nselect2 LADDEROUT 0.005153f
C57 VDD OUT 11.9877f
C58 a_4962_n5020# a_4962_n4604# 0.002207f
C59 x1.x1.nSEL1 a_4962_n4052# 7.84e-19
C60 SELECT1 a_13323_n10043# 8.84e-19
C61 x1.x3.GN3 R3R4 0.377011f
C62 R5R6 R4R5 2.29244f
C63 m2_5093_n5019# RSEL0 0.130999f
C64 RSEL1 x1.x3.GP3 0.003325f
C65 x2.x2.GN2 VRES 4.02833f
C66 x1.x4.A x2.x2.GN4 0.011047f
C67 x1.x3.GN1 x1.x5.GN 0.645006f
C68 R5R6 x1.x3.GN1 0.250515f
C69 x2.x2.GN1 VRES 2.38e-19
C70 a_4962_n4052# a_4962_n4428# 3.02e-19
C71 x2.x2.GN2 x2.x2.GP3 0.004319f
C72 a_13269_n10693# a_13269_n10869# 0.185422f
C73 VDD RSEL2 4.44873f
C74 x1.x3.GN2 RSEL2 0.001516f
C75 x2.nselect2 x1.x4.A 0.01287f
C76 x1.x3.GN3 R2R3 0.27459f
C77 x2.x1.nSEL1 SELECT1 0.275874f
C78 R5R6 R6R7 2.03637f
C79 x2.x2.GN1 x2.x2.GP3 0.002439f
C80 x1.x3.GN4 x2.x2.GN4 3.13e-20
C81 x2.x2.GN2 LADDEROUT 0.234749f
C82 x1.x1.nSEL1 RSEL0 0.169954f
C83 x1.x3.GN4 R7R8 0.13852f
C84 a_13269_n11837# SELECT1 0.02803f
C85 SELECT0 a_13269_n10181# 0.220366f
C86 x2.x2.GN1 LADDEROUT 4.69118f
C87 R4R5 x1.x3.GN3 0.123865f
C88 a_13269_n11245# SELECT1 0.254026f
C89 a_5016_n3226# x1.x3.GN4 0.001562f
C90 R1R2 R7R8 0.216753f
C91 a_4962_n4052# x1.x3.GN4 6.84e-19
C92 x2.x1.nSEL1 a_13269_n10869# 7.84e-19
C93 x1.x3.GN3 x1.x3.GN1 0.08518f
C94 x1.x3.GP3 RSEL2 1.6e-19
C95 VDD a_13269_n10181# 0.218058f
C96 m2_5093_n5019# x1.x5.GN 4e-19
C97 RSEL0 a_4962_n4428# 0.143958f
C98 a_4962_n5020# x1.x3.GN1 0.128677f
C99 x1.x3.GN3 R6R7 0.260987f
C100 a_13269_n11421# x2.x2.GN3 6.68e-19
C101 x2.x2.GN2 x1.x4.A 1.03e-20
C102 x1.x5.A R3R4 4.07e-21
C103 x2.x2.GN1 x1.x4.A 1.38e-21
C104 x2.x2.GN3 x2.x2.GN4 0.071489f
C105 a_13269_n10869# a_13269_n11245# 3.02e-19
C106 x2.x2.GN3 R7R8 0.012042f
C107 x2.x2.GN3 x2.nselect2 7.39e-21
C108 x1.x1.nSEL1 x1.x5.GN 0.10521f
C109 x1.x3.GN4 RSEL0 0.218342f
C110 LADDEROUT x1.x5.GN 0.820656f
C111 VDD SELECT0 1.59135f
C112 x2.x2.GN1 m2_13400_n11836# 0.06935f
C113 RSEL1 R7R8 4.98e-22
C114 a_4962_n5020# m2_5093_n5019# 0.01297f
C115 x1.x5.GN a_4962_n4428# 3.26e-19
C116 x1.x3.GN3 VRES 0.007817f
C117 OUT x2.x2.GN4 0.446473f
C118 RSEL1 a_5016_n3226# 8.84e-19
C119 x1.x1.nSEL0 a_4962_n4604# 0.03096f
C120 a_4962_n4052# RSEL1 0.261734f
C121 VDD x1.x3.GN2 0.70245f
C122 R4R5 x1.x5.A 4.5151f
C123 OUT R7R8 4.51509f
C124 a_5016_n4882# RSEL0 9.55e-19
C125 x1.x4.A x1.x5.GN 4.14756f
C126 R5R6 x1.x4.A 1.64e-20
C127 x1.x1.nSEL1 x1.x3.GN3 0.012418f
C128 x2.x2.GN2 x2.x2.GN3 0.067572f
C129 x2.x2.GP3 SELECT1 0.003386f
C130 x1.x5.A x1.x3.GN1 0.430802f
C131 x1.x1.nSEL1 a_4962_n5020# 0.193944f
C132 x1.x3.GN3 LADDEROUT 0.014498f
C133 x2.x2.GN1 x2.x2.GN3 0.002859f
C134 x1.x5.A R6R7 4.52052f
C135 SELECT1 LADDEROUT 0.053091f
C136 x1.x3.GN4 x1.x5.GN 9.02e-19
C137 R5R6 x1.x3.GN4 0.304696f
C138 R7R8 RSEL2 0.054741f
C139 VDD x1.x3.GP3 3.24694f
C140 x1.x3.GP3 x1.x3.GN2 0.060312f
C141 x1.x3.GN3 a_4962_n4428# 0.048646f
C142 RSEL1 RSEL0 1.99939f
C143 R3R4 m3_17234_n10416# 0.136776f
C144 a_13269_n10869# x2.x2.GP3 0.00144f
C145 a_4962_n4052# RSEL2 0.009143f
C146 x2.x2.GN2 OUT 0.429399f
C147 x1.x3.GN3 x1.x4.A 0.429865f
C148 a_5016_n4882# x1.x5.GN 1.95e-19
C149 a_13269_n10869# LADDEROUT 0.001506f
C150 x2.x2.GN1 OUT 0.430038f
C151 x1.x4.A SELECT1 0.024025f
C152 a_13269_n10181# x2.x2.GN4 0.134079f
C153 x1.x3.GN3 x1.x3.GN4 0.190989f
C154 x1.x1.nSEL0 x1.x3.GN1 0.002613f
C155 a_4962_n3876# x1.x3.GN1 1.69e-20
C156 x2.nselect2 a_13269_n10181# 9.77e-20
C157 a_13269_n10693# x2.x1.nSEL0 1.21e-20
C158 x2.x1.nSEL1 a_13295_n10741# 4.08e-19
C159 R1R2 x1.x3.GN3 4.03754f
C160 SELECT1 m2_13400_n11836# 0.183786f
C161 RSEL0 RSEL2 0.447568f
C162 R1R2 SELECT1 8.73e-20
C163 x1.x5.A LADDEROUT 4.51865f
C164 RSEL1 x1.x5.GN 0.141315f
C165 a_13269_n10869# x1.x4.A 1.34e-19
C166 a_13269_n11421# SELECT0 0.246189f
C167 x2.x2.GN4 m3_18264_n10402# 0.084813f
C168 SELECT0 x2.x2.GN4 0.218396f
C169 a_4962_n5020# a_5016_n4882# 0.006584f
C170 R7R8 m3_18264_n10402# 0.131878f
C171 x1.x1.nSEL0 m2_5093_n5019# 3.43e-19
C172 x2.x1.nSEL1 x2.x1.nSEL0 0.352716f
C173 x2.nselect2 SELECT0 1.88e-19
C174 VDD a_13269_n11421# 0.161941f
C175 x2.x2.GN2 a_13269_n10181# 7.58e-21
C176 x2.x2.GN3 SELECT1 0.272312f
C177 VDD a_4988_n4476# 5.13e-19
C178 VDD x2.x2.GN4 1.23534f
C179 a_4988_n4476# x1.x3.GN2 0.002395f
C180 x1.x5.A x1.x4.A 2.05508f
C181 VDD R7R8 3.18295f
C182 a_13269_n11837# x2.x1.nSEL0 0.081627f
C183 R7R8 x1.x3.GN2 0.260757f
C184 VDD x2.nselect2 1.22451f
C185 x1.x3.GN3 RSEL1 0.272271f
C186 a_13269_n11245# x2.x1.nSEL0 0.001174f
C187 VDD a_5016_n3226# 8.97e-19
C188 x1.x1.nSEL1 x1.x1.nSEL0 0.352716f
C189 a_4962_n5020# RSEL1 0.02803f
C190 x1.x5.GN RSEL2 3.98693f
C191 R5R6 RSEL2 2.39e-19
C192 a_5016_n3226# x1.x3.GN2 8.14e-21
C193 VDD a_4962_n4052# 0.171399f
C194 x1.x1.nSEL1 a_4962_n3876# 1.59e-19
C195 x1.x5.A x1.x3.GN4 0.446599f
C196 a_4962_n4052# x1.x3.GN2 1.61e-19
C197 a_13295_n11293# x2.x1.nSEL0 2.51e-19
C198 a_13323_n11699# SELECT0 9.55e-19
C199 a_13269_n10869# x2.x2.GN3 0.104343f
C200 m3_17234_n10416# VRES 0.003764f
C201 x2.x2.GN2 SELECT0 0.114345f
C202 x1.x3.GP3 R7R8 0.124327f
C203 x2.x2.GN1 SELECT0 0.020307f
C204 x1.x1.nSEL0 a_4962_n4428# 0.001174f
C205 VDD a_13323_n11699# 9.09e-19
C206 x2.x2.GP3 m3_17234_n10416# 0.002824f
C207 x2.x2.GN2 VDD 0.602533f
C208 a_4962_n4052# x1.x3.GP3 0.001353f
C209 x1.x3.GN3 RSEL2 0.00233f
C210 VDD RSEL0 1.15548f
C211 VDD x2.x2.GN1 1.6041f
C212 a_13295_n10741# x2.x2.GP3 4.39e-19
C213 RSEL0 x1.x3.GN2 0.114399f
C214 a_4962_n5020# RSEL2 4.33e-19
C215 SELECT1 RSEL2 9.2e-20
C216 a_13295_n10741# LADDEROUT 1.48e-19
C217 x1.x1.nSEL0 x1.x3.GN4 2.26e-20
C218 x2.x1.nSEL1 a_13269_n10693# 1.59e-19
C219 a_4962_n3876# x1.x3.GN4 0.003645f
C220 x1.x3.GP3 RSEL0 2.74e-19
C221 x1.x3.GN3 a_13269_n10181# 1.84e-20
C222 R2R3 R3R4 2.48395f
C223 SELECT1 a_13269_n10181# 0.125445f
C224 x1.x1.nSEL1 a_4988_n3924# 4.08e-19
C225 LADDEROUT x2.x1.nSEL0 9.01e-20
C226 a_13295_n10741# x1.x4.A 3.86e-20
C227 VDD x1.x5.GN 3.72608f
C228 R5R6 VDD 1.61253f
C229 x1.x3.GN2 x1.x5.GN 7.45e-19
C230 R5R6 x1.x3.GN2 0.122632f
C231 R4R5 R3R4 1.39313f
C232 a_4962_n4604# x1.x3.GN1 0.012357f
C233 x2.x1.nSEL1 a_13269_n11837# 0.193944f
C234 x2.x2.GN4 R7R8 3.97959f
C235 x2.nselect2 x2.x2.GN4 1.53e-20
C236 x1.x5.A RSEL2 5.67943f
C237 x1.x3.GN1 R3R4 3.99708f
C238 x2.x1.nSEL1 a_13269_n11245# 0.041068f
C239 x1.x1.nSEL0 RSEL1 0.137595f
C240 a_4962_n3876# RSEL1 0.127717f
C241 x2.x1.nSEL1 a_13295_n11293# 9.57e-19
C242 x1.x4.A x2.x1.nSEL0 6.2e-20
C243 SELECT0 SELECT1 1.68437f
C244 x1.x3.GP3 x1.x5.GN 3.82e-20
C245 a_4962_n4052# R7R8 7.47e-21
C246 R4R5 R2R3 7.85e-20
C247 R5R6 x1.x3.GP3 4.11452f
C248 x2.x2.GN3 m3_17234_n10416# 0.087318f
C249 VDD x1.x3.GN3 0.767502f
C250 x1.x3.GN3 x1.x3.GN2 0.175465f
C251 a_4962_n3364# x1.x3.GN4 0.134079f
C252 VDD a_4962_n5020# 0.21327f
C253 a_4962_n5020# x1.x3.GN2 0.039612f
C254 R2R3 x1.x3.GN1 2.57e-19
C255 VDD SELECT1 3.24319f
C256 x1.x3.GN4 a_4988_n3924# 3.22e-19
C257 x2.x1.nSEL0 m2_13400_n11836# 3.43e-19
C258 x2.x2.GN2 a_13269_n11421# 0.106186f
C259 x2.x2.GN3 a_13295_n10741# 0.001073f
C260 a_13269_n11421# x2.x2.GN1 0.012466f
C261 a_13269_n10869# SELECT0 0.086353f
C262 x2.x2.GN2 x2.x2.GN4 8.84e-19
C263 R4R5 x1.x3.GN1 0.334962f
C264 a_13269_n10693# x2.x2.GP3 5.21e-19
C265 x2.x2.GN2 R7R8 1.22e-19
C266 x2.x2.GN1 x2.x2.GN4 0.001074f
C267 x1.x1.nSEL0 RSEL2 0.131256f
C268 R3R4 VRES 3.1523f
C269 RSEL0 R7R8 2.25e-21
C270 x1.x3.GN3 x1.x3.GP3 5.0197f
C271 R4R5 R6R7 2.49e-19
C272 a_13269_n10693# LADDEROUT 9.74e-19
C273 a_13269_n10869# VDD 0.180589f
C274 x1.x1.nSEL1 a_4962_n4604# 0.073392f
C275 x2.x2.GP3 R3R4 4.09932f
C276 a_13323_n10043# LADDEROUT 3.17e-19
C277 a_5016_n3226# RSEL0 1.4e-19
C278 R6R7 x1.x3.GN1 0.254378f
C279 a_4962_n4052# RSEL0 0.086353f
C280 x2.x2.GN3 x2.x1.nSEL0 4.01e-20
C281 LADDEROUT R3R4 0.039417f
C282 R2R3 VRES 2.39e-19
C283 x2.x2.GN2 a_13323_n11699# 8.86e-19
C284 a_4962_n4604# a_4962_n4428# 0.185422f
C285 RSEL1 a_4962_n3364# 0.125445f
C286 x2.x2.GN1 a_13323_n11699# 0.001144f
C287 a_13269_n10693# x1.x4.A 3.32e-19
C288 VDD x1.x5.A 14.1643f
C289 x1.x5.A x1.x3.GN2 0.429382f
C290 x1.x4.A a_13323_n10043# 2.9e-19
C291 m2_5093_n5019# x1.x3.GN1 0.06935f
C292 a_4988_n4476# x1.x5.GN 1.08e-19
C293 x2.x2.GN2 x2.x2.GN1 0.065208f
C294 R2R3 LADDEROUT 0.017699f
C295 R7R8 x1.x5.GN 0.558172f
C296 R5R6 R7R8 0.318606f
C297 x2.nselect2 x1.x5.GN 4.76e-21
C298 x1.x4.A R3R4 4.53278f
C299 a_4962_n4052# x1.x5.GN 3.51e-19
C300 x1.x3.GN4 R3R4 0.237845f
C301 x1.x5.A x1.x3.GP3 0.358718f
C302 x1.x1.nSEL1 x1.x3.GN1 0.034871f
C303 x1.x3.GN1 LADDEROUT 4.27e-20
C304 R2R3 x1.x4.A 4.52053f
C305 R1R2 R3R4 0.184502f
C306 a_13269_n11421# SELECT1 0.03417f
C307 x1.x3.GN3 a_4988_n4476# 5.17e-20
C308 x1.x3.GN3 x2.x2.GN4 8.02e-21
C309 x1.x3.GN3 R7R8 0.129387f
C310 VDD x1.x1.nSEL0 0.3889f
C311 x1.x1.nSEL0 x1.x3.GN2 0.154394f
C312 SELECT1 x2.x2.GN4 0.059813f
C313 VDD a_4962_n3876# 0.262163f
C314 x2.x1.nSEL1 m2_13400_n11836# 0.00815f
C315 a_4962_n3876# x1.x3.GN2 9.62e-20
C316 R2R3 x1.x3.GN4 0.127088f
C317 a_13269_n10693# x2.x2.GN3 0.004288f
C318 x1.x3.GN1 a_4962_n4428# 1.45e-19
C319 R4R5 x1.x4.A 0.003925f
C320 x2.nselect2 SELECT1 0.001201f
C321 m3_17234_n10416# m3_18264_n10402# 0.003741f
C322 x1.x3.GN3 a_5016_n3226# 1.07e-20
C323 RSEL0 x1.x5.GN 0.136598f
C324 x1.x3.GN3 a_4962_n4052# 0.104374f
C325 x2.x2.GN3 a_13323_n10043# 1.07e-20
C326 a_13269_n11837# m2_13400_n11836# 0.01297f
C327 R1R2 R2R3 1.9897f
C328 x1.x4.A x1.x3.GN1 0.428132f
C329 x1.x1.nSEL1 m2_5093_n5019# 0.00815f
C330 x2.x2.GN3 R3R4 3.96252f
C331 R4R5 x1.x3.GN4 4.23591f
C332 x2.x2.GP3 VRES 0.050501f
C333 a_13295_n10741# SELECT0 0.001558f
C334 a_13269_n10869# x2.x2.GN4 6.84e-19
C335 RSEL1 a_4962_n4604# 0.03417f
C336 a_4962_n3876# x1.x3.GP3 4.69e-19
C337 x1.x3.GN4 x1.x3.GN1 0.142035f
C338 LADDEROUT VRES 1.8361f
C339 x2.x1.nSEL1 x2.x2.GN3 0.012418f
C340 a_13269_n10869# x2.nselect2 1.29e-19
C341 x1.x3.GN4 R6R7 0.156481f
C342 VDD a_13295_n10741# 0.001496f
C343 x2.x2.GP3 LADDEROUT 0.084041f
C344 x1.x3.GN3 RSEL0 0.254198f
C345 x2.x2.GN2 SELECT1 0.108649f
C346 a_4962_n5020# RSEL0 0.048888f
C347 OUT R3R4 4.52137f
C348 x2.x2.GN1 SELECT1 0.312198f
C349 R5R6 x1.x5.GN 7.03e-21
C350 SELECT0 x2.x1.nSEL0 0.326696f
C351 a_13269_n11245# x2.x2.GN3 0.048646f
C352 a_5016_n4882# x1.x3.GN1 0.001144f
C353 x1.x5.A R7R8 4.52065f
C354 a_13295_n11293# x2.x2.GN3 5.17e-20
C355 x1.x4.A VRES 4.51511f
C356 x1.x1.nSEL1 a_4962_n4428# 0.041068f
C357 a_4962_n4604# RSEL2 8.66e-20
C358 VDD a_4962_n3364# 0.217381f
C359 a_4962_n3364# x1.x3.GN2 7.58e-21
C360 VDD x2.x1.nSEL0 0.523674f
C361 x2.x2.GP3 x1.x4.A 0.005595f
C362 a_13269_n10869# x2.x2.GN2 1.63e-19
C363 VDD a_4988_n3924# 0.001496f
C364 a_4988_n3924# x1.x3.GN2 3.11e-20
C365 R3R4 RSEL2 2.94e-19
C366 x1.x3.GN4 VRES 4.10935f
C367 a_13269_n10869# x2.x2.GN1 6.43e-20
C368 x1.x4.A LADDEROUT 6.48818f
C369 x2.x2.GP3 x1.x3.GN4 2.78e-20
C370 RSEL1 x1.x3.GN1 0.312176f
C371 R1R2 VRES 2.31469f
C372 x1.x3.GN3 x1.x5.GN 1.63e-19
C373 R5R6 x1.x3.GN3 4.12614f
C374 a_4962_n5020# x1.x5.GN 0.001336f
C375 x2.x1.nSEL1 RSEL2 9.21e-21
C376 x1.x3.GN4 LADDEROUT 0.014367f
C377 a_13269_n10181# a_13323_n10043# 0.006584f
C378 x1.x1.nSEL0 a_4988_n4476# 2.51e-19
C379 a_4988_n3924# x1.x3.GP3 4.39e-19
C380 R1R2 LADDEROUT 0.017912f
C381 a_4962_n3876# R7R8 7.47e-21
C382 x2.x2.GN3 VRES 0.214839f
C383 R4R5 RSEL2 6.76e-20
C384 x1.x1.nSEL1 a_5016_n4882# 0.00175f
C385 a_4962_n4052# x1.x1.nSEL0 1.91e-20
C386 a_4962_n3876# a_4962_n4052# 0.185422f
C387 m2_5093_n5019# RSEL1 0.183786f
C388 x2.x2.GN3 x2.x2.GP3 2.86799f
C389 x1.x3.GN4 x1.x4.A 0.446539f
C390 a_13269_n10693# SELECT0 0.279858f
C391 x1.x3.GN1 RSEL2 0.054258f
C392 x2.x2.GN4 m3_17234_n10416# 7.07e-19
C393 x1.x3.GN3 SELECT1 7.93e-20
C394 SELECT0 a_13323_n10043# 1.4e-19
C395 R7R8 m3_17234_n10416# 0.001045f
C396 x2.x2.GN3 LADDEROUT 0.087953f
C397 R1R2 x1.x4.A 4.5214f
C398 R3R4 m3_18264_n10402# 1.46e-19
C399 a_13269_n10693# VDD 0.262214f
C400 a_13295_n10741# x2.x2.GN4 3.22e-19
C401 x1.x1.nSEL1 RSEL1 0.275603f
C402 OUT VRES 4.5205f
C403 VDD a_13323_n10043# 8.97e-19
C404 VDD a_4962_n4604# 0.164566f
C405 a_4962_n4604# x1.x3.GN2 0.106139f
C406 R1R2 x1.x3.GN4 0.628977f
C407 x1.x5.A x1.x5.GN 4.01011f
C408 R5R6 x1.x5.A 4.5214f
C409 x1.x1.nSEL0 RSEL0 0.325123f
C410 a_4962_n3876# RSEL0 0.279858f
C411 x2.x2.GP3 OUT 0.357868f
C412 x2.x1.nSEL1 SELECT0 0.168511f
C413 VDD R3R4 3.2635f
C414 x1.x3.GN2 R3R4 0.271818f
C415 m2_5093_n5019# RSEL2 4.4e-19
C416 a_13269_n10869# SELECT1 0.261734f
C417 x2.x2.GN3 x1.x4.A 8.22e-19
C418 OUT LADDEROUT 4.51998f
C419 a_13269_n11421# x2.x1.nSEL0 0.03096f
C420 a_13269_n11837# SELECT0 0.048888f
C421 RSEL1 a_4962_n4428# 0.254026f
C422 x2.x1.nSEL1 VDD 0.649185f
C423 x2.x2.GN4 x2.x1.nSEL0 2.26e-20
C424 x2.x2.GN2 m3_17234_n10416# 0.016745f
C425 a_13269_n11245# SELECT0 0.143958f
C426 x2.x2.GN3 x1.x3.GN4 1.1e-19
C427 VDD R2R3 1.6072f
C428 R2R3 x1.x3.GN2 3.9984f
C429 VDD a_13269_n11837# 0.211573f
C430 a_4962_n3364# a_5016_n3226# 0.006584f
C431 x1.x3.GP3 R3R4 0.384927f
C432 x1.x5.A x1.x3.GN3 0.429924f
C433 x1.x1.nSEL1 RSEL2 0.164995f
C434 x2.x2.GN2 a_13295_n10741# 3.11e-20
C435 LADDEROUT RSEL2 0.781024f
C436 a_13269_n11245# VDD 0.193307f
C437 a_4962_n4052# a_4988_n3924# 0.004764f
C438 RSEL1 x1.x3.GN4 0.059776f
C439 R4R5 VDD 1.56678f
C440 x1.x1.nSEL0 x1.x5.GN 0.043717f
C441 R4R5 x1.x3.GN2 0.116214f
C442 a_4962_n3876# x1.x5.GN 2.27e-19
C443 VDD a_13295_n11293# 4.32e-19
C444 VDD x1.x3.GN1 0.915728f
C445 x1.x3.GN1 x1.x3.GN2 0.143294f
C446 R2R3 x1.x3.GP3 0.115126f
C447 a_4962_n4428# RSEL2 1.67e-19
C448 VDD R6R7 1.6078f
C449 R6R7 x1.x3.GN2 4.03744f
C450 x2.x2.GN2 x2.x1.nSEL0 0.154394f
C451 x1.x4.A RSEL2 4.96785f
C452 a_4962_n3364# RSEL0 0.220366f
C453 a_13269_n10181# LADDEROUT 0.003273f
C454 x2.x2.GN1 x2.x1.nSEL0 0.004383f
C455 R4R5 x1.x3.GP3 0.346864f
C456 a_4988_n3924# RSEL0 0.001558f
C457 x1.x3.GN3 x1.x1.nSEL0 4.01e-20
C458 x1.x3.GN3 a_4962_n3876# 0.004289f
C459 x1.x3.GN4 RSEL2 5.71e-20
C460 x1.x3.GP3 x1.x3.GN1 0.075686f
C461 a_4962_n5020# x1.x1.nSEL0 0.081627f
C462 VDD m2_5093_n5019# 0.140894f
C463 x2.x2.GP3 m3_18264_n10402# 0.006132f
C464 x1.x3.GP3 R6R7 0.122655f
C465 a_13269_n10693# x2.x2.GN4 0.003699f
C466 x2.x2.GP3 SELECT0 2.82e-19
C467 x2.x2.GN3 OUT 0.429994f
C468 a_13323_n10043# x2.x2.GN4 0.001562f
C469 x1.x4.A a_13269_n10181# 0.001685f
C470 a_4962_n4604# a_4988_n4476# 0.004764f
C471 a_13269_n10693# x2.nselect2 6.01e-20
C472 VDD VRES 3.15952f
C473 SELECT0 LADDEROUT 0.022124f
C474 x2.x2.GN4 R3R4 0.269437f
C475 VDD x2.x2.GP3 1.78354f
C476 R7R8 R3R4 5.65992f
C477 a_4962_n3364# x1.x5.GN 1.19e-19
C478 VDD x1.x1.nSEL1 0.474773f
C479 x1.x1.nSEL1 x1.x3.GN2 0.209954f
C480 x2.x1.nSEL1 a_13269_n11421# 0.073392f
C481 a_4988_n3924# x1.x5.GN 9.76e-20
C482 VDD LADDEROUT 9.0607f
C483 LADDEROUT x1.x3.GN2 0.01442f
C484 R1R2 a_13269_n10181# 5.05e-21
C485 a_13269_n11421# a_13269_n11837# 0.002207f
C486 x1.x3.GP3 VRES 0.17111f
C487 x2.x1.nSEL1 x2.nselect2 0.047548f
C488 x1.x4.A SELECT0 0.001236f
C489 R2R3 R7R8 0.215077f
C490 a_13269_n11245# a_13269_n11421# 0.185422f
C491 VDD a_4962_n4428# 0.194316f
C492 x1.x3.GN2 a_4962_n4428# 0.016995f
C493 a_13269_n10693# x2.x2.GN2 5.62e-20
C494 RSEL1 RSEL2 0.460661f
C495 a_13269_n11421# a_13295_n11293# 0.004764f
C496 x2.x2.GN2 a_13323_n10043# 8.14e-21
C497 OUT VSS 12.417253f
C498 SELECT0 VSS 1.58526f
C499 SELECT1 VSS 2.059261f
C500 LADDEROUT VSS 14.893856f
C501 RSEL2 VSS 7.005585f
C502 RSEL0 VSS 1.61007f
C503 RSEL1 VSS 1.729297f
C504 VRES VSS 21.573582f
C505 VDD VSS 0.179412p
C506 m3_18264_n10402# VSS 0.066786f $ **FLOATING
C507 m3_17234_n10416# VSS 0.064102f $ **FLOATING
C508 m2_13400_n11836# VSS 0.065655f $ **FLOATING
C509 m2_5093_n5019# VSS 0.065655f $ **FLOATING
C510 a_13323_n11699# VSS 0.006505f
C511 a_13269_n11837# VSS 0.266782f
C512 x2.x1.nSEL0 VSS 0.647728f
C513 x2.x2.GN1 VSS 6.304735f
C514 a_13295_n11293# VSS 0.004461f
C515 a_13269_n11421# VSS 0.220868f
C516 x2.x1.nSEL1 VSS 0.686216f
C517 x2.x2.GN2 VSS 3.88916f
C518 a_13269_n11245# VSS 0.23458f
C519 x2.nselect2 VSS 0.451687f
C520 x2.x2.GP3 VSS 1.68642f
C521 a_13295_n10741# VSS 0.006801f
C522 x2.x2.GN3 VSS 3.65643f
C523 a_13269_n10869# VSS 0.232764f
C524 a_13269_n10693# VSS 0.249604f
C525 x2.x2.GN4 VSS 7.65266f
C526 a_13323_n10043# VSS 0.006439f
C527 a_13269_n10181# VSS 0.305716f
C528 x1.x4.A VSS 16.1289f
C529 x1.x5.A VSS 16.690754f
C530 a_5016_n4882# VSS 0.006505f
C531 a_4962_n5020# VSS 0.266782f
C532 x1.x1.nSEL0 VSS 0.650696f
C533 x1.x3.GN1 VSS 11.747699f
C534 a_4988_n4476# VSS 0.004461f
C535 a_4962_n4604# VSS 0.220868f
C536 x1.x1.nSEL1 VSS 0.682637f
C537 x1.x3.GN2 VSS 7.17674f
C538 a_4962_n4428# VSS 0.23458f
C539 x1.x5.GN VSS 5.76746f
C540 x1.x3.GP3 VSS 3.18403f
C541 a_4988_n3924# VSS 0.006801f
C542 x1.x3.GN3 VSS 6.77774f
C543 a_4962_n4052# VSS 0.232731f
C544 a_4962_n3876# VSS 0.249604f
C545 x1.x3.GN4 VSS 13.651645f
C546 a_5016_n3226# VSS 0.006583f
C547 a_4962_n3364# VSS 0.307394f
C548 R1R2 VSS 7.723106f
C549 R2R3 VSS 7.487107f
C550 R3R4 VSS 16.88881f
C551 R4R5 VSS 7.097775f
C552 R5R6 VSS 6.679734f
C553 R6R7 VSS 9.022429f
C554 R7R8 VSS 28.787964f
C555 SELECT1.t4 VSS 0.034541f
C556 SELECT1.t8 VSS 0.020355f
C557 SELECT1.t9 VSS 0.034541f
C558 SELECT1.t0 VSS 0.020355f
C559 SELECT1.n0 VSS 0.057955f
C560 SELECT1.n1 VSS 0.085627f
C561 SELECT1.n2 VSS 0.052137f
C562 SELECT1.t1 VSS 0.015983f
C563 SELECT1.t5 VSS 0.033707f
C564 SELECT1.n3 VSS 0.121038f
C565 SELECT1.n4 VSS 0.023468f
C566 SELECT1.n5 VSS 0.020215f
C567 SELECT1.t7 VSS 0.024351f
C568 SELECT1.t6 VSS 0.016734f
C569 SELECT1.n6 VSS 0.070762f
C570 SELECT1.n7 VSS 0.0163f
C571 SELECT1.n8 VSS 0.116761f
C572 SELECT1.n9 VSS 0.42291f
C573 SELECT1.t3 VSS 0.029668f
C574 SELECT1.t2 VSS 0.020145f
C575 SELECT1.n10 VSS 0.070094f
C576 SELECT1.n11 VSS 0.016777f
C577 SELECT1.n12 VSS 0.108827f
C578 SELECT1.n13 VSS 0.488144f
C579 SELECT1.n14 VSS 0.637714f
C580 R2R3.t2 VSS 0.615655f
C581 R2R3.t1 VSS 0.353436f
C582 R2R3.n0 VSS 3.42308f
C583 R2R3.t4 VSS 0.63721f
C584 R2R3.t3 VSS 0.450767f
C585 R2R3.n1 VSS 3.49982f
C586 R2R3.n2 VSS 0.553581f
C587 R2R3.n3 VSS 0.118679f
C588 R2R3.t0 VSS 0.214449f
C589 R2R3.t5 VSS 0.172939f
C590 R2R3.n4 VSS 3.41696f
C591 R2R3.n5 VSS 0.546763f
C592 R5R6.t1 VSS 0.691407f
C593 R5R6.t0 VSS 0.396924f
C594 R5R6.n0 VSS 3.84427f
C595 R5R6.t4 VSS 0.715614f
C596 R5R6.t3 VSS 0.506231f
C597 R5R6.n1 VSS 3.93045f
C598 R5R6.n2 VSS 0.621695f
C599 R5R6.n3 VSS 0.133787f
C600 R5R6.t5 VSS 0.197046f
C601 R5R6.t2 VSS 0.241304f
C602 R5R6.n4 VSS 3.70778f
C603 R5R6.n5 VSS 1.25933f
C604 x2.x2.x2.GP VSS 2.80012f
C605 x2.x1.gpo1 VSS 1.00993f
C606 x2.x2.GP2.t0 VSS 0.016198f
C607 x2.x2.GP2.t1 VSS 0.016198f
C608 x2.x2.GP2.n0 VSS 0.038624f
C609 x2.x1.x12.Y VSS 0.058789f
C610 x2.x2.GP2.n1 VSS 0.075879f
C611 x2.x2.GP2.n2 VSS 0.023609f
C612 x2.x2.GP2.t2 VSS 0.02492f
C613 x2.x2.GP2.t3 VSS 0.02492f
C614 x2.x2.GP2.n3 VSS 0.051391f
C615 x2.x2.GP2.t5 VSS 0.819753f
C616 x2.x2.GP2.t4 VSS 0.842612f
C617 x2.x2.GP2.n4 VSS 2.98946f
C618 x2.x2.GP2.n5 VSS 0.107597f
C619 x1.x3.x2.GP VSS 3.47156f
C620 x1.x2.x2.GP VSS 2.5351f
C621 x1.x1.gpo1 VSS 0.999009f
C622 x1.x3.GP2.t1 VSS 0.018287f
C623 x1.x3.GP2.t0 VSS 0.018287f
C624 x1.x3.GP2.n0 VSS 0.043605f
C625 x1.x1.x12.Y VSS 0.066371f
C626 x1.x3.GP2.n1 VSS 0.085666f
C627 x1.x3.GP2.n2 VSS 0.026654f
C628 x1.x3.GP2.t5 VSS 0.925483f
C629 x1.x3.GP2.t4 VSS 0.95129f
C630 x1.x3.GP2.n3 VSS 3.37503f
C631 x1.x3.GP2.t7 VSS 0.925483f
C632 x1.x3.GP2.t6 VSS 0.95129f
C633 x1.x3.GP2.n4 VSS 3.37503f
C634 x1.x3.GP2.n5 VSS 1.99609f
C635 x1.x3.GP2.t2 VSS 0.028134f
C636 x1.x3.GP2.t3 VSS 0.028134f
C637 x1.x3.GP2.n6 VSS 0.058019f
C638 x1.x3.GP2.n7 VSS 0.121475f
C639 x1.x3.x1.GP VSS 3.45389f
C640 x1.x2.GP1 VSS 2.34975f
C641 x1.x1.gpo0 VSS 0.786924f
C642 x1.x3.GP1.t0 VSS 0.018021f
C643 x1.x3.GP1.t1 VSS 0.018021f
C644 x1.x3.GP1.n0 VSS 0.042971f
C645 x1.x1.x11.Y VSS 0.06574f
C646 x1.x3.GP1.n1 VSS 0.084421f
C647 x1.x3.GP1.n2 VSS 0.026267f
C648 x1.x3.GP1.t6 VSS 0.912037f
C649 x1.x3.GP1.t5 VSS 0.93747f
C650 x1.x3.GP1.n3 VSS 3.31176f
C651 x1.x3.GP1.t4 VSS 0.912037f
C652 x1.x3.GP1.t7 VSS 0.93747f
C653 x1.x3.GP1.n4 VSS 3.34441f
C654 x1.x3.GP1.n5 VSS 1.76427f
C655 x1.x3.GP1.t2 VSS 0.027725f
C656 x1.x3.GP1.t3 VSS 0.027725f
C657 x1.x3.GP1.n6 VSS 0.057129f
C658 x1.x3.GP1.n7 VSS 0.121965f
C659 x2.x2.GN4.t0 VSS 0.061896f
C660 x2.x2.GN4.n0 VSS 0.071351f
C661 x2.x2.GN4.t6 VSS 0.699487f
C662 x2.x2.GN4.t5 VSS 0.68261f
C663 x2.x2.GN4.n1 VSS 3.06261f
C664 x2.x2.GN4.n2 VSS 1.5761f
C665 x2.x2.GN4.t7 VSS 0.038856f
C666 x2.x2.GN4.t3 VSS 0.022897f
C667 x2.x2.GN4.t2 VSS 0.038856f
C668 x2.x2.GN4.t4 VSS 0.022897f
C669 x2.x2.GN4.n3 VSS 0.065194f
C670 x2.x2.GN4.n4 VSS 0.096578f
C671 x2.x2.GN4.n5 VSS 0.043236f
C672 x2.x2.GN4.n6 VSS 0.35022f
C673 x2.x2.GN4.t1 VSS 0.158077f
C674 x2.x2.GN4.n7 VSS 0.028433f
C675 x2.x2.GN4.n8 VSS 0.031852f
C676 x2.x2.x1.GP VSS 2.01575f
C677 x2.x2.GP1.t1 VSS 0.012908f
C678 x2.x2.GP1.t0 VSS 0.012908f
C679 x2.x2.GP1.n0 VSS 0.030779f
C680 x2.x1.x11.Y VSS 0.047088f
C681 x2.x2.GP1.n1 VSS 0.060469f
C682 x2.x2.GP1.n2 VSS 0.018815f
C683 x2.x2.GP1.t2 VSS 0.019859f
C684 x2.x2.GP1.t3 VSS 0.019859f
C685 x2.x2.GP1.n3 VSS 0.04092f
C686 x2.x2.GP1.t5 VSS 0.653268f
C687 x2.x2.GP1.t4 VSS 0.671485f
C688 x2.x2.GP1.n4 VSS 2.37213f
C689 x2.x1.gpo0 VSS 0.636407f
C690 x2.x2.GP1.n5 VSS 0.08736f
C691 x2.x2.GN1.t0 VSS 0.030649f
C692 x2.x2.GN1.n0 VSS 0.035367f
C693 x2.x2.GN1.t6 VSS 0.346364f
C694 x2.x2.GN1.t7 VSS 0.338008f
C695 x2.x2.GN1.n1 VSS 1.51651f
C696 x2.x2.GN1.n2 VSS 0.529016f
C697 x2.x2.GN1.t3 VSS 0.01924f
C698 x2.x2.GN1.t4 VSS 0.011338f
C699 x2.x2.GN1.t5 VSS 0.01924f
C700 x2.x2.GN1.t2 VSS 0.011338f
C701 x2.x2.GN1.n3 VSS 0.032282f
C702 x2.x2.GN1.n4 VSS 0.047681f
C703 x2.x2.GN1.n5 VSS 0.046375f
C704 x2.x2.GN1.n6 VSS 0.10073f
C705 x2.x2.GN1.t1 VSS 0.078275f
C706 x2.x2.GN1.n7 VSS 0.014079f
C707 x2.x2.GN1.n8 VSS 0.015772f
C708 OUT.t7 VSS 0.326448f
C709 OUT.n0 VSS 0.487446f
C710 OUT.t1 VSS 0.333001f
C711 OUT.t5 VSS 0.4419f
C712 OUT.n1 VSS 2.22996f
C713 OUT.n2 VSS 0.754525f
C714 OUT.t2 VSS 0.430058f
C715 OUT.n3 VSS 0.534864f
C716 OUT.n4 VSS 0.670409f
C717 OUT.n5 VSS 0.349688f
C718 OUT.t8 VSS 0.326448f
C719 OUT.n6 VSS 0.487446f
C720 OUT.t9 VSS 0.333001f
C721 OUT.t3 VSS 0.4419f
C722 OUT.n7 VSS 2.22996f
C723 OUT.n8 VSS 0.754525f
C724 OUT.t6 VSS 0.430058f
C725 OUT.n9 VSS 0.534864f
C726 OUT.n10 VSS 0.659134f
C727 OUT.n11 VSS 0.291304f
C728 OUT.t14 VSS 0.326448f
C729 OUT.n12 VSS 0.487446f
C730 OUT.t15 VSS 0.333001f
C731 OUT.t11 VSS 0.4419f
C732 OUT.n13 VSS 2.22996f
C733 OUT.n14 VSS 0.754525f
C734 OUT.t10 VSS 0.430058f
C735 OUT.n15 VSS 0.534864f
C736 OUT.n16 VSS 0.657095f
C737 OUT.n17 VSS 0.299286f
C738 OUT.t0 VSS 0.326448f
C739 OUT.n18 VSS 0.487446f
C740 OUT.t4 VSS 0.333001f
C741 OUT.t13 VSS 0.4419f
C742 OUT.n19 VSS 2.22996f
C743 OUT.n20 VSS 0.754525f
C744 OUT.t12 VSS 0.430058f
C745 OUT.n21 VSS 0.534864f
C746 OUT.n22 VSS 0.679666f
C747 OUT.n23 VSS 1.00113f
C748 OUT.n24 VSS 0.948465f
C749 OUT.n25 VSS 0.561092f
C750 OUT.n26 VSS 0.007173f
C751 OUT.n27 VSS 0.004593f
C752 x2.x2.GP4.n0 VSS 0.09812f
C753 x2.x2.x4.GP VSS 2.57224f
C754 x2.x1.gpo3 VSS 1.21226f
C755 x2.x2.GP4.t2 VSS 0.012374f
C756 x2.x2.GP4.t0 VSS 0.012374f
C757 x2.x2.GP4.n1 VSS 0.029505f
C758 x2.x1.x14.Y VSS 0.106946f
C759 x2.x2.GP4.t4 VSS 0.626222f
C760 x2.x2.GP4.t5 VSS 0.643684f
C761 x2.x2.GP4.n2 VSS 2.28835f
C762 x2.x2.GP4.n3 VSS 0.018036f
C763 x2.x2.GP4.t1 VSS 0.019037f
C764 x2.x2.GP4.t3 VSS 0.019037f
C765 x2.x2.GP4.n4 VSS 0.041808f
C766 x1.x3.GN4.t0 VSS 0.055031f
C767 x1.x3.GN4.n0 VSS 0.063437f
C768 x1.x3.GN4.t7 VSS 0.621905f
C769 x1.x3.GN4.t5 VSS 0.606901f
C770 x1.x3.GN4.n1 VSS 2.72293f
C771 x1.x3.GN4.n2 VSS 1.68296f
C772 x1.x3.GN4.t2 VSS 0.621905f
C773 x1.x3.GN4.t3 VSS 0.606901f
C774 x1.x3.GN4.n3 VSS 2.72293f
C775 x1.x3.GN4.n4 VSS 2.3865f
C776 x1.x3.GN4.t4 VSS 0.034546f
C777 x1.x3.GN4.t8 VSS 0.020358f
C778 x1.x3.GN4.t6 VSS 0.034546f
C779 x1.x3.GN4.t9 VSS 0.020358f
C780 x1.x3.GN4.n5 VSS 0.057963f
C781 x1.x3.GN4.n6 VSS 0.085867f
C782 x1.x3.GN4.n7 VSS 0.038441f
C783 x1.x3.GN4.n8 VSS 0.311376f
C784 x1.x3.GN4.t1 VSS 0.140544f
C785 x1.x3.GN4.n9 VSS 0.025279f
C786 x1.x3.GN4.n10 VSS 0.028319f
C787 RSEL1.t2 VSS 0.027818f
C788 RSEL1.t5 VSS 0.016393f
C789 RSEL1.t4 VSS 0.027818f
C790 RSEL1.t1 VSS 0.016393f
C791 RSEL1.n0 VSS 0.046674f
C792 RSEL1.n1 VSS 0.06896f
C793 RSEL1.n2 VSS 0.041989f
C794 RSEL1.t7 VSS 0.012872f
C795 RSEL1.t6 VSS 0.027146f
C796 RSEL1.n3 VSS 0.097478f
C797 RSEL1.n4 VSS 0.0189f
C798 RSEL1.n5 VSS 0.01628f
C799 RSEL1.t8 VSS 0.019611f
C800 RSEL1.t0 VSS 0.013477f
C801 RSEL1.n6 VSS 0.056989f
C802 RSEL1.n7 VSS 0.013127f
C803 RSEL1.n8 VSS 0.094034f
C804 RSEL1.n9 VSS 0.340592f
C805 RSEL1.t9 VSS 0.023893f
C806 RSEL1.t3 VSS 0.016224f
C807 RSEL1.n10 VSS 0.05645f
C808 RSEL1.n11 VSS 0.013512f
C809 RSEL1.n12 VSS 0.087644f
C810 RSEL1.n13 VSS 0.393129f
C811 RSEL1.n14 VSS 0.513585f
C812 RSEL1.n15 VSS 0.158305f
C813 RSEL1.n16 VSS 0.23977f
C814 LADDEROUT.t7 VSS 0.659335f
C815 LADDEROUT.t0 VSS 0.378512f
C816 LADDEROUT.n0 VSS 3.66595f
C817 LADDEROUT.t1 VSS 0.682419f
C818 LADDEROUT.t6 VSS 0.482749f
C819 LADDEROUT.n1 VSS 3.74813f
C820 LADDEROUT.n2 VSS 0.592857f
C821 LADDEROUT.n3 VSS 0.154944f
C822 LADDEROUT.t8 VSS 0.474909f
C823 LADDEROUT.n4 VSS 0.590645f
C824 LADDEROUT.t9 VSS 0.487986f
C825 LADDEROUT.t3 VSS 0.36773f
C826 LADDEROUT.n5 VSS 2.46252f
C827 LADDEROUT.n6 VSS 0.833214f
C828 LADDEROUT.t2 VSS 0.360494f
C829 LADDEROUT.n7 VSS 0.538282f
C830 LADDEROUT.n8 VSS 0.709121f
C831 LADDEROUT.n9 VSS 0.609248f
C832 LADDEROUT.n10 VSS 3.28319f
C833 LADDEROUT.t5 VSS 0.474909f
C834 LADDEROUT.n11 VSS 0.590645f
C835 LADDEROUT.t4 VSS 0.487986f
C836 LADDEROUT.t10 VSS 0.36773f
C837 LADDEROUT.n12 VSS 2.46252f
C838 LADDEROUT.n13 VSS 0.833214f
C839 LADDEROUT.t11 VSS 0.360494f
C840 LADDEROUT.n14 VSS 0.538282f
C841 LADDEROUT.n15 VSS 0.726234f
C842 LADDEROUT.n16 VSS 0.582088f
C843 LADDEROUT.n17 VSS 1.10052f
C844 LADDEROUT.n18 VSS 0.514479f
C845 RSEL2.t1 VSS 0.600342f
C846 RSEL2.t5 VSS 0.585857f
C847 RSEL2.n0 VSS 2.65357f
C848 RSEL2.n1 VSS 0.08345f
C849 RSEL2.n2 VSS 1.60258f
C850 RSEL2.t0 VSS 0.705216f
C851 RSEL2.t4 VSS 0.724882f
C852 RSEL2.n3 VSS 2.64111f
C853 RSEL2.n4 VSS 1.7731f
C854 RSEL2.n5 VSS 4.64513f
C855 RSEL2.t2 VSS 0.033348f
C856 RSEL2.t6 VSS 0.019652f
C857 RSEL2.t3 VSS 0.033348f
C858 RSEL2.t7 VSS 0.019652f
C859 RSEL2.n6 VSS 0.055954f
C860 RSEL2.n7 VSS 0.082722f
C861 RSEL2.n8 VSS 0.082064f
C862 RSEL2.n9 VSS 1.32764f
C863 RSEL2.n10 VSS 0.236321f
C864 R3R4.t5 VSS 0.220874f
C865 R3R4.t4 VSS 0.180106f
C866 R3R4.n0 VSS 3.14849f
C867 R3R4.t7 VSS 0.639891f
C868 R3R4.t8 VSS 0.367349f
C869 R3R4.n1 VSS 3.55784f
C870 R3R4.t3 VSS 0.662294f
C871 R3R4.t2 VSS 0.468512f
C872 R3R4.n2 VSS 3.63759f
C873 R3R4.n3 VSS 0.575373f
C874 R3R4.n4 VSS 0.163342f
C875 R3R4.n5 VSS 7.10541f
C876 R3R4.n6 VSS 7.45015f
C877 R3R4.t1 VSS 0.639891f
C878 R3R4.t0 VSS 0.367349f
C879 R3R4.n7 VSS 3.55784f
C880 R3R4.t9 VSS 0.662294f
C881 R3R4.t6 VSS 0.468512f
C882 R3R4.n8 VSS 3.63759f
C883 R3R4.n9 VSS 0.575373f
C884 R3R4.n10 VSS 0.124925f
C885 x1.x3.GN1.n0 VSS 1.24311f
C886 x1.x3.GN1.t0 VSS 0.039083f
C887 x1.x3.GN1.n1 VSS 0.0451f
C888 x1.x3.GN1.t6 VSS 0.441683f
C889 x1.x3.GN1.t5 VSS 0.431027f
C890 x1.x3.GN1.n2 VSS 1.93385f
C891 x1.x3.GN1.t2 VSS 0.441683f
C892 x1.x3.GN1.t9 VSS 0.431027f
C893 x1.x3.GN1.n3 VSS 1.93385f
C894 x1.x3.GN1.n4 VSS 0.916253f
C895 x1.x3.GN1.n5 VSS 0.312185f
C896 x1.x3.GN1.t7 VSS 0.024535f
C897 x1.x3.GN1.t3 VSS 0.014458f
C898 x1.x3.GN1.t8 VSS 0.024535f
C899 x1.x3.GN1.t4 VSS 0.014458f
C900 x1.x3.GN1.n6 VSS 0.041166f
C901 x1.x3.GN1.n7 VSS 0.060803f
C902 x1.x3.GN1.n8 VSS 0.059138f
C903 x1.x3.GN1.n9 VSS 0.128451f
C904 x1.x3.GN1.t1 VSS 0.099816f
C905 x1.x3.GN1.n10 VSS 0.017954f
C906 x1.x3.GN1.n11 VSS 0.020113f
C907 VRES.t7 VSS 0.69694f
C908 VRES.t8 VSS 0.4001f
C909 VRES.n0 VSS 3.87503f
C910 VRES.t6 VSS 0.721341f
C911 VRES.t4 VSS 0.510282f
C912 VRES.n1 VSS 3.9619f
C913 VRES.n2 VSS 0.62667f
C914 VRES.n3 VSS 0.153943f
C915 VRES.t3 VSS 0.69694f
C916 VRES.t5 VSS 0.4001f
C917 VRES.n4 VSS 3.87503f
C918 VRES.t1 VSS 0.721341f
C919 VRES.t2 VSS 0.510282f
C920 VRES.n5 VSS 3.9619f
C921 VRES.n6 VSS 0.62667f
C922 VRES.n7 VSS 0.137231f
C923 VRES.t0 VSS 0.195773f
C924 VRES.n8 VSS 3.2661f
C925 VRES.n9 VSS 3.39104f
C926 R1R2.t1 VSS 0.210975f
C927 R1R2.t0 VSS 0.172971f
C928 R1R2.n0 VSS 3.23954f
C929 R1R2.t2 VSS 0.614544f
C930 R1R2.t3 VSS 0.352798f
C931 R1R2.n1 VSS 3.4169f
C932 R1R2.t4 VSS 0.63606f
C933 R1R2.t5 VSS 0.449953f
C934 R1R2.n2 VSS 3.4935f
C935 R1R2.n3 VSS 0.552582f
C936 R1R2.n4 VSS 0.118914f
C937 VDD.n0 VSS 0.057511f
C938 VDD.n1 VSS 0.255958f
C939 VDD.n2 VSS 0.12362f
C940 VDD.n3 VSS 1.04114f
C941 VDD.n4 VSS 1.04114f
C942 VDD.n5 VSS 0.171354f
C943 VDD.n6 VSS 0.125503f
C944 VDD.t84 VSS 1.38435f
C945 VDD.n9 VSS 0.125503f
C946 VDD.n10 VSS 5.32e-19
C947 VDD.n11 VSS 0.076211f
C948 VDD.n12 VSS 0.013857f
C949 VDD.n13 VSS 0.150654f
C950 VDD.n14 VSS 0.080552f
C951 VDD.n15 VSS 0.163575f
C952 VDD.n16 VSS 0.189769f
C953 VDD.n17 VSS 0.255958f
C954 VDD.n18 VSS 0.004156f
C955 VDD.n19 VSS 0.171354f
C956 VDD.n20 VSS 0.125503f
C957 VDD.t127 VSS 1.38435f
C958 VDD.n22 VSS 1.04114f
C959 VDD.n23 VSS 0.125503f
C960 VDD.n25 VSS 1.04114f
C961 VDD.n26 VSS 0.12362f
C962 VDD.n27 VSS 0.009949f
C963 VDD.n28 VSS 0.076135f
C964 VDD.n29 VSS 0.013984f
C965 VDD.n30 VSS 0.150654f
C966 VDD.n31 VSS 0.079915f
C967 VDD.n32 VSS 0.129517f
C968 VDD.n33 VSS 0.186042f
C969 VDD.n34 VSS 0.255958f
C970 VDD.n35 VSS 0.004409f
C971 VDD.n36 VSS 0.171354f
C972 VDD.n37 VSS 0.125503f
C973 VDD.t101 VSS 1.38435f
C974 VDD.n39 VSS 1.04114f
C975 VDD.n40 VSS 0.125503f
C976 VDD.n42 VSS 1.04114f
C977 VDD.n43 VSS 0.12362f
C978 VDD.n44 VSS 0.009966f
C979 VDD.n45 VSS 0.075882f
C980 VDD.n46 VSS 0.013984f
C981 VDD.n47 VSS 0.150654f
C982 VDD.n48 VSS 0.079915f
C983 VDD.n49 VSS 0.126263f
C984 VDD.n50 VSS 0.193623f
C985 VDD.n51 VSS 0.255958f
C986 VDD.n52 VSS 0.013612f
C987 VDD.n53 VSS 0.12362f
C988 VDD.n54 VSS 1.04114f
C989 VDD.n55 VSS 1.04114f
C990 VDD.n56 VSS 0.171354f
C991 VDD.n57 VSS 0.125503f
C992 VDD.t83 VSS 1.38435f
C993 VDD.n60 VSS 0.125503f
C994 VDD.n61 VSS 4.81e-19
C995 VDD.n62 VSS 0.076211f
C996 VDD.n63 VSS 0.013908f
C997 VDD.n64 VSS 0.150654f
C998 VDD.n65 VSS 0.080502f
C999 VDD.n66 VSS 0.371254f
C1000 VDD.n67 VSS 0.007798f
C1001 VDD.t124 VSS 0.015738f
C1002 VDD.n68 VSS 0.015481f
C1003 VDD.t50 VSS 0.00169f
C1004 VDD.t88 VSS 0.002567f
C1005 VDD.n69 VSS 0.004434f
C1006 VDD.t126 VSS 0.01604f
C1007 VDD.t52 VSS 0.015738f
C1008 VDD.n70 VSS 0.01499f
C1009 VDD.n71 VSS 0.007798f
C1010 VDD.n72 VSS 0.007059f
C1011 VDD.t39 VSS 0.002316f
C1012 VDD.n73 VSS 0.006573f
C1013 VDD.t116 VSS 0.009521f
C1014 VDD.n74 VSS 0.008764f
C1015 VDD.n75 VSS 0.007822f
C1016 VDD.t63 VSS 0.015742f
C1017 VDD.n76 VSS 0.001288f
C1018 VDD.t29 VSS 0.006749f
C1019 VDD.t19 VSS 0.011141f
C1020 VDD.n77 VSS 0.010984f
C1021 VDD.n78 VSS 0.013164f
C1022 VDD.t156 VSS 0.046497f
C1023 VDD.n79 VSS 0.042056f
C1024 VDD.t92 VSS 0.001261f
C1025 VDD.t122 VSS 0.003382f
C1026 VDD.n80 VSS 0.015436f
C1027 VDD.t20 VSS 0.011141f
C1028 VDD.n81 VSS 0.008152f
C1029 VDD.n82 VSS 0.030426f
C1030 VDD.n83 VSS 0.024039f
C1031 VDD.n84 VSS 0.031224f
C1032 VDD.n85 VSS 0.018029f
C1033 VDD.n86 VSS 0.013164f
C1034 VDD.n87 VSS 0.009873f
C1035 VDD.n88 VSS 0.006197f
C1036 VDD.n89 VSS 0.019524f
C1037 VDD.n90 VSS 0.030608f
C1038 VDD.t97 VSS 0.031636f
C1039 VDD.n91 VSS 0.002382f
C1040 VDD.n92 VSS 0.002432f
C1041 VDD.n93 VSS 0.009873f
C1042 VDD.n94 VSS 0.003041f
C1043 VDD.t151 VSS 0.015954f
C1044 VDD.n95 VSS 0.013093f
C1045 VDD.n96 VSS 0.007798f
C1046 VDD.t155 VSS 0.046497f
C1047 VDD.n97 VSS 0.01159f
C1048 VDD.n98 VSS 0.007798f
C1049 VDD.t37 VSS 0.001261f
C1050 VDD.t104 VSS 0.003382f
C1051 VDD.n99 VSS 0.015436f
C1052 VDD.t157 VSS 0.046497f
C1053 VDD.t114 VSS 0.006749f
C1054 VDD.n100 VSS 0.020842f
C1055 VDD.n101 VSS 0.011948f
C1056 VDD.n102 VSS 0.006197f
C1057 VDD.t13 VSS 0.011141f
C1058 VDD.n103 VSS 0.010984f
C1059 VDD.n104 VSS 0.042056f
C1060 VDD.n105 VSS 0.018029f
C1061 VDD.n106 VSS 0.031224f
C1062 VDD.t14 VSS 0.011141f
C1063 VDD.t129 VSS 0.015956f
C1064 VDD.n107 VSS 0.004507f
C1065 VDD.n108 VSS 0.005366f
C1066 VDD.t113 VSS 0.063694f
C1067 VDD.t103 VSS 0.061584f
C1068 VDD.t12 VSS 0.045556f
C1069 VDD.t36 VSS 0.065381f
C1070 VDD.t146 VSS 0.063694f
C1071 VDD.t24 VSS 0.072551f
C1072 VDD.t130 VSS 0.052726f
C1073 VDD.t53 VSS 0.028261f
C1074 VDD.t150 VSS 0.013076f
C1075 VDD.t128 VSS 0.045977f
C1076 VDD.n109 VSS 0.059997f
C1077 VDD.n110 VSS 0.041607f
C1078 VDD.n111 VSS 0.01223f
C1079 VDD.n112 VSS 0.019622f
C1080 VDD.n113 VSS 0.024039f
C1081 VDD.n114 VSS 0.008156f
C1082 VDD.n115 VSS 0.064967f
C1083 VDD.n116 VSS 0.088372f
C1084 VDD.t22 VSS 0.011141f
C1085 VDD.n117 VSS 0.021787f
C1086 VDD.n118 VSS 0.042056f
C1087 VDD.n119 VSS 0.025917f
C1088 VDD.t23 VSS 0.011141f
C1089 VDD.t79 VSS 0.016033f
C1090 VDD.n120 VSS 0.018733f
C1091 VDD.t21 VSS 0.143295f
C1092 VDD.t3 VSS 0.088033f
C1093 VDD.t45 VSS 0.036122f
C1094 VDD.t47 VSS 0.049997f
C1095 VDD.t105 VSS 0.036122f
C1096 VDD.t119 VSS 0.049997f
C1097 VDD.t81 VSS 0.036122f
C1098 VDD.t78 VSS 0.054065f
C1099 VDD.n121 VSS 0.059182f
C1100 VDD.n122 VSS 0.007798f
C1101 VDD.n123 VSS 0.003395f
C1102 VDD.t120 VSS 0.016033f
C1103 VDD.n124 VSS 0.003395f
C1104 VDD.t48 VSS 0.016033f
C1105 VDD.n125 VSS 0.22915f
C1106 VDD.n126 VSS 0.013412f
C1107 VDD.n127 VSS 0.008152f
C1108 VDD.t152 VSS 0.047225f
C1109 VDD.t4 VSS 0.011141f
C1110 VDD.n128 VSS 0.046752f
C1111 VDD.n129 VSS 0.023234f
C1112 VDD.t5 VSS 0.011141f
C1113 VDD.n130 VSS 0.030426f
C1114 VDD.n131 VSS 0.027983f
C1115 VDD.n132 VSS 0.017558f
C1116 VDD.n133 VSS 0.013702f
C1117 VDD.n134 VSS 0.013361f
C1118 VDD.t46 VSS 0.01604f
C1119 VDD.n135 VSS 0.020186f
C1120 VDD.n136 VSS 0.007798f
C1121 VDD.n137 VSS 0.013164f
C1122 VDD.n138 VSS 0.009873f
C1123 VDD.n139 VSS 0.018936f
C1124 VDD.t106 VSS 0.01604f
C1125 VDD.n140 VSS 0.02049f
C1126 VDD.n141 VSS 0.007798f
C1127 VDD.n142 VSS 0.013164f
C1128 VDD.n143 VSS 0.009873f
C1129 VDD.n144 VSS 0.018936f
C1130 VDD.t82 VSS 0.01604f
C1131 VDD.n145 VSS 0.02049f
C1132 VDD.n146 VSS 0.003395f
C1133 VDD.n147 VSS 0.013164f
C1134 VDD.n148 VSS 0.009873f
C1135 VDD.n149 VSS 0.005008f
C1136 VDD.n150 VSS 0.027358f
C1137 VDD.n151 VSS 0.01223f
C1138 VDD.n152 VSS 0.019622f
C1139 VDD.n153 VSS 0.033429f
C1140 VDD.n154 VSS 0.006654f
C1141 VDD.n155 VSS 0.06046f
C1142 VDD.n156 VSS 0.058625f
C1143 VDD.n157 VSS 0.001359f
C1144 VDD.t54 VSS 0.00169f
C1145 VDD.t131 VSS 0.002567f
C1146 VDD.n158 VSS 0.004434f
C1147 VDD.n159 VSS 0.02976f
C1148 VDD.t145 VSS 0.016033f
C1149 VDD.n160 VSS 0.018683f
C1150 VDD.t25 VSS 0.005282f
C1151 VDD.t98 VSS 0.014041f
C1152 VDD.n161 VSS 0.007965f
C1153 VDD.t147 VSS 0.015742f
C1154 VDD.n162 VSS 0.016608f
C1155 VDD.n163 VSS 0.021362f
C1156 VDD.n164 VSS 0.002813f
C1157 VDD.n165 VSS 0.013164f
C1158 VDD.n166 VSS 0.007798f
C1159 VDD.n167 VSS 0.004507f
C1160 VDD.n168 VSS 0.005008f
C1161 VDD.n169 VSS 0.026805f
C1162 VDD.n170 VSS 0.073092f
C1163 VDD.t49 VSS 0.01392f
C1164 VDD.t123 VSS 0.036276f
C1165 VDD.t125 VSS 0.040494f
C1166 VDD.t87 VSS 0.028261f
C1167 VDD.t38 VSS 0.052726f
C1168 VDD.t51 VSS 0.074239f
C1169 VDD.t62 VSS 0.036276f
C1170 VDD.t115 VSS 0.028261f
C1171 VDD.t91 VSS 0.065381f
C1172 VDD.t18 VSS 0.045556f
C1173 VDD.t121 VSS 0.061584f
C1174 VDD.t28 VSS 0.063694f
C1175 VDD.n171 VSS 0.043375f
C1176 VDD.n172 VSS 0.012601f
C1177 VDD.n173 VSS 0.00897f
C1178 VDD.n174 VSS 0.002382f
C1179 VDD.n175 VSS 0.017476f
C1180 VDD.n176 VSS 0.006665f
C1181 VDD.n177 VSS 0.013164f
C1182 VDD.n178 VSS 0.009873f
C1183 VDD.n179 VSS 0.005869f
C1184 VDD.n180 VSS 0.01995f
C1185 VDD.n181 VSS 0.014277f
C1186 VDD.n182 VSS 0.009086f
C1187 VDD.n183 VSS 0.025693f
C1188 VDD.n184 VSS 0.163422f
C1189 VDD.n185 VSS 0.083569f
C1190 VDD.n186 VSS 0.419546f
C1191 VDD.t80 VSS 0.00626f
C1192 VDD.t159 VSS 0.003689f
C1193 VDD.t77 VSS 0.00626f
C1194 VDD.t161 VSS 0.003689f
C1195 VDD.n187 VSS 0.010503f
C1196 VDD.n188 VSS 0.015528f
C1197 VDD.n189 VSS 0.015405f
C1198 VDD.n190 VSS 0.006296f
C1199 VDD.n191 VSS 0.93188f
C1200 VDD.n192 VSS 0.052382f
C1201 VDD.n193 VSS 0.078847f
C1202 VDD.n194 VSS 0.255947f
C1203 VDD.n195 VSS 0.124019f
C1204 VDD.n196 VSS 0.124019f
C1205 VDD.n197 VSS 0.123614f
C1206 VDD.n198 VSS 0.171372f
C1207 VDD.n199 VSS 0.552489f
C1208 VDD.t89 VSS 0.797375f
C1209 VDD.n200 VSS 0.769866f
C1210 VDD.t90 VSS 0.797375f
C1211 VDD.n201 VSS 0.552489f
C1212 VDD.n202 VSS 0.004857f
C1213 VDD.n203 VSS 0.135688f
C1214 VDD.n204 VSS 0.040676f
C1215 VDD.n205 VSS 0.139294f
C1216 VDD.n206 VSS 0.078847f
C1217 VDD.n207 VSS 0.255947f
C1218 VDD.n208 VSS 0.124019f
C1219 VDD.n209 VSS 0.124019f
C1220 VDD.n210 VSS 0.123614f
C1221 VDD.n211 VSS 0.171372f
C1222 VDD.n212 VSS 0.552489f
C1223 VDD.t74 VSS 0.797375f
C1224 VDD.n213 VSS 0.769866f
C1225 VDD.t55 VSS 0.797375f
C1226 VDD.n214 VSS 0.552489f
C1227 VDD.n215 VSS 0.004857f
C1228 VDD.n216 VSS 0.135688f
C1229 VDD.n217 VSS 0.040646f
C1230 VDD.n218 VSS 0.073399f
C1231 VDD.n219 VSS 0.39441f
C1232 VDD.n220 VSS 0.15613f
C1233 VDD.n221 VSS 0.255958f
C1234 VDD.n222 VSS 0.076211f
C1235 VDD.n223 VSS 1.04114f
C1236 VDD.n224 VSS 1.04114f
C1237 VDD.n225 VSS 0.12362f
C1238 VDD.n226 VSS 0.171354f
C1239 VDD.n227 VSS 0.125503f
C1240 VDD.t142 VSS 1.38435f
C1241 VDD.n230 VSS 0.125503f
C1242 VDD.n231 VSS 4.81e-19
C1243 VDD.n232 VSS 0.057511f
C1244 VDD.n233 VSS 0.255958f
C1245 VDD.n234 VSS 0.12362f
C1246 VDD.n235 VSS 1.04114f
C1247 VDD.n236 VSS 1.04114f
C1248 VDD.n237 VSS 0.171354f
C1249 VDD.n238 VSS 0.125503f
C1250 VDD.t33 VSS 1.38435f
C1251 VDD.n241 VSS 0.125503f
C1252 VDD.n242 VSS 5.32e-19
C1253 VDD.n243 VSS 0.076211f
C1254 VDD.n244 VSS 0.013857f
C1255 VDD.n245 VSS 0.150654f
C1256 VDD.n246 VSS 0.080552f
C1257 VDD.n247 VSS 0.163575f
C1258 VDD.n248 VSS 0.189769f
C1259 VDD.n249 VSS 0.255958f
C1260 VDD.n250 VSS 0.004156f
C1261 VDD.n251 VSS 0.171354f
C1262 VDD.n252 VSS 0.125503f
C1263 VDD.t134 VSS 1.38435f
C1264 VDD.n254 VSS 1.04114f
C1265 VDD.n255 VSS 0.125503f
C1266 VDD.n257 VSS 1.04114f
C1267 VDD.n258 VSS 0.12362f
C1268 VDD.n259 VSS 0.009949f
C1269 VDD.n260 VSS 0.076135f
C1270 VDD.n261 VSS 0.013984f
C1271 VDD.n262 VSS 0.150654f
C1272 VDD.n263 VSS 0.079915f
C1273 VDD.n264 VSS 0.129517f
C1274 VDD.n265 VSS 0.186042f
C1275 VDD.n266 VSS 0.255958f
C1276 VDD.n267 VSS 0.004409f
C1277 VDD.n268 VSS 0.171354f
C1278 VDD.n269 VSS 0.125503f
C1279 VDD.t35 VSS 1.38435f
C1280 VDD.n271 VSS 1.04114f
C1281 VDD.n272 VSS 0.125503f
C1282 VDD.n274 VSS 1.04114f
C1283 VDD.n275 VSS 0.12362f
C1284 VDD.n276 VSS 0.009966f
C1285 VDD.n277 VSS 0.075882f
C1286 VDD.n278 VSS 0.013984f
C1287 VDD.n279 VSS 0.150654f
C1288 VDD.n280 VSS 0.079915f
C1289 VDD.n281 VSS 0.127059f
C1290 VDD.n282 VSS 0.169406f
C1291 VDD.n283 VSS 0.013612f
C1292 VDD.n284 VSS 0.013908f
C1293 VDD.n285 VSS 0.150654f
C1294 VDD.n286 VSS 0.080502f
C1295 VDD.n287 VSS 0.144202f
C1296 VDD.n288 VSS 0.192732f
C1297 VDD.n289 VSS 0.255958f
C1298 VDD.n290 VSS 0.013648f
C1299 VDD.n291 VSS 0.12362f
C1300 VDD.n292 VSS 1.04114f
C1301 VDD.n293 VSS 1.04114f
C1302 VDD.n294 VSS 0.171354f
C1303 VDD.n295 VSS 0.125503f
C1304 VDD.t34 VSS 1.38435f
C1305 VDD.n298 VSS 0.125503f
C1306 VDD.n299 VSS 5.32e-19
C1307 VDD.n300 VSS 0.076211f
C1308 VDD.n301 VSS 0.013857f
C1309 VDD.n302 VSS 0.150654f
C1310 VDD.n303 VSS 0.080552f
C1311 VDD.n304 VSS 0.097945f
C1312 VDD.n305 VSS 0.237777f
C1313 VDD.n306 VSS 0.255958f
C1314 VDD.n307 VSS 0.004156f
C1315 VDD.n308 VSS 0.171354f
C1316 VDD.n309 VSS 0.125503f
C1317 VDD.t135 VSS 1.38435f
C1318 VDD.n311 VSS 1.04114f
C1319 VDD.n312 VSS 0.125503f
C1320 VDD.n314 VSS 1.04114f
C1321 VDD.n315 VSS 0.12362f
C1322 VDD.n316 VSS 0.009949f
C1323 VDD.n317 VSS 0.076135f
C1324 VDD.n318 VSS 0.013984f
C1325 VDD.n319 VSS 0.150654f
C1326 VDD.n320 VSS 0.079915f
C1327 VDD.n321 VSS 0.117449f
C1328 VDD.n322 VSS 0.19835f
C1329 VDD.n323 VSS 0.255958f
C1330 VDD.n324 VSS 0.004409f
C1331 VDD.n325 VSS 0.171354f
C1332 VDD.n326 VSS 0.125503f
C1333 VDD.t44 VSS 1.38435f
C1334 VDD.n328 VSS 1.04114f
C1335 VDD.n329 VSS 0.125503f
C1336 VDD.n331 VSS 1.04114f
C1337 VDD.n332 VSS 0.12362f
C1338 VDD.n333 VSS 0.010254f
C1339 VDD.n334 VSS 0.075882f
C1340 VDD.n335 VSS 0.013984f
C1341 VDD.n336 VSS 0.150654f
C1342 VDD.n337 VSS 0.079915f
C1343 VDD.n338 VSS 0.154767f
C1344 VDD.n339 VSS 0.255958f
C1345 VDD.n340 VSS 0.12362f
C1346 VDD.n341 VSS 1.04114f
C1347 VDD.n342 VSS 1.04114f
C1348 VDD.n343 VSS 0.171354f
C1349 VDD.n344 VSS 0.125503f
C1350 VDD.t32 VSS 1.38435f
C1351 VDD.n347 VSS 0.125503f
C1352 VDD.n348 VSS 4.81e-19
C1353 VDD.n349 VSS 0.076211f
C1354 VDD.n350 VSS 0.013908f
C1355 VDD.n351 VSS 0.150654f
C1356 VDD.n352 VSS 0.080502f
C1357 VDD.n353 VSS 0.153542f
C1358 VDD.n354 VSS 0.233268f
C1359 VDD.n355 VSS 1.83608f
C1360 VDD.n356 VSS 0.725969f
C1361 VDD.n357 VSS 0.217438f
C1362 VDD.n358 VSS 0.007798f
C1363 VDD.t65 VSS 0.015738f
C1364 VDD.n359 VSS 0.015481f
C1365 VDD.t59 VSS 0.00169f
C1366 VDD.t86 VSS 0.002567f
C1367 VDD.n360 VSS 0.004434f
C1368 VDD.t67 VSS 0.01604f
C1369 VDD.t27 VSS 0.015738f
C1370 VDD.n361 VSS 0.01499f
C1371 VDD.n362 VSS 0.007798f
C1372 VDD.n363 VSS 0.007059f
C1373 VDD.t69 VSS 0.002316f
C1374 VDD.n364 VSS 0.006573f
C1375 VDD.t41 VSS 0.009521f
C1376 VDD.n365 VSS 0.008764f
C1377 VDD.n366 VSS 0.007822f
C1378 VDD.t137 VSS 0.015742f
C1379 VDD.n367 VSS 0.001288f
C1380 VDD.t149 VSS 0.006749f
C1381 VDD.t16 VSS 0.011141f
C1382 VDD.n368 VSS 0.010984f
C1383 VDD.n369 VSS 0.013164f
C1384 VDD.t153 VSS 0.046497f
C1385 VDD.n370 VSS 0.042056f
C1386 VDD.t139 VSS 0.001261f
C1387 VDD.t110 VSS 0.003382f
C1388 VDD.n371 VSS 0.015436f
C1389 VDD.t17 VSS 0.011141f
C1390 VDD.n372 VSS 0.008152f
C1391 VDD.n373 VSS 0.030426f
C1392 VDD.n374 VSS 0.024039f
C1393 VDD.n375 VSS 0.031224f
C1394 VDD.n376 VSS 0.018029f
C1395 VDD.n377 VSS 0.013164f
C1396 VDD.n378 VSS 0.009873f
C1397 VDD.n379 VSS 0.006197f
C1398 VDD.n380 VSS 0.019524f
C1399 VDD.n381 VSS 0.030608f
C1400 VDD.t42 VSS 0.031636f
C1401 VDD.n382 VSS 0.002382f
C1402 VDD.n383 VSS 0.002432f
C1403 VDD.n384 VSS 0.009873f
C1404 VDD.n385 VSS 0.003041f
C1405 VDD.t108 VSS 0.015954f
C1406 VDD.n386 VSS 0.013093f
C1407 VDD.n387 VSS 0.007798f
C1408 VDD.t160 VSS 0.046497f
C1409 VDD.n388 VSS 0.01159f
C1410 VDD.n389 VSS 0.007798f
C1411 VDD.t57 VSS 0.001261f
C1412 VDD.t31 VSS 0.003382f
C1413 VDD.n390 VSS 0.015436f
C1414 VDD.t154 VSS 0.046497f
C1415 VDD.t112 VSS 0.006749f
C1416 VDD.n391 VSS 0.020842f
C1417 VDD.n392 VSS 0.011948f
C1418 VDD.n393 VSS 0.006197f
C1419 VDD.t10 VSS 0.011141f
C1420 VDD.n394 VSS 0.010984f
C1421 VDD.n395 VSS 0.042056f
C1422 VDD.n396 VSS 0.018029f
C1423 VDD.n397 VSS 0.031224f
C1424 VDD.t11 VSS 0.011141f
C1425 VDD.t61 VSS 0.015956f
C1426 VDD.n398 VSS 0.004507f
C1427 VDD.n399 VSS 0.005366f
C1428 VDD.t111 VSS 0.063694f
C1429 VDD.t30 VSS 0.061584f
C1430 VDD.t9 VSS 0.045556f
C1431 VDD.t56 VSS 0.065381f
C1432 VDD.t95 VSS 0.063694f
C1433 VDD.t93 VSS 0.072551f
C1434 VDD.t140 VSS 0.052726f
C1435 VDD.t99 VSS 0.028261f
C1436 VDD.t107 VSS 0.013076f
C1437 VDD.t60 VSS 0.045977f
C1438 VDD.n400 VSS 0.059997f
C1439 VDD.n401 VSS 0.041607f
C1440 VDD.n402 VSS 0.01223f
C1441 VDD.n403 VSS 0.019622f
C1442 VDD.n404 VSS 0.024039f
C1443 VDD.n405 VSS 0.008156f
C1444 VDD.n406 VSS 0.064967f
C1445 VDD.n407 VSS 0.088372f
C1446 VDD.t1 VSS 0.011141f
C1447 VDD.n408 VSS 0.021787f
C1448 VDD.n409 VSS 0.042056f
C1449 VDD.n410 VSS 0.025917f
C1450 VDD.t2 VSS 0.011141f
C1451 VDD.t73 VSS 0.016033f
C1452 VDD.n411 VSS 0.018733f
C1453 VDD.t0 VSS 0.143295f
C1454 VDD.t6 VSS 0.088033f
C1455 VDD.t75 VSS 0.036122f
C1456 VDD.t132 VSS 0.049997f
C1457 VDD.t117 VSS 0.036122f
C1458 VDD.t143 VSS 0.049997f
C1459 VDD.t70 VSS 0.036122f
C1460 VDD.t72 VSS 0.054065f
C1461 VDD.n412 VSS 0.059182f
C1462 VDD.n413 VSS 0.007798f
C1463 VDD.n414 VSS 0.003395f
C1464 VDD.t144 VSS 0.016033f
C1465 VDD.n415 VSS 0.003395f
C1466 VDD.t133 VSS 0.016033f
C1467 VDD.n416 VSS 0.22915f
C1468 VDD.n417 VSS 0.013412f
C1469 VDD.n418 VSS 0.008152f
C1470 VDD.t158 VSS 0.047225f
C1471 VDD.t7 VSS 0.011141f
C1472 VDD.n419 VSS 0.046752f
C1473 VDD.n420 VSS 0.023234f
C1474 VDD.t8 VSS 0.011141f
C1475 VDD.n421 VSS 0.030426f
C1476 VDD.n422 VSS 0.027983f
C1477 VDD.n423 VSS 0.017558f
C1478 VDD.n424 VSS 0.013702f
C1479 VDD.n425 VSS 0.013361f
C1480 VDD.t76 VSS 0.01604f
C1481 VDD.n426 VSS 0.020186f
C1482 VDD.n427 VSS 0.007798f
C1483 VDD.n428 VSS 0.013164f
C1484 VDD.n429 VSS 0.009873f
C1485 VDD.n430 VSS 0.018936f
C1486 VDD.t118 VSS 0.01604f
C1487 VDD.n431 VSS 0.02049f
C1488 VDD.n432 VSS 0.007798f
C1489 VDD.n433 VSS 0.013164f
C1490 VDD.n434 VSS 0.009873f
C1491 VDD.n435 VSS 0.018936f
C1492 VDD.t71 VSS 0.01604f
C1493 VDD.n436 VSS 0.02049f
C1494 VDD.n437 VSS 0.003395f
C1495 VDD.n438 VSS 0.013164f
C1496 VDD.n439 VSS 0.009873f
C1497 VDD.n440 VSS 0.005008f
C1498 VDD.n441 VSS 0.027358f
C1499 VDD.n442 VSS 0.01223f
C1500 VDD.n443 VSS 0.019622f
C1501 VDD.n444 VSS 0.033429f
C1502 VDD.n445 VSS 0.006654f
C1503 VDD.n446 VSS 0.06046f
C1504 VDD.n447 VSS 0.058625f
C1505 VDD.n448 VSS 0.001359f
C1506 VDD.t100 VSS 0.00169f
C1507 VDD.t141 VSS 0.002567f
C1508 VDD.n449 VSS 0.004434f
C1509 VDD.n450 VSS 0.02976f
C1510 VDD.t94 VSS 0.016033f
C1511 VDD.n451 VSS 0.018683f
C1512 VDD.t102 VSS 0.005282f
C1513 VDD.t43 VSS 0.014041f
C1514 VDD.n452 VSS 0.007965f
C1515 VDD.t96 VSS 0.015742f
C1516 VDD.n453 VSS 0.016608f
C1517 VDD.n454 VSS 0.021362f
C1518 VDD.n455 VSS 0.002813f
C1519 VDD.n456 VSS 0.013164f
C1520 VDD.n457 VSS 0.007798f
C1521 VDD.n458 VSS 0.004507f
C1522 VDD.n459 VSS 0.005008f
C1523 VDD.n460 VSS 0.026805f
C1524 VDD.n461 VSS 0.073092f
C1525 VDD.t58 VSS 0.01392f
C1526 VDD.t64 VSS 0.036276f
C1527 VDD.t66 VSS 0.040494f
C1528 VDD.t85 VSS 0.028261f
C1529 VDD.t68 VSS 0.052726f
C1530 VDD.t26 VSS 0.074239f
C1531 VDD.t136 VSS 0.036276f
C1532 VDD.t40 VSS 0.028261f
C1533 VDD.t138 VSS 0.065381f
C1534 VDD.t15 VSS 0.045556f
C1535 VDD.t109 VSS 0.061584f
C1536 VDD.t148 VSS 0.063694f
C1537 VDD.n462 VSS 0.043375f
C1538 VDD.n463 VSS 0.012601f
C1539 VDD.n464 VSS 0.00897f
C1540 VDD.n465 VSS 0.002382f
C1541 VDD.n466 VSS 0.017476f
C1542 VDD.n467 VSS 0.006665f
C1543 VDD.n468 VSS 0.013164f
C1544 VDD.n469 VSS 0.009873f
C1545 VDD.n470 VSS 0.005869f
C1546 VDD.n471 VSS 0.01995f
C1547 VDD.n472 VSS 0.014277f
C1548 VDD.n473 VSS 0.009086f
C1549 VDD.n474 VSS 0.025693f
C1550 VDD.n475 VSS 0.200475f
C1551 VDD.n476 VSS 0.144781f
C1552 VDD.n477 VSS 0.13208f
C1553 VDD.n478 VSS 0.20215f
C1554 R4R5.t0 VSS 0.616703f
C1555 R4R5.t1 VSS 0.354038f
C1556 R4R5.n0 VSS 3.42891f
C1557 R4R5.t2 VSS 0.638295f
C1558 R4R5.t3 VSS 0.451534f
C1559 R4R5.n1 VSS 3.50578f
C1560 R4R5.n2 VSS 0.554523f
C1561 R4R5.n3 VSS 0.121432f
C1562 R4R5.t4 VSS 0.21672f
C1563 R4R5.t5 VSS 0.173234f
C1564 R4R5.n4 VSS 3.53038f
C1565 R4R5.n5 VSS 0.592856f
C1566 x1.x5.A.n0 VSS 1.57218f
C1567 x1.x5.A.n1 VSS 1.43499f
C1568 x1.x5.A.n2 VSS 1.5115f
C1569 x1.x5.A.n3 VSS 1.43499f
C1570 x1.x5.A.n4 VSS 1.54012f
C1571 x1.x5.A.n5 VSS 1.43499f
C1572 x1.x5.A.n6 VSS 1.51409f
C1573 x1.x5.A.n7 VSS 1.43499f
C1574 x1.x5.A.n8 VSS 0.662824f
C1575 x1.x5.A.t15 VSS 0.423279f
C1576 x1.x5.A.t14 VSS 0.422273f
C1577 x1.x5.A.t17 VSS 0.560366f
C1578 x1.x5.A.n9 VSS 2.95839f
C1579 x1.x5.A.t18 VSS 0.545349f
C1580 x1.x5.A.n10 VSS 0.664947f
C1581 x1.x5.A.t1 VSS 0.423279f
C1582 x1.x5.A.t2 VSS 0.422273f
C1583 x1.x5.A.t4 VSS 0.560366f
C1584 x1.x5.A.n11 VSS 2.95839f
C1585 x1.x5.A.t3 VSS 0.545349f
C1586 x1.x5.A.n12 VSS 0.410129f
C1587 x1.x5.A.t19 VSS 0.423279f
C1588 x1.x5.A.t5 VSS 0.422273f
C1589 x1.x5.A.t16 VSS 0.560366f
C1590 x1.x5.A.n13 VSS 2.95839f
C1591 x1.x5.A.t0 VSS 0.545349f
C1592 x1.x5.A.n14 VSS 0.698266f
C1593 x1.x5.A.t7 VSS 0.783638f
C1594 x1.x5.A.t11 VSS 0.554351f
C1595 x1.x5.A.n15 VSS 4.29789f
C1596 x1.x5.A.t12 VSS 0.75713f
C1597 x1.x5.A.t13 VSS 0.434654f
C1598 x1.x5.A.n16 VSS 4.216f
C1599 x1.x5.A.n17 VSS 0.680647f
C1600 x1.x5.A.t6 VSS 0.545349f
C1601 x1.x5.A.t9 VSS 0.422273f
C1602 x1.x5.A.t10 VSS 0.560366f
C1603 x1.x5.A.n18 VSS 2.95839f
C1604 x1.x5.A.t8 VSS 0.423279f
C1605 x1.x3.GP4.n0 VSS 0.102848f
C1606 x1.x3.x4.GP VSS 2.92223f
C1607 x1.x2.x4.GP VSS 2.2958f
C1608 x1.x1.gpo3 VSS 1.43068f
C1609 x1.x3.GP4.t2 VSS 0.01297f
C1610 x1.x3.GP4.t1 VSS 0.01297f
C1611 x1.x3.GP4.n1 VSS 0.030927f
C1612 x1.x1.x14.Y VSS 0.112099f
C1613 x1.x3.GP4.t5 VSS 0.656397f
C1614 x1.x3.GP4.t7 VSS 0.674701f
C1615 x1.x3.GP4.n2 VSS 2.39862f
C1616 x1.x3.GP4.t4 VSS 0.656397f
C1617 x1.x3.GP4.t6 VSS 0.674701f
C1618 x1.x3.GP4.n3 VSS 2.39862f
C1619 x1.x3.GP4.n4 VSS 2.81741f
C1620 x1.x3.GP4.n5 VSS 0.018905f
C1621 x1.x3.GP4.t0 VSS 0.019954f
C1622 x1.x3.GP4.t3 VSS 0.019954f
C1623 x1.x3.GP4.n6 VSS 0.043823f
C1624 R6R7.t5 VSS 0.938755f
C1625 R6R7.t1 VSS 0.191596f
C1626 R6R7.n0 VSS 2.90697f
C1627 R6R7.t2 VSS 0.681991f
C1628 R6R7.t3 VSS 0.391518f
C1629 R6R7.n1 VSS 3.79192f
C1630 R6R7.t0 VSS 0.705869f
C1631 R6R7.t4 VSS 0.499337f
C1632 R6R7.n2 VSS 3.87692f
C1633 R6R7.n3 VSS 0.613229f
C1634 R6R7.n4 VSS 0.131466f
C1635 R7R8.t9 VSS 0.56478f
C1636 R7R8.t2 VSS 0.32423f
C1637 R7R8.n0 VSS 3.14022f
C1638 R7R8.t1 VSS 0.584554f
C1639 R7R8.t8 VSS 0.413518f
C1640 R7R8.n1 VSS 3.21061f
C1641 R7R8.n2 VSS 0.507836f
C1642 R7R8.n3 VSS 0.110262f
C1643 R7R8.t6 VSS 0.188087f
C1644 R7R8.t3 VSS 0.161416f
C1645 R7R8.n4 VSS 2.28338f
C1646 R7R8.t0 VSS 0.56478f
C1647 R7R8.t5 VSS 0.32423f
C1648 R7R8.n5 VSS 3.14022f
C1649 R7R8.t4 VSS 0.584554f
C1650 R7R8.t7 VSS 0.413518f
C1651 R7R8.n6 VSS 3.21061f
C1652 R7R8.n7 VSS 0.507836f
C1653 R7R8.n8 VSS 0.111208f
C1654 R7R8.n9 VSS 9.70155f
C1655 R7R8.n10 VSS 0.945745f
.ends

