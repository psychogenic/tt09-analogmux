** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sch
.subckt passgatex4 A1 GN1 GP1 Z1 A2 GN2 GP2 Z2 A3 GN3 GP3 Z3 A4 GN4 GP4 Z4 VDD VSS
*.PININFO VDD:I VSS:I GP1:I GN1:I A1:B Z1:B GP2:I GN2:I A2:B Z2:B GP3:I GN3:I A3:B Z3:B GP4:I GN4:I A4:B Z4:B
x1 A1 GN1 GP1 Z1 VDD VSS passgate
x2 A2 GN2 GP2 Z2 VDD VSS passgate
x3 A3 GN3 GP3 Z3 VDD VSS passgate
x4 A4 GN4 GP4 Z4 VDD VSS passgate
.ends

* expanding   symbol:  passgate.sym # of pins=6
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sch
.subckt passgate A GN GP Z VDD VSS
*.PININFO GN:I VDD:I VSS:I GP:I A:B Z:B
XM1 Z GN A VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 m=2
XM3 Z GP A VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=2
.ends

.end
