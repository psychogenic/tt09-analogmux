** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sch
.subckt tt_um_patdeegan_anamux ena clk rst_n ua[4] ua[5] ua[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ua[0] ua[1] ua[2] ua[3] VSS VDD
*.PININFO ena:I clk:I rst_n:I ua[4]:B ua[5]:B ua[6]:B ui_in[7]:I uio_in[0]:I uio_in[1]:I uio_in[2]:I uio_in[3]:I uio_in[4]:I
*+ uio_in[5]:I uio_in[6]:I uio_in[7]:I uio_oe[0]:O uio_oe[1]:O uio_oe[2]:O uio_oe[3]:O uio_oe[4]:O uio_oe[5]:O uio_oe[6]:O uio_oe[7]:O
*+ uio_out[0]:B uio_out[1]:B uio_out[2]:B uio_out[3]:B uio_out[4]:B uio_out[5]:B uio_out[6]:B uio_out[7]:B uo_out[0]:O uo_out[1]:O uo_out[2]:O
*+ uo_out[3]:O uo_out[4]:O uo_out[5]:O uo_out[6]:O uo_out[7]:O ui_in[0]:I ui_in[1]:I ui_in[2]:I ui_in[3]:I ui_in[4]:I ui_in[5]:I ui_in[6]:I
*+ ua[0]:B ua[1]:B ua[2]:B ua[3]:B VSS:I VDD:I
x1 ua[0] ui_in[3] VDD ui_in[4] ua[1] VSS ui_in[0] ui_in[1] ua[2] ui_in[2] ua[3] ui_in[6] ui_in[5] fulltest_userarea
.ends

* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sym # of pins=13
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sch
.subckt fulltest_userarea VRES select0 VDD select1 ring_out VSS rsel0 rsel1 muxtest_out rsel2 ladderout enable_ring
+ enable_counter
*.PININFO VDD:I VSS:I select0:I select1:I rsel0:I rsel1:I rsel2:I enable_ring:I enable_counter:I ring_out:O muxtest_out:O
*+ ladderout:O VRES:I
x1 VDD VSS VRES select0 select1 rsel0 rsel1 rsel2 muxtest_out ladderout muxtest
x2 select0 VDD select1 VSS ring_out enable_ring enable_counter ringtest
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sym # of pins=10
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sch
.subckt muxtest VDD VSS VRES SELECT0 SELECT1 RSEL0 RSEL1 RSEL2 OUT LADDEROUT
*.PININFO VSS:I VDD:I SELECT0:I SELECT1:I VRES:I RSEL0:I RSEL1:I RSEL2:I OUT:O LADDEROUT:O
x1 VDD VSS RSEL0 RSEL1 A1 A5 A6 A2 A7 A3 RSEL2 VRES A4 LADDEROUT mux8onehot
x2 SELECT1 VDD VSS A5 VRES LADDEROUT OUT OUT OUT A1 OUT SELECT0 VDD net1 mux4onehot_b
XR1 A7 VRES VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR2 A6 A7 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR3 A5 A6 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR4 A4 A5 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR5 A3 A4 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR6 A2 A3 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR7 A1 A2 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR8 VSS A1 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sym # of pins=7
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sch
.subckt ringtest select0 VDD select1 VSS mux_out enable_ring enable_counter
*.PININFO VDD:I VSS:I enable_ring:I select0:I select1:I enable_counter:I mux_out:O
x3 select1 VDD VSS counter3 drv_out ring_out mux_out mux_out mux_out counter7 mux_out select0 VDD net1 mux4onehot_b
x4 enable_counter drv_out net2 net3 net4 counter3 net5 net6 net7 counter7 net8 net9 VDD VSS simplecounter
x1 VDD VSS enable_ring ring_out ring
x2 VDD VSS ring_out drv_out driver
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sch
.subckt mux8onehot VDD VSS select0 select1 A1 A5 A6 A2 A7 A3 select2 A8 A4 Z
*.PININFO select0:I select1:I select2:I VDD:I VSS:I Z:B A1:B A2:B A3:B A4:B A5:B A6:B A7:B A8:B
x4 Z OUT_HIGH nSEL2 select2 VSS VDD passgate
x5 Z OUT_LOW select2 nSEL2 VSS VDD passgate
x2 gpo2 gpo1 gpo0 VDD gpo3 VSS A3 A2 A1 OUT_LOW OUT_LOW OUT_LOW A4 OUT_LOW gno2 gno1 gno0 gno3 passgatex4
x1 gpo0 gno0 gno1 gpo1 select0 select1 gno2 gpo2 nSEL2 select2 gno3 gpo3 VDD VSS passgatesCtrlManual
x3 gpo2 gpo1 gpo0 VDD gpo3 VSS A7 A6 A5 OUT_HIGH OUT_HIGH OUT_HIGH A8 OUT_HIGH gno2 gno1 gno0 gno3 passgatex4
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sch
.subckt mux4onehot_b select1 VDD VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 select0 select2 nselect2
*.PININFO select0:I select1:I select2:I A1:B A2:B A3:B A4:B Z1:B Z2:B Z3:B Z4:B nselect2:O VDD:I VSS:I
x2 gpo2 gpo1 gpo0 VDD gpo3 VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 gno2 gno1 gno0 gno3 passgatex4
x1 gpo0 gno0 gno1 gpo1 select0 select1 gno2 gpo2 nselect2 select2 gno3 gpo3 VDD VSS passgatesCtrlManual
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/ring.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/ring.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/ring.sch
.subckt ring VDD VSS enable out
*.PININFO VDD:B enable:I VSS:B out:O
x2 enable net18 VSS VSS VDD VDD out sky130_fd_sc_hd__nand2_2
x1 VDD VSS out net1 inverter
x3 VDD VSS net1 net2 inverter
x4 VDD VSS net2 net3 inverter
x5 VDD VSS net3 net4 inverter
x6 VDD VSS net4 net5 inverter
x7 VDD VSS net5 net6 inverter
x8 VDD VSS net6 net7 inverter
x9 VDD VSS net7 net8 inverter
x10 VDD VSS net8 net9 inverter
x11 VDD VSS net9 net10 inverter
x12 VDD VSS net10 net11 inverter
x13 VDD VSS net11 net12 inverter
x14 VDD VSS net12 net13 inverter
x15 VDD VSS net13 net14 inverter
x16 VDD VSS net14 net15 inverter
x17 VDD VSS net15 net16 inverter
x18 VDD VSS net16 net17 inverter
x19 VDD VSS net17 net18 inverter
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/driver.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/driver.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/driver.sch
.subckt driver VDD VSS in out
*.PININFO VDD:B VSS:B out:O in:I
XM9 net1 in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM10 net1 in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
XM11 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=72 nf=8 m=1
XM12 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=24 nf=8 m=1
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym # of pins=6
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sch
.subckt passgate Z A GP GN VSSBPIN VCCBPIN
*.PININFO GN:I VCCBPIN:I VSSBPIN:I GP:I A:B Z:B
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 m=2
XM3 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=2
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym # of pins=18
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sch
.subckt passgatex4 GP3 GP2 GP1 VDD GP4 VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 GN3 GN2 GN1 GN4
*.PININFO VDD:I VSS:I GP1:I GN1:I A1:B Z1:B GP2:I GN2:I A2:B Z2:B GP3:I GN3:I A3:B Z3:B GP4:I GN4:I A4:B Z4:B
x1 Z1 A1 GP1 GN1 VSS VDD passgate
x2 Z2 A2 GP2 GN2 VSS VDD passgate
x3 Z3 A3 GP3 GN3 VSS VDD passgate
x4 Z4 A4 GP4 GN4 VSS VDD passgate
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sch
.subckt passgatesCtrlManual gpo0 gno0 gno1 gpo1 SEL0 SEL1 gno2 gpo2 nSEL2 SEL2 gno3 gpo3 VDD VSS
*.PININFO SEL0:I SEL1:I SEL2:I gno0:O gpo0:O gno1:O gpo1:O gno2:O gpo2:O gno3:O gpo3:O nSEL2:O VDD:I VSS:I
x1 SEL0 VSS VSS VDD VDD nSEL0 sky130_fd_sc_hd__inv_2
x2 SEL1 VSS VSS VDD VDD nSEL1 sky130_fd_sc_hd__inv_2
x7 nSEL0 nSEL1 VSS VSS VDD VDD gno0 sky130_fd_sc_hd__and2_1
x10 SEL1 SEL0 VSS VSS VDD VDD gno3 sky130_fd_sc_hd__and2_1
x11 gno0 VSS VSS VDD VDD gpo0 sky130_fd_sc_hd__inv_2
x12 gno1 VSS VSS VDD VDD gpo1 sky130_fd_sc_hd__inv_2
x13 gno2 VSS VSS VDD VDD gpo2 sky130_fd_sc_hd__inv_2
x14 gno3 VSS VSS VDD VDD gpo3 sky130_fd_sc_hd__inv_2
x15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x16 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x17 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x8 SEL1 SEL0 VSS VSS VDD VDD gno1 sky130_fd_sc_hd__and2b_1
x9 SEL0 SEL1 VSS VSS VDD VDD gno2 sky130_fd_sc_hd__and2b_1
x18 SEL2 VSS VSS VDD VDD nSEL2 sky130_fd_sc_hd__inv_2
x19 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/inverter.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/inverter.sch
.subckt inverter VDD VSS in out
*.PININFO out:O VDD:B VSS:B in:I
x1 in VSS VSS VDD VDD out sky130_fd_sc_hd__inv_2
.ends

.end
