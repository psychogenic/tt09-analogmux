* NGSPICE file created from tt_um_patdeegan_anamux_parax.ext - technology: sky130A

.subckt tt_um_patdeegan_anamux_parax clk ena rst_n ua[4] ua[5] ua[6] ua[7] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ ui_in[5] ua[0] ua[3] ui_in[1] ua[1] ui_in[4] ui_in[2] ui_in[6] ui_in[0] ua[2] ui_in[3]
+ VGND VDPWR
X0 a_21007_3867# ringtest_0.x4.net2.t2 VGND.t926 VGND.t925 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X1 VGND.t899 VDPWR.t1166 VGND.t898 VGND.t897 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X2 VGND.t901 VDPWR.t1167 VGND.t900 VGND.t671 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X3 a_24527_5340# a_24361_5340# VGND.t165 VGND.t164 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X4 ua[2].t3 muxtest_0.x2.x2.GP1.t4 ua[3].t4 VDPWR.t314 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X5 ringtest_0.x4.clknet_0_clk.t15 a_23879_6940# VGND.t642 VGND.t641 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X6 a_24135_3867# ringtest_0.x4.net6.t2 VDPWR.t160 VDPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X7 VGND.t1093 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t15 VGND.t1092 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X8 VDPWR.t1046 ui_in[1].t0 muxtest_0.x1.x1.nSEL1 VDPWR.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X9 a_22399_8976# a_21852_8720# a_22052_8875# VDPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=2310,139
X10 muxtest_0.x1.x3.GP1.t3 muxtest_0.x1.x3.GN1 VDPWR.t73 VDPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X11 a_27491_4566# ringtest_0.x4._23_ ringtest_0.x4._09_ VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=3510,184
X12 VGND.t550 a_27065_5156# a_27233_5058# VGND.t549 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X13 VDPWR.t1135 ringtest_0.x4._05_ a_24883_6800# VDPWR.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=4368,272
X14 VDPWR.t1039 a_16579_11759# ringtest_0.x3.x2.GN3 VDPWR.t1038 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X15 VDPWR.t754 VGND.t1127 VDPWR.t753 VDPWR.t752 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X16 a_25309_5334# a_24527_5340# a_25225_5334# VDPWR.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X17 a_12019_24012# muxtest_0.x2.x1.nSEL1 VGND.t548 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X18 a_26913_4566# ringtest_0.x4._15_ a_26817_4566# VGND.t575 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4160,194
X19 VGND.t579 ringtest_0.x4._21_ a_24545_5878# VGND.t578 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X20 muxtest_0.x1.x3.GP4.t3 muxtest_0.x1.x3.GN4 VDPWR.t1011 VDPWR.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X21 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR.t77 VDPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X22 VDPWR.t361 ringtest_0.x4._15_ a_25925_6788# VDPWR.t360 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X23 a_24004_6128# ringtest_0.x4._17_ a_23932_6128# VDPWR.t1143 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6600,266
X24 VGND.t904 VDPWR.t1168 VGND.t903 VGND.t902 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X25 a_23467_4818# ringtest_0.x4._11_.t4 a_23381_4818# VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X26 a_19114_31955# a_19290_32287# a_19242_32347# VGND.t967 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X27 VGND.t906 VDPWR.t1169 VGND.t905 VGND.t85 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X28 ringtest_0.x4.clknet_1_1__leaf_clk.t14 a_25364_5878# VGND.t1091 VGND.t1090 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X29 VDPWR.t963 a_21375_3867# ringtest_0.x4.counter[1] VDPWR.t962 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X30 VDPWR.t129 ringtest_0.x4.net5 a_22486_4246# VDPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=11200,512
X31 muxtest_0.x1.x1.nSEL0 ui_in[0].t0 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X32 VDPWR.t849 a_19842_32287# a_19666_31955# VDPWR.t848 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X33 muxtest_0.R3R4.t9 muxtest_0.x2.x2.GN3 ua[2].t11 VGND.t947 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X34 VDPWR.t751 VGND.t1128 VDPWR.t750 VDPWR.t749 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X35 a_12473_23980# ui_in[4].t0 VDPWR.t789 VDPWR.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X36 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP3 muxtest_0.R1R2.t1 VDPWR.t123 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X37 a_16579_11759# a_16755_12091# a_16707_12151# VGND.t929 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X38 VDPWR.t5 a_13501_23906# muxtest_0.x2.x2.GN4 VDPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X39 VDPWR.t219 a_19289_13081.t2 ringtest_0.drv_out.t18 VDPWR.t218 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X40 VGND.t5 a_21465_9294# ringtest_0.x4.net2.t0 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X41 ringtest_0.x4.clknet_0_clk.t31 a_23879_6940# VDPWR.t425 VDPWR.t424 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X42 VDPWR.t249 a_22021_4220# ringtest_0.x4._03_ VDPWR.t248 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=7430,283
X43 VGND.t304 ringtest_0.x4.net5 a_23467_4584# VGND.t303 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X44 muxtest_0.x2.nselect2 VDPWR.t951 VDPWR.t953 VDPWR.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X45 a_16707_12151# ui_in[4].t1 VGND.t114 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X46 VGND.t909 VDPWR.t1170 VGND.t908 VGND.t907 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X47 VDPWR.t748 VGND.t1129 VDPWR.t747 VDPWR.t613 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X48 ringtest_0.x4._15_ a_23381_4584# VGND.t829 VGND.t828 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X49 a_23899_5334# ringtest_0.x4._15_ VDPWR.t359 VDPWR.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0 ps=0 w=1 l=0.15
**devattr s=6900,269 d=6400,264
X50 VDPWR.t330 a_27065_5156# a_27233_5058# VDPWR.t320 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X51 muxtest_0.x1.x3.GP3 muxtest_0.x1.x3.GN3 VDPWR.t852 VDPWR.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X52 VGND.t912 VDPWR.t1171 VGND.t911 VGND.t910 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X53 VGND.t993 ringtest_0.x4.net3.t2 ringtest_0.x4._12_ VGND.t992 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X54 VGND.t11 a_25975_3867# ringtest_0.x4.counter[6] VGND.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X55 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk.t32 VDPWR.t1159 VDPWR.t1158 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X56 muxtest_0.x1.x5.A ui_in[2].t0 ua[3].t8 VDPWR.t772 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X57 ua[1].t1 ringtest_0.x3.x2.GP4.t4 ringtest_0.counter7.t1 VDPWR.t1094 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X58 a_22392_5990# a_22224_6244# VDPWR.t921 VDPWR.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0 ps=0 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X59 ringtest_0.x4.clknet_1_0__leaf_clk.t31 a_21395_6940# VDPWR.t1086 VDPWR.t1085 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X60 VGND.t1017 ringtest_0.x4._22_ a_26913_4566# VGND.t1016 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.104 ps=0.97 w=0.65 l=0.15
**devattr s=4160,194 d=4485,199
X61 a_26640_5334# a_26367_5340# a_26555_5334# VDPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X62 ringtest_0.x4.clknet_1_1__leaf_clk.t31 a_25364_5878# VDPWR.t1131 VDPWR.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X63 VDPWR.t746 VGND.t1130 VDPWR.t745 VDPWR.t744 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X64 VGND.t39 VDPWR.t1172 VGND.t38 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X65 a_21785_8054# ringtest_0.x4.net3.t3 VDPWR.t1018 VDPWR.t1017 sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X66 ringtest_0.x4._17_ a_25925_6788# VGND.t479 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X67 VGND.t359 a_19114_31955# muxtest_0.x1.x3.GN2 VGND.t358 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X68 VDPWR.t183 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR.t182 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X69 VDPWR.t950 VDPWR.t948 ringtest_0.x3.nselect2 VDPWR.t949 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X70 VDPWR.t423 a_23879_6940# ringtest_0.x4.clknet_0_clk.t30 VDPWR.t422 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X71 VGND.t856 ringtest_0.x4.net4 ringtest_0.x4._13_ VGND.t855 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X72 a_24317_4942# ringtest_0.x4.net6.t3 a_24551_4790# VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=4368,272
X73 VGND.t723 ringtest_0.x4.clknet_0_clk.t32 a_25364_5878# VGND.t722 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X74 VGND.t127 a_22111_10993# ringtest_0.x4.net1 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X75 VGND.t42 VDPWR.t1173 VGND.t41 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X76 VDPWR.t141 a_27815_3867# ringtest_0.x4.counter[8] VDPWR.t140 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X77 ringtest_0.x4._00_ a_21425_9686# a_21675_9686# VDPWR.t857 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X78 VDPWR.t743 VGND.t1131 VDPWR.t742 VDPWR.t602 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X79 VDPWR.t741 VGND.t1132 VDPWR.t740 VDPWR.t739 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X80 VDPWR.t841 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR.t840 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X81 VDPWR.t175 ringtest_0.x4._00_ a_22399_9142# VDPWR.t174 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=4368,272
X82 VGND.t640 a_23879_6940# ringtest_0.x4.clknet_0_clk.t14 VGND.t639 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X83 a_21675_4790# a_21509_4790# VGND.t557 VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X84 VGND.t1055 ui_in[0].t1 a_19842_32287# VGND.t1054 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X85 VGND.t45 VDPWR.t1174 VGND.t44 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X86 VDPWR.t1084 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t30 VDPWR.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X87 VGND.t136 a_23399_3867# ringtest_0.counter3.t2 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X88 VDPWR.t286 a_18662_32213# muxtest_0.x1.x3.GN1 VDPWR.t285 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X89 VDPWR.t941 ringtest_0.x4.net2.t3 a_21507_9686# VDPWR.t940 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X90 VDPWR.t738 VGND.t1133 VDPWR.t737 VDPWR.t736 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X91 a_27659_4246# ringtest_0.x4.net11 VDPWR.t809 VDPWR.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X92 a_22390_4566# ringtest_0.x4.net5 VGND.t302 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6890,366
X93 ringtest_0.x3.x1.nSEL1 ui_in[4].t2 VGND.t116 VGND.t115 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X94 ringtest_0.x4.clknet_1_0__leaf_clk.t15 a_21395_6940# VGND.t1051 VGND.t1050 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X95 a_22649_6244# a_21785_5878# a_22392_5990# VDPWR.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X96 muxtest_0.x1.x3.GP2.t3 muxtest_0.x1.x3.GN2 VDPWR.t179 VDPWR.t178 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X97 ua[3].t9 ui_in[2].t1 muxtest_0.x1.x4.A VGND.t662 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X98 muxtest_0.R5R6.t5 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A VGND.t838 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X99 VGND.t965 a_24329_6640# a_24336_6544# VGND.t964 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X100 a_27303_4246# a_27273_4220# ringtest_0.x4._09_ VDPWR.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.3 ps=2.6 w=1 l=0.15
**devattr s=12000,520 d=10400,504
X101 VDPWR.t735 VGND.t1134 VDPWR.t734 VDPWR.t733 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X102 ringtest_0.x4.clknet_1_0__leaf_clk.t29 a_21395_6940# VDPWR.t1082 VDPWR.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X103 VGND.t924 ringtest_0.x4.net2.t4 a_21425_9686# VGND.t923 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X104 a_19666_31955# a_19842_32287# a_19794_32347# VGND.t830 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X105 muxtest_0.R3R4.t1 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A VGND.t155 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X106 VDPWR.t885 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR.t884 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X107 a_21845_8816# ringtest_0.x4.clknet_1_0__leaf_clk.t32 VDPWR.t1014 VDPWR.t1013 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X108 VGND.t1049 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t14 VGND.t1048 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X109 a_21672_5334# a_21399_5340# a_21587_5334# VDPWR.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X110 ringtest_0.x4.clknet_1_1__leaf_clk.t30 a_25364_5878# VDPWR.t1129 VDPWR.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X111 VDPWR.t732 VGND.t1135 VDPWR.t731 VDPWR.t730 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X112 a_18662_32213# muxtest_0.x1.x1.nSEL0 a_18836_32319# VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X113 a_16203_12091# ui_in[4].t3 VDPWR.t113 VDPWR.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X114 a_19794_32347# ui_in[1].t1 VGND.t752 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X115 VDPWR.t729 VGND.t1136 VDPWR.t728 VDPWR.t727 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X116 VDPWR.t813 a_22817_6146# a_22733_6244# VDPWR.t812 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X117 VDPWR.t207 a_17231_12017# ringtest_0.x3.x2.GN4 VDPWR.t206 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X118 VDPWR.t421 a_23879_6940# ringtest_0.x4.clknet_0_clk.t29 VDPWR.t420 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X119 VGND.t1089 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t13 VGND.t1088 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X120 ringtest_0.x3.nselect2 VDPWR.t945 VDPWR.t947 VDPWR.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X121 a_25925_6788# ringtest_0.x4.net6.t4 VDPWR.t162 VDPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X122 a_25975_3867# ringtest_0.x4.net8 VDPWR.t802 VDPWR.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X123 ringtest_0.x4.net10 a_27233_5308# VDPWR.t832 VDPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X124 a_11845_23906# muxtest_0.x2.x1.nSEL1 VDPWR.t329 VDPWR.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X125 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VGND.t514 VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X126 VDPWR.t276 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR.t275 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X127 a_21939_8054# ringtest_0.x4.net3.t4 a_21867_8054# VGND.t994 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X128 a_26721_4246# ringtest_0.x4.net10 a_26627_4246# VDPWR.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.32 ps=2.64 w=1 l=0.15
**devattr s=12800,528 d=6600,266
X129 a_22116_4902# a_21948_5156# VGND.t847 VGND.t846 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X130 VDPWR.t1080 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t28 VDPWR.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X131 a_25149_4220# ringtest_0.x4.net7 VDPWR.t228 VDPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0 ps=0 w=0.42 l=0.15
**devattr s=3108,158 d=2940,154
X132 VDPWR.t891 a_21840_5308# a_21767_5334# VDPWR.t890 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X133 VGND.t48 VDPWR.t1175 VGND.t47 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X134 VGND.t51 VDPWR.t1176 VGND.t50 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X135 VDPWR.t173 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR.t172 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X136 VDPWR.t726 VGND.t1137 VDPWR.t725 VDPWR.t724 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X137 a_24627_6200# ringtest_0.x4._21_ VDPWR.t365 VDPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X138 VGND.t658 ringtest_0.x4._16_.t2 a_24986_5878# VGND.t657 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2646,147 d=3945,196
X139 VGND.t54 VDPWR.t1177 VGND.t53 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X140 VDPWR.t349 a_22245_8054# ringtest_0.x4._11_.t3 VDPWR.t348 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X141 a_25977_4220# ringtest_0.x4._11_.t5 VDPWR.t1041 VDPWR.t1040 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0 ps=0 w=0.42 l=0.15
**devattr s=3108,158 d=2940,154
X142 VGND.t57 VDPWR.t1178 VGND.t56 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X143 a_26367_4790# a_26201_4790# VGND.t321 VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X144 VDPWR.t723 VGND.t1138 VDPWR.t722 VDPWR.t624 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X145 a_25677_5156# a_24895_4790# a_25593_5156# VDPWR.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X146 VDPWR.t1142 ringtest_0.x4._17_ a_23349_6422# VDPWR.t1141 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X147 VDPWR.t357 ringtest_0.x4._15_ a_25977_4220# VDPWR.t356 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=3108,158
X148 VDPWR.t721 VGND.t1139 VDPWR.t720 VDPWR.t498 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X149 VDPWR.t187 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2.t3 VDPWR.t186 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X150 VDPWR.t309 a_24070_5852# a_24004_6128# VDPWR.t308 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=12000,520
X151 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP2.t4 muxtest_0.R6R7.t1 VDPWR.t13 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X152 ua[0].t1 muxtest_0.x2.x2.GN2 ua[2].t1 VGND.t357 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X153 VGND.t587 a_25977_4220# ringtest_0.x4._23_ VGND.t586 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=7851,266
X154 VDPWR.t719 VGND.t1140 VDPWR.t718 VDPWR.t717 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X155 VDPWR.t716 VGND.t1141 VDPWR.t715 VDPWR.t714 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X156 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X157 VDPWR.t87 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X158 a_21425_9686# ringtest_0.x4.net1 VGND.t134 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X159 VGND.t721 a_24317_4942# ringtest_0.x4._20_ VGND.t720 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=5266,228
X160 muxtest_0.x1.x1.nSEL1 ui_in[1].t2 VDPWR.t815 VDPWR.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X161 a_21465_8830# a_21561_8830# VGND.t970 VGND.t881 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X162 ringtest_0.x4.clknet_0_clk.t13 a_23879_6940# VGND.t638 VGND.t637 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X163 a_22295_3867# ringtest_0.x4.net4 VDPWR.t875 VDPWR.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X164 muxtest_0.R7R8.t9 muxtest_0.R6R7.t5 VGND.t643 sky130_fd_pr__res_high_po_1p41 l=1.75
X165 VDPWR.t713 VGND.t1142 VDPWR.t712 VDPWR.t711 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X166 a_26808_4902# a_26640_5156# VDPWR.t199 VDPWR.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0 ps=0 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X167 VGND.t60 VDPWR.t1179 VGND.t59 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X168 ringtest_0.x4.clknet_1_1__leaf_clk.t29 a_25364_5878# VDPWR.t1127 VDPWR.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X169 VGND.t731 a_26808_5308# a_26766_5712# VGND.t730 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X170 a_25351_5712# a_24361_5340# a_25225_5334# VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X171 VGND.t1047 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t13 VGND.t1046 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X172 VGND.t63 VDPWR.t1180 VGND.t62 VGND.t61 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X173 muxtest_0.R7R8.t8 muxtest_0.x2.x2.GN4 ua[2].t13 VGND.t961 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X174 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VGND.t776 VGND.t503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X175 VGND.t66 VDPWR.t1181 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X176 a_21007_3867# ringtest_0.x4.net2.t5 VDPWR.t939 VDPWR.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X177 ringtest_0.x4.net4 a_22265_5308# VDPWR.t215 VDPWR.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X178 VDPWR.t895 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR.t894 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X179 VGND.t391 a_19289_13081.t3 ringtest_0.drv_out.t10 VGND.t390 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X180 a_22373_5156# a_21509_4790# a_22116_4902# VDPWR.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X181 VDPWR.t710 VGND.t1143 VDPWR.t709 VDPWR.t565 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X182 a_26895_3867# ringtest_0.x4.net9 VGND.t522 VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X183 a_27191_4790# a_26201_4790# a_27065_5156# VGND.t319 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X184 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR.t845 VDPWR.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X185 VDPWR.t708 VGND.t1144 VDPWR.t707 VDPWR.t489 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X186 VGND.t69 VDPWR.t1182 VGND.t68 VGND.t67 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X187 a_22116_4902# a_21948_5156# VDPWR.t863 VDPWR.t862 sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0 ps=0 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X188 VGND.t738 ringtest_0.x4.net8 a_23837_5878# VGND.t737 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=6890,366 d=3510,184
X189 VDPWR.t1078 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t27 VDPWR.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X190 a_16755_12091# ui_in[3].t0 VDPWR.t131 VDPWR.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X191 VDPWR.t1125 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t28 VDPWR.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X192 VDPWR.t1138 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 VDPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X193 ringtest_0.x4.clknet_1_0__leaf_clk.t12 a_21395_6940# VGND.t1045 VGND.t1044 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X194 VGND.t72 VDPWR.t1183 VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X195 VGND.t161 a_21007_3867# ringtest_0.x4.counter[0] VGND.t160 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X196 a_22181_5334# a_21399_5340# a_22097_5334# VDPWR.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X197 a_20318_32213# ui_in[1].t3 a_20492_32319# VGND.t288 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X198 VGND.t339 ringtest_0.x4._00_ a_22399_9142# VGND.t338 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.087554 ps=0.893846 w=0.42 l=0.15
**devattr s=3252,166 d=4368,272
X199 a_22224_6244# a_21951_5878# a_22139_5878# VDPWR.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X200 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VGND.t535 VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X201 VGND.t532 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1.t1 VGND.t531 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X202 VDPWR.t127 ringtest_0.x4.net5 a_23381_4584# VDPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X203 a_26555_5334# ringtest_0.x4._08_ VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X204 ua[2].t5 muxtest_0.x2.x2.GP3 muxtest_0.R3R4.t3 VDPWR.t282 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X205 a_16027_11759# ui_in[3].t1 VDPWR.t56 VDPWR.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X206 VDPWR.t205 a_22541_5058# a_22457_5156# VDPWR.t204 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X207 ringtest_0.x4.clknet_1_1__leaf_clk.t12 a_25364_5878# VGND.t1087 VGND.t1086 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X208 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VGND.t866 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X209 ringtest_0.x4._19_ a_23529_6422# VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X210 a_26569_6422# ringtest_0.x4._23_ VGND.t607 VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X211 a_24895_4790# a_24729_4790# VDPWR.t144 VDPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X212 VDPWR.t313 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR.t312 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X213 ringtest_0.ring_out.t4 ringtest_0.x3.x2.GN1 ua[1].t9 VGND.t530 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X214 ringtest_0.drv_out.t9 a_19289_13081.t4 VGND.t393 VGND.t392 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X215 a_23899_5334# ringtest_0.x4.net6.t5 VDPWR.t1026 VDPWR.t1025 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0 ps=0 w=1 l=0.15
**devattr s=6600,266 d=6600,266
X216 VDPWR.t706 VGND.t1145 VDPWR.t705 VDPWR.t704 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X217 a_24045_6654# a_24336_6544# a_24287_6422# VDPWR.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=2268,138
X218 a_24800_5334# a_24527_5340# a_24715_5334# VDPWR.t816 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X219 muxtest_0.R7R8.t1 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A VGND.t154 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X220 muxtest_0.x2.x2.GP3 muxtest_0.x2.x2.GN3 VGND.t946 VGND.t945 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X221 VGND.t75 VDPWR.t1184 VGND.t74 VGND.t73 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X222 a_25925_6788# ringtest_0.x4._11_.t6 VDPWR.t1043 VDPWR.t1042 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0 ps=0 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X223 ringtest_0.x4.net10 a_27233_5308# VGND.t769 VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X224 VGND.t870 a_21840_5308# a_21798_5712# VGND.t869 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X225 VGND.t140 ui_in[3].t2 muxtest_0.x2.x1.nSEL0 VGND.t139 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X226 VDPWR.t703 VGND.t1146 VDPWR.t702 VDPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X227 VDPWR.t1054 a_22392_5990# a_22319_6244# VDPWR.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X228 VGND.t78 VDPWR.t1185 VGND.t77 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X229 VGND.t477 a_15575_12017# ringtest_0.x3.x2.GN1 VGND.t476 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X230 a_22201_9142# a_21981_9142# VGND.t335 VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.074954 pd=0.823846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4838,217 d=2784,153
X231 ringtest_0.counter7.t3 ringtest_0.x3.x2.GN4 ua[1].t6 VGND.t383 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X232 VDPWR.t226 ringtest_0.x4.net7 a_25925_6788# VDPWR.t225 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X233 VDPWR.t8 a_25975_3867# ringtest_0.x4.counter[6] VDPWR.t7 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X234 VGND.t725 ringtest_0.x4.clknet_0_clk.t33 a_25364_5878# VGND.t724 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X235 VDPWR.t701 VGND.t1147 VDPWR.t700 VDPWR.t699 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X236 VGND.t727 ringtest_0.x4.clknet_0_clk.t34 a_21395_6940# VGND.t726 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X237 a_19114_31955# ui_in[0].t2 VDPWR.t1090 VDPWR.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X238 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VGND.t466 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X239 VDPWR.t698 VGND.t1148 VDPWR.t697 VDPWR.t696 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X240 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR.t893 VDPWR.t892 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X241 VDPWR.t881 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2.t3 VDPWR.t880 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X242 VDPWR.t1016 ringtest_0.x4.clknet_1_0__leaf_clk.t33 a_21509_4790# VDPWR.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X243 VDPWR.t695 VGND.t1149 VDPWR.t694 VDPWR.t616 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X244 a_21803_9508# a_21465_9294# VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=3528,168
X245 a_22052_9116# a_21852_9416# a_22201_9142# VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.064246 ps=0.706154 w=0.36 l=0.15
**devattr s=2784,153 d=2484,141
X246 VGND.t81 VDPWR.t1186 VGND.t80 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X247 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VGND.t504 VGND.t503 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X248 ringtest_0.x4._12_ ringtest_0.x4.net2.t6 a_21132_8918# VGND.t922 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
**devattr s=3835,189 d=3640,186
X249 a_22052_8875# a_21852_8720# a_22201_8964# VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.064246 ps=0.706154 w=0.36 l=0.15
**devattr s=2784,153 d=2484,141
X250 a_27065_5156# a_26201_4790# a_26808_4902# VDPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X251 ringtest_0.x4.clknet_1_0__leaf_clk.t11 a_21395_6940# VGND.t1043 VGND.t1042 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X252 a_21587_5334# ringtest_0.x4._02_ VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X253 VGND.t1057 ui_in[0].t3 muxtest_0.x1.x1.nSEL0 VGND.t1056 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X254 VGND.t84 VDPWR.t1187 VGND.t83 VGND.t82 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X255 VDPWR.t1 a_21465_9294# ringtest_0.x4.net2.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X256 ringtest_0.x4._25_ a_26749_6422# VDPWR.t268 VDPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X257 VDPWR.t52 a_23399_3867# ringtest_0.counter3.t3 VDPWR.t51 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X258 VDPWR.t1123 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t27 VDPWR.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X259 muxtest_0.x2.x2.GP2.t1 muxtest_0.x2.x2.GN2 VGND.t356 VGND.t355 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X260 ringtest_0.x3.x2.GP1.t0 ringtest_0.x3.x2.GN1 VGND.t529 VGND.t528 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X261 VGND.t87 VDPWR.t1188 VGND.t86 VGND.t85 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X262 VDPWR.t693 VGND.t1150 VDPWR.t692 VDPWR.t583 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X263 a_26817_4566# ringtest_0.x4._11_.t7 a_26627_4246# VGND.t1012 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X264 a_22649_6244# a_21951_5878# a_22392_5990# VGND.t740 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X265 VDPWR.t850 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 VDPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X266 VDPWR.t691 VGND.t1151 VDPWR.t690 VDPWR.t536 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X267 VGND.t331 a_21845_9116# a_21852_9416# VGND.t306 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X268 a_21591_6128# ringtest_0.x4._11_.t8 ringtest_0.x4._13_ VDPWR.t1044 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X269 VDPWR.t355 ringtest_0.x4._15_ a_23381_4818# VDPWR.t354 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X270 a_21981_9142# a_21845_9116# a_21561_9116# VDPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.078615 pd=0.771795 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4380,215
X271 VDPWR.t689 VGND.t1152 VDPWR.t688 VDPWR.t687 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X272 VGND.t1085 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t11 VGND.t1084 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X273 VGND.t153 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1.t1 VGND.t152 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X274 muxtest_0.R6R7.t3 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A VGND.t347 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X275 VDPWR.t686 VGND.t1153 VDPWR.t685 VDPWR.t684 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X276 ringtest_0.x4.clknet_0_clk.t12 a_23879_6940# VGND.t636 VGND.t635 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X277 VDPWR.t1145 a_27233_5058# a_27149_5156# VDPWR.t829 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X278 VDPWR.t683 VGND.t1154 VDPWR.t682 VDPWR.t681 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X279 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VGND.t177 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X280 VDPWR.t680 VGND.t1155 VDPWR.t679 VDPWR.t678 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X281 ringtest_0.x4.clknet_1_1__leaf_clk.t26 a_25364_5878# VDPWR.t1121 VDPWR.t1120 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X282 a_26839_6788# a_26569_6422# a_26749_6422# VGND.t850 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X283 VGND.t90 VDPWR.t1189 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X284 VGND.t1041 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t10 VGND.t1040 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X285 VGND.t673 VDPWR.t1190 VGND.t672 VGND.t671 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X286 ringtest_0.x4.net8 a_25393_5308# VDPWR.t384 VDPWR.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X287 VGND.t991 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP4.t1 VGND.t990 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X288 a_24479_4790# ringtest_0.x4.net8 VGND.t736 VGND.t735 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0 ps=0 w=0.42 l=0.15
**devattr s=5266,228 d=1764,126
X289 ringtest_0.x4.net9 a_25761_5058# VGND.t539 VGND.t538 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X290 a_27191_5712# a_26201_5340# a_27065_5334# VGND.t656 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X291 VGND.t605 ringtest_0.x4._23_ a_27273_4220# VGND.t604 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X292 a_25593_5156# a_24895_4790# a_25336_4902# VGND.t650 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X293 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR.t171 VDPWR.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X294 VGND.t746 ringtest_0.x4.net11 a_27489_3702# VGND.t745 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X295 ringtest_0.drv_out.t8 a_19289_13081.t5 VGND.t395 VGND.t394 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X296 ringtest_0.x3.x2.GP3 ringtest_0.x3.x2.GN3 VGND.t1102 VGND.t1101 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X297 VGND.t676 VDPWR.t1191 VGND.t675 VGND.t674 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X298 ringtest_0.counter3.t5 ringtest_0.x3.x2.GN3 ua[1].t14 VGND.t1100 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X299 ringtest_0.x4.clknet_0_clk.t28 a_23879_6940# VDPWR.t419 VDPWR.t418 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X300 a_24699_6200# ringtest_0.x4.net9 a_24627_6200# VDPWR.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2688,148
X301 VGND.t679 VDPWR.t1192 VGND.t678 VGND.t677 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X302 VDPWR.t677 VGND.t1156 VDPWR.t676 VDPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X303 VGND.t681 VDPWR.t1193 muxtest_0.x2.nselect2 VGND.t680 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X304 ringtest_0.x4.clknet_1_0__leaf_clk.t9 a_21395_6940# VGND.t1039 VGND.t1038 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
X305 a_24264_6788# a_23949_6654# VGND.t593 VGND.t592 sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X306 VGND.t146 a_24135_3867# ringtest_0.x4.counter[4] VGND.t145 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X307 VGND.t684 VDPWR.t1194 VGND.t683 VGND.t682 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X308 VDPWR.t784 ringtest_0.x4.clknet_1_1__leaf_clk.t33 a_26201_4790# VDPWR.t783 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X309 a_21465_8830# a_21561_8830# VDPWR.t993 VDPWR.t992 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X310 a_19666_31955# ui_in[1].t4 VDPWR.t105 VDPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X311 VDPWR.t177 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2.t2 VDPWR.t176 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X312 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP2.t5 muxtest_0.R6R7.t0 VDPWR.t67 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X313 ua[0].t8 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A VGND.t989 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X314 ringtest_0.x4.net5 a_22541_5058# VGND.t375 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X315 VGND.t944 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 VGND.t943 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X316 VDPWR.t217 a_16027_11759# ringtest_0.x3.x2.GN2 VDPWR.t216 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X317 VDPWR.t1119 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t25 VDPWR.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X318 VGND.t687 VDPWR.t1195 VGND.t686 VGND.t685 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X319 a_21395_6940# ringtest_0.x4.clknet_0_clk.t35 VGND.t664 VGND.t663 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X320 a_23949_6654# a_24045_6654# VDPWR.t54 VDPWR.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X321 VDPWR.t786 ringtest_0.x4.clknet_1_1__leaf_clk.t34 a_24361_5340# VDPWR.t785 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X322 VDPWR.t193 a_23770_5308# ringtest_0.x4._18_ VDPWR.t192 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6900,269
X323 VGND.t976 a_22765_4478# ringtest_0.x4._14_ VGND.t975 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X324 VDPWR.t369 ringtest_0.ring_out.t10 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR.t368 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X325 VGND.t981 ringtest_0.x4._10_ a_22245_8054# VGND.t980 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=2730,149
X326 a_21675_10006# ringtest_0.x4.net2.t7 VGND.t921 VGND.t920 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X327 VGND.t147 a_22052_8875# a_21981_8976# VGND.t102 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.126592 ps=1.2736 w=0.64 l=0.15
**devattr s=3956,199 d=4838,217
X328 ringtest_0.x4.net9 a_25761_5058# VDPWR.t319 VDPWR.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X329 VDPWR.t675 VGND.t1157 VDPWR.t674 VDPWR.t673 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X330 VGND.t758 a_19289_13081.t6 ringtest_0.drv_out.t7 VGND.t757 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=37200,1324
X331 VGND.t978 a_24968_5308# a_24926_5712# VGND.t977 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X332 VGND.t290 ui_in[1].t5 muxtest_0.x1.x1.nSEL1 VGND.t289 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X333 muxtest_0.x1.x3.GP1.t0 muxtest_0.x1.x3.GN1 VGND.t151 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X334 a_16027_11759# a_16203_12091# a_16155_12151# VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X335 ringtest_0.x4.clknet_0_clk.t11 a_23879_6940# VGND.t634 VGND.t633 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X336 VDPWR.t48 ringtest_0.x4.net1 a_21049_8598# VDPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=10600,506 d=5900,259
X337 VDPWR.t672 VGND.t1158 VDPWR.t671 VDPWR.t670 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
**devattr d=9048,452
X338 VGND.t690 VDPWR.t1196 VGND.t689 VGND.t688 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X339 VGND.t526 a_20318_32213# muxtest_0.x1.x3.GN4 VGND.t525 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X340 muxtest_0.x2.x1.nSEL0 ui_in[3].t3 VDPWR.t58 VDPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X341 a_16155_12151# ui_in[3].t4 VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X342 a_26269_4612# ringtest_0.x4._15_ a_26173_4612# VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3192,160
X343 VDPWR.t669 VGND.t1159 VDPWR.t668 VDPWR.t667 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X344 VDPWR.t666 VGND.t1160 VDPWR.t665 VDPWR.t664 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X345 VGND.t1037 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t8 VGND.t1036 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X346 a_25149_4220# ringtest_0.x4.net9 VDPWR.t298 VDPWR.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0 ps=0 w=0.42 l=0.15
**devattr s=12498,336 d=2352,140
X347 a_22223_5712# a_21233_5340# a_22097_5334# VGND.t951 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X348 muxtest_0.x1.x3.GP4.t0 muxtest_0.x1.x3.GN4 VGND.t988 VGND.t987 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X349 VGND.t692 VDPWR.t1197 VGND.t691 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X350 VGND.t695 VDPWR.t1198 VGND.t694 VGND.t693 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X351 ringtest_0.x4.net5 a_22541_5058# VDPWR.t203 VDPWR.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X352 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR.t85 VDPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X353 VGND.t698 VDPWR.t1199 VGND.t697 VGND.t696 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X354 VGND.t287 ringtest_0.x4._11_.t9 ringtest_0.x4._01_ VGND.t286 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X355 a_22765_5308# ringtest_0.x4._16_.t3 a_23151_5334# VDPWR.t771 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X356 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP1.t4 muxtest_0.R7R8.t4 VDPWR.t1035 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X357 a_25977_4220# ringtest_0.x4._22_ VDPWR.t1052 VDPWR.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0 ps=0 w=0.42 l=0.15
**devattr s=12498,336 d=2352,140
X358 a_25083_4790# ringtest_0.x4._07_ VDPWR.t1161 VDPWR.t1160 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X359 VGND.t701 VDPWR.t1200 VGND.t700 VGND.t699 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X360 VDPWR.t663 VGND.t1161 VDPWR.t662 VDPWR.t661 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X361 a_22983_5654# ringtest_0.x4._16_.t4 ringtest_0.x4._04_ VGND.t659 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=3510,184
X362 VGND.t704 VDPWR.t1201 VGND.t703 VGND.t702 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X363 VDPWR.t60 ui_in[3].t5 ringtest_0.x3.x1.nSEL0 VDPWR.t59 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X364 a_23879_6940# ringtest_0.drv_out.t20 VDPWR.t1020 VDPWR.t1019 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X365 a_22164_4362# ringtest_0.x4._16_.t5 VGND.t1114 VGND.t1113 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=4010,197 d=4368,272
X366 a_25168_5156# a_24729_4790# a_25083_4790# VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X367 VDPWR.t660 VGND.t1162 VDPWR.t659 VDPWR.t658 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X368 VGND.t1019 a_22392_5990# a_22350_5878# VGND.t1018 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X369 VDPWR.t756 ringtest_0.x4._20_ a_23809_4790# VDPWR.t755 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X370 muxtest_0.x2.nselect2 VDPWR.t1202 VGND.t706 VGND.t705 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X371 a_21780_8964# a_21465_8830# VGND.t972 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X372 ringtest_0.x4._11_.t1 a_22245_8054# VGND.t567 VGND.t566 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2730,149 d=2268,138
X373 a_26895_3867# ringtest_0.x4.net9 VDPWR.t296 VDPWR.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X374 a_24715_5334# ringtest_0.x4._06_ VGND.t120 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X375 VGND.t708 VDPWR.t1203 VGND.t707 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X376 VDPWR.t99 ringtest_0.x4._11_.t10 a_23899_5334# VDPWR.t98 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6400,264 d=6600,266
X377 VDPWR.t1117 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t24 VDPWR.t1116 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X378 VDPWR.t332 a_25421_6641# ringtest_0.x4._05_ VDPWR.t331 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X379 muxtest_0.x1.x3.GP3 muxtest_0.x1.x3.GN3 VGND.t837 VGND.t836 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X380 muxtest_0.x1.x4.A muxtest_0.x1.x5.GN ua[3].t3 VDPWR.t119 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X381 ua[2].t2 muxtest_0.x2.x2.GP1.t5 ua[3].t5 VDPWR.t315 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X382 ua[0].t0 muxtest_0.x2.x2.GN2 ua[2].t0 VGND.t354 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X383 a_25294_4790# a_24895_4790# a_25168_5156# VGND.t649 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X384 a_21863_4790# ringtest_0.x4._03_ VDPWR.t251 VDPWR.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X385 VDPWR.t657 VGND.t1163 VDPWR.t656 VDPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X386 VDPWR.t79 a_21007_3867# ringtest_0.x4.counter[0] VDPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X387 VGND.t711 VDPWR.t1204 VGND.t710 VGND.t709 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X388 a_21948_5156# a_21509_4790# a_21863_4790# VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X389 VGND.t714 VDPWR.t1205 VGND.t713 VGND.t712 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X390 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.ring_out.t11 VDPWR.t371 VDPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X391 VGND.t744 ringtest_0.x4.net11 a_27491_4566# VGND.t743 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X392 ringtest_0.x4.net11 a_27233_5058# VGND.t1112 VGND.t1111 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X393 ringtest_0.x4._21_ a_23809_4790# VDPWR.t33 VDPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X394 VGND.t349 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VGND.t348 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X395 VGND.t716 VDPWR.t1206 ringtest_0.x3.nselect2 VGND.t715 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X396 VDPWR.t919 ringtest_0.x4._01_ a_22399_8976# VDPWR.t918 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=4368,272
X397 VDPWR.t417 a_23879_6940# ringtest_0.x4.clknet_0_clk.t27 VDPWR.t416 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X398 a_25149_4220# ringtest_0.x4.net6.t6 a_25547_4612# VGND.t1000 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=4368,272
X399 ringtest_0.x4.net8 a_25393_5308# VGND.t603 VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X400 VGND.t844 a_21425_9686# ringtest_0.x4._00_ VGND.t843 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X401 VGND.t589 a_25336_4902# a_25294_4790# VGND.t588 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X402 VDPWR.t415 a_23879_6940# ringtest_0.x4.clknet_0_clk.t26 VDPWR.t414 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X403 ua[2].t8 muxtest_0.x2.x2.GP4.t4 muxtest_0.R7R8.t5 VDPWR.t762 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X404 a_22139_5878# ringtest_0.x4._04_ VGND.t955 VGND.t954 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X405 ringtest_0.x3.x2.GP2.t2 ringtest_0.x3.x2.GN2 VDPWR.t879 VDPWR.t878 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X406 ringtest_0.x4.clknet_0_clk.t10 a_23879_6940# VGND.t632 VGND.t631 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X407 a_25977_4220# ringtest_0.x4.net10 a_26375_4612# VGND.t774 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=4368,272
X408 VGND.t719 VDPWR.t1207 VGND.t718 VGND.t717 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X409 VGND.t553 a_25421_6641# ringtest_0.x4._05_ VGND.t552 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X410 VDPWR.t969 ringtest_0.x4._24_ a_26749_6422# VDPWR.t968 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X411 VGND.t610 ringtest_0.x4.clknet_1_0__leaf_clk.t34 a_21785_5878# VGND.t609 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X412 VGND.t775 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VGND.t501 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X413 VDPWR.t820 a_19289_13081.t7 ringtest_0.drv_out.t17 VDPWR.t819 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X414 a_22021_4220# a_22164_4362# VDPWR.t266 VDPWR.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
**devattr s=12000,520 d=6600,266
X415 VDPWR.t843 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR.t842 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X416 VGND.t781 VDPWR.t1208 VGND.t780 VGND.t779 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X417 VDPWR.t101 ringtest_0.x4._11_.t11 a_23809_4790# VDPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X418 ua[3].t11 muxtest_0.x2.x2.GN1 ua[2].t15 VGND.t1126 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X419 VDPWR.t655 VGND.t1164 VDPWR.t654 VDPWR.t653 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X420 a_19242_32347# ui_in[0].t4 VGND.t1059 VGND.t1058 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X421 muxtest_0.x1.x3.GP2.t1 muxtest_0.x1.x3.GN2 VGND.t346 VGND.t345 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X422 ringtest_0.x4.clknet_1_0__leaf_clk.t7 a_21395_6940# VGND.t1035 VGND.t1034 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X423 VGND.t941 ringtest_0.x4._24_ a_26839_6788# VGND.t940 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X424 VDPWR.t391 ringtest_0.x4.clknet_1_0__leaf_clk.t35 a_21785_5878# VDPWR.t390 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X425 VGND.t760 a_19289_13081.t8 ringtest_0.drv_out.t6 VGND.t759 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X426 VDPWR.t652 VGND.t1165 VDPWR.t651 VDPWR.t650 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X427 ringtest_0.x4.net11 a_27233_5058# VDPWR.t1144 VDPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X428 muxtest_0.x2.x1.nSEL1 ui_in[4].t4 VDPWR.t115 VDPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X429 a_15575_12017# ringtest_0.x3.x1.nSEL0 a_15749_12123# VGND.t966 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X430 a_25083_4790# ringtest_0.x4._07_ VGND.t1120 VGND.t1119 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X431 VDPWR.t111 a_19666_31955# muxtest_0.x1.x3.GN3 VDPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X432 VGND.t939 ringtest_0.x4._14_ ringtest_0.x4._02_ VGND.t938 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X433 muxtest_0.R1R2.t2 ua[0].t4 VGND.t467 sky130_fd_pr__res_high_po_1p41 l=1.75
X434 VGND.t784 VDPWR.t1209 VGND.t783 VGND.t782 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X435 VGND.t630 a_23879_6940# ringtest_0.x4.clknet_0_clk.t9 VGND.t629 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X436 VGND.t670 ringtest_0.x4.clknet_1_1__leaf_clk.t35 a_24729_4790# VGND.t669 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X437 a_26808_5308# a_26640_5334# VGND.t756 VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X438 VDPWR.t1115 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t23 VDPWR.t1114 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X439 VDPWR.t649 VGND.t1166 VDPWR.t648 VDPWR.t450 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X440 VDPWR.t647 VGND.t1167 VDPWR.t646 VDPWR.t456 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X441 VGND.t787 VDPWR.t1210 VGND.t786 VGND.t785 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X442 VGND.t790 VDPWR.t1211 VGND.t789 VGND.t788 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X443 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP4.t4 muxtest_0.R4R5.t2 VDPWR.t956 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X444 VDPWR.t873 ringtest_0.x4.net4 a_21591_6128# VDPWR.t872 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X445 a_21055_5334# ringtest_0.x4._13_ VDPWR.t877 VDPWR.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X446 VDPWR.t288 a_11845_23906# muxtest_0.x2.x2.GN1 VDPWR.t287 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X447 VGND.t865 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VGND.t174 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X448 VDPWR.t645 VGND.t1168 VDPWR.t644 VDPWR.t643 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X449 a_21395_6940# ringtest_0.x4.clknet_0_clk.t36 VGND.t666 VGND.t665 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X450 VDPWR.t800 ringtest_0.x4.net8 a_25149_4220# VDPWR.t799 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=3108,158
X451 ringtest_0.drv_out.t16 a_19289_13081.t9 VDPWR.t822 VDPWR.t821 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X452 VDPWR.t889 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR.t888 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X453 VDPWR.t642 VGND.t1169 VDPWR.t641 VDPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X454 a_25168_5156# a_24895_4790# a_25083_4790# VDPWR.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X455 VDPWR.t787 ringtest_0.x4.clknet_1_1__leaf_clk.t36 a_26201_5340# VDPWR.t783 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X456 VDPWR.t1028 ringtest_0.x4.net6.t7 a_22795_5334# VDPWR.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X457 a_25364_5878# ringtest_0.x4.clknet_0_clk.t37 VDPWR.t782 VDPWR.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X458 a_21863_4790# ringtest_0.x4._03_ VGND.t471 VGND.t470 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X459 ringtest_0.x3.nselect2 VDPWR.t1212 VGND.t792 VGND.t791 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X460 a_23949_6654# a_24045_6654# VGND.t138 VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X461 a_23529_6422# a_23349_6422# VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X462 a_25055_3867# ringtest_0.x4.net7 VGND.t402 VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X463 a_26555_4790# ringtest_0.x4._09_ VDPWR.t264 VDPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X464 a_22795_5334# a_22765_5308# ringtest_0.x4._04_ VDPWR.t991 sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.3 ps=2.6 w=1 l=0.15
**devattr s=12000,520 d=10400,504
X465 VDPWR.t982 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP4.t3 VDPWR.t981 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X466 VGND.t795 VDPWR.t1213 VGND.t794 VGND.t793 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X467 VDPWR.t255 ringtest_0.drv_out.t21 a_23879_6940# VDPWR.t254 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X468 ringtest_0.x4._24_ a_26627_4246# VGND.t98 VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0 ps=0 w=0.65 l=0.15
**devattr s=4485,199 d=6890,366
X469 a_26640_5156# a_26201_4790# a_26555_4790# VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X470 a_21675_9686# ringtest_0.x4.net2.t8 VDPWR.t937 VDPWR.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X471 VDPWR.t27 a_22052_9116# a_21981_9142# VDPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.140385 ps=1.378205 w=0.75 l=0.15
**devattr s=4380,215 d=7155,252
X472 VDPWR.t899 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR.t898 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X473 VGND.t465 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VGND.t348 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X474 VDPWR.t639 VGND.t1170 VDPWR.t638 VDPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
**devattr d=9048,452
X475 a_27303_4246# ringtest_0.x4._23_ VDPWR.t389 VDPWR.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X476 a_21948_5156# a_21675_4790# a_21863_4790# VDPWR.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X477 a_13675_24012# ui_in[3].t6 VGND.t1005 VGND.t1004 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X478 VGND.t798 VDPWR.t1214 VGND.t797 VGND.t796 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X479 VGND.t801 VDPWR.t1215 VGND.t800 VGND.t799 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X480 VGND.t804 VDPWR.t1216 VGND.t803 VGND.t802 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X481 a_26766_4790# a_26367_4790# a_26640_5156# VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X482 VGND.t337 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VGND.t158 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X483 VDPWR.t636 VGND.t1171 VDPWR.t635 VDPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X484 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk.t37 VGND.t483 VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X485 VDPWR.t1097 ui_in[2].t2 muxtest_0.x1.x5.GN VDPWR.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X486 a_26721_4246# ringtest_0.x4._15_ VDPWR.t353 VDPWR.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0 ps=0 w=1 l=0.15
**devattr s=6600,266 d=6400,264
X487 VGND.t125 a_22295_3867# ringtest_0.x4.counter[2] VGND.t124 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X488 VGND.t485 ringtest_0.x4.clknet_1_1__leaf_clk.t38 a_24361_5340# VGND.t484 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X489 VGND.t502 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VGND.t501 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X490 VGND.t1096 ringtest_0.x4._05_ a_24883_6800# VGND.t1095 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.087554 ps=0.893846 w=0.42 l=0.15
**devattr s=3252,166 d=4368,272
X491 VDPWR.t376 a_25336_4902# a_25263_5156# VDPWR.t375 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X492 a_20318_32213# ui_in[0].t5 VDPWR.t1092 VDPWR.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X493 VGND.t1011 a_16579_11759# ringtest_0.x3.x2.GN3 VGND.t1010 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X494 ringtest_0.counter7.t2 ringtest_0.x3.x2.GN4 ua[1].t5 VGND.t382 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X495 VDPWR.t634 VGND.t1172 VDPWR.t633 VDPWR.t429 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X496 a_23879_6940# ringtest_0.drv_out.t22 VDPWR.t257 VDPWR.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X497 a_26808_5308# a_26640_5334# VDPWR.t818 VDPWR.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0 ps=0 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X498 ringtest_0.x4.clknet_1_1__leaf_clk.t10 a_25364_5878# VGND.t1083 VGND.t1082 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X499 a_26095_6788# ringtest_0.x4.net7 a_26007_6788# VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X500 ringtest_0.x4._07_ a_24699_6200# VDPWR.t367 VDPWR.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5830,267 d=10400,504
X501 a_21840_5308# a_21672_5334# VGND.t496 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X502 a_15749_12123# ringtest_0.x3.x1.nSEL1 VGND.t729 VGND.t728 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X503 VGND.t807 VDPWR.t1217 VGND.t806 VGND.t805 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X504 VGND.t573 ringtest_0.x4._15_ a_26201_6788# VGND.t572 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X505 VDPWR.t808 ringtest_0.x4.net11 a_27489_3702# VDPWR.t807 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X506 VGND.t370 a_26808_4902# a_26766_4790# VGND.t369 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X507 VDPWR.t632 VGND.t1173 VDPWR.t631 VDPWR.t630 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X508 a_25263_5156# a_24729_4790# a_25168_5156# VDPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X509 VGND.t353 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2.t0 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X510 ua[2].t9 muxtest_0.x2.x2.GP4.t5 muxtest_0.R7R8.t6 VDPWR.t763 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X511 VGND.t628 a_23879_6940# ringtest_0.x4.clknet_0_clk.t8 VGND.t627 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X512 VGND.t809 VDPWR.t1218 VGND.t808 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X513 a_21375_3867# ringtest_0.x4.net3.t5 VGND.t647 VGND.t646 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X514 VDPWR.t292 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR.t291 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X515 VGND.t812 VDPWR.t1219 VGND.t811 VGND.t810 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X516 ringtest_0.x4._15_ a_23381_4584# VDPWR.t847 VDPWR.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X517 VDPWR.t64 a_24135_3867# ringtest_0.x4.counter[4] VDPWR.t63 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X518 VDPWR.t393 ringtest_0.x4.clknet_1_0__leaf_clk.t36 a_21233_5340# VDPWR.t392 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X519 muxtest_0.x1.x1.nSEL1 ui_in[1].t6 VGND.t292 VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X520 ringtest_0.ring_out.t3 ringtest_0.x3.x2.GN1 ua[1].t8 VGND.t527 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X521 ringtest_0.x4._10_ a_21785_8054# VDPWR.t95 VDPWR.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X522 ua[1].t3 ringtest_0.x3.x2.GP3 ringtest_0.counter3.t1 VDPWR.t50 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X523 a_22164_4362# ringtest_0.x4._16_.t6 VDPWR.t1147 VDPWR.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
**devattr s=7430,283 d=4704,280
X524 a_23467_4584# ringtest_0.x4.net4 a_23381_4584# VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X525 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP2.t6 muxtest_0.R2R3.t1 VDPWR.t68 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X526 VGND.t668 ringtest_0.x4.clknet_0_clk.t38 a_21395_6940# VGND.t667 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X527 VDPWR.t629 VGND.t1174 VDPWR.t628 VDPWR.t627 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X528 VGND.t175 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VGND.t174 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X529 a_24685_6788# a_24465_6800# VGND.t406 VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.074954 pd=0.823846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4838,217 d=2784,153
X530 VDPWR.t626 VGND.t1175 VDPWR.t625 VDPWR.t624 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X531 VDPWR.t859 ui_in[6].t0 ringtest_0.ring_out.t7 VDPWR.t858 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X532 VGND.t814 VDPWR.t1220 VGND.t813 VGND.t233 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X533 VGND.t817 VDPWR.t1221 VGND.t816 VGND.t815 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X534 VGND.t1033 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t6 VGND.t1032 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X535 VDPWR.t1050 ringtest_0.x4._22_ a_26721_4246# VDPWR.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6400,264 d=6900,269
X536 VGND.t645 ringtest_0.x4._20_ a_23963_4790# VGND.t644 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X537 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP1.t5 muxtest_0.R7R8.t3 VDPWR.t1036 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X538 a_22695_8304# ringtest_0.x4._12_ ringtest_0.x4._01_ VDPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X539 ringtest_0.x4._17_ a_25925_6788# VDPWR.t263 VDPWR.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X540 muxtest_0.x2.x2.GP4.t2 muxtest_0.x2.x2.GN4 VDPWR.t980 VDPWR.t979 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X541 ringtest_0.x4.clknet_0_clk.t7 a_23879_6940# VGND.t626 VGND.t625 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
X542 a_26555_4790# ringtest_0.x4._09_ VGND.t481 VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X543 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VGND.t778 VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X544 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR.t897 VDPWR.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X545 ringtest_0.x4.clknet_1_1__leaf_clk.t22 a_25364_5878# VDPWR.t1113 VDPWR.t1112 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X546 VDPWR.t935 ringtest_0.x4.net2.t9 a_21785_8054# VDPWR.t934 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X547 a_27169_6641# ringtest_0.x4._25_ VDPWR.t901 VDPWR.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X548 a_24317_4942# ringtest_0.x4.net8 VDPWR.t798 VDPWR.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0 ps=0 w=0.42 l=0.15
**devattr s=5689,267 d=2646,147
X549 ringtest_0.x4._16_.t0 a_23381_4818# VGND.t1094 VGND.t828 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X550 ringtest_0.drv_out.t15 a_19289_13081.t10 VDPWR.t824 VDPWR.t823 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X551 muxtest_0.R5R6.t4 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A VGND.t835 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X552 muxtest_0.R4R5.t0 muxtest_0.R3R4.t4 VGND.t371 sky130_fd_pr__res_high_po_1p41 l=1.75
X553 VGND.t1099 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X554 a_21845_8816# ringtest_0.x4.clknet_1_0__leaf_clk.t37 VGND.t761 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X555 a_27815_3867# ringtest_0.x4.net10 VGND.t773 VGND.t772 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X556 a_21561_9116# a_21845_9116# a_21780_9142# VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2736,148
X557 a_21840_5308# a_21672_5334# VDPWR.t272 VDPWR.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0 ps=0 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X558 muxtest_0.x1.x5.GN ui_in[2].t3 VDPWR.t1099 VDPWR.t1098 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X559 VGND.t933 a_12297_23648# muxtest_0.x2.x2.GN2 VGND.t932 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X560 VDPWR.t988 ringtest_0.x3.x1.nSEL0 a_15575_12017# VDPWR.t987 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X561 ringtest_0.x4.clknet_1_0__leaf_clk.t5 a_21395_6940# VGND.t1031 VGND.t1030 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X562 VGND.t404 a_25149_4220# ringtest_0.x4._22_ VGND.t403 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=7851,266
X563 VDPWR.t211 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP4.t3 VDPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X564 VDPWR.t623 VGND.t1176 VDPWR.t622 VDPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X565 a_21561_8830# a_21845_8816# a_21780_8964# VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2736,148
X566 VDPWR.t621 VGND.t1177 VDPWR.t620 VDPWR.t619 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X567 VGND.t819 VDPWR.t1222 VGND.t818 VGND.t810 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X568 VDPWR.t618 VGND.t1178 VDPWR.t617 VDPWR.t616 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X569 VGND.t159 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VGND.t158 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X570 VGND.t508 a_18662_32213# muxtest_0.x1.x3.GN1 VGND.t507 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X571 VDPWR.t1165 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1.t3 VDPWR.t1164 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X572 VDPWR.t615 VGND.t1179 VDPWR.t614 VDPWR.t613 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X573 VGND.t822 VDPWR.t1223 VGND.t821 VGND.t820 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X574 VDPWR.t31 a_13025_23980# a_12849_23648# VDPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X575 a_21507_9686# ringtest_0.x4.net1 a_21425_9686# VDPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X576 VDPWR.t612 VGND.t1180 VDPWR.t611 VDPWR.t610 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X577 VGND.t825 VDPWR.t1224 VGND.t824 VGND.t823 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X578 a_24045_6654# a_24329_6640# a_24264_6788# VGND.t963 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2736,148
X579 VGND.t937 ringtest_0.x4._14_ a_22390_4566# VGND.t936 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=4290,196 d=3510,184
X580 a_25719_4790# a_24729_4790# a_25593_5156# VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X581 a_17405_12123# ui_in[3].t7 VGND.t1007 VGND.t1006 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X582 VDPWR.t609 VGND.t1181 VDPWR.t608 VDPWR.t459 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X583 ringtest_0.counter3.t4 ringtest_0.x3.x2.GN3 ua[1].t15 VGND.t1097 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X584 a_27169_6641# ringtest_0.x4._25_ VGND.t878 VGND.t877 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X585 ringtest_0.drv_out.t5 a_19289_13081.t11 VGND.t561 VGND.t560 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=37200,1324 d=19800,666
X586 ringtest_0.x3.x1.nSEL0 ui_in[3].t8 VDPWR.t1032 VDPWR.t1031 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X587 VGND.t827 VDPWR.t1225 VGND.t826 VGND.t815 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X588 VDPWR.t413 a_23879_6940# ringtest_0.x4.clknet_0_clk.t25 VDPWR.t412 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X589 VGND.t235 VDPWR.t1226 VGND.t234 VGND.t233 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X590 ringtest_0.x4._00_ ringtest_0.x4.net1 a_21675_10006# VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X591 VDPWR.t1149 ringtest_0.x4._16_.t7 a_24763_6143# VDPWR.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.129 ps=1.18 w=0.42 l=0.15
**devattr s=5160,236 d=5830,267
X592 VGND.t238 VDPWR.t1227 VGND.t237 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X593 a_21803_8598# a_21465_8830# VDPWR.t997 VDPWR.t996 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=3528,168
X594 a_22457_5156# a_21675_4790# a_22373_5156# VDPWR.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X595 a_18836_32319# muxtest_0.x1.x1.nSEL1 VGND.t144 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X596 VGND.t241 VDPWR.t1228 VGND.t240 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X597 VDPWR.t607 VGND.t1182 VDPWR.t606 VDPWR.t605 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X598 a_25364_5878# ringtest_0.x4.clknet_0_clk.t39 VDPWR.t774 VDPWR.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0 ps=0 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X599 VDPWR.t340 a_19289_13081.t12 ringtest_0.drv_out.t14 VDPWR.t339 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=111600,3724
X600 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP3 muxtest_0.R5R6.t1 VDPWR.t122 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X601 muxtest_0.R4R5.t5 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A VGND.t986 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X602 ringtest_0.x4.net6.t0 a_22817_6146# VGND.t750 VGND.t749 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X603 a_24986_5878# ringtest_0.x4._22_ a_24763_6143# VGND.t1015 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2646,147
X604 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP4.t5 muxtest_0.R4R5.t1 VDPWR.t957 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X605 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk.t38 VDPWR.t826 VDPWR.t825 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X606 a_24287_6422# a_23949_6654# VDPWR.t380 VDPWR.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=3528,168
X607 VDPWR.t201 a_26808_4902# a_26735_5156# VDPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X608 a_26640_5334# a_26201_5340# a_26555_5334# VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X609 VGND.t864 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2.t1 VGND.t863 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X610 VDPWR.t259 ringtest_0.drv_out.t23 a_23879_6940# VDPWR.t258 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X611 a_23837_5878# ringtest_0.x4._17_ VGND.t1108 VGND.t1107 sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=4290,196
X612 ringtest_0.ring_out.t8 ui_in[6].t1 VDPWR.t861 VDPWR.t860 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X613 VDPWR.t137 a_21845_8816# a_21852_8720# VDPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X614 ringtest_0.x4.net4 a_22265_5308# VGND.t387 VGND.t386 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X615 VGND.t1009 ui_in[3].t9 a_13025_23980# VGND.t1008 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X616 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP4.t6 ua[0].t6 VDPWR.t958 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X617 VDPWR.t604 VGND.t1183 VDPWR.t603 VDPWR.t602 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X618 VDPWR.t601 VGND.t1184 VDPWR.t600 VDPWR.t599 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X619 a_13501_23906# ui_in[3].t10 VDPWR.t1034 VDPWR.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X620 VGND.t244 VDPWR.t1229 VGND.t243 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X621 a_26735_5156# a_26201_4790# a_26640_5156# VDPWR.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X622 VGND.t247 VDPWR.t1230 VGND.t246 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X623 VDPWR.t598 VGND.t1185 VDPWR.t597 VDPWR.t596 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X624 VGND.t377 a_17231_12017# ringtest_0.x3.x2.GN4 VGND.t376 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X625 ringtest_0.x4.clknet_0_clk.t6 a_23879_6940# VGND.t624 VGND.t623 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X626 VGND.t250 VDPWR.t1231 VGND.t249 VGND.t248 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X627 a_26766_5712# a_26367_5340# a_26640_5334# VGND.t974 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X628 VDPWR.t595 VGND.t1186 VDPWR.t594 VDPWR.t474 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X629 a_21981_8976# a_21845_8816# a_21561_8830# VDPWR.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.078615 pd=0.771795 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4380,215
X630 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VGND.t500 VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X631 a_26007_6788# ringtest_0.x4.net6.t8 a_25925_6788# VGND.t1001 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X632 VDPWR.t593 VGND.t1187 VDPWR.t592 VDPWR.t513 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X633 VDPWR.t363 ringtest_0.x4._21_ a_24070_5852# VDPWR.t362 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=7430,283
X634 VGND.t537 a_25761_5058# a_25719_4790# VGND.t536 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X635 VDPWR.t19 a_12473_23980# a_12297_23648# VDPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X636 a_15575_12017# ringtest_0.x3.x1.nSEL1 VDPWR.t793 VDPWR.t792 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X637 ringtest_0.x4.clknet_0_clk.t24 a_23879_6940# VDPWR.t411 VDPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X638 VGND.t253 VDPWR.t1232 VGND.t252 VGND.t251 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X639 a_24465_6800# a_24329_6640# a_24045_6654# VDPWR.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.078615 pd=0.771795 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4380,215
X640 VGND.t487 ringtest_0.x4.clknet_1_1__leaf_clk.t39 a_26201_5340# VGND.t486 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X641 VDPWR.t1111 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t21 VDPWR.t1110 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X642 VDPWR.t591 VGND.t1188 VDPWR.t590 VDPWR.t589 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X643 ringtest_0.x4._06_ a_24004_6128# VGND.t983 VGND.t982 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X644 VDPWR.t588 VGND.t1189 VDPWR.t587 VDPWR.t586 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
**devattr d=9048,452
X645 ringtest_0.x4.net6.t1 a_22817_6146# VDPWR.t811 VDPWR.t810 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X646 VGND.t834 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 VGND.t833 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X647 VGND.t255 VDPWR.t1233 VGND.t254 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X648 ringtest_0.x4.clknet_1_0__leaf_clk.t4 a_21395_6940# VGND.t1029 VGND.t1028 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X649 ringtest_0.x4.clknet_1_1__leaf_clk.t9 a_25364_5878# VGND.t1081 VGND.t1080 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X650 muxtest_0.x2.x2.GP1.t2 muxtest_0.x2.x2.GN1 VDPWR.t1163 VDPWR.t1162 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X651 VGND.t622 a_23879_6940# ringtest_0.x4.clknet_0_clk.t5 VGND.t621 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X652 VDPWR.t905 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR.t904 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X653 muxtest_0.R1R2.t5 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A VGND.t832 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X654 VGND.t258 VDPWR.t1234 VGND.t257 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X655 a_27065_5334# a_26201_5340# a_26808_5308# VDPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X656 VGND.t107 a_12849_23648# muxtest_0.x2.x2.GN3 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X657 VDPWR.t374 a_25977_4220# ringtest_0.x4._23_ VDPWR.t7 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=12498,336
X658 VDPWR.t765 muxtest_0.x1.x1.nSEL0 a_18662_32213# VDPWR.t764 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X659 a_23349_6422# ringtest_0.x4._17_ VGND.t1106 VGND.t1105 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X660 ringtest_0.x4.clknet_1_1__leaf_clk.t20 a_25364_5878# VDPWR.t1109 VDPWR.t1108 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X661 a_21675_4790# a_21509_4790# VDPWR.t335 VDPWR.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X662 a_21672_5334# a_21233_5340# a_21587_5334# VGND.t950 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X663 a_22765_4478# ringtest_0.x4.net4 a_22939_4584# VGND.t853 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X664 VGND.t296 ui_in[4].t5 a_12473_23980# VGND.t295 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X665 VGND.t1027 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t3 VGND.t1026 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X666 VDPWR.t585 VGND.t1190 VDPWR.t584 VDPWR.t583 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X667 a_25441_4612# ringtest_0.x4.net8 a_25345_4612# VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3192,160
X668 a_27149_5156# a_26367_4790# a_27065_5156# VDPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X669 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VGND.t336 VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X670 VGND.t971 a_21465_8830# ringtest_0.x4.net3.t0 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X671 muxtest_0.R2R3.t3 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A VGND.t344 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X672 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR.t887 VDPWR.t886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X673 a_22224_6244# a_21785_5878# a_22139_5878# VGND.t327 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X674 a_25055_3867# ringtest_0.x4.net7 VDPWR.t224 VDPWR.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X675 VGND.t601 a_25393_5308# a_25351_5712# VGND.t600 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X676 a_21798_5712# a_21399_5340# a_21672_5334# VGND.t516 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X677 muxtest_0.R7R8.t0 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A VGND.t149 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X678 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP2.t7 muxtest_0.R2R3.t0 VDPWR.t69 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X679 VDPWR.t582 VGND.t1191 VDPWR.t581 VDPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X680 VDPWR.t93 a_24763_6143# a_24699_6200# VDPWR.t92 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0672 ps=0.74 w=0.42 l=0.15
**devattr s=2688,148 d=8370,269
X681 VDPWR.t191 a_24536_6699# a_24465_6800# VDPWR.t190 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.140385 ps=1.378205 w=0.75 l=0.15
**devattr s=4380,215 d=7155,252
X682 VDPWR.t830 a_27233_5308# a_27149_5334# VDPWR.t829 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X683 VGND.t261 VDPWR.t1235 VGND.t260 VGND.t259 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X684 VGND.t343 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2.t0 VGND.t342 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X685 VDPWR.t342 a_19289_13081.t13 ringtest_0.drv_out.t13 VDPWR.t341 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X686 a_22350_5878# a_21951_5878# a_22224_6244# VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X687 VGND.t399 ringtest_0.x4.net7 a_23770_5308# VGND.t398 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=8320,388
X688 VGND.t763 ringtest_0.x4.clknet_1_0__leaf_clk.t39 a_21233_5340# VGND.t762 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X689 ringtest_0.x4.clknet_1_0__leaf_clk.t2 a_21395_6940# VGND.t1025 VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X690 VDPWR.t117 ui_in[4].t6 muxtest_0.x2.x1.nSEL1 VDPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X691 a_19289_13081.t0 ringtest_0.ring_out.t12 VGND.t583 VGND.t582 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=34800,1316 d=34800,1316
X692 VDPWR.t579 VGND.t1192 VDPWR.t578 VDPWR.t577 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X693 VDPWR.t776 ringtest_0.x4.clknet_0_clk.t40 a_25364_5878# VDPWR.t775 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X694 ringtest_0.x4.counter[9] a_27489_3702# VGND.t285 VGND.t284 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X695 ringtest_0.x4.clknet_1_1__leaf_clk.t8 a_25364_5878# VGND.t1079 VGND.t1078 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X696 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR.t311 VDPWR.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X697 a_17231_12017# ui_in[3].t11 VDPWR.t909 VDPWR.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X698 VDPWR.t576 VGND.t1193 VDPWR.t575 VDPWR.t574 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X699 VGND.t263 VDPWR.t1236 VGND.t262 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X700 VDPWR.t39 a_22295_3867# ringtest_0.x4.counter[2] VDPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X701 VDPWR.t573 VGND.t1194 VDPWR.t572 VDPWR.t571 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X702 a_22765_5308# ringtest_0.x4.net6.t9 VGND.t1003 VGND.t1002 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X703 ua[3].t1 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A VGND.t298 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X704 VGND.t620 a_23879_6940# ringtest_0.x4.clknet_0_clk.t4 VGND.t619 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X705 ua[2].t7 muxtest_0.x2.x2.GP2.t4 ua[0].t3 VDPWR.t761 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X706 a_22097_5334# a_21233_5340# a_21840_5308# VDPWR.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X707 muxtest_0.R3R4.t8 muxtest_0.x2.x2.GN3 ua[2].t10 VGND.t942 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X708 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR.t903 VDPWR.t902 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X709 VGND.t266 VDPWR.t1237 VGND.t265 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X710 VDPWR.t409 a_23879_6940# ringtest_0.x4.clknet_0_clk.t23 VDPWR.t408 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X711 ringtest_0.x4._19_ a_23529_6422# VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X712 a_23381_4584# ringtest_0.x4.net4 VDPWR.t871 VDPWR.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X713 VGND.t652 a_25593_5156# a_25761_5058# VGND.t651 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X714 a_22139_5878# ringtest_0.x4._04_ VDPWR.t978 VDPWR.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X715 muxtest_0.x2.x1.nSEL0 ui_in[3].t12 VGND.t884 VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X716 VGND.t269 VDPWR.t1238 VGND.t268 VGND.t267 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X717 a_21375_3867# ringtest_0.x4.net3.t6 VDPWR.t758 VDPWR.t757 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X718 a_24317_4942# ringtest_0.x4.net6.t10 VDPWR.t1030 VDPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X719 VDPWR.t197 a_16203_12091# a_16027_11759# VDPWR.t196 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X720 VDPWR.t103 ringtest_0.x4._11_.t12 a_22695_8304# VDPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X721 ringtest_0.x4.clknet_1_0__leaf_clk.t26 a_21395_6940# VDPWR.t1076 VDPWR.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X722 VGND.t272 VDPWR.t1239 VGND.t271 VGND.t270 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X723 VGND.t524 a_26895_3867# ringtest_0.counter7.t4 VGND.t523 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X724 ua[1].t2 ringtest_0.x3.x2.GP3 ringtest_0.counter3.t0 VDPWR.t49 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X725 VGND.t275 VDPWR.t1240 VGND.t274 VGND.t273 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X726 VGND.t1023 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t1 VGND.t1022 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X727 ua[2].t4 muxtest_0.x2.x2.GP3 muxtest_0.R3R4.t2 VDPWR.t281 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X728 VDPWR.t570 VGND.t1195 VDPWR.t569 VDPWR.t568 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X729 VDPWR.t567 VGND.t1196 VDPWR.t566 VDPWR.t565 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X730 VGND.t278 VDPWR.t1241 VGND.t277 VGND.t276 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X731 a_26367_4790# a_26201_4790# VDPWR.t148 VDPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X732 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR.t247 VDPWR.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X733 a_24545_5878# ringtest_0.x4.net9 VGND.t520 VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X734 muxtest_0.R6R7.t2 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A VGND.t341 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X735 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP3 muxtest_0.R5R6.t0 VDPWR.t121 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X736 a_24968_5308# a_24800_5334# VGND.t310 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X737 VDPWR.t213 a_22265_5308# a_22181_5334# VDPWR.t212 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X738 a_13501_23906# ui_in[4].t7 a_13675_24012# VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X739 VGND.t886 ui_in[3].t13 ringtest_0.x3.x1.nSEL0 VGND.t885 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X740 VDPWR.t378 a_23949_6654# ringtest_0.x4.net7 VDPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X741 VGND.t280 VDPWR.t1242 VGND.t279 VGND.t251 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X742 VDPWR.t564 VGND.t1197 VDPWR.t563 VDPWR.t562 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X743 VGND.t571 ringtest_0.x4._15_ a_23467_4818# VGND.t303 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X744 VDPWR.t1074 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t25 VDPWR.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X745 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VGND.t157 VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X746 VGND.t996 ui_in[4].t8 a_16203_12091# VGND.t995 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X747 VDPWR.t561 VGND.t1198 VDPWR.t560 VDPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X748 VGND.t283 VDPWR.t1243 VGND.t282 VGND.t281 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X749 VDPWR.t107 ui_in[1].t7 a_20318_32213# VDPWR.t106 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X750 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP4.t7 ua[0].t5 VDPWR.t959 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X751 a_24004_6128# a_24070_5852# a_23837_5878# VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=4290,196 d=6760,364
X752 VDPWR.t769 a_25593_5156# a_25761_5058# VDPWR.t768 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X753 a_22373_5156# a_21675_4790# a_22116_4902# VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X754 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR.t280 VDPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X755 a_21465_9294# a_21561_9116# VGND.t882 VGND.t881 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X756 VDPWR.t1107 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t19 VDPWR.t1106 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X757 ua[3].t0 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A VGND.t298 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X758 a_23932_6128# ringtest_0.x4.net8 VDPWR.t796 VDPWR.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0 ps=0 w=1 l=0.15
**devattr s=11200,512 d=4200,242
X759 a_23399_3867# ringtest_0.x4.net5 VGND.t300 VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X760 a_27815_3867# ringtest_0.x4.net10 VDPWR.t836 VDPWR.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X761 ringtest_0.x4.clknet_1_1__leaf_clk.t7 a_25364_5878# VGND.t1077 VGND.t1076 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X762 VGND.t7 a_13501_23906# muxtest_0.x2.x2.GN4 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X763 VDPWR.t66 a_22052_8875# a_21981_8976# VDPWR.t65 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.140385 ps=1.378205 w=0.75 l=0.15
**devattr s=4380,215 d=7155,252
X764 VDPWR.t558 VGND.t1199 VDPWR.t557 VDPWR.t556 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X765 ringtest_0.x3.x2.GP4.t2 ringtest_0.x3.x2.GN4 VDPWR.t209 VDPWR.t208 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X766 VDPWR.t913 ringtest_0.x4._11_.t13 a_26721_4246# VDPWR.t912 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6600,266 d=6600,266
X767 a_23899_5654# ringtest_0.x4._15_ VGND.t570 VGND.t569 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0 ps=0 w=0.65 l=0.15
**devattr s=4485,199 d=4160,194
X768 ringtest_0.x3.x2.GP2.t0 ringtest_0.x3.x2.GN2 VGND.t862 VGND.t861 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X769 VDPWR.t189 a_19114_31955# muxtest_0.x1.x3.GN2 VDPWR.t188 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X770 VDPWR.t243 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.ring_out.t2 VDPWR.t242 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X771 VDPWR.t1022 ui_in[4].t9 ringtest_0.x3.x1.nSEL1 VDPWR.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X772 VDPWR.t555 VGND.t1200 VDPWR.t554 VDPWR.t553 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
**devattr d=9048,452
X773 a_24800_5334# a_24361_5340# a_24715_5334# VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X774 VGND.t409 VDPWR.t1244 VGND.t408 VGND.t407 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X775 VGND.t1021 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t0 VGND.t1020 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X776 a_23381_4818# ringtest_0.x4._11_.t14 VDPWR.t915 VDPWR.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X777 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR.t91 VDPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X778 a_21561_9116# a_21852_9416# a_21803_9508# VDPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=2268,138
X779 VGND.t777 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VGND.t497 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X780 VGND.t1075 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t6 VGND.t1074 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X781 a_24968_5308# a_24800_5334# VDPWR.t139 VDPWR.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0 ps=0 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X782 a_24926_5712# a_24527_5340# a_24800_5334# VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X783 VDPWR.t552 VGND.t1201 VDPWR.t551 VDPWR.t550 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X784 VGND.t565 a_22245_8054# ringtest_0.x4._11_.t0 VGND.t564 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X785 a_21132_8918# ringtest_0.x4.net1 VGND.t131 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0 ps=0 w=0.65 l=0.15
**devattr s=6890,366 d=3835,189
X786 ringtest_0.x4._09_ a_27273_4220# VGND.t333 VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0 ps=0 w=0.65 l=0.15
**devattr s=8320,388 d=10010,284
X787 a_24551_4790# ringtest_0.x4.net7 a_24479_4790# VGND.t397 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X788 VGND.t412 VDPWR.t1245 VGND.t411 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X789 muxtest_0.x2.x1.nSEL1 ui_in[4].t10 VGND.t998 VGND.t997 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X790 ua[0].t7 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A VGND.t985 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X791 VDPWR.t961 a_16755_12091# a_16579_11759# VDPWR.t960 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X792 a_27273_4220# ringtest_0.x4._23_ a_27659_4246# VDPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X793 VDPWR.t791 a_24317_4942# ringtest_0.x4._20_ VDPWR.t790 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5689,267
X794 VGND.t767 a_27233_5308# a_27191_5712# VGND.t766 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X795 ua[2].t6 muxtest_0.x2.x2.GP2.t5 ua[0].t2 VDPWR.t760 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X796 VGND.t415 VDPWR.t1246 VGND.t414 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X797 ringtest_0.x4.clknet_0_clk.t22 a_23879_6940# VDPWR.t407 VDPWR.t406 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X798 a_22733_6244# a_21951_5878# a_22649_6244# VDPWR.t803 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X799 VDPWR.t549 VGND.t1202 VDPWR.t548 VDPWR.t426 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X800 VDPWR.t547 VGND.t1203 VDPWR.t546 VDPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X801 a_27273_4220# ringtest_0.x4.net11 VGND.t742 VGND.t741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X802 VDPWR.t1140 a_25225_5334# a_25393_5308# VDPWR.t1139 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X803 a_25225_5334# a_24527_5340# a_24968_5308# VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X804 a_22111_10993# ui_in[5].t0 VDPWR.t1088 VDPWR.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X805 VDPWR.t1072 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t24 VDPWR.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X806 VDPWR.t544 VGND.t1204 VDPWR.t543 VDPWR.t542 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X807 VDPWR.t45 ringtest_0.x4.net1 a_21785_8054# VDPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X808 a_27065_5156# a_26367_4790# a_26808_4902# VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X809 VGND.t868 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VGND.t172 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X810 a_17231_12017# ui_in[4].t11 a_17405_12123# VGND.t999 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X811 ringtest_0.x4._12_ ringtest_0.x4.net3.t7 a_21049_8598# VDPWR.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X812 a_25225_5334# a_24361_5340# a_24968_5308# VDPWR.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X813 VDPWR.t541 VGND.t1205 VDPWR.t540 VDPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X814 VDPWR.t538 VGND.t1206 VDPWR.t537 VDPWR.t536 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X815 VDPWR.t995 a_21465_8830# ringtest_0.x4.net3.t1 VDPWR.t994 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X816 VGND.t418 VDPWR.t1247 VGND.t417 VGND.t416 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X817 muxtest_0.R5R6.t3 muxtest_0.R4R5.t3 VGND.t643 sky130_fd_pr__res_high_po_1p41 l=1.75
X818 ringtest_0.drv_out.t12 a_19289_13081.t14 VDPWR.t344 VDPWR.t343 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=111600,3724 d=59400,1866
X819 VDPWR.t999 a_22765_4478# ringtest_0.x4._14_ VDPWR.t998 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X820 VGND.t389 a_16027_11759# ringtest_0.x3.x2.GN2 VGND.t388 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X821 VGND.t888 ui_in[3].t14 a_16755_12091# VGND.t887 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X822 VGND.t421 VDPWR.t1248 VGND.t420 VGND.t419 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X823 VGND.t960 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP4.t1 VGND.t959 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X824 VDPWR.t869 ringtest_0.x4.net4 a_22765_4478# VDPWR.t868 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X825 a_22074_4790# a_21675_4790# a_21948_5156# VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X826 a_21780_9142# a_21465_9294# VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X827 a_24763_6143# ringtest_0.x4._22_ VDPWR.t1048 VDPWR.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0 ps=0 w=0.42 l=0.15
**devattr s=8370,269 d=5160,236
X828 VGND.t424 VDPWR.t1249 VGND.t423 VGND.t422 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X829 ringtest_0.x4.clknet_1_0__leaf_clk.t23 a_21395_6940# VDPWR.t1070 VDPWR.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X830 ringtest_0.ring_out.t1 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR.t241 VDPWR.t240 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X831 VGND.t876 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VGND.t873 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X832 a_23809_4790# ringtest_0.x4._15_ VDPWR.t351 VDPWR.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X833 VDPWR.t535 VGND.t1207 VDPWR.t534 VDPWR.t441 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X834 VGND.t427 VDPWR.t1250 VGND.t426 VGND.t425 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X835 VGND.t458 muxtest_0.R7R8.t2 VGND.t457 sky130_fd_pr__res_high_po_1p41 l=1.75
X836 VGND.t429 VDPWR.t1251 VGND.t428 VGND.t193 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X837 VDPWR.t533 VGND.t1208 VDPWR.t532 VDPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X838 a_22052_9116# a_21845_9116# a_22228_9508# VDPWR.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=2730,149
X839 a_22939_4584# ringtest_0.x4._11_.t15 VGND.t890 VGND.t889 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X840 VGND.t849 a_22116_4902# a_22074_4790# VGND.t848 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X841 ringtest_0.x4.clknet_1_1__leaf_clk.t18 a_25364_5878# VDPWR.t1105 VDPWR.t1104 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X842 VDPWR.t1024 ui_in[4].t12 a_13501_23906# VDPWR.t1023 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X843 a_22228_9508# a_21981_9142# VDPWR.t169 VDPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0 ps=0 w=0.42 l=0.15
**devattr s=7155,252 d=3066,157
X844 VGND.t1061 ui_in[2].t4 muxtest_0.x1.x5.GN VGND.t1060 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X845 VDPWR.t382 a_25393_5308# a_25309_5334# VDPWR.t381 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X846 a_24895_4790# a_24729_4790# VGND.t314 VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X847 VGND.t385 a_22265_5308# a_22223_5712# VGND.t384 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X848 VGND.t1073 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t5 VGND.t1072 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X849 VGND.t432 VDPWR.t1252 VGND.t431 VGND.t430 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X850 VDPWR.t985 a_24329_6640# a_24336_6544# VDPWR.t984 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X851 VGND.t434 VDPWR.t1253 VGND.t433 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X852 muxtest_0.R7R8.t7 muxtest_0.x2.x2.GN4 ua[2].t12 VGND.t958 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X853 a_26555_5334# ringtest_0.x4._08_ VDPWR.t12 VDPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X854 a_19290_32287# ui_in[1].t8 VDPWR.t109 VDPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X855 muxtest_0.R6R7.t4 muxtest_0.R5R6.t2 VGND.t371 sky130_fd_pr__res_high_po_1p41 l=1.75
X856 VGND.t498 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VGND.t497 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X857 VDPWR.t530 VGND.t1209 VDPWR.t529 VDPWR.t528 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X858 a_26627_4246# ringtest_0.x4.net10 VGND.t771 VGND.t770 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0 ps=0 w=0.65 l=0.15
**devattr s=8320,388 d=4290,196
X859 VGND.t436 VDPWR.t1254 VGND.t435 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X860 a_22775_5878# a_21785_5878# a_22649_6244# VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X861 VGND.t439 VDPWR.t1255 VGND.t438 VGND.t437 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X862 a_22795_5334# ringtest_0.x4._16_.t8 VDPWR.t1151 VDPWR.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X863 ringtest_0.x4._13_ ringtest_0.x4._11_.t16 VGND.t892 VGND.t891 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X864 VGND.t512 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VGND.t511 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X865 VGND.t591 a_23949_6654# ringtest_0.x4.net7 VGND.t590 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X866 VDPWR.t778 ringtest_0.x4.clknet_0_clk.t41 a_25364_5878# VDPWR.t777 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X867 a_26367_5340# a_26201_5340# VDPWR.t770 VDPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X868 VDPWR.t780 ringtest_0.x4.clknet_0_clk.t42 a_21395_6940# VDPWR.t779 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X869 ringtest_0.drv_out.t4 a_19289_13081.t15 VGND.t563 VGND.t562 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X870 ua[1].t12 ringtest_0.x3.x2.GP1.t4 ringtest_0.ring_out.t6 VDPWR.t1012 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X871 VGND.t365 ringtest_0.x4._18_ a_23619_6788# VGND.t364 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X872 VGND.t441 VDPWR.t1256 VGND.t440 VGND.t419 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X873 a_12849_23648# ui_in[4].t13 VDPWR.t925 VDPWR.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X874 ringtest_0.x4.clknet_1_1__leaf_clk.t4 a_25364_5878# VGND.t1071 VGND.t1070 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
X875 VDPWR.t527 VGND.t1210 VDPWR.t526 VDPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X876 a_26640_5156# a_26367_4790# a_26555_4790# VDPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X877 muxtest_0.R3R4.t0 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A VGND.t148 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X878 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP1.t6 muxtest_0.R3R4.t6 VDPWR.t1037 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X879 VGND.t444 VDPWR.t1257 VGND.t443 VGND.t442 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X880 VGND.t447 VDPWR.t1258 VGND.t446 VGND.t445 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X881 VDPWR.t524 VGND.t1211 VDPWR.t523 VDPWR.t522 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X882 a_22399_9142# a_21852_9416# a_22052_9116# VDPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=2310,139
X883 VDPWR.t43 ringtest_0.x4.net1 a_21675_9686# VDPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X884 ringtest_0.x4.counter[9] a_27489_3702# VDPWR.t97 VDPWR.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X885 VGND.t110 ringtest_0.x4.clknet_1_0__leaf_clk.t40 a_21509_4790# VGND.t109 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X886 a_22392_5990# a_22224_6244# VGND.t914 VGND.t913 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X887 muxtest_0.x1.x1.nSEL0 ui_in[0].t6 VDPWR.t234 VDPWR.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X888 a_17377_14114# ui_in[6].t2 ringtest_0.ring_out.t9 VGND.t845 sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X889 ua[1].t13 ringtest_0.x3.x2.GP2.t4 ringtest_0.drv_out.t19 VDPWR.t1093 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X890 VDPWR.t806 ringtest_0.x4.net11 a_27303_4246# VDPWR.t805 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X891 muxtest_0.x2.x2.GP4.t0 muxtest_0.x2.x2.GN4 VGND.t957 VGND.t956 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X892 muxtest_0.R2R3.t4 muxtest_0.R1R2.t3 VGND.t551 sky130_fd_pr__res_high_po_1p41 l=1.75
X893 VGND.t173 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VGND.t172 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X894 ringtest_0.x4.clknet_1_0__leaf_clk.t22 a_21395_6940# VDPWR.t1068 VDPWR.t1067 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X895 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VGND.t875 VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X896 ringtest_0.x4.clknet_0_clk.t3 a_23879_6940# VGND.t618 VGND.t617 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X897 VDPWR.t222 ringtest_0.x4.net7 a_24317_4942# VDPWR.t221 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=2268,138
X898 VGND.t748 a_22817_6146# a_22775_5878# VGND.t747 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X899 VGND.t450 VDPWR.t1259 VGND.t449 VGND.t448 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X900 VDPWR.t301 a_26895_3867# ringtest_0.counter7.t5 VDPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X901 VGND.t874 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VGND.t873 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X902 VDPWR.t521 VGND.t1212 VDPWR.t520 VDPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X903 VDPWR.t1005 ringtest_0.x4._10_ a_22245_8054# VDPWR.t1004 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6500,265
X904 VGND.t1104 a_25225_5334# a_25393_5308# VGND.t1103 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X905 a_21587_5334# ringtest_0.x4._02_ VDPWR.t10 VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X906 muxtest_0.x1.x5.GN ui_in[2].t5 VGND.t661 VGND.t660 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X907 a_25336_4902# a_25168_5156# VGND.t506 VGND.t505 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X908 VGND.t1069 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t3 VGND.t1068 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X909 VGND.t381 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP4.t1 VGND.t380 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X910 VDPWR.t1103 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t17 VDPWR.t1102 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X911 VGND.t453 VDPWR.t1260 VGND.t452 VGND.t451 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X912 ringtest_0.x4.clknet_0_clk.t21 a_23879_6940# VDPWR.t405 VDPWR.t404 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X913 VGND.t1125 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1.t1 VGND.t1124 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X914 ringtest_0.drv_out.t2 ringtest_0.x3.x2.GN2 ua[1].t11 VGND.t860 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X915 VGND.t129 ringtest_0.x4.net1 a_21939_8054# VGND.t128 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X916 a_21399_5340# a_21233_5340# VDPWR.t975 VDPWR.t974 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X917 muxtest_0.x1.x5.A ui_in[2].t6 ua[3].t6 VDPWR.t772 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X918 a_19289_13081.t1 ringtest_0.ring_out.t13 VDPWR.t373 VDPWR.t372 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=104400,3716 d=104400,3716
X919 VDPWR.t518 VGND.t1213 VDPWR.t517 VDPWR.t516 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X920 a_12297_23648# ui_in[3].t15 VDPWR.t911 VDPWR.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X921 a_25345_4612# ringtest_0.x4.net9 VGND.t518 VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0 ps=0 w=0.42 l=0.15
**devattr s=7851,266 d=2772,150
X922 VGND.t456 VDPWR.t1261 VGND.t455 VGND.t454 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X923 VGND.t183 VDPWR.t1262 VGND.t182 VGND.t181 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X924 VDPWR.t1066 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t21 VDPWR.t1065 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X925 VGND.t186 VDPWR.t1263 VGND.t185 VGND.t184 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X926 ringtest_0.x3.x1.nSEL0 ui_in[3].t16 VGND.t840 VGND.t839 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X927 a_25547_4612# ringtest_0.x4.net7 a_25441_4612# VGND.t396 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2436,142
X928 VDPWR.t865 a_22116_4902# a_22043_5156# VDPWR.t864 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X929 VDPWR.t927 ui_in[4].t14 a_17231_12017# VDPWR.t926 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X930 VDPWR.t386 ringtest_0.x4._23_ a_26569_6422# VDPWR.t385 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X931 VDPWR.t321 a_27065_5334# a_27233_5308# VDPWR.t320 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X932 a_27065_5334# a_26367_5340# a_26808_5308# VGND.t973 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X933 ringtest_0.x4._02_ ringtest_0.x4._14_ a_21055_5334# VDPWR.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X934 VDPWR.t515 VGND.t1214 VDPWR.t514 VDPWR.t513 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X935 a_26173_4612# ringtest_0.x4._22_ VGND.t1014 VGND.t1013 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0 ps=0 w=0.42 l=0.15
**devattr s=7851,266 d=2772,150
X936 VGND.t294 a_19666_31955# muxtest_0.x1.x3.GN3 VGND.t293 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X937 ringtest_0.x3.x1.nSEL1 ui_in[4].t15 VDPWR.t929 VDPWR.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X938 a_26375_4612# ringtest_0.x4._11_.t17 a_26269_4612# VGND.t893 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2436,142
X939 VGND.t189 VDPWR.t1264 VGND.t188 VGND.t187 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X940 VGND.t192 VDPWR.t1265 VGND.t191 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X941 a_22043_5156# a_21509_4790# a_21948_5156# VDPWR.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X942 VGND.t534 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VGND.t511 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X943 a_26749_6422# a_26569_6422# VDPWR.t867 VDPWR.t866 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X944 a_23770_5308# ringtest_0.x4.net6.t11 a_23993_5654# VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X945 VGND.t103 a_22052_9116# a_21981_9142# VGND.t102 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.126592 ps=1.2736 w=0.64 l=0.15
**devattr s=3956,199 d=4838,217
X946 a_23399_3867# ringtest_0.x4.net5 VDPWR.t125 VDPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X947 VGND.t195 VDPWR.t1266 VGND.t194 VGND.t193 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X948 ringtest_0.ring_out.t0 ui_in[6].t3 a_17377_14114# VGND.t123 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X949 VDPWR.t261 a_15575_12017# ringtest_0.x3.x2.GN1 VDPWR.t260 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X950 ringtest_0.x4._11_.t2 a_22245_8054# VDPWR.t347 VDPWR.t346 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=6500,265 d=5400,254
X951 ringtest_0.x4._02_ ringtest_0.x4._13_ VGND.t858 VGND.t857 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X952 ringtest_0.x4.clknet_1_0__leaf_clk.t20 a_21395_6940# VDPWR.t1064 VDPWR.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X953 muxtest_0.x1.x4.A muxtest_0.x1.x5.GN ua[3].t2 VDPWR.t119 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X954 VGND.t469 a_22021_4220# ringtest_0.x4._03_ VGND.t468 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4010,197
X955 VGND.t489 ringtest_0.x4.clknet_1_1__leaf_clk.t40 a_26201_4790# VGND.t488 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X956 VDPWR.t512 VGND.t1215 VDPWR.t511 VDPWR.t510 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X957 VDPWR.t509 VGND.t1216 VDPWR.t508 VDPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X958 VDPWR.t506 VGND.t1217 VDPWR.t505 VDPWR.t504 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X959 a_23879_6940# ringtest_0.drv_out.t24 VGND.t475 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X960 ringtest_0.x4._24_ a_26627_4246# VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0 ps=0 w=1 l=0.15
**devattr s=6900,269 d=10600,506
X961 a_25593_5156# a_24729_4790# a_25336_4902# VDPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X962 a_22111_10993# ui_in[5].t1 VGND.t1053 VGND.t1052 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X963 a_21395_6940# ringtest_0.x4.clknet_0_clk.t43 VDPWR.t1153 VDPWR.t1152 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X964 VDPWR.t245 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR.t244 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X965 ua[3].t10 muxtest_0.x2.x2.GN1 ua[2].t14 VGND.t1123 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X966 ringtest_0.drv_out.t1 ringtest_0.x3.x2.GN2 ua[1].t10 VGND.t859 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X967 VGND.t896 ringtest_0.x4._01_ a_22399_8976# VGND.t338 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.087554 ps=0.893846 w=0.42 l=0.15
**devattr s=3252,166 d=4368,272
X968 a_25336_4902# a_25168_5156# VDPWR.t284 VDPWR.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0 ps=0 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X969 VGND.t1067 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t2 VGND.t1066 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X970 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VGND.t872 VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X971 VGND.t198 VDPWR.t1267 VGND.t197 VGND.t196 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X972 VDPWR.t794 a_26808_5308# a_26735_5334# VDPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X973 ringtest_0.x4.clknet_0_clk.t20 a_23879_6940# VDPWR.t403 VDPWR.t402 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X974 VDPWR.t278 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR.t277 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X975 VDPWR.t503 VGND.t1218 VDPWR.t502 VDPWR.t501 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X976 muxtest_0.x2.x2.GP1.t0 muxtest_0.x2.x2.GN1 VGND.t1122 VGND.t1121 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X977 a_21465_9294# a_21561_9116# VDPWR.t907 VDPWR.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X978 VDPWR.t500 VGND.t1219 VDPWR.t499 VDPWR.t498 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X979 ringtest_0.x4._21_ a_23809_4790# VGND.t118 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X980 VGND.t880 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VGND.t584 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X981 VGND.t201 VDPWR.t1268 VGND.t200 VGND.t199 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X982 VGND.t616 a_23879_6940# ringtest_0.x4.clknet_0_clk.t2 VGND.t615 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X983 muxtest_0.R3R4.t7 muxtest_0.R2R3.t5 VGND.t643 sky130_fd_pr__res_high_po_1p41 l=1.75
X984 VDPWR.t1062 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t19 VDPWR.t1061 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X985 a_23891_4790# ringtest_0.x4._11_.t18 a_23809_4790# VGND.t894 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X986 VDPWR.t497 VGND.t1220 VDPWR.t496 VDPWR.t495 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X987 VDPWR.t37 a_22097_5334# a_22265_5308# VDPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X988 a_22097_5334# a_21399_5340# a_21840_5308# VGND.t515 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X989 ua[3].t7 ui_in[2].t7 muxtest_0.x1.x4.A VGND.t662 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X990 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR.t290 VDPWR.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X991 VGND.t916 a_25055_3867# ringtest_0.x4.counter[5] VGND.t915 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X992 VGND.t204 VDPWR.t1269 VGND.t203 VGND.t202 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X993 VDPWR.t317 a_25761_5058# a_25677_5156# VDPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X994 a_26735_5334# a_26201_5340# a_26640_5334# VDPWR.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X995 ua[1].t4 ringtest_0.x3.x2.GP1.t5 ringtest_0.ring_out.t5 VDPWR.t118 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X996 VGND.t614 a_23879_6940# ringtest_0.x4.clknet_0_clk.t1 VGND.t613 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X997 ringtest_0.x4._25_ a_26749_6422# VGND.t492 VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X998 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk.t41 VGND.t112 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X999 VGND.t473 a_19289_13081.t16 ringtest_0.drv_out.t3 VGND.t472 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X1000 VDPWR.t494 VGND.t1221 VDPWR.t493 VDPWR.t492 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X1001 a_22201_8964# a_21981_8976# VGND.t979 VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.074954 pd=0.823846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4838,217 d=2784,153
X1002 VGND.t207 VDPWR.t1270 VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X1003 VGND.t210 VDPWR.t1271 VGND.t209 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X1004 VGND.t213 VDPWR.t1272 VGND.t212 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X1005 a_24135_3867# ringtest_0.x4.net6.t12 VGND.t544 VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X1006 a_26808_4902# a_26640_5156# VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X1007 a_22499_4790# a_21509_4790# a_22373_5156# VGND.t554 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X1008 a_12849_23648# a_13025_23980# a_12977_24040# VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X1009 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VGND.t867 VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1010 VDPWR.t89 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1011 a_22765_4478# ringtest_0.x4._11_.t19 VDPWR.t917 VDPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X1012 VDPWR.t491 VGND.t1222 VDPWR.t490 VDPWR.t489 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1013 a_19842_32287# ui_in[0].t7 VDPWR.t236 VDPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X1014 a_11845_23906# muxtest_0.x2.x1.nSEL0 a_12019_24012# VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X1015 VDPWR.t488 VGND.t1223 VDPWR.t487 VDPWR.t486 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1016 VDPWR.t485 VGND.t1224 VDPWR.t484 VDPWR.t483 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X1017 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR.t181 VDPWR.t180 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1018 VDPWR.t482 VGND.t1225 VDPWR.t481 VDPWR.t480 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
**devattr d=9048,452
X1019 VDPWR.t323 ringtest_0.x4.clknet_1_1__leaf_clk.t41 a_24729_4790# VDPWR.t322 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X1020 a_26367_5340# a_26201_5340# VGND.t654 VGND.t653 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1021 VDPWR.t479 VGND.t1226 VDPWR.t478 VDPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X1022 a_24715_5334# ringtest_0.x4._06_ VDPWR.t35 VDPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X1023 muxtest_0.R4R5.t4 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A VGND.t984 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X1024 a_23619_6788# a_23349_6422# a_23529_6422# VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X1025 VGND.t1065 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t1 VGND.t1064 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X1026 VGND.t918 ui_in[4].t16 muxtest_0.x2.x1.nSEL1 VGND.t917 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1027 a_21049_8598# ringtest_0.x4.net2.t10 VDPWR.t933 VDPWR.t932 sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0 ps=0 w=1 l=0.15
**devattr s=5900,259 d=5600,256
X1028 VGND.t216 VDPWR.t1273 VGND.t215 VGND.t214 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X1029 VGND.t931 a_21375_3867# ringtest_0.x4.counter[1] VGND.t930 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X1030 VGND.t219 VDPWR.t1274 VGND.t218 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X1031 VGND.t541 a_27065_5334# a_27233_5308# VGND.t540 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1032 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR.t839 VDPWR.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1033 VGND.t577 ringtest_0.x4._21_ a_24070_5852# VGND.t576 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4010,197
X1034 a_24527_5340# a_24361_5340# VDPWR.t82 VDPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X1035 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP1.t7 muxtest_0.R3R4.t5 VDPWR.t345 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X1036 VDPWR.t965 a_12297_23648# muxtest_0.x2.x2.GN2 VDPWR.t964 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X1037 a_27149_5334# a_26367_5340# a_27065_5334# VDPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X1038 VDPWR.t230 a_25149_4220# ringtest_0.x4._22_ VDPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=12498,336
X1039 a_21767_5334# a_21233_5340# a_21672_5334# VDPWR.t973 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X1040 VGND.t307 a_21845_8816# a_21852_8720# VGND.t306 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1041 VGND.t222 VDPWR.t1275 VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X1042 ringtest_0.x4.clknet_0_clk.t19 a_23879_6940# VDPWR.t401 VDPWR.t400 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1043 a_25364_5878# ringtest_0.x4.clknet_0_clk.t44 VGND.t1118 VGND.t1117 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X1044 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VGND.t879 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1045 VDPWR.t325 ringtest_0.x4.net6.t13 a_25149_4220# VDPWR.t324 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=4368,272
X1046 VDPWR.t75 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1047 VGND.t225 VDPWR.t1276 VGND.t224 VGND.t223 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X1048 VGND.t373 a_22541_5058# a_22499_4790# VGND.t372 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X1049 VDPWR.t476 VGND.t1227 VDPWR.t475 VDPWR.t474 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1050 VGND.t595 ringtest_0.drv_out.t25 a_23879_6940# VGND.t594 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X1051 a_22486_4246# ringtest_0.x4._14_ a_22021_4220# VDPWR.t966 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=4200,242
X1052 VGND.t363 a_23770_5308# ringtest_0.x4._18_ VGND.t362 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=4485,199
X1053 VDPWR.t834 ringtest_0.x4.net10 a_25977_4220# VDPWR.t833 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=4368,272
X1054 a_12297_23648# a_12473_23980# a_12425_24040# VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X1055 VGND.t585 ringtest_0.ring_out.t14 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VGND.t584 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1056 ua[1].t0 ringtest_0.x3.x2.GP4.t5 ringtest_0.counter7.t0 VDPWR.t1095 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X1057 VDPWR.t307 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1.t3 VDPWR.t306 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1058 ringtest_0.x4.clknet_1_0__leaf_clk.t18 a_21395_6940# VDPWR.t1060 VDPWR.t1059 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1059 a_24536_6699# a_24336_6544# a_24685_6788# VGND.t765 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.064246 ps=0.706154 w=0.36 l=0.15
**devattr s=2784,153 d=2484,141
X1060 VDPWR.t473 VGND.t1228 VDPWR.t472 VDPWR.t471 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
**devattr d=9048,452
X1061 VGND.t227 VDPWR.t1277 VGND.t226 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X1062 a_12425_24040# ui_in[3].t17 VGND.t842 VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X1063 VDPWR.t955 a_27169_6641# ringtest_0.x4._08_ VDPWR.t954 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1064 VDPWR.t303 a_20318_32213# muxtest_0.x1.x3.GN4 VDPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X1065 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR.t883 VDPWR.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1066 VDPWR.t399 a_23879_6940# ringtest_0.x4.clknet_0_clk.t18 VDPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X1067 a_24536_6699# a_24329_6640# a_24712_6422# VDPWR.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=2730,149
X1068 VGND.t312 a_27815_3867# ringtest_0.x4.counter[8] VGND.t311 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X1069 muxtest_0.R1R2.t4 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A VGND.t831 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X1070 ua[1].t7 ringtest_0.x3.x2.GP2.t5 ringtest_0.drv_out.t0 VDPWR.t239 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X1071 a_25421_6641# ringtest_0.x4._19_ VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X1072 VDPWR.t470 VGND.t1229 VDPWR.t469 VDPWR.t468 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X1073 a_23879_6940# ringtest_0.drv_out.t26 VGND.t597 VGND.t596 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X1074 a_21399_5340# a_21233_5340# VGND.t949 VGND.t948 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1075 VGND.t361 a_24536_6699# a_24465_6800# VGND.t360 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.126592 ps=1.2736 w=0.64 l=0.15
**devattr s=3956,199 d=4838,217
X1076 a_24883_6800# a_24329_6640# a_24536_6699# VGND.t962 sky130_fd_pr__nfet_01v8 ad=0.075046 pd=0.766154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=3252,166
X1077 muxtest_0.x2.x2.GP3 muxtest_0.x2.x2.GN3 VDPWR.t972 VDPWR.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1078 a_21395_6940# ringtest_0.x4.clknet_0_clk.t45 VDPWR.t1155 VDPWR.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1079 a_26201_6788# ringtest_0.x4._11_.t20 a_26095_6788# VGND.t895 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X1080 VGND.t329 a_22649_6244# a_22817_6146# VGND.t328 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1081 VGND.t229 VDPWR.t1278 VGND.t228 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X1082 ringtest_0.x4._07_ a_24699_6200# VGND.t581 VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3945,196 d=6760,364
X1083 VDPWR.t164 a_21845_9116# a_21852_9416# VDPWR.t163 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X1084 a_24712_6422# a_24465_6800# VDPWR.t232 VDPWR.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0 ps=0 w=0.42 l=0.15
**devattr s=7155,252 d=3066,157
X1085 VDPWR.t854 ui_in[3].t18 muxtest_0.x2.x1.nSEL0 VDPWR.t853 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1086 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VGND.t171 VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1087 VGND.t1116 ringtest_0.x4._16_.t9 a_22765_5308# VGND.t1115 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1088 VGND.t122 a_22097_5334# a_22265_5308# VGND.t121 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1089 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP3 muxtest_0.R1R2.t0 VDPWR.t120 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X1090 a_16579_11759# ui_in[4].t17 VDPWR.t931 VDPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X1091 VDPWR.t467 VGND.t1230 VDPWR.t466 VDPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X1092 VGND.t928 a_27169_6641# ringtest_0.x4._08_ VGND.t927 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X1093 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR.t274 VDPWR.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1094 muxtest_0.R2R3.t2 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A VGND.t340 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X1095 a_25421_6641# ringtest_0.x4._19_ VGND.t95 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X1096 VDPWR.t41 a_22111_10993# ringtest_0.x4.net1 VDPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1097 ringtest_0.drv_out.t11 a_19289_13081.t17 VDPWR.t253 VDPWR.t252 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X1098 ringtest_0.x3.x2.GP4.t0 ringtest_0.x3.x2.GN4 VGND.t379 VGND.t378 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1099 a_21561_8830# a_21852_8720# a_21803_8598# VDPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=2268,138
X1100 VDPWR.t464 VGND.t1231 VDPWR.t463 VDPWR.t462 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
**devattr d=9048,452
X1101 a_23993_5654# ringtest_0.x4._11_.t21 a_23899_5654# VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
**devattr s=4160,194 d=4290,196
X1102 VDPWR.t461 VGND.t1232 VDPWR.t460 VDPWR.t459 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X1103 VGND.t935 ui_in[1].t9 a_19290_32287# VGND.t934 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X1104 a_17377_14114# ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VGND.t464 VGND.t463 sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1105 VGND.t167 ui_in[4].t18 ringtest_0.x3.x1.nSEL1 VGND.t166 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1106 a_24883_6800# a_24336_6544# a_24536_6699# VDPWR.t827 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=2310,139
X1107 VDPWR.t238 ui_in[0].t8 muxtest_0.x1.x1.nSEL0 VDPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1108 a_18662_32213# muxtest_0.x1.x1.nSEL1 VDPWR.t62 VDPWR.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X1109 VDPWR.t458 VGND.t1233 VDPWR.t457 VDPWR.t456 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1110 VDPWR.t455 VGND.t1234 VDPWR.t454 VDPWR.t453 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X1111 VDPWR.t158 a_22649_6244# a_22817_6146# VDPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X1112 VDPWR.t452 VGND.t1235 VDPWR.t451 VDPWR.t450 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1113 VGND.t1110 a_27233_5058# a_27191_4790# VGND.t1109 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X1114 VDPWR.t29 a_12849_23648# muxtest_0.x2.x2.GN3 VDPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X1115 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.ring_out.t15 VGND.t105 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1116 ringtest_0.x4.clknet_1_1__leaf_clk.t0 a_25364_5878# VGND.t1063 VGND.t1062 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X1117 a_24699_6200# a_24763_6143# a_24545_5878# VGND.t178 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1118 muxtest_0.x2.x2.GP2.t2 muxtest_0.x2.x2.GN2 VDPWR.t185 VDPWR.t184 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1119 ringtest_0.x3.x2.GP1.t2 ringtest_0.x3.x2.GN1 VDPWR.t305 VDPWR.t304 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1120 ringtest_0.x4.clknet_1_1__leaf_clk.t16 a_25364_5878# VDPWR.t1101 VDPWR.t1100 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1121 VDPWR.t146 muxtest_0.x2.x1.nSEL0 a_11845_23906# VDPWR.t145 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X1122 a_21951_5878# a_21785_5878# VGND.t325 VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1123 VGND.t494 a_22373_5156# a_22541_5058# VGND.t493 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1124 VDPWR.t449 VGND.t1236 VDPWR.t448 VDPWR.t447 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
**devattr d=9048,452
X1125 a_25975_3867# ringtest_0.x4.net8 VGND.t733 VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X1126 a_21981_9142# a_21852_9416# a_21561_9116# VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.071208 pd=0.7164 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=3956,199
X1127 VGND.t232 VDPWR.t1279 VGND.t231 VGND.t230 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X1128 VDPWR.t397 a_23879_6940# ringtest_0.x4.clknet_0_clk.t17 VDPWR.t396 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1129 VGND.t18 VDPWR.t1280 VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X1130 a_21981_8976# a_21852_8720# a_21561_8830# VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.071208 pd=0.7164 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=3956,199
X1131 VDPWR.t446 VGND.t1237 VDPWR.t445 VDPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1132 a_22319_6244# a_21785_5878# a_22224_6244# VDPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X1133 VDPWR.t71 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1.t2 VDPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1134 VGND.t21 VDPWR.t1281 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X1135 VDPWR.t990 a_19290_32287# a_19114_31955# VDPWR.t989 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X1136 VGND.t24 VDPWR.t1282 VGND.t23 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X1137 VDPWR.t443 VGND.t1238 VDPWR.t442 VDPWR.t441 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1138 VGND.t27 VDPWR.t1283 VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X1139 a_21951_5878# a_21785_5878# VDPWR.t154 VDPWR.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X1140 ringtest_0.x4._06_ a_24004_6128# VDPWR.t1007 VDPWR.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=7430,283 d=10400,504
X1141 VDPWR.t1001 a_24968_5308# a_24895_5334# VDPWR.t1000 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X1142 a_24465_6800# a_24336_6544# a_24045_6654# VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.071208 pd=0.7164 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=3956,199
X1143 VDPWR.t440 VGND.t1239 VDPWR.t439 VDPWR.t438 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X1144 a_22390_4566# a_22164_4362# a_22021_4220# VGND.t490 sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X1145 VDPWR.t1157 ringtest_0.x4.clknet_0_clk.t46 a_21395_6940# VDPWR.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X1146 VDPWR.t195 ringtest_0.x4._18_ a_23529_6422# VDPWR.t194 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X1147 VDPWR.t1009 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP4.t2 VDPWR.t1008 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1148 a_12977_24040# ui_in[4].t19 VGND.t169 VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X1149 VDPWR.t437 VGND.t1240 VDPWR.t436 VDPWR.t435 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
**devattr d=9048,452
X1150 ringtest_0.x4._10_ a_21785_8054# VGND.t180 VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X1151 VGND.t612 a_23879_6940# ringtest_0.x4.clknet_0_clk.t0 VGND.t611 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X1152 a_23963_4790# ringtest_0.x4._15_ a_23891_4790# VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X1153 VDPWR.t1058 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t17 VDPWR.t1057 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1154 VGND.t30 VDPWR.t1284 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X1155 a_24895_5334# a_24361_5340# a_24800_5334# VDPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X1156 a_23770_5308# ringtest_0.x4.net7 a_23899_5334# VDPWR.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6600,266 d=12800,528
X1157 a_22399_9142# a_21845_9116# a_22052_9116# VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.075046 pd=0.766154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=3252,166
X1158 a_21867_8054# ringtest_0.x4.net2.t11 a_21785_8054# VGND.t919 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X1159 VDPWR.t434 VGND.t1241 VDPWR.t433 VDPWR.t432 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X1160 ringtest_0.x4._04_ a_22765_5308# VGND.t969 VGND.t968 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0 ps=0 w=0.65 l=0.15
**devattr s=8320,388 d=10010,284
X1161 VGND.t33 VDPWR.t1285 VGND.t32 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X1162 ringtest_0.x4.clknet_0_clk.t16 a_23879_6940# VDPWR.t395 VDPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X1163 a_25364_5878# ringtest_0.x4.clknet_0_clk.t47 VGND.t546 VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X1164 a_22399_8976# a_21845_8816# a_22052_8875# VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.075046 pd=0.766154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=3252,166
X1165 a_20492_32319# ui_in[0].t9 VGND.t460 VGND.t459 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X1166 ringtest_0.x3.x2.GP3 ringtest_0.x3.x2.GN3 VDPWR.t1137 VDPWR.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1167 VDPWR.t270 a_22373_5156# a_22541_5058# VDPWR.t269 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X1168 VDPWR.t431 VGND.t1242 VDPWR.t430 VDPWR.t429 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1169 a_22052_8875# a_21845_8816# a_22228_8598# VDPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=2730,149
X1170 a_22228_8598# a_21981_8976# VDPWR.t1003 VDPWR.t1002 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0 ps=0 w=0.42 l=0.15
**devattr s=7155,252 d=3066,157
X1171 ringtest_0.x4._01_ ringtest_0.x4._12_ VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1172 VGND.t599 ringtest_0.drv_out.t27 a_23879_6940# VGND.t598 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X1173 ringtest_0.x4._16_.t1 a_23381_4818# VDPWR.t1133 VDPWR.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X1174 a_23151_5334# ringtest_0.x4.net6.t14 VDPWR.t327 VDPWR.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1175 VDPWR.t944 VDPWR.t942 muxtest_0.x2.nselect2 VDPWR.t943 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1176 VGND.t510 a_11845_23906# muxtest_0.x2.x2.GN1 VGND.t509 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X1177 a_22295_3867# ringtest_0.x4.net4 VGND.t852 VGND.t851 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X1178 VDPWR.t428 VGND.t1243 VDPWR.t427 VDPWR.t426 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X1179 a_13025_23980# ui_in[3].t19 VDPWR.t856 VDPWR.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X1180 VGND.t462 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B a_17377_14114# VGND.t461 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1181 VGND.t36 VDPWR.t1286 VGND.t35 VGND.t34 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X1182 VDPWR.t923 a_25055_3867# ringtest_0.x4.counter[5] VDPWR.t922 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1183 VGND.t953 ringtest_0.x4.net6.t15 a_22983_5654# VGND.t952 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1184 VDPWR.t970 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 VDPWR.t924 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1185 ringtest_0.x4.clknet_1_0__leaf_clk.t16 a_21395_6940# VDPWR.t1056 VDPWR.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
R0 ringtest_0.x4.net2.n14 ringtest_0.x4.net2.t1 315.034
R1 ringtest_0.x4.net2.t0 ringtest_0.x4.net2.n14 265.769
R2 ringtest_0.x4.net2 ringtest_0.x4.net2.t0 262.318
R3 ringtest_0.x4.net2.n4 ringtest_0.x4.net2.t5 260.322
R4 ringtest_0.x4.net2.n9 ringtest_0.x4.net2.t10 241.536
R5 ringtest_0.x4.net2.n0 ringtest_0.x4.net2.t8 212.081
R6 ringtest_0.x4.net2.n1 ringtest_0.x4.net2.t3 212.081
R7 ringtest_0.x4.net2.n6 ringtest_0.x4.net2.t9 183.505
R8 ringtest_0.x4.net2.n4 ringtest_0.x4.net2.t2 175.169
R9 ringtest_0.x4.net2.n9 ringtest_0.x4.net2.t6 169.237
R10 ringtest_0.x4.net2.n10 ringtest_0.x4.net2.n9 159.952
R11 ringtest_0.x4.net2.n7 ringtest_0.x4.net2.n6 153.863
R12 ringtest_0.x4.net2.n3 ringtest_0.x4.net2.n2 152.698
R13 ringtest_0.x4.net2.n5 ringtest_0.x4.net2.n4 152
R14 ringtest_0.x4.net2.n0 ringtest_0.x4.net2.t7 139.78
R15 ringtest_0.x4.net2.n1 ringtest_0.x4.net2.t4 139.78
R16 ringtest_0.x4.net2.n6 ringtest_0.x4.net2.t11 114.532
R17 ringtest_0.x4.net2.n2 ringtest_0.x4.net2.n0 37.246
R18 ringtest_0.x4.net2.n8 ringtest_0.x4.net2.n5 34.4715
R19 ringtest_0.x4.net2.n2 ringtest_0.x4.net2.n1 24.1005
R20 ringtest_0.x4.net2.n12 ringtest_0.x4.net2.n3 18.9449
R21 ringtest_0.x4.net2.n13 ringtest_0.x4.net2.n12 14.916
R22 ringtest_0.x4.net2.n11 ringtest_0.x4.net2.n10 13.8005
R23 ringtest_0.x4.net2 ringtest_0.x4.net2.n7 10.8927
R24 ringtest_0.x4.net2.n14 ringtest_0.x4.net2.n13 8.72777
R25 ringtest_0.x4.net2.n8 ringtest_0.x4.net2 6.07742
R26 ringtest_0.x4.net2.n10 ringtest_0.x4.net2 3.33963
R27 ringtest_0.x4.net2.n10 ringtest_0.x4.net2 3.29747
R28 ringtest_0.x4.net2 ringtest_0.x4.net2.n13 3.29747
R29 ringtest_0.x4.net2.n11 ringtest_0.x4.net2.n8 3.19006
R30 ringtest_0.x4.net2.n3 ringtest_0.x4.net2 1.97868
R31 ringtest_0.x4.net2.n7 ringtest_0.x4.net2 1.97868
R32 ringtest_0.x4.net2.n5 ringtest_0.x4.net2 1.55726
R33 ringtest_0.x4.net2.n12 ringtest_0.x4.net2.n11 1.38649
R34 VGND.n3406 VGND.n64 4.7454e+06
R35 VGND.n318 VGND.n65 4.7454e+06
R36 VGND.n3406 VGND.n65 3.52e+06
R37 VGND.n360 VGND.n64 3.52e+06
R38 VGND.n3212 VGND.n173 3.3176e+06
R39 VGND.n3281 VGND.n3280 3.3176e+06
R40 VGND.n378 VGND.n376 2.347e+06
R41 VGND.n376 VGND.n64 2.3386e+06
R42 VGND.n3191 VGND.n173 2.3386e+06
R43 VGND.n3281 VGND.n3250 2.3386e+06
R44 VGND.n321 VGND.n66 2.15447e+06
R45 VGND.n3250 VGND.n3249 2.1446e+06
R46 VGND.n3192 VGND.n3191 2.1446e+06
R47 VGND.n3283 VGND.n3234 1.86572e+06
R48 VGND.n303 VGND.n65 1.2338e+06
R49 VGND.n334 VGND.n65 1.18072e+06
R50 VGND.n310 VGND.n309 1.1798e+06
R51 VGND.n3284 VGND.n3232 1.1798e+06
R52 VGND.n3229 VGND.n176 1.1798e+06
R53 VGND.n311 VGND.n310 1.17976e+06
R54 VGND.n3284 VGND.n3233 1.17976e+06
R55 VGND.n3229 VGND.n3228 1.17976e+06
R56 VGND.n376 VGND.t152 1.17724e+06
R57 VGND.n3250 VGND.t378 1.17707e+06
R58 VGND.n3191 VGND.t956 1.17707e+06
R59 VGND.n3405 VGND.t845 1.0027e+06
R60 VGND.n3077 VGND.n224 573621
R61 VGND.n323 VGND.n318 396385
R62 VGND.n362 VGND.n360 396385
R63 VGND.n3214 VGND.n3212 396385
R64 VGND.n3280 VGND.n3279 396385
R65 VGND.n318 VGND.n317 391216
R66 VGND.n360 VGND.n359 391216
R67 VGND.n3280 VGND.n3251 391216
R68 VGND.n3212 VGND.n3211 391216
R69 VGND.n3283 VGND.n3282 293853
R70 VGND.n3405 VGND.n66 291597
R71 VGND.n3290 VGND.n3289 86912.4
R72 VGND.n3290 VGND.n66 81673.6
R73 VGND.n3235 VGND.n67 72143.6
R74 VGND.n310 VGND.n172 66245.4
R75 VGND.n3061 VGND.n224 61252.6
R76 VGND.n3081 VGND.n172 52488.3
R77 VGND.n3289 VGND.n3288 52128.6
R78 VGND.n3394 VGND.n3393 38301.6
R79 VGND VGND.n175 35992.3
R80 VGND.n3407 VGND.n63 35421.6
R81 VGND.n3395 VGND.n3394 29605.7
R82 VGND.n3288 VGND.n173 29419.1
R83 VGND.n3288 VGND.n172 29145.5
R84 VGND.n399 VGND 25742.3
R85 VGND.n2394 VGND 23608
R86 VGND.n3404 VGND.n67 18854
R87 VGND.n3288 VGND.n3287 17410.5
R88 VGND.n341 VGND.n222 16580.9
R89 VGND.n2394 VGND.t757 13977.5
R90 VGND VGND.n173 13964.9
R91 VGND.n3231 VGND.n174 13854.2
R92 VGND.n369 VGND.n341 13333.2
R93 VGND.n3289 VGND.n74 13232.9
R94 VGND.n379 VGND.n371 11744.7
R95 VGND.n383 VGND.n371 11744.7
R96 VGND.n379 VGND.n372 11744.7
R97 VGND.n383 VGND.n372 11744.7
R98 VGND.n358 VGND.n346 11744.7
R99 VGND.n354 VGND.n346 11744.7
R100 VGND.n358 VGND.n348 11744.7
R101 VGND.n354 VGND.n348 11744.7
R102 VGND.n396 VGND.n282 11744.7
R103 VGND.n396 VGND.n388 11744.7
R104 VGND.n388 VGND.n280 11744.7
R105 VGND.n282 VGND.n280 11744.7
R106 VGND.n335 VGND.n284 11744.7
R107 VGND.n339 VGND.n284 11744.7
R108 VGND.n335 VGND.n285 11744.7
R109 VGND.n339 VGND.n285 11744.7
R110 VGND.n316 VGND.n293 11744.7
R111 VGND.n312 VGND.n293 11744.7
R112 VGND.n316 VGND.n294 11744.7
R113 VGND.n312 VGND.n294 11744.7
R114 VGND.n304 VGND.n298 11744.7
R115 VGND.n308 VGND.n298 11744.7
R116 VGND.n304 VGND.n299 11744.7
R117 VGND.n308 VGND.n299 11744.7
R118 VGND.n320 VGND.n291 11744.7
R119 VGND.n320 VGND.n292 11744.7
R120 VGND.n324 VGND.n292 11744.7
R121 VGND.n324 VGND.n291 11744.7
R122 VGND.n363 VGND.n342 11744.7
R123 VGND.n367 VGND.n342 11744.7
R124 VGND.n363 VGND.n343 11744.7
R125 VGND.n367 VGND.n343 11744.7
R126 VGND.n3248 VGND.n3236 11744.7
R127 VGND.n3243 VGND.n3236 11744.7
R128 VGND.n3248 VGND.n3238 11744.7
R129 VGND.n3243 VGND.n3238 11744.7
R130 VGND.n3266 VGND.n3263 11744.7
R131 VGND.n3266 VGND.n3264 11744.7
R132 VGND.n3268 VGND.n3263 11744.7
R133 VGND.n3268 VGND.n3264 11744.7
R134 VGND.n206 VGND.n197 11744.7
R135 VGND.n206 VGND.n199 11744.7
R136 VGND.n199 VGND.n196 11744.7
R137 VGND.n197 VGND.n196 11744.7
R138 VGND.n3210 VGND.n177 11744.7
R139 VGND.n3227 VGND.n177 11744.7
R140 VGND.n3210 VGND.n178 11744.7
R141 VGND.n3227 VGND.n178 11744.7
R142 VGND.n3194 VGND.n185 11744.7
R143 VGND.n3194 VGND.n186 11744.7
R144 VGND.n3196 VGND.n185 11744.7
R145 VGND.n3196 VGND.n186 11744.7
R146 VGND.n3215 VGND.n3204 11744.7
R147 VGND.n3215 VGND.n3208 11744.7
R148 VGND.n3205 VGND.n3204 11744.7
R149 VGND.n3208 VGND.n3205 11744.7
R150 VGND.n3391 VGND.n75 11744.7
R151 VGND.n3391 VGND.n76 11744.7
R152 VGND.n75 VGND.n73 11744.7
R153 VGND.n76 VGND.n73 11744.7
R154 VGND.n3278 VGND.n3252 11744.7
R155 VGND.n3278 VGND.n3254 11744.7
R156 VGND.n3257 VGND.n3252 11744.7
R157 VGND.n3257 VGND.n3254 11744.7
R158 VGND.n3076 VGND.n225 11744.7
R159 VGND.n3072 VGND.n226 11744.7
R160 VGND.n3076 VGND.n226 11744.7
R161 VGND.n3059 VGND.n3057 11744.7
R162 VGND.n3063 VGND.n3057 11744.7
R163 VGND.n3060 VGND.n3059 11744.7
R164 VGND.n3063 VGND.n3060 11744.7
R165 VGND.n370 VGND.n369 9554.71
R166 VGND.n3396 VGND.n3395 9243.96
R167 VGND.n3082 VGND.n3081 8452.32
R168 VGND.n3078 VGND.n222 7337.33
R169 VGND.n323 VGND.t989 7088.89
R170 VGND.t985 VGND.n321 7088.89
R171 VGND.n362 VGND.t984 7088.89
R172 VGND.n368 VGND.t986 7088.89
R173 VGND.n3214 VGND.t958 7088.89
R174 VGND.t961 VGND.n174 7088.89
R175 VGND.n3279 VGND.t382 7088.89
R176 VGND.t383 VGND.n3234 7088.89
R177 VGND.n303 VGND.t340 6925.66
R178 VGND.n309 VGND.t344 6925.66
R179 VGND.n317 VGND.t831 6925.66
R180 VGND.n311 VGND.t832 6925.66
R181 VGND.n3249 VGND.t860 6925.66
R182 VGND.t859 VGND.n3232 6925.66
R183 VGND.t1097 VGND.n3251 6925.66
R184 VGND.t1100 VGND.n3233 6925.66
R185 VGND.t357 VGND.n3192 6925.66
R186 VGND.t354 VGND.n176 6925.66
R187 VGND.n3211 VGND.t942 6925.66
R188 VGND.n3228 VGND.t947 6925.66
R189 VGND.n359 VGND.t838 6925.66
R190 VGND.t835 VGND.n283 6925.66
R191 VGND.n378 VGND.t341 6925.66
R192 VGND.n384 VGND.t347 6925.66
R193 VGND.n3081 VGND.t959 6843.4
R194 VGND.t989 VGND.n322 6733.33
R195 VGND.n322 VGND.t985 6733.33
R196 VGND.t984 VGND.n361 6733.33
R197 VGND.n361 VGND.t986 6733.33
R198 VGND.t958 VGND.n3213 6733.33
R199 VGND.n3213 VGND.t961 6733.33
R200 VGND.n3253 VGND.t382 6733.33
R201 VGND.n3253 VGND.t383 6733.33
R202 VGND.t340 VGND.n302 6578.29
R203 VGND.n302 VGND.t344 6578.29
R204 VGND.n297 VGND.t831 6578.29
R205 VGND.t832 VGND.n297 6578.29
R206 VGND.n3237 VGND.t860 6578.29
R207 VGND.n3237 VGND.t859 6578.29
R208 VGND.n3267 VGND.t1097 6578.29
R209 VGND.n3267 VGND.t1100 6578.29
R210 VGND.n3195 VGND.t357 6578.29
R211 VGND.n3195 VGND.t354 6578.29
R212 VGND.t942 VGND.n3209 6578.29
R213 VGND.n3209 VGND.t947 6578.29
R214 VGND.n347 VGND.t838 6578.29
R215 VGND.n347 VGND.t835 6578.29
R216 VGND.t341 VGND.n377 6578.29
R217 VGND.n377 VGND.t347 6578.29
R218 VGND.n334 VGND.t155 6418.9
R219 VGND.n340 VGND.t148 6418.9
R220 VGND.t155 VGND.n333 6096.95
R221 VGND.n333 VGND.t148 6096.95
R222 VGND.n386 VGND.n385 5782.24
R223 VGND.n385 VGND.n370 5742.37
R224 VGND.n479 VGND.n423 5452.27
R225 VGND.n479 VGND.n470 5452.27
R226 VGND.n423 VGND.n421 5452.27
R227 VGND.n470 VGND.n421 5452.27
R228 VGND.n467 VGND.n428 5452.27
R229 VGND.n459 VGND.n428 5452.27
R230 VGND.n467 VGND.n429 5452.27
R231 VGND.n459 VGND.n429 5452.27
R232 VGND.n489 VGND.n402 5452.27
R233 VGND.n419 VGND.n402 5452.27
R234 VGND.n489 VGND.n403 5452.27
R235 VGND.n419 VGND.n403 5452.27
R236 VGND.n434 VGND.n425 5452.27
R237 VGND.n461 VGND.n434 5452.27
R238 VGND.n437 VGND.n425 5452.27
R239 VGND.n461 VGND.n437 5452.27
R240 VGND.n413 VGND.n400 5452.27
R241 VGND.n416 VGND.n413 5452.27
R242 VGND.n414 VGND.n400 5452.27
R243 VGND.n416 VGND.n414 5452.27
R244 VGND.n439 VGND.n427 5452.27
R245 VGND.n458 VGND.n439 5452.27
R246 VGND.n440 VGND.n427 5452.27
R247 VGND.n458 VGND.n440 5452.27
R248 VGND.n481 VGND.n410 5452.27
R249 VGND.n411 VGND.n410 5452.27
R250 VGND.n481 VGND.n480 5452.27
R251 VGND.n480 VGND.n411 5452.27
R252 VGND.n451 VGND.n449 5452.27
R253 VGND.n453 VGND.n449 5452.27
R254 VGND.n452 VGND.n451 5452.27
R255 VGND.n453 VGND.n452 5452.27
R256 VGND.n2392 VGND.n1001 5434.88
R257 VGND.n2392 VGND.n1003 5434.88
R258 VGND.n1003 VGND.n1000 5434.88
R259 VGND.n1001 VGND.n1000 5434.88
R260 VGND.n3230 VGND.n3229 5417.76
R261 VGND.n3082 VGND.n3080 5047.41
R262 VGND VGND.t810 4888.89
R263 VGND.n3080 VGND.n3079 4736.53
R264 VGND.t810 VGND 4408.43
R265 VGND.n385 VGND.n384 4081.58
R266 VGND.n370 VGND.n283 4038.16
R267 VGND.t46 VGND.t37 3877.39
R268 VGND.t820 VGND.t43 3877.39
R269 VGND.n310 VGND.n222 3666.67
R270 VGND.n1010 VGND.n1007 3464.88
R271 VGND.n1013 VGND.n1007 3464.88
R272 VGND.n1010 VGND.n1008 3464.88
R273 VGND.n1013 VGND.n1008 3464.88
R274 VGND.n3230 VGND.n175 3363.82
R275 VGND VGND.t696 3346.36
R276 VGND.t430 VGND 3346.36
R277 VGND.t902 VGND 3346.36
R278 VGND.t276 VGND 3346.36
R279 VGND VGND.t281 3346.36
R280 VGND VGND.t208 3346.36
R281 VGND VGND.t73 3346.36
R282 VGND.n3062 VGND.n3061 3340.87
R283 VGND.n3078 VGND.n3077 3323.88
R284 VGND.n198 VGND.n175 3119.26
R285 VGND.t845 VGND.n3404 3111.89
R286 VGND.t34 VGND.t793 3101.92
R287 VGND.t451 VGND.t779 3101.92
R288 VGND.t782 VGND.t823 3101.92
R289 VGND.n386 VGND.n224 2996.82
R290 VGND.n2031 VGND 2973.14
R291 VGND.n3284 VGND.n3283 2937.79
R292 VGND.n172 VGND.n66 2904
R293 VGND.n369 VGND.n368 2881.39
R294 VGND VGND.t259 2857.47
R295 VGND VGND.t52 2857.47
R296 VGND.t422 VGND 2857.47
R297 VGND.t25 VGND 2857.47
R298 VGND.t40 VGND 2857.47
R299 VGND VGND.t688 2857.47
R300 VGND.n3285 VGND.n3284 2647.82
R301 VGND.n341 VGND.n340 2595.64
R302 VGND.n399 VGND.n398 2555.51
R303 VGND.n1222 VGND 2552.48
R304 VGND.t1024 VGND.t28 2495.02
R305 VGND.n2037 VGND 2469.73
R306 VGND VGND.t58 2452.87
R307 VGND VGND.t217 2452.87
R308 VGND.t815 VGND.t236 2326.44
R309 VGND.t79 VGND.t193 2326.44
R310 VGND.t242 VGND.t85 2326.44
R311 VGND VGND.t248 2081.99
R312 VGND.t425 VGND 2081.99
R313 VGND.n3079 VGND.n223 2065.3
R314 VGND.n198 VGND.t1123 2053.05
R315 VGND.n3285 VGND.n3231 2012.27
R316 VGND.n207 VGND.t1123 1950.07
R317 VGND.n2036 VGND.t64 1938.7
R318 VGND.t1126 VGND.n207 1926.65
R319 VGND.n2035 VGND.n1222 1896.67
R320 VGND.n2035 VGND.n2034 1896.67
R321 VGND.n2034 VGND.n2033 1896.67
R322 VGND.n2033 VGND.n2032 1896.67
R323 VGND.n2032 VGND.n2031 1896.67
R324 VGND.t248 VGND 1812.26
R325 VGND VGND.t34 1795.4
R326 VGND.t779 VGND 1795.4
R327 VGND VGND.t782 1795.4
R328 VGND VGND.t410 1795.4
R329 VGND.n3406 VGND.n3405 1791.03
R330 VGND VGND.t897 1786.97
R331 VGND.t245 VGND 1786.97
R332 VGND VGND.t205 1786.97
R333 VGND VGND.t70 1702.68
R334 VGND VGND.n1368 1677.39
R335 VGND.t2 VGND.t881 1593.1
R336 VGND.t766 VGND.t540 1593.1
R337 VGND.t493 VGND.t372 1593.1
R338 VGND.t306 VGND.t338 1584.67
R339 VGND.t491 VGND.t927 1584.67
R340 VGND.t117 VGND.t187 1567.82
R341 VGND.t696 VGND.t211 1550.96
R342 VGND.t259 VGND.t430 1550.96
R343 VGND.t52 VGND.t902 1550.96
R344 VGND.t843 VGND.t132 1550.96
R345 VGND.t413 VGND.t276 1550.96
R346 VGND.t281 VGND.t785 1550.96
R347 VGND.t208 VGND.t25 1550.96
R348 VGND.t73 VGND.t40 1550.96
R349 VGND.t688 VGND.t245 1550.96
R350 VGND.n3084 VGND.t6 1550.96
R351 VGND.n3083 VGND.n3080 1530.43
R352 VGND VGND.t442 1502.01
R353 VGND.n491 VGND.n399 1445.53
R354 VGND.t332 VGND.t549 1416.09
R355 VGND VGND.t233 1407.66
R356 VGND.t256 VGND 1407.66
R357 VGND VGND.t671 1407.66
R358 VGND.t31 VGND 1407.66
R359 VGND.t828 VGND 1407.66
R360 VGND VGND.t419 1407.66
R361 VGND VGND.t251 1399.23
R362 VGND.t572 VGND.t478 1399.23
R363 VGND.t4 VGND 1390.8
R364 VGND.t211 VGND 1306.51
R365 VGND.t793 VGND 1306.51
R366 VGND VGND.t88 1306.51
R367 VGND.t897 VGND 1306.51
R368 VGND VGND.t413 1306.51
R369 VGND VGND.t451 1306.51
R370 VGND.t64 VGND 1306.51
R371 VGND.t264 VGND 1306.51
R372 VGND.t785 VGND 1306.51
R373 VGND.t823 VGND 1306.51
R374 VGND.t273 VGND 1306.51
R375 VGND VGND.t220 1306.51
R376 VGND.t28 VGND 1306.51
R377 VGND VGND.t49 1306.51
R378 VGND.t205 VGND 1306.51
R379 VGND.n2938 VGND.n522 1294.86
R380 VGND.t1054 VGND 1289.66
R381 VGND VGND.t887 1289.66
R382 VGND.t1008 VGND 1289.66
R383 VGND VGND.t1119 1272.8
R384 VGND.n3463 VGND.t525 1229.99
R385 VGND.n3421 VGND.n3408 1198.25
R386 VGND.n3462 VGND.n3461 1198.25
R387 VGND.n3368 VGND.n86 1198.25
R388 VGND.n113 VGND.n112 1198.25
R389 VGND.n71 VGND.n68 1198.25
R390 VGND.n3403 VGND.n3402 1198.25
R391 VGND.n1420 VGND.n1419 1198.25
R392 VGND.n1931 VGND.n1917 1198.25
R393 VGND.n2030 VGND.n2029 1198.25
R394 VGND.n2498 VGND.n2395 1198.25
R395 VGND.n2986 VGND.n2985 1198.25
R396 VGND.n2988 VGND.n2987 1198.25
R397 VGND.n2036 VGND.n581 1196.22
R398 VGND.n2038 VGND.n2037 1196.22
R399 VGND.n3464 VGND.n3463 1194.5
R400 VGND.n3190 VGND.n3189 1194.5
R401 VGND.n3094 VGND.n219 1194.5
R402 VGND.n3085 VGND.n3084 1194.5
R403 VGND.n3316 VGND.n72 1194.5
R404 VGND.n2236 VGND.n2225 1194.5
R405 VGND.n2224 VGND.n2223 1194.5
R406 VGND.n2725 VGND.n731 1194.5
R407 VGND.n2790 VGND.n693 1194.5
R408 VGND.n1500 VGND.n1368 1194.5
R409 VGND.n2594 VGND.n842 1194.5
R410 VGND.n1661 VGND.n1581 1194.5
R411 VGND.n1916 VGND.n1915 1194.5
R412 VGND.t576 VGND.t398 1188.51
R413 VGND.n3446 VGND.n38 1171.32
R414 VGND.n3175 VGND.n208 1171.32
R415 VGND.n95 VGND.n94 1171.32
R416 VGND.n1916 VGND.t651 1146.36
R417 VGND VGND.t843 1137.93
R418 VGND.n3393 VGND.n3392 1105.32
R419 VGND.t768 VGND 1104.21
R420 VGND.t948 VGND 1078.93
R421 VGND.t720 VGND.t735 1078.93
R422 VGND.t644 VGND.t117 1078.93
R423 VGND.t286 VGND 1070.5
R424 VGND.t179 VGND 1036.78
R425 VGND.t478 VGND 1036.78
R426 VGND.n491 VGND.n490 1032.02
R427 VGND VGND.t422 1019.92
R428 VGND VGND.t46 1019.92
R429 VGND VGND.t820 1019.92
R430 VGND.t220 VGND 1019.92
R431 VGND.t334 VGND.t102 1003.07
R432 VGND.t606 VGND 1003.07
R433 VGND.t846 VGND.t848 1003.07
R434 VGND.n2173 VGND.n2172 999.607
R435 VGND.n2142 VGND.n2141 999.607
R436 VGND.n2680 VGND.n2679 999.607
R437 VGND.t92 VGND.t617 960.92
R438 VGND.t747 VGND.t659 952.49
R439 VGND.t338 VGND.t305 944.062
R440 VGND.t480 VGND.t318 944.062
R441 VGND.t555 VGND.t470 944.062
R442 VGND VGND.n2224 927.203
R443 VGND.n731 VGND 927.203
R444 VGND.n3463 VGND 918.774
R445 VGND VGND.t507 918.774
R446 VGND VGND.n70 918.774
R447 VGND.t236 VGND 918.774
R448 VGND.n2225 VGND 918.774
R449 VGND.t233 VGND 918.774
R450 VGND VGND.t79 918.774
R451 VGND.t251 VGND 918.774
R452 VGND.t85 VGND 918.774
R453 VGND VGND.n693 918.774
R454 VGND VGND.t256 918.774
R455 VGND.t671 VGND 918.774
R456 VGND VGND.t31 918.774
R457 VGND.t190 VGND 918.774
R458 VGND.t419 VGND 918.774
R459 VGND VGND.n72 918.774
R460 VGND.t476 VGND 918.774
R461 VGND.n3084 VGND 918.774
R462 VGND.t509 VGND 918.774
R463 VGND.t303 VGND.t828 910.346
R464 VGND.t6 VGND.t1004 910.346
R465 VGND.n1419 VGND 901.917
R466 VGND.n1917 VGND 901.917
R467 VGND.t100 VGND.t308 893.487
R468 VGND.t740 VGND.t326 893.487
R469 VGND.n1432 VGND.n1431 870.4
R470 VGND.n1222 VGND 851.341
R471 VGND VGND.n2035 851.341
R472 VGND.t102 VGND.t100 851.341
R473 VGND.n2034 VGND 851.341
R474 VGND.n2033 VGND 851.341
R475 VGND.n2032 VGND 851.341
R476 VGND.t495 VGND.t515 851.341
R477 VGND.n2031 VGND 851.341
R478 VGND VGND.t854 851.341
R479 VGND VGND.n3082 851.341
R480 VGND.t578 VGND.t164 842.913
R481 VGND.n3080 VGND.n222 839.237
R482 VGND.t305 VGND.t101 834.484
R483 VGND.t101 VGND.t334 834.484
R484 VGND.t754 VGND.t162 834.484
R485 VGND.t569 VGND.t362 834.484
R486 VGND.t739 VGND.t1018 834.484
R487 VGND.t950 VGND.t516 834.484
R488 VGND.t316 VGND.t649 834.484
R489 VGND.t293 VGND.t751 826.054
R490 VGND.t358 VGND.t1058 826.054
R491 VGND.t940 VGND.t491 826.054
R492 VGND.t214 VGND.t99 826.054
R493 VGND.t490 VGND.t846 826.054
R494 VGND.t113 VGND.t1010 826.054
R495 VGND.t141 VGND.t388 826.054
R496 VGND.t168 VGND.t106 826.054
R497 VGND.t841 VGND.t932 826.054
R498 VGND.t895 VGND.t572 809.196
R499 VGND.t1119 VGND.t403 809.196
R500 VGND.n314 VGND.n313 807.013
R501 VGND.n307 VGND.n306 807.013
R502 VGND.n319 VGND.n290 807.013
R503 VGND.n338 VGND.n337 807.013
R504 VGND.n382 VGND.n381 807.013
R505 VGND.n356 VGND.n355 807.013
R506 VGND.n366 VGND.n365 807.013
R507 VGND.n204 VGND.n203 807.013
R508 VGND.t796 VGND 805.538
R509 VGND.t308 VGND.t2 800.766
R510 VGND.t980 VGND.t566 800.766
R511 VGND.t656 VGND.t766 800.766
R512 VGND.t319 VGND.t1109 800.766
R513 VGND.t289 VGND.t934 792.337
R514 VGND.t564 VGND.t802 792.337
R515 VGND.t400 VGND.t230 792.337
R516 VGND.t995 VGND.t166 792.337
R517 VGND.t295 VGND.t917 792.337
R518 VGND.n315 VGND.n314 785.722
R519 VGND.n306 VGND.n305 785.722
R520 VGND.n325 VGND.n290 785.722
R521 VGND.n337 VGND.n336 785.722
R522 VGND.n381 VGND.n380 785.722
R523 VGND.n357 VGND.n356 785.722
R524 VGND.n365 VGND.n364 785.722
R525 VGND.n203 VGND.n202 785.722
R526 VGND.t936 VGND.t559 783.909
R527 VGND.t410 VGND.t425 775.48
R528 VGND.n3074 VGND.n3073 767.294
R529 VGND.n3058 VGND.n3056 767.294
R530 VGND.n313 VGND.n296 763.106
R531 VGND.n307 VGND.n300 763.106
R532 VGND.n319 VGND.n289 763.106
R533 VGND.n338 VGND.n286 763.106
R534 VGND.n382 VGND.n373 763.106
R535 VGND.n355 VGND.n353 763.106
R536 VGND.n366 VGND.n344 763.106
R537 VGND.n205 VGND.n204 763.106
R538 VGND.n3073 VGND.n3070 763.106
R539 VGND.n3058 VGND.n3055 763.106
R540 VGND.n394 VGND.n393 763.09
R541 VGND.n3245 VGND.n3244 763.09
R542 VGND.n3269 VGND.n3262 763.09
R543 VGND.n3226 VGND.n3225 763.09
R544 VGND.n3207 VGND.n3206 763.09
R545 VGND.n3197 VGND.n184 763.09
R546 VGND.n3389 VGND.n3388 763.09
R547 VGND.n3259 VGND.n3258 763.09
R548 VGND.t1105 VGND.t214 758.621
R549 VGND.t1113 VGND.t558 758.621
R550 VGND.t922 VGND.t130 750.192
R551 VGND.n296 VGND.n295 748.977
R552 VGND.n301 VGND.n300 748.977
R553 VGND.n332 VGND.n286 748.977
R554 VGND.n345 VGND.n344 748.977
R555 VGND.n326 VGND.n289 748.977
R556 VGND.n375 VGND.n373 748.977
R557 VGND.n353 VGND.n352 748.977
R558 VGND.n205 VGND.n201 748.977
R559 VGND.t927 VGND.t877 741.763
R560 VGND.t1001 VGND.t400 741.763
R561 VGND.t1068 VGND.t973 741.763
R562 VGND.t893 VGND.t774 741.763
R563 VGND.n393 VGND.n392 732.236
R564 VGND.n3246 VGND.n3245 732.236
R565 VGND.n3270 VGND.n3269 732.236
R566 VGND.n3225 VGND.n3224 732.236
R567 VGND.n3207 VGND.n3202 732.236
R568 VGND.n3198 VGND.n3197 732.236
R569 VGND.n3388 VGND.n3387 732.236
R570 VGND.n3276 VGND.n3259 732.236
R571 VGND.t992 VGND.t922 724.904
R572 VGND.t474 VGND.t594 724.904
R573 VGND.t619 VGND.t641 724.904
R574 VGND.t625 VGND.t621 724.904
R575 VGND.t639 VGND.t637 724.904
R576 VGND.t635 VGND.t639 724.904
R577 VGND.t667 VGND.t663 724.904
R578 VGND.t663 VGND.t726 724.904
R579 VGND.t726 VGND.t665 724.904
R580 VGND.t665 VGND.t1036 724.904
R581 VGND.t1036 VGND.t1042 724.904
R582 VGND.t1046 VGND.t1050 724.904
R583 VGND.t1050 VGND.t1040 724.904
R584 VGND.t1040 VGND.t1044 724.904
R585 VGND.t1044 VGND.t1048 724.904
R586 VGND.t1048 VGND.t1038 724.904
R587 VGND.t1022 VGND.t1028 724.904
R588 VGND.t1028 VGND.t1032 724.904
R589 VGND.t1032 VGND.t1034 724.904
R590 VGND.t1034 VGND.t1026 724.904
R591 VGND.t1026 VGND.t1030 724.904
R592 VGND.t1030 VGND.t1020 724.904
R593 VGND.t1076 VGND.t1072 724.904
R594 VGND.t1070 VGND.t1066 724.904
R595 VGND.t1082 VGND.t1084 724.904
R596 VGND.t724 VGND.t1117 724.904
R597 VGND.t1117 VGND.t722 724.904
R598 VGND.t538 VGND.t1013 724.904
R599 VGND.t598 VGND.t552 716.476
R600 VGND.t1092 VGND.t196 716.476
R601 VGND.t398 VGND.t533 716.476
R602 VGND.t542 VGND.t1107 716.476
R603 VGND.n3392 VGND.n74 709.47
R604 VGND.t660 VGND.t1060 708.047
R605 VGND.t291 VGND.t289 708.047
R606 VGND.t0 VGND.t1056 708.047
R607 VGND.t143 VGND.t648 708.047
R608 VGND.n3395 VGND.n70 708.047
R609 VGND.t104 VGND.t584 708.047
R610 VGND.t156 VGND.t158 708.047
R611 VGND.t350 VGND.t348 708.047
R612 VGND.t170 VGND.t172 708.047
R613 VGND.t176 VGND.t174 708.047
R614 VGND.t513 VGND.t511 708.047
R615 VGND.t499 VGND.t497 708.047
R616 VGND.t503 VGND.t501 708.047
R617 VGND.t871 VGND.t873 708.047
R618 VGND.n3291 VGND.n3290 708.047
R619 VGND.t132 VGND.t920 708.047
R620 VGND.t920 VGND.t923 708.047
R621 VGND.t923 VGND.t133 708.047
R622 VGND.t111 VGND.t306 708.047
R623 VGND.t881 VGND.t4 708.047
R624 VGND.t8 VGND.t286 708.047
R625 VGND.t566 VGND.t564 708.047
R626 VGND.t519 VGND.t578 708.047
R627 VGND.t1002 VGND.t1115 708.047
R628 VGND.t954 VGND.t951 708.047
R629 VGND.t891 VGND.t855 708.047
R630 VGND.t762 VGND.t948 708.047
R631 VGND.t857 VGND.t938 708.047
R632 VGND.t743 VGND.t741 708.047
R633 VGND.t488 VGND.t320 708.047
R634 VGND.t669 VGND.t313 708.047
R635 VGND.t854 VGND.t303 708.047
R636 VGND.t556 VGND.t109 708.047
R637 VGND.n3394 VGND.n72 708.047
R638 VGND.t715 VGND.t791 708.047
R639 VGND.t166 VGND.t115 708.047
R640 VGND.t885 VGND.t839 708.047
R641 VGND.t966 VGND.t728 708.047
R642 VGND.t680 VGND.t705 708.047
R643 VGND.t917 VGND.t997 708.047
R644 VGND.t139 VGND.t883 708.047
R645 VGND.t317 VGND.t547 708.047
R646 VGND.t405 VGND.t631 699.617
R647 VGND.t617 VGND.t590 691.188
R648 VGND.t709 VGND.t768 691.188
R649 VGND.t600 VGND.t545 691.188
R650 VGND.t468 VGND 682.76
R651 VGND.n208 VGND.t717 681.482
R652 VGND.n94 VGND.t805 681.482
R653 VGND.t613 VGND.t137 674.331
R654 VGND.t1084 VGND 674.331
R655 VGND.t178 VGND.t119 674.331
R656 VGND.t586 VGND.t538 674.331
R657 VGND.t850 VGND.t940 657.471
R658 VGND.t99 VGND.t364 657.471
R659 VGND.t386 VGND.t740 657.471
R660 VGND.t1016 VGND.t322 657.471
R661 VGND VGND.t61 649.043
R662 VGND.t952 VGND.t749 640.614
R663 VGND.t659 VGND.t328 640.614
R664 VGND.n3291 VGND 632.184
R665 VGND VGND.t815 632.184
R666 VGND.n2224 VGND 632.184
R667 VGND.n2225 VGND 632.184
R668 VGND.t193 VGND 632.184
R669 VGND.n2037 VGND 632.184
R670 VGND VGND.n2036 632.184
R671 VGND VGND.t242 632.184
R672 VGND VGND.n731 632.184
R673 VGND VGND.n693 632.184
R674 VGND.t70 VGND 632.184
R675 VGND.n1368 VGND 632.184
R676 VGND.t592 VGND.t611 632.184
R677 VGND.n1419 VGND 632.184
R678 VGND.t58 VGND 632.184
R679 VGND.t1088 VGND.t602 632.184
R680 VGND VGND.n842 632.184
R681 VGND.t217 VGND 632.184
R682 VGND.n1917 VGND 632.184
R683 VGND.t1066 VGND.t14 623.755
R684 VGND.t1062 VGND.t755 615.327
R685 VGND.n1581 VGND.t1088 615.327
R686 VGND.t1090 VGND.t1103 615.327
R687 VGND.t91 VGND.t737 615.327
R688 VGND.t994 VGND.t128 606.898
R689 VGND.t919 VGND.t994 606.898
R690 VGND.t82 VGND.t1024 606.898
R691 VGND.t655 VGND.t1080 606.898
R692 VGND.t397 VGND.t330 606.898
R693 VGND.t735 VGND.t397 606.898
R694 VGND.t568 VGND.t644 606.898
R695 VGND.t894 VGND.t568 606.898
R696 VGND.t889 VGND.t374 606.898
R697 VGND.t239 VGND.n38 606.351
R698 VGND.n70 VGND.n69 599.125
R699 VGND.n3292 VGND.n3291 599.125
R700 VGND.t641 VGND.t964 598.467
R701 VGND.t968 VGND.t747 598.467
R702 VGND.t575 VGND.t367 598.467
R703 VGND.t734 VGND.t505 598.467
R704 VGND.t301 VGND.t554 598.467
R705 VGND.t765 VGND.t627 590.038
R706 VGND VGND.t850 581.61
R707 VGND.t615 VGND.t482 581.61
R708 VGND VGND.t857 581.61
R709 VGND.t608 VGND.t1111 573.181
R710 VGND.n3061 VGND.n175 570.136
R711 VGND VGND.t660 564.751
R712 VGND VGND.t0 564.751
R713 VGND.t648 VGND 564.751
R714 VGND.n398 VGND 564.751
R715 VGND VGND.t104 564.751
R716 VGND VGND.t156 564.751
R717 VGND VGND.t350 564.751
R718 VGND VGND.t170 564.751
R719 VGND VGND.t176 564.751
R720 VGND VGND.t513 564.751
R721 VGND VGND.t499 564.751
R722 VGND VGND.t503 564.751
R723 VGND VGND.t871 564.751
R724 VGND.n2394 VGND 564.751
R725 VGND.n2394 VGND 564.751
R726 VGND.t128 VGND 564.751
R727 VGND.n2394 VGND 564.751
R728 VGND.n2394 VGND 564.751
R729 VGND.t327 VGND.t384 564.751
R730 VGND.n2394 VGND 564.751
R731 VGND VGND.t853 564.751
R732 VGND.n2394 VGND 564.751
R733 VGND.t791 VGND 564.751
R734 VGND.t839 VGND 564.751
R735 VGND VGND.t966 564.751
R736 VGND.n3393 VGND 564.751
R737 VGND.t297 VGND 564.751
R738 VGND.t705 VGND 564.751
R739 VGND.t883 VGND 564.751
R740 VGND VGND.t317 564.751
R741 VGND.t459 VGND.t525 563.702
R742 VGND VGND.t980 556.322
R743 VGND.t963 VGND.t633 556.322
R744 VGND.t396 VGND.t650 556.322
R745 VGND VGND.t919 547.894
R746 VGND VGND.t606 547.894
R747 VGND VGND.t1001 547.894
R748 VGND VGND.t1105 547.894
R749 VGND.t309 VGND.t657 547.894
R750 VGND.t362 VGND 547.894
R751 VGND.t324 VGND.t495 547.894
R752 VGND VGND.t894 547.894
R753 VGND VGND.t8 539.465
R754 VGND VGND.t416 539.465
R755 VGND.t907 VGND 531.034
R756 VGND.t37 VGND 531.034
R757 VGND.t43 VGND 531.034
R758 VGND VGND.t223 531.034
R759 VGND.t685 VGND.t126 526.468
R760 VGND.t184 VGND.t143 522.606
R761 VGND VGND.t92 522.606
R762 VGND.t1086 VGND 522.606
R763 VGND.t728 VGND.t799 522.606
R764 VGND.n3083 VGND.t297 522.606
R765 VGND.t547 VGND.t712 522.606
R766 VGND VGND.t179 514.177
R767 VGND.t121 VGND.t913 514.177
R768 VGND VGND.t480 514.177
R769 VGND.t1015 VGND.t754 505.748
R770 VGND VGND.t12 505.748
R771 VGND.t55 VGND.t1046 497.318
R772 VGND.t974 VGND.t1064 497.318
R773 VGND VGND.t889 497.318
R774 VGND.t1018 VGND.t121 488.889
R775 VGND VGND.t967 480.461
R776 VGND.t962 VGND.t623 480.461
R777 VGND.t1074 VGND.t653 480.461
R778 VGND.t164 VGND 480.461
R779 VGND VGND.t536 480.461
R780 VGND.t366 VGND 480.461
R781 VGND.t96 VGND 480.461
R782 VGND VGND.t677 473.495
R783 VGND VGND.t19 473.495
R784 VGND VGND.t674 473.495
R785 VGND.n2395 VGND.t693 465.17
R786 VGND VGND.t598 463.603
R787 VGND.t623 VGND.t1095 463.603
R788 VGND.t629 VGND.t360 463.603
R789 VGND.t717 VGND 459.26
R790 VGND.t805 VGND 459.26
R791 VGND.t657 VGND.t977 455.173
R792 VGND.t869 VGND.t324 455.173
R793 VGND VGND.t319 455.173
R794 VGND.t318 VGND.t770 455.173
R795 VGND VGND.t656 446.743
R796 VGND.t973 VGND 446.743
R797 VGND VGND.t753 446.743
R798 VGND VGND.t604 446.743
R799 VGND.t536 VGND.n1916 446.743
R800 VGND VGND.t315 446.743
R801 VGND.t288 VGND.t459 438.435
R802 VGND VGND.t576 438.315
R803 VGND VGND.t1022 429.885
R804 VGND.t323 VGND.t1012 429.885
R805 VGND.t649 VGND.t517 429.885
R806 VGND.t677 VGND 426.228
R807 VGND.t19 VGND 426.228
R808 VGND.t674 VGND 426.228
R809 VGND VGND.t685 426.228
R810 VGND.n3231 VGND.n3230 406.803
R811 VGND VGND.t486 404.599
R812 VGND VGND.t609 404.599
R813 VGND VGND.t762 404.599
R814 VGND.t369 VGND.t575 404.599
R815 VGND.t1012 VGND.t369 404.599
R816 VGND.t588 VGND.t734 404.599
R817 VGND.t517 VGND.t588 404.599
R818 VGND VGND.t669 404.599
R819 VGND.t975 VGND.t493 404.599
R820 VGND.t109 VGND 404.599
R821 VGND.t530 VGND.n74 403.983
R822 VGND.t507 VGND.t184 387.74
R823 VGND.t764 VGND.t629 387.74
R824 VGND.t730 VGND.t1062 387.74
R825 VGND.t799 VGND.t476 387.74
R826 VGND.t712 VGND.t509 387.74
R827 VGND.n281 VGND 384.901
R828 VGND.t693 VGND 380.899
R829 VGND.t770 VGND.t323 379.31
R830 VGND.t1013 VGND 379.31
R831 VGND.t470 VGND.t190 370.882
R832 VGND VGND.t943 370.37
R833 VGND.t1124 VGND 370.37
R834 VGND VGND.t1098 370.37
R835 VGND.t531 VGND 370.37
R836 VGND.n2030 VGND.t437 361.798
R837 VGND.n415 VGND.n407 354.26
R838 VGND.n415 VGND.n406 354.26
R839 VGND.n418 VGND.n405 354.26
R840 VGND.n418 VGND.n417 354.26
R841 VGND.n478 VGND.n477 354.26
R842 VGND.n477 VGND.n476 354.26
R843 VGND.n445 VGND.n408 354.26
R844 VGND.n466 VGND.n430 354.26
R845 VGND.n466 VGND.n465 354.26
R846 VGND.n435 VGND.n432 354.26
R847 VGND.n436 VGND.n435 354.26
R848 VGND.n443 VGND.n442 354.26
R849 VGND.n444 VGND.n443 354.26
R850 VGND.n2391 VGND.n1004 353.13
R851 VGND.n2391 VGND.n2390 353.13
R852 VGND.n2539 VGND.n947 352
R853 VGND VGND.t288 349.704
R854 VGND VGND.t682 341.574
R855 VGND VGND.t67 341.574
R856 VGND VGND.t448 341.574
R857 VGND.t830 VGND.n3462 337.166
R858 VGND.t633 VGND.t764 337.166
R859 VGND.t1064 VGND.t730 337.166
R860 VGND.t753 VGND 337.166
R861 VGND.n112 VGND.t929 337.166
R862 VGND.t108 VGND.n219 337.166
R863 VGND.n3190 VGND.n187 334.815
R864 VGND.n93 VGND.n86 334.815
R865 VGND.n2390 VGND.n2389 330.486
R866 VGND.t977 VGND.t1015 328.736
R867 VGND.t1115 VGND 328.736
R868 VGND.t604 VGND 328.736
R869 VGND.n3075 VGND.n3074 325.502
R870 VGND.n3064 VGND.n3056 325.502
R871 VGND.t910 VGND 325.171
R872 VGND.n2388 VGND.n1004 324.425
R873 VGND VGND.t270 323.541
R874 VGND.n3462 VGND.t751 320.307
R875 VGND.t315 VGND 320.307
R876 VGND.n112 VGND.t113 320.307
R877 VGND.n219 VGND.t168 320.307
R878 VGND.t313 VGND 311.877
R879 VGND.n3075 VGND.n3069 308.137
R880 VGND.n3065 VGND.n3064 308.137
R881 VGND.n3206 VGND.n3203 304.553
R882 VGND.n3258 VGND.n3256 304.553
R883 VGND.n395 VGND.n394 304.553
R884 VGND.n3244 VGND.n3242 304.553
R885 VGND.n3265 VGND.n3262 304.553
R886 VGND.n3193 VGND.n184 304.553
R887 VGND.n3226 VGND.n179 304.553
R888 VGND.n3390 VGND.n3389 304.553
R889 VGND.t364 VGND 303.449
R890 VGND.t163 VGND 303.449
R891 VGND.t374 VGND.t975 303.449
R892 VGND.n3287 VGND.n3286 299.892
R893 VGND VGND.t830 295.019
R894 VGND.t505 VGND.t396 295.019
R895 VGND VGND.t556 295.019
R896 VGND.t929 VGND 295.019
R897 VGND VGND.t108 295.019
R898 VGND.n1008 VGND.n1005 292.5
R899 VGND.t582 VGND.n1008 292.5
R900 VGND.n1007 VGND.n1006 292.5
R901 VGND.t582 VGND.n1007 292.5
R902 VGND VGND.t992 286.591
R903 VGND.t1038 VGND 286.591
R904 VGND VGND.t574 286.591
R905 VGND.n637 VGND.t993 281.25
R906 VGND.t584 VGND 278.161
R907 VGND.t158 VGND 278.161
R908 VGND.t348 VGND 278.161
R909 VGND.t172 VGND 278.161
R910 VGND.t174 VGND 278.161
R911 VGND.t511 VGND 278.161
R912 VGND.t497 VGND 278.161
R913 VGND.t501 VGND 278.161
R914 VGND.t873 VGND 278.161
R915 VGND.n387 VGND.t154 277.575
R916 VGND.t682 VGND 277.529
R917 VGND.t437 VGND 277.529
R918 VGND.t67 VGND 277.529
R919 VGND.t448 VGND 277.529
R920 VGND.n1168 VGND.t1211 276.531
R921 VGND.n1204 VGND.t1191 276.531
R922 VGND.n747 VGND.t1192 276.531
R923 VGND.t270 VGND 276.274
R924 VGND VGND.t910 276.274
R925 VGND.n533 VGND.t134 275.293
R926 VGND.n2593 VGND.t1116 275.293
R927 VGND.n1845 VGND.t605 275.293
R928 VGND VGND.t667 269.733
R929 VGND.t162 VGND.t178 269.733
R930 VGND.t384 VGND.t739 269.733
R931 VGND.n2105 VGND.t1201 269.488
R932 VGND.n2889 VGND.t1162 269.445
R933 VGND.n395 VGND.n389 266.349
R934 VGND.n3242 VGND.n3239 266.349
R935 VGND.n3265 VGND.n3260 266.349
R936 VGND.n3193 VGND.n182 266.349
R937 VGND.n3222 VGND.n179 266.349
R938 VGND.n3217 VGND.n3203 266.349
R939 VGND.n3390 VGND.n77 266.349
R940 VGND.n3256 VGND.n3255 266.349
R941 VGND.n561 VGND.t1232 265.317
R942 VGND.n819 VGND.t1152 265.317
R943 VGND.n1152 VGND.t1157 265.298
R944 VGND.n732 VGND.t1203 265.298
R945 VGND.t149 VGND.n397 263.652
R946 VGND.n397 VGND.t154 263.652
R947 VGND.n1172 VGND.t1167 262.784
R948 VGND.n1173 VGND.t1151 262.784
R949 VGND.n1175 VGND.t1172 262.784
R950 VGND.n2171 VGND.t1212 262.784
R951 VGND.n548 VGND.t1166 262.784
R952 VGND.n549 VGND.t1131 262.784
R953 VGND.n1185 VGND.t1206 262.784
R954 VGND.n1187 VGND.t1238 262.784
R955 VGND.n1188 VGND.t1146 262.784
R956 VGND.n1197 VGND.t1178 262.784
R957 VGND.n612 VGND.t1183 262.784
R958 VGND.n613 VGND.t1214 262.784
R959 VGND.n2842 VGND.t1187 262.784
R960 VGND.n2844 VGND.t1190 262.784
R961 VGND.n751 VGND.t1207 262.784
R962 VGND.n752 VGND.t1210 262.784
R963 VGND.n754 VGND.t1149 262.784
R964 VGND.n2678 VGND.t1155 262.784
R965 VGND.n1320 VGND.t1171 262.784
R966 VGND.n1321 VGND.t1175 262.784
R967 VGND.n806 VGND.t1150 262.784
R968 VGND.n807 VGND.t1156 262.784
R969 VGND.n1538 VGND.t1138 262.784
R970 VGND.n1540 VGND.t1144 262.784
R971 VGND.n883 VGND.t1237 262.784
R972 VGND.n884 VGND.t1243 262.784
R973 VGND.n1292 VGND.t1222 262.784
R974 VGND.n1837 VGND.t1227 262.784
R975 VGND.n966 VGND.t1202 262.784
R976 VGND.n967 VGND.t1208 262.784
R977 VGND.n2207 VGND.t1229 262.719
R978 VGND.n2269 VGND.t1196 262.719
R979 VGND.n1132 VGND.t1180 262.719
R980 VGND.n1150 VGND.t1230 262.719
R981 VGND.n2241 VGND.t1193 262.719
R982 VGND.n2945 VGND.t1234 262.719
R983 VGND.n2945 VGND.t1164 262.719
R984 VGND.n1220 VGND.t1198 262.719
R985 VGND.n2075 VGND.t1127 262.719
R986 VGND.n2063 VGND.t1160 262.719
R987 VGND.n2898 VGND.t1165 262.719
R988 VGND.n2840 VGND.t1188 262.719
R989 VGND.n2817 VGND.t1173 262.719
R990 VGND.n2714 VGND.t1169 262.719
R991 VGND.n712 VGND.t1128 262.719
R992 VGND.n2754 VGND.t1241 262.719
R993 VGND.n696 VGND.t1168 262.719
R994 VGND.n2784 VGND.t1133 262.719
R995 VGND.n2635 VGND.t1141 262.719
R996 VGND.n1353 VGND.t1221 262.719
R997 VGND.n1502 VGND.t1145 262.719
R998 VGND.n1251 VGND.t1215 262.719
R999 VGND.n2349 VGND.t1181 262.719
R1000 VGND.n497 VGND.t1176 262.719
R1001 VGND.n1104 VGND.t1143 262.719
R1002 VGND.n275 VGND.t1177 262.719
R1003 VGND.t934 VGND 261.303
R1004 VGND VGND.t111 261.303
R1005 VGND.t94 VGND 261.303
R1006 VGND.t1095 VGND.t619 261.303
R1007 VGND.t49 VGND 261.303
R1008 VGND.t580 VGND.t309 261.303
R1009 VGND.t223 VGND 261.303
R1010 VGND.t741 VGND 261.303
R1011 VGND.t97 VGND 261.303
R1012 VGND.t774 VGND 261.303
R1013 VGND.t1000 VGND 261.303
R1014 VGND.t330 VGND 261.303
R1015 VGND VGND.t995 261.303
R1016 VGND VGND.t295 261.303
R1017 VGND.t160 VGND.t76 260.675
R1018 VGND.n1664 VGND.t1220 259.082
R1019 VGND.n1926 VGND.t1135 259.082
R1020 VGND.n2542 VGND.t1216 259.082
R1021 VGND.n1745 VGND.t1186 259.082
R1022 VGND.n2438 VGND.t1163 259.082
R1023 VGND.n2354 VGND.t1235 259.082
R1024 VGND.n1061 VGND.t1223 259.082
R1025 VGND.n3037 VGND.t1242 259.082
R1026 VGND.n245 VGND.t1233 259.082
R1027 VGND.n447 VGND.n446 255.839
R1028 VGND.n446 VGND.n445 253.365
R1029 VGND.t802 VGND 252.875
R1030 VGND.t360 VGND.t625 252.875
R1031 VGND VGND.t580 252.875
R1032 VGND.t609 VGND.t869 252.875
R1033 VGND.t938 VGND 252.875
R1034 VGND.n648 VGND.t3 251
R1035 VGND.n648 VGND.t972 251
R1036 VGND.n2587 VGND.t748 251
R1037 VGND.n916 VGND.t385 251
R1038 VGND.n1286 VGND.t1110 251
R1039 VGND.n2559 VGND.t373 251
R1040 VGND.t943 VGND.t945 248.889
R1041 VGND.t355 VGND.t352 248.889
R1042 VGND.t1121 VGND.t1124 248.889
R1043 VGND.t1098 VGND.t1101 248.889
R1044 VGND.t861 VGND.t863 248.889
R1045 VGND.t528 VGND.t531 248.889
R1046 VGND.n1460 VGND.t593 245.82
R1047 VGND.n1704 VGND.t767 245.82
R1048 VGND.n1599 VGND.t601 245.82
R1049 VGND.n1914 VGND.t537 245.82
R1050 VGND VGND.t702 244.445
R1051 VGND.t88 VGND 244.445
R1052 VGND VGND.t273 244.445
R1053 VGND.t267 VGND 244.445
R1054 VGND.t627 VGND.t962 244.445
R1055 VGND.t416 VGND 244.445
R1056 VGND.t22 VGND 244.445
R1057 VGND VGND.t454 244.445
R1058 VGND.n663 VGND.t339 243.028
R1059 VGND.n663 VGND.t896 243.028
R1060 VGND.n1631 VGND.t120 243.028
R1061 VGND.n911 VGND.t955 243.028
R1062 VGND.n1242 VGND.t1120 243.028
R1063 VGND.n1882 VGND.t481 243.028
R1064 VGND.n1447 VGND.t618 242.067
R1065 VGND.n1556 VGND.t1069 242.067
R1066 VGND VGND.t202 241.573
R1067 VGND.n1495 VGND.t595 240.948
R1068 VGND.n1642 VGND.t546 240.948
R1069 VGND.n16 VGND.t935 240.575
R1070 VGND.n110 VGND.t996 240.575
R1071 VGND.n1393 VGND.t1096 238.675
R1072 VGND.n1678 VGND.t15 238.675
R1073 VGND.n875 VGND.t13 238.675
R1074 VGND.n2543 VGND.t471 238.675
R1075 VGND.n803 VGND.t1025 238.44
R1076 VGND VGND.t16 238.202
R1077 VGND.n7 VGND.t1055 237.327
R1078 VGND.n3098 VGND.t296 237.327
R1079 VGND.n3088 VGND.t1009 237.327
R1080 VGND.n3320 VGND.t888 237.327
R1081 VGND.n1438 VGND.t1106 237.327
R1082 VGND.n1515 VGND.t607 237.327
R1083 VGND.t653 VGND.t1070 236.016
R1084 VGND.t982 VGND 236.016
R1085 VGND.t951 VGND.t327 236.016
R1086 VGND.n2816 VGND.t565 235.607
R1087 VGND.n1971 VGND.n1970 234.667
R1088 VGND.n1624 VGND.t399 230.977
R1089 VGND.n1866 VGND.t771 230.977
R1090 VGND.n621 VGND.t131 229.833
R1091 VGND.n1612 VGND.n1611 228.294
R1092 VGND.n943 VGND.n942 228.294
R1093 VGND.t788 VGND 228.09
R1094 VGND.t1042 VGND.t55 227.587
R1095 VGND.t1080 VGND.t974 227.587
R1096 VGND.t486 VGND.t1074 227.587
R1097 VGND VGND.t484 227.587
R1098 VGND.n2043 VGND.t47 227.256
R1099 VGND.n1431 VGND.t668 226.708
R1100 VGND.n3144 VGND.t797 225.427
R1101 VGND.n3169 VGND.t718 225.427
R1102 VGND.n3089 VGND.t455 225.427
R1103 VGND.n3108 VGND.t713 225.427
R1104 VGND.n1014 VGND.n1006 225.13
R1105 VGND.n1009 VGND.n1006 225.13
R1106 VGND.t445 VGND.t181 224.931
R1107 VGND.n1715 VGND.t1139 224.196
R1108 VGND.n1124 VGND.t1137 224.102
R1109 VGND.n717 VGND.t1197 224.102
R1110 VGND.n2791 VGND.t42 223.282
R1111 VGND.n1449 VGND.n1413 222.691
R1112 VGND VGND.n3190 222.222
R1113 VGND.n208 VGND 222.222
R1114 VGND VGND.n86 222.222
R1115 VGND.n94 VGND 222.222
R1116 VGND.n690 VGND.t1132 221.972
R1117 VGND.n845 VGND.n843 221.804
R1118 VGND.t152 VGND.t150 221.451
R1119 VGND.n839 VGND.t1218 220.952
R1120 VGND.n840 VGND.t1224 220.952
R1121 VGND.n692 VGND.t221 219.972
R1122 VGND.n628 VGND.n626 218.506
R1123 VGND.n628 VGND.n627 218.506
R1124 VGND.n1709 VGND.n1551 218.506
R1125 VGND.n1656 VGND.n1585 218.506
R1126 VGND.n918 VGND.n853 218.506
R1127 VGND.n1853 VGND.n1288 218.506
R1128 VGND.n1891 VGND.n1890 218.506
R1129 VGND.n934 VGND.n933 218.506
R1130 VGND.n57 VGND.t1184 218.308
R1131 VGND.n3436 VGND.t1205 218.308
R1132 VGND.n25 VGND.t1240 218.308
R1133 VGND.n9 VGND.t1185 218.308
R1134 VGND.n212 VGND.t1159 218.308
R1135 VGND.n3167 VGND.t1154 218.308
R1136 VGND.n221 VGND.t1147 218.308
R1137 VGND.n3107 VGND.t1213 218.308
R1138 VGND.n3302 VGND.t1209 218.308
R1139 VGND.n98 VGND.t1161 218.308
R1140 VGND.n3322 VGND.t1142 218.308
R1141 VGND.n3346 VGND.t1195 218.308
R1142 VGND.n555 VGND.t1129 218.308
R1143 VGND.n619 VGND.t1179 218.308
R1144 VGND.n2883 VGND.t1130 218.308
R1145 VGND.n813 VGND.t1148 218.308
R1146 VGND.n1440 VGND.t1136 218.308
R1147 VGND.n1844 VGND.t1219 218.308
R1148 VGND.n1811 VGND.t1239 218.308
R1149 VGND.n996 VGND.t1134 218.308
R1150 VGND.n1604 VGND.n1603 218.13
R1151 VGND.n1133 VGND.t903 217.977
R1152 VGND.n1123 VGND.t431 217.977
R1153 VGND.n2761 VGND.t74 217.977
R1154 VGND.n2740 VGND.t209 217.977
R1155 VGND.n2217 VGND.t795 217.953
R1156 VGND.n730 VGND.t825 217.953
R1157 VGND.n2261 VGND.t261 217.892
R1158 VGND.n2759 VGND.t27 217.892
R1159 VGND.n212 VGND.t798 217.78
R1160 VGND.n3167 VGND.t719 217.78
R1161 VGND.n221 VGND.t456 217.78
R1162 VGND.n3107 VGND.t714 217.78
R1163 VGND.n1340 VGND.t249 216.933
R1164 VGND.n1125 VGND.t89 216.589
R1165 VGND.n718 VGND.t274 216.589
R1166 VGND.n2802 VGND.t803 216.579
R1167 VGND.n1549 VGND.t710 215.992
R1168 VGND.n1124 VGND.t90 214.487
R1169 VGND.n717 VGND.t275 214.487
R1170 VGND.n8 VGND.t704 214.456
R1171 VGND.n3 VGND.t703 214.456
R1172 VGND.n58 VGND.t701 214.456
R1173 VGND.n42 VGND.t700 214.456
R1174 VGND.n3437 VGND.t241 214.456
R1175 VGND.n40 VGND.t240 214.456
R1176 VGND.n26 VGND.t186 214.456
R1177 VGND.n32 VGND.t185 214.456
R1178 VGND.n81 VGND.t201 214.456
R1179 VGND.n3305 VGND.t200 214.456
R1180 VGND.n99 VGND.t807 214.456
R1181 VGND.n97 VGND.t806 214.456
R1182 VGND.n3345 VGND.t801 214.456
R1183 VGND.n3341 VGND.t800 214.456
R1184 VGND.n3323 VGND.t24 214.456
R1185 VGND.n115 VGND.t23 214.456
R1186 VGND.n554 VGND.t909 214.456
R1187 VGND.n554 VGND.t899 214.456
R1188 VGND.n546 VGND.t898 214.456
R1189 VGND.n525 VGND.t908 214.456
R1190 VGND.n521 VGND.t819 214.456
R1191 VGND.n2227 VGND.t818 214.456
R1192 VGND.n521 VGND.t812 214.456
R1193 VGND.n2227 VGND.t811 214.456
R1194 VGND.n2226 VGND.t54 214.456
R1195 VGND.n1151 VGND.t904 214.456
R1196 VGND.n1140 VGND.t53 214.456
R1197 VGND.n2263 VGND.t432 214.456
R1198 VGND.n2277 VGND.t260 214.456
R1199 VGND.n1157 VGND.t794 214.456
R1200 VGND.n2214 VGND.t36 214.456
R1201 VGND.n1158 VGND.t213 214.456
R1202 VGND.n2185 VGND.t35 214.456
R1203 VGND.n2178 VGND.t698 214.456
R1204 VGND.n1171 VGND.t212 214.456
R1205 VGND.n1171 VGND.t697 214.456
R1206 VGND.n1172 VGND.t827 214.456
R1207 VGND.n1172 VGND.t826 214.456
R1208 VGND.n1173 VGND.t817 214.456
R1209 VGND.n1173 VGND.t816 214.456
R1210 VGND.n1175 VGND.t255 214.456
R1211 VGND.n1175 VGND.t254 214.456
R1212 VGND.n2171 VGND.t238 214.456
R1213 VGND.n2171 VGND.t237 214.456
R1214 VGND.n548 VGND.t235 214.456
R1215 VGND.n548 VGND.t234 214.456
R1216 VGND.n549 VGND.t814 214.456
R1217 VGND.n549 VGND.t813 214.456
R1218 VGND.n2892 VGND.t822 214.456
R1219 VGND.n577 VGND.t44 214.456
R1220 VGND.n2064 VGND.t821 214.456
R1221 VGND.n576 VGND.t39 214.456
R1222 VGND.n2069 VGND.t48 214.456
R1223 VGND.n2060 VGND.t38 214.456
R1224 VGND.n2082 VGND.t424 214.456
R1225 VGND.n2099 VGND.t453 214.456
R1226 VGND.n2039 VGND.t423 214.456
R1227 VGND.n2117 VGND.t452 214.456
R1228 VGND.n1221 VGND.t781 214.456
R1229 VGND.n1216 VGND.t415 214.456
R1230 VGND.n2131 VGND.t780 214.456
R1231 VGND.n1200 VGND.t278 214.456
R1232 VGND.n1198 VGND.t414 214.456
R1233 VGND.n1198 VGND.t277 214.456
R1234 VGND.n1185 VGND.t195 214.456
R1235 VGND.n1185 VGND.t194 214.456
R1236 VGND.n1187 VGND.t429 214.456
R1237 VGND.n1187 VGND.t428 214.456
R1238 VGND.n1188 VGND.t692 214.456
R1239 VGND.n1188 VGND.t691 214.456
R1240 VGND.n1197 VGND.t81 214.456
R1241 VGND.n1197 VGND.t80 214.456
R1242 VGND.n2882 VGND.t66 214.456
R1243 VGND.n582 VGND.t65 214.456
R1244 VGND.n2882 VGND.t45 214.456
R1245 VGND.n618 VGND.t266 214.456
R1246 VGND.n610 VGND.t265 214.456
R1247 VGND.n612 VGND.t280 214.456
R1248 VGND.n612 VGND.t279 214.456
R1249 VGND.n613 VGND.t253 214.456
R1250 VGND.n613 VGND.t252 214.456
R1251 VGND.n2785 VGND.t75 214.456
R1252 VGND.n2764 VGND.t41 214.456
R1253 VGND.n690 VGND.t222 214.456
R1254 VGND.n680 VGND.t804 214.456
R1255 VGND.n2829 VGND.t246 214.456
R1256 VGND.n2841 VGND.t690 214.456
R1257 VGND.n2836 VGND.t689 214.456
R1258 VGND.n2841 VGND.t247 214.456
R1259 VGND.n2842 VGND.t708 214.456
R1260 VGND.n2842 VGND.t707 214.456
R1261 VGND.n2844 VGND.t258 214.456
R1262 VGND.n2844 VGND.t257 214.456
R1263 VGND.n710 VGND.t210 214.456
R1264 VGND.n2742 VGND.t26 214.456
R1265 VGND.n736 VGND.t824 214.456
R1266 VGND.n2721 VGND.t784 214.456
R1267 VGND.n737 VGND.t787 214.456
R1268 VGND.n2692 VGND.t783 214.456
R1269 VGND.n2685 VGND.t283 214.456
R1270 VGND.n750 VGND.t786 214.456
R1271 VGND.n750 VGND.t282 214.456
R1272 VGND.n751 VGND.t244 214.456
R1273 VGND.n751 VGND.t243 214.456
R1274 VGND.n752 VGND.t436 214.456
R1275 VGND.n752 VGND.t435 214.456
R1276 VGND.n754 VGND.t906 214.456
R1277 VGND.n754 VGND.t905 214.456
R1278 VGND.n2678 VGND.t87 214.456
R1279 VGND.n2678 VGND.t86 214.456
R1280 VGND.n1320 VGND.t72 214.456
R1281 VGND.n1320 VGND.t71 214.456
R1282 VGND.n1321 VGND.t809 214.456
R1283 VGND.n1321 VGND.t808 214.456
R1284 VGND.n1439 VGND.t216 214.456
R1285 VGND.n1418 VGND.t215 214.456
R1286 VGND.n2628 VGND.t57 214.456
R1287 VGND.n1429 VGND.t56 214.456
R1288 VGND.n781 VGND.t83 214.456
R1289 VGND.n812 VGND.t30 214.456
R1290 VGND.n804 VGND.t29 214.456
R1291 VGND.n812 VGND.t84 214.456
R1292 VGND.n806 VGND.t901 214.456
R1293 VGND.n806 VGND.t900 214.456
R1294 VGND.n807 VGND.t673 214.456
R1295 VGND.n807 VGND.t672 214.456
R1296 VGND.n1370 VGND.t232 214.456
R1297 VGND.n1516 VGND.t231 214.456
R1298 VGND.n1361 VGND.t269 214.456
R1299 VGND.n1313 VGND.t268 214.456
R1300 VGND.n1346 VGND.t250 214.456
R1301 VGND.n879 VGND.t418 214.456
R1302 VGND.n877 VGND.t417 214.456
R1303 VGND.n1663 VGND.t198 214.456
R1304 VGND.n1578 VGND.t197 214.456
R1305 VGND.n1700 VGND.t711 214.456
R1306 VGND.n1715 VGND.t51 214.456
R1307 VGND.n1541 VGND.t50 214.456
R1308 VGND.n1538 VGND.t227 214.456
R1309 VGND.n1538 VGND.t226 214.456
R1310 VGND.n1540 VGND.t60 214.456
R1311 VGND.n1540 VGND.t59 214.456
R1312 VGND.n839 VGND.t263 214.456
R1313 VGND.n839 VGND.t262 214.456
R1314 VGND.n840 VGND.t207 214.456
R1315 VGND.n840 VGND.t206 214.456
R1316 VGND.n883 VGND.t434 214.456
R1317 VGND.n883 VGND.t433 214.456
R1318 VGND.n884 VGND.t33 214.456
R1319 VGND.n884 VGND.t32 214.456
R1320 VGND.n971 VGND.t427 214.456
R1321 VGND.n963 VGND.t426 214.456
R1322 VGND.n971 VGND.t412 214.456
R1323 VGND.n960 VGND.t411 214.456
R1324 VGND.n2541 VGND.t192 214.456
R1325 VGND.n944 VGND.t191 214.456
R1326 VGND.n1925 VGND.t63 214.456
R1327 VGND.n1918 VGND.t62 214.456
R1328 VGND.n1945 VGND.t189 214.456
R1329 VGND.n1968 VGND.t188 214.456
R1330 VGND.n1843 VGND.t225 214.456
R1331 VGND.n1290 VGND.t224 214.456
R1332 VGND.n1292 VGND.t229 214.456
R1333 VGND.n1292 VGND.t228 214.456
R1334 VGND.n1837 VGND.t219 214.456
R1335 VGND.n1837 VGND.t218 214.456
R1336 VGND.n966 VGND.t441 214.456
R1337 VGND.n966 VGND.t440 214.456
R1338 VGND.n967 VGND.t421 214.456
R1339 VGND.n967 VGND.t420 214.456
R1340 VGND.n2437 VGND.t78 214.456
R1341 VGND.n2435 VGND.t77 214.456
R1342 VGND.n2417 VGND.t450 214.456
R1343 VGND.n2416 VGND.t449 214.456
R1344 VGND.n2474 VGND.t695 214.456
R1345 VGND.n2397 VGND.t694 214.456
R1346 VGND.n997 VGND.t18 214.456
R1347 VGND.n2509 VGND.t17 214.456
R1348 VGND.n1996 VGND.t69 214.456
R1349 VGND.n1995 VGND.t68 214.456
R1350 VGND.n1227 VGND.t439 214.456
R1351 VGND.n1225 VGND.t438 214.456
R1352 VGND.n1781 VGND.t684 214.456
R1353 VGND.n1780 VGND.t683 214.456
R1354 VGND.n1810 VGND.t204 214.456
R1355 VGND.n1763 VGND.t203 214.456
R1356 VGND.n1741 VGND.t790 214.456
R1357 VGND.n1746 VGND.t789 214.456
R1358 VGND.n240 VGND.t447 214.456
R1359 VGND.n246 VGND.t446 214.456
R1360 VGND.n3036 VGND.t183 214.456
R1361 VGND.n3039 VGND.t182 214.456
R1362 VGND.n258 VGND.t271 214.456
R1363 VGND.n3021 VGND.t272 214.456
R1364 VGND.n277 VGND.t679 214.456
R1365 VGND.n271 VGND.t678 214.456
R1366 VGND.n1060 VGND.t409 214.456
R1367 VGND.n1059 VGND.t408 214.456
R1368 VGND.n1098 VGND.t21 214.456
R1369 VGND.n1075 VGND.t20 214.456
R1370 VGND.n495 VGND.t676 214.456
R1371 VGND.n1080 VGND.t675 214.456
R1372 VGND.n1039 VGND.t911 214.456
R1373 VGND.n1032 VGND.t912 214.456
R1374 VGND.n2350 VGND.t687 214.456
R1375 VGND.n2338 VGND.t686 214.456
R1376 VGND.n2353 VGND.t444 214.456
R1377 VGND.n2351 VGND.t443 214.456
R1378 VGND.n1009 VGND.n1005 214.409
R1379 VGND.n1015 VGND.n1014 213.911
R1380 VGND.n3401 VGND.n3400 212.78
R1381 VGND.n1631 VGND.n1608 212.317
R1382 VGND.t311 VGND.t284 211.237
R1383 VGND.t853 VGND 210.728
R1384 VGND.n3287 VGND.t530 209.996
R1385 VGND.n2601 VGND.n836 207.965
R1386 VGND.n937 VGND.n936 207.965
R1387 VGND.n1373 VGND.n1372 206.909
R1388 VGND.n3286 VGND.n3285 206.876
R1389 VGND.n1671 VGND.n1670 205.971
R1390 VGND.n1466 VGND.n1396 205.899
R1391 VGND.n1469 VGND.n1468 205.899
R1392 VGND.n1398 VGND.n1397 205.481
R1393 VGND.n1572 VGND.n1571 205.481
R1394 VGND.n2626 VGND.n2625 205.385
R1395 VGND.n1449 VGND.n1412 204.692
R1396 VGND.n1476 VGND.n1475 204.692
R1397 VGND.n48 VGND.n44 204.457
R1398 VGND.n3310 VGND.n3309 204.457
R1399 VGND.n1939 VGND.n1937 204.457
R1400 VGND.n1939 VGND.n1938 204.457
R1401 VGND.n1921 VGND.n1919 204.457
R1402 VGND.n2823 VGND.n2822 204.201
R1403 VGND.n1249 VGND.n1248 204.201
R1404 VGND.n1263 VGND.n1262 204.201
R1405 VGND.n1425 VGND.n1422 202.724
R1406 VGND.n772 VGND.n771 202.724
R1407 VGND.n1484 VGND.n1387 202.724
R1408 VGND.n1655 VGND.n1586 202.724
R1409 VGND.n1598 VGND.n1597 202.724
R1410 VGND VGND.t1092 202.299
R1411 VGND.t326 VGND.t968 202.299
R1412 VGND.t855 VGND.t950 202.299
R1413 VGND.t372 VGND.t301 202.299
R1414 VGND.n780 VGND.n779 201.458
R1415 VGND.n1575 VGND.n1574 201.458
R1416 VGND.n1459 VGND.n1400 201.129
R1417 VGND.n2618 VGND.n784 201.129
R1418 VGND.n2620 VGND.n783 201.129
R1419 VGND.n1680 VGND.n1573 201.129
R1420 VGND.n2084 VGND.n2083 200.692
R1421 VGND.n1702 VGND.n1701 200.692
R1422 VGND.n2479 VGND.n2478 200.692
R1423 VGND.n3023 VGND.n3022 200.692
R1424 VGND.n2327 VGND.n2326 200.692
R1425 VGND.n2599 VGND.n838 200.516
R1426 VGND.n1285 VGND.n1284 200.516
R1427 VGND.n793 VGND.n792 200.508
R1428 VGND.n774 VGND.n773 200.508
R1429 VGND.n2634 VGND.n776 200.508
R1430 VGND.n1392 VGND.n1391 200.508
R1431 VGND.n1560 VGND.n1559 200.508
R1432 VGND.n1665 VGND.n1580 200.508
R1433 VGND.n1583 VGND.n1582 200.508
R1434 VGND.n3460 VGND.n15 200.231
R1435 VGND.n3452 VGND.n21 200.231
R1436 VGND.n3329 VGND.n3328 200.231
R1437 VGND.n108 VGND.n107 200.231
R1438 VGND.n1446 VGND.n1416 200.231
R1439 VGND.n845 VGND.n844 200.127
R1440 VGND.n1851 VGND.n1850 200.127
R1441 VGND.n30 VGND.n24 200.105
R1442 VGND.n3109 VGND.n3106 200.105
R1443 VGND.n3138 VGND.n214 200.105
R1444 VGND.n3348 VGND.n3343 200.105
R1445 VGND.n599 VGND.n597 199.739
R1446 VGND.n599 VGND.n598 199.739
R1447 VGND.n1494 VGND.n1374 199.739
R1448 VGND.n1629 VGND.n1610 199.739
R1449 VGND.n1272 VGND.n1271 199.739
R1450 VGND.n1823 VGND.n1758 199.739
R1451 VGND.n1818 VGND.n1762 199.739
R1452 VGND.n1805 VGND.n1767 199.739
R1453 VGND.n1784 VGND.n1783 199.739
R1454 VGND.n1992 VGND.n1991 199.739
R1455 VGND.n2519 VGND.n990 199.739
R1456 VGND.n999 VGND.n998 199.739
R1457 VGND.n2413 VGND.n2412 199.739
R1458 VGND.n2421 VGND.n2420 199.739
R1459 VGND.n2444 VGND.n2434 199.739
R1460 VGND.n1031 VGND.n1030 199.739
R1461 VGND.n682 VGND.n681 199.662
R1462 VGND.n657 VGND.n655 199.53
R1463 VGND.n657 VGND.n656 199.53
R1464 VGND.n1470 VGND.n1467 199.53
R1465 VGND.n1637 VGND.n1605 199.53
R1466 VGND.n917 VGND.n854 199.53
R1467 VGND.n1241 VGND.n1240 199.53
R1468 VGND.n1865 VGND.n1864 199.53
R1469 VGND.n940 VGND.n939 199.53
R1470 VGND.t956 VGND 198.519
R1471 VGND.t945 VGND 198.519
R1472 VGND VGND.t355 198.519
R1473 VGND VGND.t1121 198.519
R1474 VGND.t378 VGND 198.519
R1475 VGND.t1101 VGND 198.519
R1476 VGND VGND.t861 198.519
R1477 VGND VGND.t528 198.519
R1478 VGND VGND.n38 197.724
R1479 VGND.n3101 VGND.n3100 197.476
R1480 VGND.n3095 VGND.n218 197.476
R1481 VGND.n1359 VGND.n1307 197.476
R1482 VGND.n536 VGND.n535 196.831
R1483 VGND.n1694 VGND.n1558 196.589
R1484 VGND.n909 VGND.n859 196.589
R1485 VGND.n1352 VGND.n1310 196.442
R1486 VGND.n1483 VGND.n1388 196.442
R1487 VGND.n1673 VGND.n1577 196.442
R1488 VGND.n861 VGND.n860 196.442
R1489 VGND.n890 VGND.n878 196.442
R1490 VGND.n308 VGND.n307 195
R1491 VGND.n309 VGND.n308 195
R1492 VGND.n305 VGND.n304 195
R1493 VGND.n304 VGND.n303 195
R1494 VGND.n313 VGND.n312 195
R1495 VGND.n312 VGND.n311 195
R1496 VGND.n316 VGND.n315 195
R1497 VGND.n317 VGND.n316 195
R1498 VGND.n320 VGND.n319 195
R1499 VGND.n321 VGND.n320 195
R1500 VGND.n325 VGND.n324 195
R1501 VGND.n324 VGND.n323 195
R1502 VGND.n367 VGND.n366 195
R1503 VGND.n368 VGND.n367 195
R1504 VGND.n364 VGND.n363 195
R1505 VGND.n363 VGND.n362 195
R1506 VGND.n339 VGND.n338 195
R1507 VGND.n340 VGND.n339 195
R1508 VGND.n336 VGND.n335 195
R1509 VGND.n335 VGND.n334 195
R1510 VGND.n391 VGND.n282 195
R1511 VGND.n282 VGND.n281 195
R1512 VGND.n3244 VGND.n3243 195
R1513 VGND.n3243 VGND.n3232 195
R1514 VGND.n3248 VGND.n3247 195
R1515 VGND.n3249 VGND.n3248 195
R1516 VGND.n3264 VGND.n3262 195
R1517 VGND.n3264 VGND.n3233 195
R1518 VGND.n3263 VGND.n3261 195
R1519 VGND.n3263 VGND.n3251 195
R1520 VGND.n3206 VGND.n3205 195
R1521 VGND.n3205 VGND.n174 195
R1522 VGND.n3216 VGND.n3215 195
R1523 VGND.n3215 VGND.n3214 195
R1524 VGND.n186 VGND.n184 195
R1525 VGND.n186 VGND.n176 195
R1526 VGND.n185 VGND.n183 195
R1527 VGND.n3192 VGND.n185 195
R1528 VGND.n3227 VGND.n3226 195
R1529 VGND.n3228 VGND.n3227 195
R1530 VGND.n3210 VGND.n180 195
R1531 VGND.n3211 VGND.n3210 195
R1532 VGND.n3389 VGND.n76 195
R1533 VGND.n3286 VGND.n76 195
R1534 VGND.n202 VGND.n197 195
R1535 VGND.n197 VGND.n187 195
R1536 VGND.n204 VGND.n199 195
R1537 VGND.n199 VGND.n198 195
R1538 VGND.n3258 VGND.n3257 195
R1539 VGND.n3257 VGND.n3234 195
R1540 VGND.n3278 VGND.n3277 195
R1541 VGND.n3279 VGND.n3278 195
R1542 VGND.n3386 VGND.n75 195
R1543 VGND.n93 VGND.n75 195
R1544 VGND.n355 VGND.n354 195
R1545 VGND.n354 VGND.n283 195
R1546 VGND.n358 VGND.n357 195
R1547 VGND.n359 VGND.n358 195
R1548 VGND.n383 VGND.n382 195
R1549 VGND.n384 VGND.n383 195
R1550 VGND.n380 VGND.n379 195
R1551 VGND.n379 VGND.n378 195
R1552 VGND.n394 VGND.n388 195
R1553 VGND.n388 VGND.n387 195
R1554 VGND.n3074 VGND.n226 195
R1555 VGND.n226 VGND.t298 195
R1556 VGND.n3070 VGND.n225 195
R1557 VGND.n3060 VGND.n3056 195
R1558 VGND.t662 VGND.n3060 195
R1559 VGND.n3057 VGND.n3055 195
R1560 VGND.t662 VGND.n3057 195
R1561 VGND.n398 VGND.t149 194.406
R1562 VGND.t913 VGND.t386 193.87
R1563 VGND.t367 VGND.t1016 193.87
R1564 VGND.n2057 VGND.n2055 190.399
R1565 VGND.n1555 VGND.n1552 190.399
R1566 VGND.n2477 VGND.n2476 190.399
R1567 VGND.n263 VGND.n261 190.399
R1568 VGND.n2325 VGND.n2324 190.399
R1569 VGND.n1970 VGND.n1244 189.268
R1570 VGND.n947 VGND.n946 189.201
R1571 VGND.n3071 VGND.n225 188.968
R1572 VGND.t515 VGND.t954 185.441
R1573 VGND.t650 VGND.t1000 185.441
R1574 VGND.t1004 VGND.n3083 185.441
R1575 VGND.n438 VGND.t699 179.556
R1576 VGND.t523 VGND 177.529
R1577 VGND.t915 VGND 177.529
R1578 VGND.t145 VGND 177.529
R1579 VGND.t124 VGND 177.529
R1580 VGND.t930 VGND 177.529
R1581 VGND.t1058 VGND 177.012
R1582 VGND.t737 VGND.t569 177.012
R1583 VGND.t1109 VGND.t332 177.012
R1584 VGND.t322 VGND.t97 177.012
R1585 VGND VGND.t141 177.012
R1586 VGND VGND.t841 177.012
R1587 VGND.t150 VGND 176.633
R1588 VGND.n398 VGND 176.633
R1589 VGND.n3072 VGND.n3071 174.41
R1590 VGND.t202 VGND 174.157
R1591 VGND.t16 VGND 174.157
R1592 VGND.t611 VGND.t963 168.583
R1593 VGND.t484 VGND.t982 168.583
R1594 VGND.n387 VGND.n386 163.297
R1595 VGND.n3429 VGND.t991 162.471
R1596 VGND.n3424 VGND.t834 162.471
R1597 VGND.n3420 VGND.t343 162.471
R1598 VGND.n3415 VGND.t153 162.471
R1599 VGND.n3455 VGND.t290 162.471
R1600 VGND.n3376 VGND.t381 162.471
R1601 VGND.n3371 VGND.t1099 162.471
R1602 VGND.n3367 VGND.t864 162.471
R1603 VGND.n3362 VGND.t532 162.471
R1604 VGND.n3334 VGND.t167 162.471
R1605 VGND.n2986 VGND 162.179
R1606 VGND.n127 VGND.t880 162.022
R1607 VGND.n132 VGND.t337 162.022
R1608 VGND.n137 VGND.t349 162.022
R1609 VGND.n142 VGND.t868 162.022
R1610 VGND.n147 VGND.t865 162.022
R1611 VGND.n152 VGND.t512 162.022
R1612 VGND.n157 VGND.t777 162.022
R1613 VGND.n162 VGND.t775 162.022
R1614 VGND.n167 VGND.t876 162.022
R1615 VGND.n131 VGND.t105 162.022
R1616 VGND.n136 VGND.t157 162.022
R1617 VGND.n141 VGND.t466 162.022
R1618 VGND.n146 VGND.t171 162.022
R1619 VGND.n151 VGND.t177 162.022
R1620 VGND.n156 VGND.t535 162.022
R1621 VGND.n161 VGND.t500 162.022
R1622 VGND.n166 VGND.t504 162.022
R1623 VGND.n171 VGND.t872 162.022
R1624 VGND.n3460 VGND.t1061 160.046
R1625 VGND.n3452 VGND.t1057 160.046
R1626 VGND.n3329 VGND.t716 160.046
R1627 VGND.n108 VGND.t886 160.046
R1628 VGND.n127 VGND.t585 160.017
R1629 VGND.n132 VGND.t159 160.017
R1630 VGND.n137 VGND.t465 160.017
R1631 VGND.n142 VGND.t173 160.017
R1632 VGND.n147 VGND.t175 160.017
R1633 VGND.n152 VGND.t534 160.017
R1634 VGND.n157 VGND.t498 160.017
R1635 VGND.n162 VGND.t502 160.017
R1636 VGND.n167 VGND.t874 160.017
R1637 VGND.n60 VGND.t988 160.017
R1638 VGND.n3422 VGND.t837 160.017
R1639 VGND.n3411 VGND.t346 160.017
R1640 VGND.n39 VGND.t151 160.017
R1641 VGND.n3453 VGND.t292 160.017
R1642 VGND.n22 VGND.t1 160.017
R1643 VGND.n83 VGND.t379 160.017
R1644 VGND.n3369 VGND.t1102 160.017
R1645 VGND.n89 VGND.t862 160.017
R1646 VGND.n3360 VGND.t529 160.017
R1647 VGND.n3336 VGND.t116 160.017
R1648 VGND.n3353 VGND.t840 160.017
R1649 VGND.n131 VGND.t879 160.017
R1650 VGND.n136 VGND.t336 160.017
R1651 VGND.n141 VGND.t351 160.017
R1652 VGND.n146 VGND.t867 160.017
R1653 VGND.n151 VGND.t866 160.017
R1654 VGND.n156 VGND.t514 160.017
R1655 VGND.n161 VGND.t778 160.017
R1656 VGND.n166 VGND.t776 160.017
R1657 VGND.n171 VGND.t875 160.017
R1658 VGND.n16 VGND.t661 158.534
R1659 VGND.n110 VGND.t792 158.534
R1660 VGND.t10 VGND.n2030 157.304
R1661 VGND.n2395 VGND.t135 157.304
R1662 VGND.n3146 VGND.t960 157.291
R1663 VGND.n3148 VGND.t944 157.291
R1664 VGND.n191 VGND.t353 157.291
R1665 VGND.n192 VGND.t1125 157.291
R1666 VGND.n3097 VGND.t681 157.291
R1667 VGND.n3124 VGND.t918 157.291
R1668 VGND.n3117 VGND.t140 157.291
R1669 VGND.n3156 VGND.t957 155.286
R1670 VGND.n3150 VGND.t946 155.286
R1671 VGND.n3184 VGND.t356 155.286
R1672 VGND.n3178 VGND.t1122 155.286
R1673 VGND.n3129 VGND.t706 155.286
R1674 VGND.n3122 VGND.t998 155.286
R1675 VGND.n3115 VGND.t884 155.286
R1676 VGND.n904 VGND.t856 154.131
R1677 VGND.n2814 VGND.t9 152.381
R1678 VGND.n874 VGND.t892 152.381
R1679 VGND.n882 VGND.t939 152.381
R1680 VGND.n2085 VGND.n2084 152
R1681 VGND.n1703 VGND.n1702 152
R1682 VGND.n2478 VGND.n2411 152
R1683 VGND.n2326 VGND.n1034 152
R1684 VGND.n3024 VGND.n3023 152
R1685 VGND.n2803 VGND.t287 150.101
R1686 VGND.n882 VGND.t858 150.101
R1687 VGND.n2987 VGND.t407 149.954
R1688 VGND VGND.n3403 144.951
R1689 VGND.n848 VGND.t969 144.886
R1690 VGND.n1858 VGND.t333 144.886
R1691 VGND.t482 VGND.t596 143.296
R1692 VGND VGND.n842 143.296
R1693 VGND.t61 VGND 143.296
R1694 VGND.n474 VGND.n473 139.727
R1695 VGND.t662 VGND.n223 137.912
R1696 VGND.n3062 VGND.t662 137.912
R1697 VGND.t123 VGND 135.415
R1698 VGND.t631 VGND.t765 134.867
R1699 VGND.t1111 VGND.t743 134.867
R1700 VGND.t549 VGND.t608 134.867
R1701 VGND.t403 VGND.t316 134.867
R1702 VGND.n71 VGND.t376 133.507
R1703 VGND.t964 VGND.t615 126.438
R1704 VGND.n522 VGND.t844 124.688
R1705 VGND.n431 VGND.n430 123.882
R1706 VGND.t76 VGND 122.472
R1707 VGND.n879 VGND.t1231 121.927
R1708 VGND.n2417 VGND.t1228 121.927
R1709 VGND.n1996 VGND.t1158 121.927
R1710 VGND.n1227 VGND.t1225 121.927
R1711 VGND.n1781 VGND.t1170 121.927
R1712 VGND VGND.t1126 121.481
R1713 VGND VGND.t527 121.481
R1714 VGND.n3079 VGND.n3078 120.984
R1715 VGND.n3077 VGND.n3076 118.285
R1716 VGND.t596 VGND 118.008
R1717 VGND.t1020 VGND.t82 118.008
R1718 VGND.t1072 VGND.t655 118.008
R1719 VGND.t574 VGND.t488 118.008
R1720 VGND.n452 VGND.n448 117.001
R1721 VGND.n452 VGND.t467 117.001
R1722 VGND.n449 VGND.n447 117.001
R1723 VGND.n449 VGND.t467 117.001
R1724 VGND.n480 VGND.n412 117.001
R1725 VGND.n480 VGND.t551 117.001
R1726 VGND.n410 VGND.n408 117.001
R1727 VGND.t551 VGND.n410 117.001
R1728 VGND.n444 VGND.n440 117.001
R1729 VGND.n440 VGND.t643 117.001
R1730 VGND.n442 VGND.n439 117.001
R1731 VGND.t643 VGND.n439 117.001
R1732 VGND.n414 VGND.n407 117.001
R1733 VGND.n414 VGND.t371 117.001
R1734 VGND.n413 VGND.n406 117.001
R1735 VGND.n413 VGND.t371 117.001
R1736 VGND.n437 VGND.n436 117.001
R1737 VGND.t643 VGND.n437 117.001
R1738 VGND.n434 VGND.n432 117.001
R1739 VGND.t643 VGND.n434 117.001
R1740 VGND.n405 VGND.n403 117.001
R1741 VGND.t371 VGND.n403 117.001
R1742 VGND.n417 VGND.n402 117.001
R1743 VGND.t371 VGND.n402 117.001
R1744 VGND.n465 VGND.n429 117.001
R1745 VGND.t643 VGND.n429 117.001
R1746 VGND.n430 VGND.n428 117.001
R1747 VGND.t643 VGND.n428 117.001
R1748 VGND.n476 VGND.n421 117.001
R1749 VGND.t457 VGND.n421 117.001
R1750 VGND.n479 VGND.n478 117.001
R1751 VGND.t457 VGND.n479 117.001
R1752 VGND.n972 VGND.t1200 116.734
R1753 VGND.n1347 VGND.t1189 116.734
R1754 VGND.n1978 VGND.n1977 114.377
R1755 VGND.n1509 VGND.n1365 110.349
R1756 VGND.n1889 VGND.n1270 110.349
R1757 VGND.t755 VGND.t1068 109.579
R1758 VGND.n1581 VGND.t1086 109.579
R1759 VGND.t1103 VGND.t724 109.579
R1760 VGND.t545 VGND.t163 109.579
R1761 VGND.t554 VGND.t936 109.579
R1762 VGND.n1365 VGND.t573 108.505
R1763 VGND.n1977 VGND.t518 108.505
R1764 VGND.n1270 VGND.t1014 108.505
R1765 VGND VGND.t380 106.942
R1766 VGND.t463 VGND.t999 102.992
R1767 VGND.t461 VGND.t1006 102.992
R1768 VGND.n2178 VGND.t1140 102.353
R1769 VGND.n1200 VGND.t1226 102.353
R1770 VGND.n2685 VGND.t1199 102.353
R1771 VGND.n2822 VGND.t129 101.43
R1772 VGND.n1248 VGND.t736 101.43
R1773 VGND.n1262 VGND.t645 101.43
R1774 VGND.t230 VGND.t895 101.15
R1775 VGND.t14 VGND.t1076 101.15
R1776 VGND.n2850 VGND.t1182 99.7825
R1777 VGND.n964 VGND.t1204 99.7825
R1778 VGND.t772 VGND.t311 98.8769
R1779 VGND.t284 VGND.t745 98.8769
R1780 VGND.t521 VGND.t523 98.8769
R1781 VGND.t732 VGND.t10 98.8769
R1782 VGND.t401 VGND.t915 98.8769
R1783 VGND.t543 VGND.t145 98.8769
R1784 VGND.t299 VGND.t135 98.8769
R1785 VGND.t851 VGND.t124 98.8769
R1786 VGND.t646 VGND.t930 98.8769
R1787 VGND.t925 VGND.t160 98.8769
R1788 VGND.t637 VGND.t592 92.7208
R1789 VGND.t1078 VGND 92.7208
R1790 VGND.t602 VGND.t1090 92.7208
R1791 VGND.t533 VGND.t542 92.7208
R1792 VGND.t1107 VGND.t91 92.7208
R1793 VGND VGND.t555 92.7208
R1794 VGND.n476 VGND.n475 89.224
R1795 VGND.n465 VGND.n464 89.224
R1796 VGND.n463 VGND.n432 89.224
R1797 VGND.n436 VGND.n433 89.224
R1798 VGND.n442 VGND.n441 89.224
R1799 VGND.n456 VGND.n444 89.224
R1800 VGND.t181 VGND 88.8318
R1801 VGND.t407 VGND 88.8318
R1802 VGND.n455 VGND.n447 88.4711
R1803 VGND.t352 VGND.n187 85.9264
R1804 VGND.t863 VGND.n93 85.9264
R1805 VGND.n483 VGND.n408 84.7064
R1806 VGND.t967 VGND.t291 84.2917
R1807 VGND.t133 VGND.t907 84.2917
R1808 VGND.t115 VGND.t366 84.2917
R1809 VGND.t997 VGND.t96 84.2917
R1810 VGND VGND.t788 84.2702
R1811 VGND.n3282 VGND 83.8426
R1812 VGND.n484 VGND.n407 80.1887
R1813 VGND.n486 VGND.n406 80.1887
R1814 VGND.n487 VGND.n405 80.1887
R1815 VGND.n417 VGND.n404 80.1887
R1816 VGND.n2394 VGND 76.6073
R1817 VGND.t848 VGND.t1113 75.8626
R1818 VGND VGND.n2394 75.2814
R1819 VGND.n655 VGND.t103 74.8666
R1820 VGND.n656 VGND.t147 74.8666
R1821 VGND.n1467 VGND.t361 74.8666
R1822 VGND.n1558 VGND.t756 74.8666
R1823 VGND.n1605 VGND.t310 74.8666
R1824 VGND.n854 VGND.t914 74.8666
R1825 VGND.n859 VGND.t496 74.8666
R1826 VGND.n1240 VGND.t506 74.8666
R1827 VGND.n1864 VGND.t368 74.8666
R1828 VGND.n939 VGND.t847 74.8666
R1829 VGND.n24 VGND.t144 72.8576
R1830 VGND.n44 VGND.t460 72.8576
R1831 VGND.n3106 VGND.t548 72.8576
R1832 VGND.n214 VGND.t1005 72.8576
R1833 VGND.n3309 VGND.t1007 72.8576
R1834 VGND.n3343 VGND.t729 72.8576
R1835 VGND.n1937 VGND.t571 72.8576
R1836 VGND.n1938 VGND.t304 72.8576
R1837 VGND.n1919 VGND.t890 72.8576
R1838 VGND.t643 VGND.n426 72.7469
R1839 VGND.n460 VGND.t467 72.7469
R1840 VGND.t126 VGND.t1052 71.7175
R1841 VGND.t745 VGND 70.787
R1842 VGND.t959 VGND.t796 67.6928
R1843 VGND.t749 VGND.t1002 67.4335
R1844 VGND.t328 VGND.t952 67.4335
R1845 VGND.t320 VGND.t893 67.4335
R1846 VGND.n422 VGND.t371 66.396
R1847 VGND.t457 VGND.n420 66.396
R1848 VGND.n482 VGND.n409 64.8307
R1849 VGND.n3077 VGND.t298 61.6916
R1850 VGND VGND.t445 61.1229
R1851 VGND VGND.n2986 61.1229
R1852 VGND.n1002 VGND.n63 59.6152
R1853 VGND.n1011 VGND.n63 59.6152
R1854 VGND.t558 VGND.t468 59.0043
R1855 VGND.n451 VGND.n450 58.7133
R1856 VGND.n15 VGND.t752 58.5719
R1857 VGND.n21 VGND.t1059 58.5719
R1858 VGND.n3100 VGND.t842 58.5719
R1859 VGND.n218 VGND.t169 58.5719
R1860 VGND.n3328 VGND.t114 58.5719
R1861 VGND.n107 VGND.t142 58.5719
R1862 VGND.n1416 VGND.t365 58.5719
R1863 VGND.n1307 VGND.t941 58.5719
R1864 VGND.n3404 VGND.t123 57.2177
R1865 VGND.t999 VGND.t461 57.2177
R1866 VGND.n3394 VGND.n71 57.2177
R1867 VGND VGND.n492 56.2331
R1868 VGND.n391 VGND.n389 54.2123
R1869 VGND.n3247 VGND.n3239 54.2123
R1870 VGND.n3261 VGND.n3260 54.2123
R1871 VGND.n3222 VGND.n180 54.2123
R1872 VGND.n3217 VGND.n3216 54.2123
R1873 VGND.n183 VGND.n182 54.2123
R1874 VGND.n3386 VGND.n77 54.2123
R1875 VGND.n3277 VGND.n3255 54.2123
R1876 VGND.n1004 VGND.n1001 53.1823
R1877 VGND.n1001 VGND.t757 53.1823
R1878 VGND.n2390 VGND.n1003 53.1823
R1879 VGND.n1003 VGND.n1002 53.1823
R1880 VGND.n1014 VGND.n1013 53.1823
R1881 VGND.n1013 VGND.n1012 53.1823
R1882 VGND.n1010 VGND.n1009 53.1823
R1883 VGND.n1011 VGND.n1010 53.1823
R1884 VGND.n681 VGND.t567 52.8576
R1885 VGND.n454 VGND.n448 51.7522
R1886 VGND.t1060 VGND.t293 50.5752
R1887 VGND.t1056 VGND.t358 50.5752
R1888 VGND.t137 VGND.t635 50.5752
R1889 VGND VGND.t1078 50.5752
R1890 VGND.t1010 VGND.t715 50.5752
R1891 VGND.t388 VGND.t885 50.5752
R1892 VGND.t106 VGND.t680 50.5752
R1893 VGND.t932 VGND.t139 50.5752
R1894 VGND.n1002 VGND.t560 50.3004
R1895 VGND.t582 VGND.n1011 49.0584
R1896 VGND.n1012 VGND.t582 49.0584
R1897 VGND.n2389 VGND.n1000 48.7505
R1898 VGND.n2393 VGND.n1000 48.7505
R1899 VGND.n2392 VGND.n2391 48.7505
R1900 VGND.n2393 VGND.n2392 48.7505
R1901 VGND.n1603 VGND.t658 48.5719
R1902 VGND.t380 VGND.n3281 47.9103
R1903 VGND.n1611 VGND.t577 47.1434
R1904 VGND.n942 VGND.t1114 47.1434
R1905 VGND.t699 VGND 44.7453
R1906 VGND.n50 VGND 43.9579
R1907 VGND.n3140 VGND 43.9579
R1908 VGND.n3308 VGND 43.9579
R1909 VGND.n475 VGND.n474 42.1089
R1910 VGND.n488 VGND.n404 42.1089
R1911 VGND.n488 VGND.n487 42.1089
R1912 VGND.n486 VGND.n485 42.1089
R1913 VGND.n485 VGND.n484 42.1089
R1914 VGND.n483 VGND.n482 42.1089
R1915 VGND.n3403 VGND.t376 41.9598
R1916 VGND.n655 VGND.t335 40.0005
R1917 VGND.n656 VGND.t979 40.0005
R1918 VGND.n681 VGND.t981 40.0005
R1919 VGND.n1400 VGND.t638 40.0005
R1920 VGND.n1400 VGND.t640 40.0005
R1921 VGND.n784 VGND.t1035 40.0005
R1922 VGND.n784 VGND.t1027 40.0005
R1923 VGND.n783 VGND.t1029 40.0005
R1924 VGND.n783 VGND.t1033 40.0005
R1925 VGND.n792 VGND.t1031 40.0005
R1926 VGND.n792 VGND.t1021 40.0005
R1927 VGND.n1422 VGND.t664 40.0005
R1928 VGND.n1422 VGND.t727 40.0005
R1929 VGND.n771 VGND.t666 40.0005
R1930 VGND.n771 VGND.t1037 40.0005
R1931 VGND.n773 VGND.t1043 40.0005
R1932 VGND.n773 VGND.t1047 40.0005
R1933 VGND.n776 VGND.t1051 40.0005
R1934 VGND.n776 VGND.t1041 40.0005
R1935 VGND.n779 VGND.t1045 40.0005
R1936 VGND.n779 VGND.t1049 40.0005
R1937 VGND.n2625 VGND.t1039 40.0005
R1938 VGND.n1396 VGND.t626 40.0005
R1939 VGND.n1397 VGND.t634 40.0005
R1940 VGND.n1397 VGND.t612 40.0005
R1941 VGND.n1412 VGND.t636 40.0005
R1942 VGND.n1412 VGND.t614 40.0005
R1943 VGND.n1467 VGND.t406 40.0005
R1944 VGND.n1468 VGND.t632 40.0005
R1945 VGND.n1468 VGND.t622 40.0005
R1946 VGND.n1475 VGND.t624 40.0005
R1947 VGND.n1475 VGND.t628 40.0005
R1948 VGND.n1391 VGND.t642 40.0005
R1949 VGND.n1391 VGND.t620 40.0005
R1950 VGND.n1387 VGND.t597 40.0005
R1951 VGND.n1387 VGND.t616 40.0005
R1952 VGND.n1372 VGND.t475 40.0005
R1953 VGND.n1372 VGND.t599 40.0005
R1954 VGND.n1559 VGND.t1063 40.0005
R1955 VGND.n1559 VGND.t1065 40.0005
R1956 VGND.n1558 VGND.t731 40.0005
R1957 VGND.n1571 VGND.t1081 40.0005
R1958 VGND.n1571 VGND.t1073 40.0005
R1959 VGND.n1573 VGND.t1077 40.0005
R1960 VGND.n1573 VGND.t1067 40.0005
R1961 VGND.n1574 VGND.t1075 40.0005
R1962 VGND.n1670 VGND.t1079 40.0005
R1963 VGND.n1670 VGND.t1085 40.0005
R1964 VGND.n1580 VGND.t1083 40.0005
R1965 VGND.n1580 VGND.t1093 40.0005
R1966 VGND.n1582 VGND.t1087 40.0005
R1967 VGND.n1582 VGND.t1089 40.0005
R1968 VGND.n1586 VGND.t1091 40.0005
R1969 VGND.n1586 VGND.t725 40.0005
R1970 VGND.n1597 VGND.t1118 40.0005
R1971 VGND.n1597 VGND.t723 40.0005
R1972 VGND.n1605 VGND.t978 40.0005
R1973 VGND.n854 VGND.t1019 40.0005
R1974 VGND.n859 VGND.t870 40.0005
R1975 VGND.n1240 VGND.t589 40.0005
R1976 VGND.n1864 VGND.t370 40.0005
R1977 VGND.n939 VGND.t849 40.0005
R1978 VGND.n484 VGND.n483 39.4771
R1979 VGND.n1365 VGND.t479 38.7697
R1980 VGND.n838 VGND.t363 38.7697
R1981 VGND.n1977 VGND.t404 38.7697
R1982 VGND.n1284 VGND.t98 38.7697
R1983 VGND.n1270 VGND.t587 38.7697
R1984 VGND.n597 VGND.t112 38.5719
R1985 VGND.n597 VGND.t331 38.5719
R1986 VGND.n598 VGND.t761 38.5719
R1987 VGND.n598 VGND.t307 38.5719
R1988 VGND.n2625 VGND.t1023 38.5719
R1989 VGND.n1396 VGND.t630 38.5719
R1990 VGND.n1388 VGND.t483 38.5719
R1991 VGND.n1388 VGND.t965 38.5719
R1992 VGND.n1574 VGND.t1071 38.5719
R1993 VGND.n1577 VGND.t654 38.5719
R1994 VGND.n1577 VGND.t487 38.5719
R1995 VGND.n1608 VGND.t520 38.5719
R1996 VGND.n1608 VGND.t579 38.5719
R1997 VGND.n1610 VGND.t165 38.5719
R1998 VGND.n1610 VGND.t485 38.5719
R1999 VGND.n860 VGND.t325 38.5719
R2000 VGND.n860 VGND.t610 38.5719
R2001 VGND.n878 VGND.t949 38.5719
R2002 VGND.n878 VGND.t763 38.5719
R2003 VGND.n1244 VGND.t314 38.5719
R2004 VGND.n1244 VGND.t670 38.5719
R2005 VGND.n1271 VGND.t321 38.5719
R2006 VGND.n1271 VGND.t489 38.5719
R2007 VGND.n946 VGND.t557 38.5719
R2008 VGND.n946 VGND.t110 38.5719
R2009 VGND.n3407 VGND.t342 38.3944
R2010 VGND VGND.t990 36.085
R2011 VGND VGND.t833 36.085
R2012 VGND.n1611 VGND.t983 35.4291
R2013 VGND.n942 VGND.t469 35.4291
R2014 VGND.n487 VGND.n486 35.2902
R2015 VGND.n464 VGND.n431 34.659
R2016 VGND.n463 VGND.n462 34.659
R2017 VGND.n462 VGND.n433 34.659
R2018 VGND.n457 VGND.n441 34.659
R2019 VGND.n457 VGND.n456 34.659
R2020 VGND.n455 VGND.n454 34.659
R2021 VGND.n1478 VGND.n1477 34.6358
R2022 VGND.n50 VGND.n49 34.6358
R2023 VGND.n47 VGND.n2 34.6358
R2024 VGND.n3161 VGND.n3145 34.6358
R2025 VGND.n3161 VGND.n3160 34.6358
R2026 VGND.n3155 VGND.n3154 34.6358
R2027 VGND.n3189 VGND.n188 34.6358
R2028 VGND.n3189 VGND.n189 34.6358
R2029 VGND.n3183 VGND.n3182 34.6358
R2030 VGND.n3177 VGND.n3176 34.6358
R2031 VGND.n3176 VGND.n195 34.6358
R2032 VGND.n3170 VGND.n195 34.6358
R2033 VGND.n3140 VGND.n3139 34.6358
R2034 VGND.n3137 VGND.n215 34.6358
R2035 VGND.n3085 VGND.n215 34.6358
R2036 VGND.n3087 VGND.n3085 34.6358
R2037 VGND.n3090 VGND.n220 34.6358
R2038 VGND.n3094 VGND.n220 34.6358
R2039 VGND.n3114 VGND.n3103 34.6358
R2040 VGND.n3110 VGND.n3103 34.6358
R2041 VGND.n3311 VGND.n3308 34.6358
R2042 VGND.n3315 VGND.n3299 34.6358
R2043 VGND.n636 VGND.n629 34.6358
R2044 VGND.n654 VGND.n602 34.6358
R2045 VGND.n650 VGND.n602 34.6358
R2046 VGND.n650 VGND.n649 34.6358
R2047 VGND.n662 VGND.n600 34.6358
R2048 VGND.n658 VGND.n600 34.6358
R2049 VGND.n1459 VGND.n1401 34.6358
R2050 VGND.n1474 VGND.n1394 34.6358
R2051 VGND.n1482 VGND.n1389 34.6358
R2052 VGND.n1658 VGND.n1657 34.6358
R2053 VGND.n1654 VGND.n1587 34.6358
R2054 VGND.n1641 VGND.n1601 34.6358
R2055 VGND.n1636 VGND.n1635 34.6358
R2056 VGND.n1635 VGND.n1606 34.6358
R2057 VGND.n2602 VGND.n835 34.6358
R2058 VGND.n920 VGND.n919 34.6358
R2059 VGND.n915 VGND.n857 34.6358
R2060 VGND.n903 VGND.n863 34.6358
R2061 VGND.n1936 VGND.n1935 34.6358
R2062 VGND.n1935 VGND.n1267 34.6358
R2063 VGND.n1940 VGND.n1265 34.6358
R2064 VGND.n1913 VGND.n1896 34.6358
R2065 VGND.n1904 VGND.n1896 34.6358
R2066 VGND.n1905 VGND.n1904 34.6358
R2067 VGND.n1888 VGND.n1887 34.6358
R2068 VGND.n1915 VGND.n1268 34.6358
R2069 VGND.n2555 VGND.n2554 34.6358
R2070 VGND.n2554 VGND.n2553 34.6358
R2071 VGND.n2549 VGND.n2548 34.6358
R2072 VGND.n1822 VGND.n1760 34.6358
R2073 VGND.n1804 VGND.n1768 34.6358
R2074 VGND.n2007 VGND.n2006 34.6358
R2075 VGND.n2518 VGND.n991 34.6358
R2076 VGND.n2468 VGND.n2467 34.6358
R2077 VGND.n2449 VGND.n2448 34.6358
R2078 VGND.n2448 VGND.n2432 34.6358
R2079 VGND.n1042 VGND.n493 34.6358
R2080 VGND.n2057 VGND.t1236 34.2973
R2081 VGND.n1555 VGND.t1194 34.2973
R2082 VGND.n2477 VGND.t1174 34.2973
R2083 VGND.n263 VGND.t1217 34.2973
R2084 VGND.n2325 VGND.t1153 34.2973
R2085 VGND.n3157 VGND.n3156 33.8829
R2086 VGND.n3151 VGND.n3150 33.8829
R2087 VGND.n3185 VGND.n3184 33.8829
R2088 VGND.n3179 VGND.n3178 33.8829
R2089 VGND.n3130 VGND.n3129 33.8829
R2090 VGND.n3123 VGND.n3122 33.8829
R2091 VGND.n3116 VGND.n3115 33.8829
R2092 VGND.n1673 VGND.n1672 33.8829
R2093 VGND.n905 VGND.n861 33.8829
R2094 VGND.t590 VGND.t613 33.717
R2095 VGND.t722 VGND.t600 33.717
R2096 VGND.t119 VGND.t519 33.717
R2097 VGND.t516 VGND 33.717
R2098 VGND.t12 VGND.t891 33.717
R2099 VGND.t651 VGND.t586 33.717
R2100 VGND.n1310 VGND.t878 33.462
R2101 VGND.n1310 VGND.t928 33.462
R2102 VGND.n1374 VGND.t95 33.462
R2103 VGND.n1374 VGND.t553 33.462
R2104 VGND.n1758 VGND.t773 33.462
R2105 VGND.n1758 VGND.t312 33.462
R2106 VGND.n1762 VGND.t285 33.462
R2107 VGND.n1762 VGND.t746 33.462
R2108 VGND.n1767 VGND.t522 33.462
R2109 VGND.n1767 VGND.t524 33.462
R2110 VGND.n1783 VGND.t733 33.462
R2111 VGND.n1783 VGND.t11 33.462
R2112 VGND.n1991 VGND.t402 33.462
R2113 VGND.n1991 VGND.t916 33.462
R2114 VGND.n990 VGND.t544 33.462
R2115 VGND.n990 VGND.t146 33.462
R2116 VGND.n998 VGND.t300 33.462
R2117 VGND.n998 VGND.t136 33.462
R2118 VGND.n2412 VGND.t852 33.462
R2119 VGND.n2412 VGND.t125 33.462
R2120 VGND.n2420 VGND.t647 33.462
R2121 VGND.n2420 VGND.t931 33.462
R2122 VGND.n2434 VGND.t926 33.462
R2123 VGND.n2434 VGND.t161 33.462
R2124 VGND.n1030 VGND.t1053 33.462
R2125 VGND.n1030 VGND.t127 33.462
R2126 VGND.n3157 VGND.n3146 33.1299
R2127 VGND.n3151 VGND.n3148 33.1299
R2128 VGND.n3185 VGND.n191 33.1299
R2129 VGND.n3179 VGND.n192 33.1299
R2130 VGND.n3095 VGND.n3094 33.1299
R2131 VGND.n3130 VGND.n3097 33.1299
R2132 VGND.n3124 VGND.n3123 33.1299
R2133 VGND.n3121 VGND.n3101 33.1299
R2134 VGND.n3117 VGND.n3116 33.1299
R2135 VGND.n492 VGND.n491 32.9096
R2136 VGND.n2383 VGND.t561 32.8043
R2137 VGND.n1018 VGND.t758 32.8043
R2138 VGND VGND.t772 32.5848
R2139 VGND VGND.t521 32.5848
R2140 VGND VGND.t732 32.5848
R2141 VGND VGND.t401 32.5848
R2142 VGND VGND.t543 32.5848
R2143 VGND VGND.t299 32.5848
R2144 VGND VGND.t851 32.5848
R2145 VGND VGND.t646 32.5848
R2146 VGND VGND.t925 32.5848
R2147 VGND.n1603 VGND.t581 32.5719
R2148 VGND.n454 VGND.n453 32.5005
R2149 VGND.n453 VGND.n438 32.5005
R2150 VGND.n451 VGND.n426 32.5005
R2151 VGND.n445 VGND.n411 32.5005
R2152 VGND.n424 VGND.n411 32.5005
R2153 VGND.n482 VGND.n481 32.5005
R2154 VGND.n481 VGND.n401 32.5005
R2155 VGND.n458 VGND.n457 32.5005
R2156 VGND.n460 VGND.n458 32.5005
R2157 VGND.n443 VGND.n427 32.5005
R2158 VGND.n468 VGND.n427 32.5005
R2159 VGND.n416 VGND.n415 32.5005
R2160 VGND.n420 VGND.n416 32.5005
R2161 VGND.n485 VGND.n400 32.5005
R2162 VGND.n490 VGND.n400 32.5005
R2163 VGND.n462 VGND.n461 32.5005
R2164 VGND.n461 VGND.n460 32.5005
R2165 VGND.n435 VGND.n425 32.5005
R2166 VGND.n468 VGND.n425 32.5005
R2167 VGND.n419 VGND.n418 32.5005
R2168 VGND.n420 VGND.n419 32.5005
R2169 VGND.n489 VGND.n488 32.5005
R2170 VGND.n490 VGND.n489 32.5005
R2171 VGND.n459 VGND.n431 32.5005
R2172 VGND.n460 VGND.n459 32.5005
R2173 VGND.n467 VGND.n466 32.5005
R2174 VGND.n468 VGND.n467 32.5005
R2175 VGND.n477 VGND.n470 32.5005
R2176 VGND.n470 VGND.n469 32.5005
R2177 VGND.n474 VGND.n423 32.5005
R2178 VGND.n423 VGND.n422 32.5005
R2179 VGND.n441 VGND.n433 32.4928
R2180 VGND.n3125 VGND.n3098 32.377
R2181 VGND.n628 VGND.n604 32.377
R2182 VGND.n1854 VGND.n1853 32.377
R2183 VGND.n1891 VGND.n1268 32.377
R2184 VGND.n2560 VGND.n934 32.377
R2185 VGND.n1678 VGND.n1677 32.377
R2186 VGND.n1889 VGND.n1888 31.624
R2187 VGND.n648 VGND.n604 31.2476
R2188 VGND.n2588 VGND.n2587 31.2476
R2189 VGND.n1854 VGND.n1286 31.2476
R2190 VGND.n2560 VGND.n2559 31.2476
R2191 VGND.n456 VGND.n455 30.9174
R2192 VGND.n478 VGND.n473 30.8711
R2193 VGND.n392 VGND.n391 30.8711
R2194 VGND.n3247 VGND.n3246 30.8711
R2195 VGND.n3270 VGND.n3261 30.8711
R2196 VGND.n3224 VGND.n180 30.8711
R2197 VGND.n3216 VGND.n3202 30.8711
R2198 VGND.n3198 VGND.n183 30.8711
R2199 VGND.n3387 VGND.n3386 30.8711
R2200 VGND.n3277 VGND.n3276 30.8711
R2201 VGND.n658 VGND.n657 30.8711
R2202 VGND.n1637 VGND.n1636 30.8711
R2203 VGND.n1979 VGND.n1241 30.8711
R2204 VGND.n1867 VGND.n1865 30.8711
R2205 VGND.n475 VGND.n404 30.7444
R2206 VGND.n1570 VGND.n1560 30.4946
R2207 VGND.n1624 VGND.n835 30.4946
R2208 VGND.n1867 VGND.n1866 30.4946
R2209 VGND.n2377 VGND.t583 30.3424
R2210 VGND.n1461 VGND.n1460 30.1181
R2211 VGND.n1681 VGND.n1680 30.1181
R2212 VGND.n1600 VGND.n1599 30.1181
R2213 VGND.n1914 VGND.n1913 30.1181
R2214 VGND.n3402 VGND.n3401 29.8168
R2215 VGND.t392 VGND.t472 29.8079
R2216 VGND.t472 VGND.t562 29.8079
R2217 VGND.t394 VGND.t759 29.8079
R2218 VGND.t390 VGND.t394 29.8079
R2219 VGND.t560 VGND.t390 29.8079
R2220 VGND.n1465 VGND.n1398 29.7417
R2221 VGND.n2593 VGND.n2592 29.3652
R2222 VGND.n1449 VGND.n1448 28.9887
R2223 VGND.n464 VGND.n463 28.259
R2224 VGND.n1485 VGND.n1484 27.8593
R2225 VGND.n1655 VGND.n1654 27.8593
R2226 VGND.n663 VGND.n662 27.4829
R2227 VGND.n1631 VGND.n1606 27.4829
R2228 VGND.n2599 VGND.n2598 27.4829
R2229 VGND.n917 VGND.n916 27.4829
R2230 VGND.n911 VGND.n857 27.4829
R2231 VGND.n1978 VGND.n1976 27.4829
R2232 VGND.n1976 VGND.n1242 27.4829
R2233 VGND.n1859 VGND.n1285 27.4829
R2234 VGND.n1882 VGND.n1273 27.4829
R2235 VGND.n1485 VGND.n1373 27.1064
R2236 VGND.n3446 VGND.n3445 26.9246
R2237 VGND.n3359 VGND.n95 26.9246
R2238 VGND.n1625 VGND.n1612 26.7299
R2239 VGND.n2337 VGND.n2336 26.6009
R2240 VGND.n1944 VGND.n1265 26.314
R2241 VGND.n2383 VGND.n2382 26.1653
R2242 VGND.n2385 VGND.n2384 26.1653
R2243 VGND.n1018 VGND.n1017 26.1653
R2244 VGND.n469 VGND.n468 25.9813
R2245 VGND.n2822 VGND.t180 25.9346
R2246 VGND.n1248 VGND.t721 25.9346
R2247 VGND.n1262 VGND.t118 25.9346
R2248 VGND.n3235 VGND.t199 25.8199
R2249 VGND.n1662 VGND.n1661 25.7355
R2250 VGND.n1924 VGND.n1922 25.7355
R2251 VGND.n2548 VGND.n2547 25.7355
R2252 VGND.n1824 VGND.n1757 25.7355
R2253 VGND.n2443 VGND.n2442 25.7355
R2254 VGND.n3464 VGND.n2 25.6926
R2255 VGND.n3316 VGND.n3315 25.6926
R2256 VGND.n1817 VGND.n1816 25.6926
R2257 VGND.n1809 VGND.n1765 25.6926
R2258 VGND.n1779 VGND.n1768 25.6926
R2259 VGND.n2006 VGND.n1993 25.6926
R2260 VGND.n2510 VGND.n991 25.6926
R2261 VGND.n2504 VGND.n2503 25.6926
R2262 VGND.n2467 VGND.n2414 25.6926
R2263 VGND.n1043 VGND.n1042 25.6926
R2264 VGND.n637 VGND.n636 25.6005
R2265 VGND.n1677 VGND.n1575 25.6005
R2266 VGND.n15 VGND.t294 25.4291
R2267 VGND.n21 VGND.t359 25.4291
R2268 VGND.n3100 VGND.t933 25.4291
R2269 VGND.n218 VGND.t107 25.4291
R2270 VGND.n3328 VGND.t1011 25.4291
R2271 VGND.n107 VGND.t389 25.4291
R2272 VGND.n1416 VGND.t93 25.4291
R2273 VGND.n1307 VGND.t492 25.4291
R2274 VGND.t130 VGND.t264 25.2879
R2275 VGND.t621 VGND.t405 25.2879
R2276 VGND.t559 VGND.t490 25.2879
R2277 VGND.n3429 VGND.n3428 25.224
R2278 VGND.n3428 VGND.n60 25.224
R2279 VGND.n3424 VGND.n3423 25.224
R2280 VGND.n3423 VGND.n3422 25.224
R2281 VGND.n3420 VGND.n3419 25.224
R2282 VGND.n3419 VGND.n3411 25.224
R2283 VGND.n3415 VGND.n3414 25.224
R2284 VGND.n3414 VGND.n39 25.224
R2285 VGND.n3455 VGND.n3454 25.224
R2286 VGND.n3454 VGND.n3453 25.224
R2287 VGND.n3451 VGND.n22 25.224
R2288 VGND.n3376 VGND.n3375 25.224
R2289 VGND.n3375 VGND.n83 25.224
R2290 VGND.n3371 VGND.n3370 25.224
R2291 VGND.n3370 VGND.n3369 25.224
R2292 VGND.n3367 VGND.n3366 25.224
R2293 VGND.n3366 VGND.n89 25.224
R2294 VGND.n3362 VGND.n3361 25.224
R2295 VGND.n3361 VGND.n3360 25.224
R2296 VGND.n3335 VGND.n3334 25.224
R2297 VGND.n3336 VGND.n3335 25.224
R2298 VGND.n3353 VGND.n3340 25.224
R2299 VGND.n127 VGND.n125 25.224
R2300 VGND.n131 VGND.n125 25.224
R2301 VGND.n132 VGND.n124 25.224
R2302 VGND.n136 VGND.n124 25.224
R2303 VGND.n137 VGND.n123 25.224
R2304 VGND.n141 VGND.n123 25.224
R2305 VGND.n142 VGND.n122 25.224
R2306 VGND.n146 VGND.n122 25.224
R2307 VGND.n147 VGND.n121 25.224
R2308 VGND.n151 VGND.n121 25.224
R2309 VGND.n152 VGND.n120 25.224
R2310 VGND.n156 VGND.n120 25.224
R2311 VGND.n157 VGND.n119 25.224
R2312 VGND.n161 VGND.n119 25.224
R2313 VGND.n162 VGND.n118 25.224
R2314 VGND.n166 VGND.n118 25.224
R2315 VGND.n167 VGND.n117 25.224
R2316 VGND.n171 VGND.n117 25.224
R2317 VGND.n1572 VGND.n1570 25.224
R2318 VGND.n1681 VGND.n1572 25.224
R2319 VGND.n2473 VGND.n2472 24.9894
R2320 VGND.n2332 VGND.n2331 24.9894
R2321 VGND.n3144 VGND.n3143 24.9767
R2322 VGND.n3169 VGND.n3168 24.9767
R2323 VGND.n3108 VGND.n3105 24.9767
R2324 VGND.n2881 VGND.n585 24.968
R2325 VGND.n3400 VGND.t464 24.9236
R2326 VGND.n3400 VGND.t462 24.9236
R2327 VGND.n535 VGND.t921 24.9236
R2328 VGND.n535 VGND.t924 24.9236
R2329 VGND.n627 VGND.t970 24.9236
R2330 VGND.n627 VGND.t971 24.9236
R2331 VGND.n626 VGND.t882 24.9236
R2332 VGND.n626 VGND.t5 24.9236
R2333 VGND.n1413 VGND.t138 24.9236
R2334 VGND.n1413 VGND.t591 24.9236
R2335 VGND.n1551 VGND.t769 24.9236
R2336 VGND.n1551 VGND.t541 24.9236
R2337 VGND.n1585 VGND.t603 24.9236
R2338 VGND.n1585 VGND.t1104 24.9236
R2339 VGND.n836 VGND.t1108 24.9236
R2340 VGND.n836 VGND.t738 24.9236
R2341 VGND.n838 VGND.t570 24.9236
R2342 VGND.n844 VGND.t1003 24.9236
R2343 VGND.n844 VGND.t953 24.9236
R2344 VGND.n843 VGND.t750 24.9236
R2345 VGND.n843 VGND.t329 24.9236
R2346 VGND.n853 VGND.t387 24.9236
R2347 VGND.n853 VGND.t122 24.9236
R2348 VGND.n1850 VGND.t742 24.9236
R2349 VGND.n1850 VGND.t744 24.9236
R2350 VGND.n1288 VGND.t1112 24.9236
R2351 VGND.n1288 VGND.t550 24.9236
R2352 VGND.n1284 VGND.t1017 24.9236
R2353 VGND.n1890 VGND.t539 24.9236
R2354 VGND.n1890 VGND.t652 24.9236
R2355 VGND.n933 VGND.t375 24.9236
R2356 VGND.n933 VGND.t494 24.9236
R2357 VGND.n936 VGND.t302 24.9236
R2358 VGND.n936 VGND.t937 24.9236
R2359 VGND VGND.t463 24.7946
R2360 VGND.n1695 VGND.n1694 24.4711
R2361 VGND.n910 VGND.n909 24.4711
R2362 VGND.n2602 VGND.n2601 24.4711
R2363 VGND.n905 VGND.n904 24.4711
R2364 VGND.n904 VGND.n903 24.4711
R2365 VGND.n2555 VGND.n937 24.4711
R2366 VGND.t990 VGND.t987 24.2493
R2367 VGND.t833 VGND.t836 24.2493
R2368 VGND.t342 VGND.t345 24.2493
R2369 VGND.n3459 VGND.n16 24.0946
R2370 VGND.n3330 VGND.n110 24.0946
R2371 VGND.n281 VGND.t239 23.7273
R2372 VGND.n2594 VGND.n841 23.7181
R2373 VGND.n1328 VGND.n1314 23.7181
R2374 VGND.n1339 VGND.n1314 23.7181
R2375 VGND.n1433 VGND.n1420 23.7181
R2376 VGND.n1433 VGND.n1432 23.7181
R2377 VGND.n1642 VGND.n1641 23.7181
R2378 VGND.n2598 VGND.n841 23.7181
R2379 VGND.n2586 VGND.n848 23.7181
R2380 VGND.n920 VGND.n848 23.7181
R2381 VGND.n1931 VGND.n1267 23.7181
R2382 VGND.n1859 VGND.n1858 23.7181
R2383 VGND.n1789 VGND.n1788 23.7181
R2384 VGND.n2029 VGND.n1223 23.7181
R2385 VGND.n2012 VGND.n2011 23.7181
R2386 VGND.n1999 VGND.n989 23.7181
R2387 VGND.n2499 VGND.n2498 23.7181
R2388 VGND.n2460 VGND.n2459 23.7181
R2389 VGND.n2985 VGND.n493 23.7181
R2390 VGND.t1052 VGND 23.6345
R2391 VGND.n876 VGND.n875 23.4338
R2392 VGND.n1392 VGND.n1389 23.3417
R2393 VGND.n1658 VGND.n1583 23.3417
R2394 VGND.n450 VGND.n448 23.2076
R2395 VGND.n3176 VGND.n3175 23.1729
R2396 VGND.n664 VGND.n599 22.9652
R2397 VGND.n664 VGND.n663 22.9652
R2398 VGND.n1631 VGND.n1630 22.9652
R2399 VGND.n1630 VGND.n1629 22.9652
R2400 VGND.n2588 VGND.n845 22.9652
R2401 VGND.n911 VGND.n910 22.9652
R2402 VGND.n1972 VGND.n1242 22.9652
R2403 VGND.n1972 VGND.n1971 22.9652
R2404 VGND.n1852 VGND.n1851 22.9652
R2405 VGND.n1883 VGND.n1882 22.9652
R2406 VGND.n1883 VGND.n1272 22.9652
R2407 VGND.n943 VGND.n940 22.9652
R2408 VGND.n3282 VGND.n3235 22.9387
R2409 VGND.n3393 VGND.t527 22.8805
R2410 VGND.n1642 VGND.n1600 22.5887
R2411 VGND.n24 VGND.t508 22.3257
R2412 VGND.n44 VGND.t526 22.3257
R2413 VGND.n3106 VGND.t510 22.3257
R2414 VGND.n214 VGND.t7 22.3257
R2415 VGND.n3309 VGND.t377 22.3257
R2416 VGND.n3343 VGND.t477 22.3257
R2417 VGND.n1937 VGND.t1094 22.3257
R2418 VGND.n1938 VGND.t829 22.3257
R2419 VGND.n1919 VGND.t976 22.3257
R2420 VGND.n649 VGND.n648 22.2123
R2421 VGND.n2587 VGND.n2586 22.2123
R2422 VGND.n916 VGND.n915 22.2123
R2423 VGND.n2559 VGND.n2558 22.2123
R2424 VGND.n1824 VGND.n1823 22.2123
R2425 VGND.n1823 VGND.n1822 22.2123
R2426 VGND.n1818 VGND.n1760 22.2123
R2427 VGND.n1818 VGND.n1817 22.2123
R2428 VGND.n1805 VGND.n1765 22.2123
R2429 VGND.n1805 VGND.n1804 22.2123
R2430 VGND.n1788 VGND.n1784 22.2123
R2431 VGND.n1784 VGND.n1223 22.2123
R2432 VGND.n2011 VGND.n1992 22.2123
R2433 VGND.n2007 VGND.n1992 22.2123
R2434 VGND.n2519 VGND.n989 22.2123
R2435 VGND.n2519 VGND.n2518 22.2123
R2436 VGND.n2503 VGND.n999 22.2123
R2437 VGND.n2499 VGND.n999 22.2123
R2438 VGND.n2472 VGND.n2413 22.2123
R2439 VGND.n2468 VGND.n2413 22.2123
R2440 VGND.n2459 VGND.n2421 22.2123
R2441 VGND.n2449 VGND.n2421 22.2123
R2442 VGND.n2444 VGND.n2432 22.2123
R2443 VGND.n2444 VGND.n2443 22.2123
R2444 VGND.n2336 VGND.n1031 22.2123
R2445 VGND.n2332 VGND.n1031 22.2123
R2446 VGND.n446 VGND.n412 21.6752
R2447 VGND.n3408 VGND 21.6512
R2448 VGND.n3460 VGND.n3459 21.4593
R2449 VGND.n3452 VGND.n3451 21.4593
R2450 VGND.n3330 VGND.n3329 21.4593
R2451 VGND.n3340 VGND.n108 21.4593
R2452 VGND.n599 VGND.n585 21.4593
R2453 VGND.n1629 VGND.n1628 21.4593
R2454 VGND.n2592 VGND.n845 21.4593
R2455 VGND.n1979 VGND.n1978 21.4593
R2456 VGND.n1887 VGND.n1272 21.4593
R2457 VGND.n1699 VGND.n1556 20.8482
R2458 VGND.n1461 VGND.n1398 20.7064
R2459 VGND.n1449 VGND.n1401 20.7064
R2460 VGND.n3424 VGND.n60 20.3299
R2461 VGND.n3415 VGND.n3411 20.3299
R2462 VGND.n3371 VGND.n83 20.3299
R2463 VGND.n3362 VGND.n89 20.3299
R2464 VGND.t987 VGND 19.3418
R2465 VGND.t836 VGND 19.3418
R2466 VGND.t345 VGND 19.3418
R2467 VGND.n3430 VGND.n3429 19.2926
R2468 VGND.n3377 VGND.n3376 19.2926
R2469 VGND.n2394 VGND.t392 19.2511
R2470 VGND.t1006 VGND 19.0729
R2471 VGND.n3138 VGND.n3137 18.824
R2472 VGND.n132 VGND.n131 18.824
R2473 VGND.n137 VGND.n136 18.824
R2474 VGND.n142 VGND.n141 18.824
R2475 VGND.n147 VGND.n146 18.824
R2476 VGND.n152 VGND.n151 18.824
R2477 VGND.n157 VGND.n156 18.824
R2478 VGND.n162 VGND.n161 18.824
R2479 VGND.n167 VGND.n166 18.824
R2480 VGND.n2828 VGND.n2827 18.2791
R2481 VGND.n1517 VGND.n1362 18.2791
R2482 VGND.n1097 VGND.n1096 18.2791
R2483 VGND.n33 VGND.n22 17.7867
R2484 VGND.n3353 VGND.n3352 17.7867
R2485 VGND.n1074 VGND.n1055 17.7007
R2486 VGND.n2359 VGND.n2358 17.4137
R2487 VGND.n3421 VGND.n3420 17.3181
R2488 VGND.n3145 VGND.n3144 17.3181
R2489 VGND.n3170 VGND.n3169 17.3181
R2490 VGND.n3090 VGND.n3089 17.3181
R2491 VGND.n3368 VGND.n3367 17.3181
R2492 VGND.n1447 VGND.n1446 17.3181
R2493 VGND.n2233 VGND.n2232 17.195
R2494 VGND.n2792 VGND.n692 16.9936
R2495 VGND.n3020 VGND.n264 16.9545
R2496 VGND.n2600 VGND.n2599 16.9417
R2497 VGND.n1863 VGND.n1285 16.9417
R2498 VGND.t702 VGND.t1054 16.8587
R2499 VGND.t877 VGND.t267 16.8587
R2500 VGND.t540 VGND.t709 16.8587
R2501 VGND.t187 VGND.t720 16.8587
R2502 VGND.t887 VGND.t22 16.8587
R2503 VGND.t454 VGND.t1008 16.8587
R2504 VGND.n3040 VGND.n255 16.8353
R2505 VGND.n3035 VGND.n256 16.7924
R2506 VGND.n523 VGND.n522 16.763
R2507 VGND.n1012 VGND.n67 16.4566
R2508 VGND.n1466 VGND.n1465 16.1887
R2509 VGND.n1448 VGND.n1447 16.1887
R2510 VGND.n1695 VGND.n1556 16.1887
R2511 VGND.n3422 VGND.n3421 15.8123
R2512 VGND.n3445 VGND.n39 15.8123
R2513 VGND.n3139 VGND.n3138 15.8123
R2514 VGND.n3110 VGND.n3109 15.8123
R2515 VGND.n3369 VGND.n3368 15.8123
R2516 VGND.n3360 VGND.n3359 15.8123
R2517 VGND.n127 VGND.n69 15.8123
R2518 VGND.n3292 VGND.n171 15.8123
R2519 VGND.n1496 VGND.n1495 15.3963
R2520 VGND.n2985 VGND.n2984 15.3963
R2521 VGND.n2989 VGND.n2988 15.3963
R2522 VGND.n3089 VGND.n3088 15.0593
R2523 VGND.t562 VGND.n2393 14.9042
R2524 VGND.n2393 VGND.t759 14.9042
R2525 VGND.n1931 VGND.n1930 14.8179
R2526 VGND.n2988 VGND.n278 14.8179
R2527 VGND.n3445 VGND.n3444 14.775
R2528 VGND.n3461 VGND.n4 14.775
R2529 VGND.n3359 VGND.n92 14.775
R2530 VGND.n3324 VGND.n113 14.775
R2531 VGND.n617 VGND.n614 14.775
R2532 VGND.n1437 VGND.n1420 14.775
R2533 VGND.n1721 VGND.n1720 14.775
R2534 VGND.n1839 VGND.n1838 14.775
R2535 VGND.n2029 VGND.n2028 14.775
R2536 VGND.n2498 VGND.n2497 14.775
R2537 VGND.n2939 VGND.n2938 14.2735
R2538 VGND.n2540 VGND.n2539 14.065
R2539 VGND.n553 VGND.n550 14.0503
R2540 VGND.n2846 VGND.n2845 14.0503
R2541 VGND.n811 VGND.n808 14.0503
R2542 VGND.n1625 VGND.n1624 13.9299
R2543 VGND.n1866 VGND.n1273 13.9299
R2544 VGND.n970 VGND.n969 13.8859
R2545 VGND.n3455 VGND.n16 13.5534
R2546 VGND.n3334 VGND.n110 13.5534
R2547 VGND.n3396 VGND.n69 12.8005
R2548 VGND.n3396 VGND.n68 12.8005
R2549 VGND.n3402 VGND.n68 12.8005
R2550 VGND.n2172 VGND.n1174 12.8005
R2551 VGND.n2143 VGND.n2142 12.8005
R2552 VGND.n2679 VGND.n753 12.8005
R2553 VGND.n887 VGND.n886 12.8005
R2554 VGND.n1851 VGND.n1289 12.5161
R2555 VGND.n3070 VGND.n3069 12.424
R2556 VGND.n3065 VGND.n3055 12.424
R2557 VGND.n2792 VGND.n2791 12.1384
R2558 VGND.n1672 VGND.n1671 11.9309
R2559 VGND.n3143 VGND.n3142 11.3835
R2560 VGND.n1661 VGND.n1583 11.2946
R2561 VGND.n1858 VGND.n1286 11.2946
R2562 VGND.n53 VGND.n52 11.2844
R2563 VGND.n3307 VGND.n3306 11.2844
R2564 VGND.n306 VGND.n299 11.0382
R2565 VGND.n302 VGND.n299 11.0382
R2566 VGND.n300 VGND.n298 11.0382
R2567 VGND.n302 VGND.n298 11.0382
R2568 VGND.n314 VGND.n294 11.0382
R2569 VGND.n297 VGND.n294 11.0382
R2570 VGND.n296 VGND.n293 11.0382
R2571 VGND.n297 VGND.n293 11.0382
R2572 VGND.n291 VGND.n289 11.0382
R2573 VGND.n322 VGND.n291 11.0382
R2574 VGND.n292 VGND.n290 11.0382
R2575 VGND.n322 VGND.n292 11.0382
R2576 VGND.n365 VGND.n343 11.0382
R2577 VGND.n361 VGND.n343 11.0382
R2578 VGND.n344 VGND.n342 11.0382
R2579 VGND.n361 VGND.n342 11.0382
R2580 VGND.n337 VGND.n285 11.0382
R2581 VGND.n333 VGND.n285 11.0382
R2582 VGND.n286 VGND.n284 11.0382
R2583 VGND.n333 VGND.n284 11.0382
R2584 VGND.n3245 VGND.n3238 11.0382
R2585 VGND.n3238 VGND.n3237 11.0382
R2586 VGND.n3242 VGND.n3236 11.0382
R2587 VGND.n3237 VGND.n3236 11.0382
R2588 VGND.n3269 VGND.n3268 11.0382
R2589 VGND.n3268 VGND.n3267 11.0382
R2590 VGND.n3266 VGND.n3265 11.0382
R2591 VGND.n3267 VGND.n3266 11.0382
R2592 VGND.n3208 VGND.n3207 11.0382
R2593 VGND.n3213 VGND.n3208 11.0382
R2594 VGND.n3204 VGND.n3203 11.0382
R2595 VGND.n3213 VGND.n3204 11.0382
R2596 VGND.n3197 VGND.n3196 11.0382
R2597 VGND.n3196 VGND.n3195 11.0382
R2598 VGND.n3194 VGND.n3193 11.0382
R2599 VGND.n3195 VGND.n3194 11.0382
R2600 VGND.n3225 VGND.n178 11.0382
R2601 VGND.n3209 VGND.n178 11.0382
R2602 VGND.n179 VGND.n177 11.0382
R2603 VGND.n3209 VGND.n177 11.0382
R2604 VGND.n203 VGND.n196 11.0382
R2605 VGND.n207 VGND.n196 11.0382
R2606 VGND.n206 VGND.n205 11.0382
R2607 VGND.n207 VGND.n206 11.0382
R2608 VGND.n3259 VGND.n3254 11.0382
R2609 VGND.n3254 VGND.n3253 11.0382
R2610 VGND.n3256 VGND.n3252 11.0382
R2611 VGND.n3253 VGND.n3252 11.0382
R2612 VGND.n3388 VGND.n73 11.0382
R2613 VGND.n3392 VGND.n73 11.0382
R2614 VGND.n3391 VGND.n3390 11.0382
R2615 VGND.n3392 VGND.n3391 11.0382
R2616 VGND.n356 VGND.n348 11.0382
R2617 VGND.n348 VGND.n347 11.0382
R2618 VGND.n353 VGND.n346 11.0382
R2619 VGND.n347 VGND.n346 11.0382
R2620 VGND.n381 VGND.n372 11.0382
R2621 VGND.n377 VGND.n372 11.0382
R2622 VGND.n373 VGND.n371 11.0382
R2623 VGND.n377 VGND.n371 11.0382
R2624 VGND.n393 VGND.n280 11.0382
R2625 VGND.n397 VGND.n280 11.0382
R2626 VGND.n396 VGND.n395 11.0382
R2627 VGND.n397 VGND.n396 11.0382
R2628 VGND.n3076 VGND.n3075 11.0382
R2629 VGND.n3073 VGND.n3072 11.0382
R2630 VGND.n3064 VGND.n3063 11.0382
R2631 VGND.n3063 VGND.n3062 11.0382
R2632 VGND.n3059 VGND.n3058 11.0382
R2633 VGND.n3059 VGND.n223 11.0382
R2634 VGND.n2098 VGND.n2042 10.9091
R2635 VGND.n1431 VGND.n1430 10.8805
R2636 VGND.n471 VGND.t458 10.6509
R2637 VGND.n3066 VGND.n3065 10.6195
R2638 VGND.n3069 VGND.n3068 10.6189
R2639 VGND.n1340 VGND.n1339 10.5983
R2640 VGND.n657 VGND.n654 10.5417
R2641 VGND.n1470 VGND.n1466 10.5417
R2642 VGND.n1905 VGND.n1241 10.5417
R2643 VGND.n1865 VGND.n1863 10.5417
R2644 VGND.n2553 VGND.n940 10.5417
R2645 VGND.n392 VGND.n390 10.4476
R2646 VGND.n3246 VGND.n3241 10.4476
R2647 VGND.n3271 VGND.n3270 10.4476
R2648 VGND.n3224 VGND.n3223 10.4476
R2649 VGND.n3218 VGND.n3202 10.4476
R2650 VGND.n3199 VGND.n3198 10.4476
R2651 VGND.n3387 VGND.n3385 10.4476
R2652 VGND.n3276 VGND.n3275 10.4476
R2653 VGND.n3453 VGND.n3452 10.1652
R2654 VGND.n3336 VGND.n108 10.1652
R2655 VGND.n1495 VGND.n1494 10.1652
R2656 VGND.n1494 VGND.n1373 10.1652
R2657 VGND.n1694 VGND.n1693 10.1652
R2658 VGND.n2601 VGND.n2600 10.1652
R2659 VGND.n909 VGND.n908 10.1652
R2660 VGND.n2558 VGND.n937 10.1652
R2661 VGND.n637 VGND.n625 9.88085
R2662 VGND.n1747 VGND.n1746 9.7205
R2663 VGND.n247 VGND.n246 9.7205
R2664 VGND.n2437 VGND.n2436 9.71789
R2665 VGND.n2353 VGND.n2352 9.71789
R2666 VGND.n53 VGND.n42 9.70901
R2667 VGND.n3438 VGND.n3437 9.70901
R2668 VGND.n27 VGND.n26 9.70901
R2669 VGND.n3306 VGND.n3305 9.70901
R2670 VGND.n100 VGND.n99 9.70901
R2671 VGND.n3345 VGND.n3344 9.70901
R2672 VGND.n48 VGND.n47 9.41227
R2673 VGND.n3310 VGND.n3299 9.41227
R2674 VGND.n1637 VGND.n1604 9.41227
R2675 VGND.n1940 VGND.n1939 9.41227
R2676 VGND.n1921 VGND.n1920 9.41227
R2677 VGND.n2153 VGND.n1174 9.3031
R2678 VGND.n2143 VGND.n1182 9.3031
R2679 VGND.n2661 VGND.n753 9.3031
R2680 VGND.n1328 VGND.n1327 9.3031
R2681 VGND.n1721 VGND.n1535 9.3031
R2682 VGND.n1838 VGND.n1836 9.3031
R2683 VGND.n3447 VGND.n3446 9.3005
R2684 VGND.n3440 VGND.n3439 9.3005
R2685 VGND.n3442 VGND.n3441 9.3005
R2686 VGND.n3444 VGND.n3443 9.3005
R2687 VGND.n3445 VGND.n36 9.3005
R2688 VGND.n55 VGND.n54 9.3005
R2689 VGND.n56 VGND.n41 9.3005
R2690 VGND.n3431 VGND.n3430 9.3005
R2691 VGND.n3429 VGND.n59 9.3005
R2692 VGND.n3428 VGND.n3427 9.3005
R2693 VGND.n3426 VGND.n60 9.3005
R2694 VGND.n3425 VGND.n3424 9.3005
R2695 VGND.n3423 VGND.n61 9.3005
R2696 VGND.n3422 VGND.n62 9.3005
R2697 VGND.n3421 VGND.n3409 9.3005
R2698 VGND.n3420 VGND.n3410 9.3005
R2699 VGND.n3419 VGND.n3418 9.3005
R2700 VGND.n3417 VGND.n3411 9.3005
R2701 VGND.n3416 VGND.n3415 9.3005
R2702 VGND.n3414 VGND.n3413 9.3005
R2703 VGND.n3412 VGND.n39 9.3005
R2704 VGND.n29 VGND.n28 9.3005
R2705 VGND.n31 VGND.n23 9.3005
R2706 VGND.n34 VGND.n33 9.3005
R2707 VGND.n3461 VGND.n13 9.3005
R2708 VGND.n3460 VGND.n14 9.3005
R2709 VGND.n3459 VGND.n3458 9.3005
R2710 VGND.n3457 VGND.n16 9.3005
R2711 VGND.n3456 VGND.n3455 9.3005
R2712 VGND.n3454 VGND.n18 9.3005
R2713 VGND.n3453 VGND.n19 9.3005
R2714 VGND.n3452 VGND.n20 9.3005
R2715 VGND.n3451 VGND.n3450 9.3005
R2716 VGND.n35 VGND.n22 9.3005
R2717 VGND.n51 VGND.n50 9.3005
R2718 VGND.n49 VGND.n43 9.3005
R2719 VGND.n47 VGND.n46 9.3005
R2720 VGND.n45 VGND.n2 9.3005
R2721 VGND.n3465 VGND.n3464 9.3005
R2722 VGND.n6 VGND.n5 9.3005
R2723 VGND.n11 VGND.n10 9.3005
R2724 VGND.n12 VGND.n4 9.3005
R2725 VGND.n3111 VGND.n3110 9.3005
R2726 VGND.n3112 VGND.n3103 9.3005
R2727 VGND.n3141 VGND.n3140 9.3005
R2728 VGND.n3139 VGND.n213 9.3005
R2729 VGND.n3137 VGND.n3136 9.3005
R2730 VGND.n3135 VGND.n215 9.3005
R2731 VGND.n3085 VGND.n216 9.3005
R2732 VGND.n3087 VGND.n3086 9.3005
R2733 VGND.n3091 VGND.n3090 9.3005
R2734 VGND.n3092 VGND.n220 9.3005
R2735 VGND.n3094 VGND.n3093 9.3005
R2736 VGND.n3096 VGND.n217 9.3005
R2737 VGND.n3131 VGND.n3130 9.3005
R2738 VGND.n3128 VGND.n3127 9.3005
R2739 VGND.n3126 VGND.n3125 9.3005
R2740 VGND.n3123 VGND.n3099 9.3005
R2741 VGND.n3121 VGND.n3120 9.3005
R2742 VGND.n3119 VGND.n3118 9.3005
R2743 VGND.n3116 VGND.n3102 9.3005
R2744 VGND.n3114 VGND.n3113 9.3005
R2745 VGND.n3175 VGND.n3174 9.3005
R2746 VGND.n3171 VGND.n3170 9.3005
R2747 VGND.n3172 VGND.n195 9.3005
R2748 VGND.n3176 VGND.n194 9.3005
R2749 VGND.n3145 VGND.n211 9.3005
R2750 VGND.n3162 VGND.n3161 9.3005
R2751 VGND.n3160 VGND.n3159 9.3005
R2752 VGND.n3158 VGND.n3157 9.3005
R2753 VGND.n3155 VGND.n3147 9.3005
R2754 VGND.n3154 VGND.n3153 9.3005
R2755 VGND.n3152 VGND.n3151 9.3005
R2756 VGND.n3149 VGND.n188 9.3005
R2757 VGND.n3189 VGND.n3188 9.3005
R2758 VGND.n3187 VGND.n189 9.3005
R2759 VGND.n3186 VGND.n3185 9.3005
R2760 VGND.n3183 VGND.n190 9.3005
R2761 VGND.n3182 VGND.n3181 9.3005
R2762 VGND.n3180 VGND.n3179 9.3005
R2763 VGND.n3177 VGND.n193 9.3005
R2764 VGND.n3356 VGND.n95 9.3005
R2765 VGND.n102 VGND.n101 9.3005
R2766 VGND.n104 VGND.n103 9.3005
R2767 VGND.n105 VGND.n92 9.3005
R2768 VGND.n3359 VGND.n3358 9.3005
R2769 VGND.n3304 VGND.n3301 9.3005
R2770 VGND.n3303 VGND.n80 9.3005
R2771 VGND.n3378 VGND.n3377 9.3005
R2772 VGND.n3376 VGND.n82 9.3005
R2773 VGND.n3375 VGND.n3374 9.3005
R2774 VGND.n3373 VGND.n83 9.3005
R2775 VGND.n3372 VGND.n3371 9.3005
R2776 VGND.n3370 VGND.n84 9.3005
R2777 VGND.n3369 VGND.n85 9.3005
R2778 VGND.n3368 VGND.n87 9.3005
R2779 VGND.n3367 VGND.n88 9.3005
R2780 VGND.n3366 VGND.n3365 9.3005
R2781 VGND.n3364 VGND.n89 9.3005
R2782 VGND.n3363 VGND.n3362 9.3005
R2783 VGND.n3361 VGND.n90 9.3005
R2784 VGND.n3360 VGND.n91 9.3005
R2785 VGND.n3347 VGND.n3342 9.3005
R2786 VGND.n3350 VGND.n3349 9.3005
R2787 VGND.n3352 VGND.n3351 9.3005
R2788 VGND.n3308 VGND.n3300 9.3005
R2789 VGND.n3312 VGND.n3311 9.3005
R2790 VGND.n3313 VGND.n3299 9.3005
R2791 VGND.n3315 VGND.n3314 9.3005
R2792 VGND.n3317 VGND.n3316 9.3005
R2793 VGND.n3319 VGND.n3318 9.3005
R2794 VGND.n3321 VGND.n114 9.3005
R2795 VGND.n3325 VGND.n3324 9.3005
R2796 VGND.n3326 VGND.n113 9.3005
R2797 VGND.n3329 VGND.n3327 9.3005
R2798 VGND.n3331 VGND.n3330 9.3005
R2799 VGND.n3332 VGND.n110 9.3005
R2800 VGND.n3334 VGND.n3333 9.3005
R2801 VGND.n3335 VGND.n109 9.3005
R2802 VGND.n3337 VGND.n3336 9.3005
R2803 VGND.n3338 VGND.n108 9.3005
R2804 VGND.n3340 VGND.n3339 9.3005
R2805 VGND.n3354 VGND.n3353 9.3005
R2806 VGND.n3293 VGND.n3292 9.3005
R2807 VGND.n171 VGND.n170 9.3005
R2808 VGND.n3402 VGND.n3399 9.3005
R2809 VGND.n3398 VGND.n68 9.3005
R2810 VGND.n3397 VGND.n3396 9.3005
R2811 VGND.n126 VGND.n69 9.3005
R2812 VGND.n128 VGND.n127 9.3005
R2813 VGND.n129 VGND.n125 9.3005
R2814 VGND.n131 VGND.n130 9.3005
R2815 VGND.n133 VGND.n132 9.3005
R2816 VGND.n134 VGND.n124 9.3005
R2817 VGND.n136 VGND.n135 9.3005
R2818 VGND.n138 VGND.n137 9.3005
R2819 VGND.n139 VGND.n123 9.3005
R2820 VGND.n141 VGND.n140 9.3005
R2821 VGND.n143 VGND.n142 9.3005
R2822 VGND.n144 VGND.n122 9.3005
R2823 VGND.n146 VGND.n145 9.3005
R2824 VGND.n148 VGND.n147 9.3005
R2825 VGND.n149 VGND.n121 9.3005
R2826 VGND.n151 VGND.n150 9.3005
R2827 VGND.n153 VGND.n152 9.3005
R2828 VGND.n154 VGND.n120 9.3005
R2829 VGND.n156 VGND.n155 9.3005
R2830 VGND.n158 VGND.n157 9.3005
R2831 VGND.n159 VGND.n119 9.3005
R2832 VGND.n161 VGND.n160 9.3005
R2833 VGND.n163 VGND.n162 9.3005
R2834 VGND.n164 VGND.n118 9.3005
R2835 VGND.n166 VGND.n165 9.3005
R2836 VGND.n168 VGND.n167 9.3005
R2837 VGND.n169 VGND.n117 9.3005
R2838 VGND.n553 VGND.n552 9.3005
R2839 VGND.n556 VGND.n547 9.3005
R2840 VGND.n558 VGND.n557 9.3005
R2841 VGND.n560 VGND.n559 9.3005
R2842 VGND.n563 VGND.n562 9.3005
R2843 VGND.n545 VGND.n544 9.3005
R2844 VGND.n538 VGND.n537 9.3005
R2845 VGND.n527 VGND.n526 9.3005
R2846 VGND.n2932 VGND.n2931 9.3005
R2847 VGND.n2933 VGND.n524 9.3005
R2848 VGND.n2935 VGND.n2934 9.3005
R2849 VGND.n2937 VGND.n2936 9.3005
R2850 VGND.n2160 VGND.n1174 9.3005
R2851 VGND.n2156 VGND.n1174 9.3005
R2852 VGND.n2174 VGND.n2173 9.3005
R2853 VGND.n2176 VGND.n2175 9.3005
R2854 VGND.n2177 VGND.n1170 9.3005
R2855 VGND.n2181 VGND.n2180 9.3005
R2856 VGND.n2184 VGND.n2183 9.3005
R2857 VGND.n2186 VGND.n1167 9.3005
R2858 VGND.n2188 VGND.n2187 9.3005
R2859 VGND.n2201 VGND.n2200 9.3005
R2860 VGND.n2203 VGND.n2202 9.3005
R2861 VGND.n2205 VGND.n2204 9.3005
R2862 VGND.n2206 VGND.n1156 9.3005
R2863 VGND.n2209 VGND.n2208 9.3005
R2864 VGND.n2210 VGND.n1155 9.3005
R2865 VGND.n2212 VGND.n2211 9.3005
R2866 VGND.n2213 VGND.n1154 9.3005
R2867 VGND.n2216 VGND.n2215 9.3005
R2868 VGND.n2223 VGND.n2222 9.3005
R2869 VGND.n2221 VGND.n1153 9.3005
R2870 VGND.n2220 VGND.n2219 9.3005
R2871 VGND.n2219 VGND.n2218 9.3005
R2872 VGND.n2287 VGND.n2286 9.3005
R2873 VGND.n2286 VGND.n2285 9.3005
R2874 VGND.n2279 VGND.n2278 9.3005
R2875 VGND.n2276 VGND.n1127 9.3005
R2876 VGND.n2275 VGND.n2274 9.3005
R2877 VGND.n2273 VGND.n1128 9.3005
R2878 VGND.n2272 VGND.n2271 9.3005
R2879 VGND.n2270 VGND.n1129 9.3005
R2880 VGND.n2268 VGND.n2267 9.3005
R2881 VGND.n2266 VGND.n1130 9.3005
R2882 VGND.n2265 VGND.n2264 9.3005
R2883 VGND.n2262 VGND.n1131 9.3005
R2884 VGND.n1143 VGND.n1142 9.3005
R2885 VGND.n1147 VGND.n1146 9.3005
R2886 VGND.n2250 VGND.n2249 9.3005
R2887 VGND.n2248 VGND.n1139 9.3005
R2888 VGND.n2247 VGND.n2246 9.3005
R2889 VGND.n2245 VGND.n1148 9.3005
R2890 VGND.n2244 VGND.n2243 9.3005
R2891 VGND.n2242 VGND.n1149 9.3005
R2892 VGND.n2240 VGND.n2239 9.3005
R2893 VGND.n2238 VGND.n2237 9.3005
R2894 VGND.n2236 VGND.n2235 9.3005
R2895 VGND.n2234 VGND.n2233 9.3005
R2896 VGND.n2232 VGND.n2231 9.3005
R2897 VGND.n2230 VGND.n2229 9.3005
R2898 VGND.n2228 VGND.n513 9.3005
R2899 VGND.n517 VGND.n514 9.3005
R2900 VGND.n2952 VGND.n2951 9.3005
R2901 VGND.n2950 VGND.n2949 9.3005
R2902 VGND.n2948 VGND.n518 9.3005
R2903 VGND.n2947 VGND.n2946 9.3005
R2904 VGND.n2944 VGND.n519 9.3005
R2905 VGND.n2943 VGND.n2942 9.3005
R2906 VGND.n2941 VGND.n520 9.3005
R2907 VGND.n2940 VGND.n2939 9.3005
R2908 VGND.n2891 VGND.n580 9.3005
R2909 VGND.n2894 VGND.n2893 9.3005
R2910 VGND.n2895 VGND.n579 9.3005
R2911 VGND.n2897 VGND.n2896 9.3005
R2912 VGND.n2899 VGND.n578 9.3005
R2913 VGND.n2901 VGND.n2900 9.3005
R2914 VGND.n2903 VGND.n2902 9.3005
R2915 VGND.n583 VGND.n581 9.3005
R2916 VGND.n2888 VGND.n2887 9.3005
R2917 VGND.n2886 VGND.n2885 9.3005
R2918 VGND.n2884 VGND.n584 9.3005
R2919 VGND.n2881 VGND.n2880 9.3005
R2920 VGND.n599 VGND.n595 9.3005
R2921 VGND.n663 VGND.n596 9.3005
R2922 VGND.n638 VGND.n637 9.3005
R2923 VGND.n620 VGND.n611 9.3005
R2924 VGND.n617 VGND.n616 9.3005
R2925 VGND.n623 VGND.n622 9.3005
R2926 VGND.n625 VGND.n624 9.3005
R2927 VGND.n636 VGND.n635 9.3005
R2928 VGND.n631 VGND.n629 9.3005
R2929 VGND.n605 VGND.n604 9.3005
R2930 VGND.n648 VGND.n647 9.3005
R2931 VGND.n649 VGND.n603 9.3005
R2932 VGND.n651 VGND.n650 9.3005
R2933 VGND.n652 VGND.n602 9.3005
R2934 VGND.n654 VGND.n653 9.3005
R2935 VGND.n657 VGND.n601 9.3005
R2936 VGND.n659 VGND.n658 9.3005
R2937 VGND.n660 VGND.n600 9.3005
R2938 VGND.n662 VGND.n661 9.3005
R2939 VGND.n665 VGND.n664 9.3005
R2940 VGND.n593 VGND.n585 9.3005
R2941 VGND.n2905 VGND.n2904 9.3005
R2942 VGND.n2914 VGND.n2913 9.3005
R2943 VGND.n2916 VGND.n2915 9.3005
R2944 VGND.n2065 VGND.n575 9.3005
R2945 VGND.n2067 VGND.n2066 9.3005
R2946 VGND.n2144 VGND.n2143 9.3005
R2947 VGND.n2143 VGND.n1186 9.3005
R2948 VGND.n2141 VGND.n2140 9.3005
R2949 VGND.n2139 VGND.n2138 9.3005
R2950 VGND.n2137 VGND.n1199 9.3005
R2951 VGND.n2136 VGND.n2135 9.3005
R2952 VGND.n2133 VGND.n2132 9.3005
R2953 VGND.n2130 VGND.n2129 9.3005
R2954 VGND.n1212 VGND.n1205 9.3005
R2955 VGND.n1217 VGND.n1214 9.3005
R2956 VGND.n2119 VGND.n2118 9.3005
R2957 VGND.n2116 VGND.n1215 9.3005
R2958 VGND.n2115 VGND.n2114 9.3005
R2959 VGND.n2113 VGND.n1218 9.3005
R2960 VGND.n2112 VGND.n2111 9.3005
R2961 VGND.n2110 VGND.n1219 9.3005
R2962 VGND.n2109 VGND.n2108 9.3005
R2963 VGND.n2107 VGND.n2106 9.3005
R2964 VGND.n2040 VGND.n2038 9.3005
R2965 VGND.n2103 VGND.n2102 9.3005
R2966 VGND.n2101 VGND.n2100 9.3005
R2967 VGND.n2098 VGND.n2097 9.3005
R2968 VGND.n2044 VGND.n2043 9.3005
R2969 VGND.n2054 VGND.n2052 9.3005
R2970 VGND.n2087 VGND.n2086 9.3005
R2971 VGND.n2056 VGND.n2053 9.3005
R2972 VGND.n2081 VGND.n2080 9.3005
R2973 VGND.n2079 VGND.n2058 9.3005
R2974 VGND.n2078 VGND.n2077 9.3005
R2975 VGND.n2076 VGND.n2059 9.3005
R2976 VGND.n2074 VGND.n2073 9.3005
R2977 VGND.n2072 VGND.n2061 9.3005
R2978 VGND.n2071 VGND.n2070 9.3005
R2979 VGND.n2068 VGND.n2062 9.3005
R2980 VGND.n2788 VGND.n694 9.3005
R2981 VGND.n2787 VGND.n2786 9.3005
R2982 VGND.n2783 VGND.n695 9.3005
R2983 VGND.n2782 VGND.n2781 9.3005
R2984 VGND.n2780 VGND.n2779 9.3005
R2985 VGND.n2778 VGND.n697 9.3005
R2986 VGND.n2777 VGND.n2776 9.3005
R2987 VGND.n2775 VGND.n698 9.3005
R2988 VGND.n2763 VGND.n2762 9.3005
R2989 VGND.n2766 VGND.n2765 9.3005
R2990 VGND.n2790 VGND.n2789 9.3005
R2991 VGND.n2793 VGND.n2792 9.3005
R2992 VGND.n2801 VGND.n2800 9.3005
R2993 VGND.n2804 VGND.n2803 9.3005
R2994 VGND.n685 VGND.n684 9.3005
R2995 VGND.n2813 VGND.n2812 9.3005
R2996 VGND.n2815 VGND.n683 9.3005
R2997 VGND.n2819 VGND.n2818 9.3005
R2998 VGND.n2820 VGND.n682 9.3005
R2999 VGND.n2821 VGND 9.3005
R3000 VGND.n2825 VGND.n2824 9.3005
R3001 VGND.n2827 VGND.n2826 9.3005
R3002 VGND.n2828 VGND.n679 9.3005
R3003 VGND.n2831 VGND.n2830 9.3005
R3004 VGND.n2832 VGND.n678 9.3005
R3005 VGND.n2834 VGND.n2833 9.3005
R3006 VGND.n2835 VGND.n676 9.3005
R3007 VGND.n2864 VGND.n2863 9.3005
R3008 VGND.n2862 VGND.n2861 9.3005
R3009 VGND.n2854 VGND.n2837 9.3005
R3010 VGND.n2853 VGND.n2852 9.3005
R3011 VGND.n2851 VGND.n2839 9.3005
R3012 VGND.n2849 VGND.n2848 9.3005
R3013 VGND.n2847 VGND.n2846 9.3005
R3014 VGND.n2668 VGND.n753 9.3005
R3015 VGND.n2664 VGND.n753 9.3005
R3016 VGND.n2681 VGND.n2680 9.3005
R3017 VGND.n2683 VGND.n2682 9.3005
R3018 VGND.n2684 VGND.n749 9.3005
R3019 VGND.n2688 VGND.n2687 9.3005
R3020 VGND.n2691 VGND.n2690 9.3005
R3021 VGND.n2693 VGND.n746 9.3005
R3022 VGND.n2695 VGND.n2694 9.3005
R3023 VGND.n2708 VGND.n2707 9.3005
R3024 VGND.n2710 VGND.n2709 9.3005
R3025 VGND.n2712 VGND.n2711 9.3005
R3026 VGND.n2713 VGND.n735 9.3005
R3027 VGND.n2716 VGND.n2715 9.3005
R3028 VGND.n2717 VGND.n734 9.3005
R3029 VGND.n2719 VGND.n2718 9.3005
R3030 VGND.n2720 VGND.n733 9.3005
R3031 VGND.n2723 VGND.n2722 9.3005
R3032 VGND.n2725 VGND.n2724 9.3005
R3033 VGND.n2727 VGND.n2726 9.3005
R3034 VGND.n2729 VGND.n2728 9.3005
R3035 VGND.n2730 VGND.n2729 9.3005
R3036 VGND.n2739 VGND.n716 9.3005
R3037 VGND.n2739 VGND.n2738 9.3005
R3038 VGND.n2741 VGND.n715 9.3005
R3039 VGND.n2744 VGND.n2743 9.3005
R3040 VGND.n2745 VGND.n714 9.3005
R3041 VGND.n2747 VGND.n2746 9.3005
R3042 VGND.n2748 VGND.n713 9.3005
R3043 VGND.n2750 VGND.n2749 9.3005
R3044 VGND.n2752 VGND.n2751 9.3005
R3045 VGND.n2753 VGND.n711 9.3005
R3046 VGND.n2756 VGND.n2755 9.3005
R3047 VGND.n2758 VGND.n2757 9.3005
R3048 VGND.n1494 VGND.n1493 9.3005
R3049 VGND.n1482 VGND.n1481 9.3005
R3050 VGND.n1479 VGND.n1478 9.3005
R3051 VGND.n1446 VGND.n1445 9.3005
R3052 VGND.n1437 VGND.n1436 9.3005
R3053 VGND.n1426 VGND.n1421 9.3005
R3054 VGND.n1428 VGND.n1427 9.3005
R3055 VGND.n1424 VGND.n767 9.3005
R3056 VGND.n1423 VGND.n768 9.3005
R3057 VGND.n2642 VGND.n2641 9.3005
R3058 VGND.n2640 VGND.n2639 9.3005
R3059 VGND.n2638 VGND.n2637 9.3005
R3060 VGND.n2636 VGND.n775 9.3005
R3061 VGND.n2633 VGND.n2632 9.3005
R3062 VGND.n2631 VGND.n777 9.3005
R3063 VGND.n2630 VGND.n2629 9.3005
R3064 VGND.n2627 VGND.n778 9.3005
R3065 VGND.n2624 VGND.n2623 9.3005
R3066 VGND.n2622 VGND.n2621 9.3005
R3067 VGND.n2619 VGND.n782 9.3005
R3068 VGND.n2618 VGND.n2617 9.3005
R3069 VGND.n786 VGND.n785 9.3005
R3070 VGND.n801 VGND.n800 9.3005
R3071 VGND.n802 VGND.n791 9.3005
R3072 VGND.n821 VGND.n820 9.3005
R3073 VGND.n818 VGND.n817 9.3005
R3074 VGND.n816 VGND.n815 9.3005
R3075 VGND.n814 VGND.n805 9.3005
R3076 VGND.n811 VGND.n810 9.3005
R3077 VGND.n1434 VGND.n1433 9.3005
R3078 VGND.n1435 VGND.n1420 9.3005
R3079 VGND.n1441 VGND.n1417 9.3005
R3080 VGND.n1443 VGND.n1442 9.3005
R3081 VGND.n1444 VGND.n1415 9.3005
R3082 VGND.n1447 VGND.n1414 9.3005
R3083 VGND.n1448 VGND.n1411 9.3005
R3084 VGND.n1450 VGND.n1449 9.3005
R3085 VGND.n1403 VGND.n1401 9.3005
R3086 VGND.n1459 VGND.n1458 9.3005
R3087 VGND.n1462 VGND.n1461 9.3005
R3088 VGND.n1463 VGND.n1398 9.3005
R3089 VGND.n1465 VGND.n1464 9.3005
R3090 VGND.n1466 VGND.n1395 9.3005
R3091 VGND.n1471 VGND.n1470 9.3005
R3092 VGND.n1472 VGND.n1394 9.3005
R3093 VGND.n1474 VGND.n1473 9.3005
R3094 VGND.n1477 VGND.n1390 9.3005
R3095 VGND.n1480 VGND.n1389 9.3005
R3096 VGND.n1486 VGND.n1485 9.3005
R3097 VGND.n1386 VGND.n1373 9.3005
R3098 VGND.n1495 VGND.n1371 9.3005
R3099 VGND.n1497 VGND.n1496 9.3005
R3100 VGND.n1498 VGND.n1369 9.3005
R3101 VGND.n1500 VGND.n1499 9.3005
R3102 VGND.n1501 VGND.n1367 9.3005
R3103 VGND.n1504 VGND.n1503 9.3005
R3104 VGND.n1505 VGND.n1366 9.3005
R3105 VGND.n1507 VGND.n1506 9.3005
R3106 VGND.n1508 VGND.n1364 9.3005
R3107 VGND.n1511 VGND.n1510 9.3005
R3108 VGND.n1512 VGND.n1363 9.3005
R3109 VGND.n1514 VGND.n1513 9.3005
R3110 VGND.n1518 VGND.n1517 9.3005
R3111 VGND.n1328 VGND.n1318 9.3005
R3112 VGND.n1329 VGND.n1328 9.3005
R3113 VGND.n1337 VGND.n1314 9.3005
R3114 VGND.n1339 VGND.n1338 9.3005
R3115 VGND.n1342 VGND.n1341 9.3005
R3116 VGND.n1344 VGND.n1343 9.3005
R3117 VGND.n1345 VGND.n1312 9.3005
R3118 VGND.n1348 VGND.n1347 9.3005
R3119 VGND.n1349 VGND.n1311 9.3005
R3120 VGND.n1351 VGND.n1350 9.3005
R3121 VGND.n1352 VGND.n1309 9.3005
R3122 VGND.n1355 VGND.n1354 9.3005
R3123 VGND.n1356 VGND.n1308 9.3005
R3124 VGND.n1358 VGND.n1357 9.3005
R3125 VGND.n1360 VGND.n1303 9.3005
R3126 VGND.n1362 VGND.n1304 9.3005
R3127 VGND.n1722 VGND.n1721 9.3005
R3128 VGND.n1721 VGND.n1539 9.3005
R3129 VGND.n1720 VGND.n1719 9.3005
R3130 VGND.n1718 VGND.n1717 9.3005
R3131 VGND.n1712 VGND.n1711 9.3005
R3132 VGND.n1710 VGND.n1550 9.3005
R3133 VGND.n1708 VGND.n1707 9.3005
R3134 VGND.n1706 VGND.n1705 9.3005
R3135 VGND.n1554 VGND.n1553 9.3005
R3136 VGND.n1699 VGND.n1698 9.3005
R3137 VGND.n1697 VGND.n1556 9.3005
R3138 VGND.n1696 VGND.n1695 9.3005
R3139 VGND.n1693 VGND.n1692 9.3005
R3140 VGND.n1570 VGND.n1569 9.3005
R3141 VGND.n1572 VGND.n1566 9.3005
R3142 VGND.n1682 VGND.n1681 9.3005
R3143 VGND.n1679 VGND.n1567 9.3005
R3144 VGND.n1677 VGND.n1676 9.3005
R3145 VGND.n1675 VGND.n1674 9.3005
R3146 VGND.n1672 VGND.n1576 9.3005
R3147 VGND.n1669 VGND.n1668 9.3005
R3148 VGND.n1667 VGND.n1666 9.3005
R3149 VGND.n1662 VGND.n1579 9.3005
R3150 VGND.n1661 VGND.n1660 9.3005
R3151 VGND.n1659 VGND.n1658 9.3005
R3152 VGND.n1657 VGND.n1584 9.3005
R3153 VGND.n1654 VGND.n1653 9.3005
R3154 VGND.n1589 VGND.n1587 9.3005
R3155 VGND.n1600 VGND.n1596 9.3005
R3156 VGND.n1643 VGND.n1642 9.3005
R3157 VGND.n1641 VGND.n1640 9.3005
R3158 VGND.n1639 VGND.n1601 9.3005
R3159 VGND.n1638 VGND.n1637 9.3005
R3160 VGND.n1636 VGND.n1602 9.3005
R3161 VGND.n1635 VGND.n1634 9.3005
R3162 VGND.n1633 VGND.n1606 9.3005
R3163 VGND.n1632 VGND.n1631 9.3005
R3164 VGND.n1630 VGND.n1607 9.3005
R3165 VGND.n1629 VGND.n1609 9.3005
R3166 VGND.n1628 VGND.n1627 9.3005
R3167 VGND.n1626 VGND.n1625 9.3005
R3168 VGND.n1624 VGND.n1623 9.3005
R3169 VGND.n1615 VGND.n835 9.3005
R3170 VGND.n2603 VGND.n2602 9.3005
R3171 VGND.n2600 VGND.n834 9.3005
R3172 VGND.n2599 VGND.n837 9.3005
R3173 VGND.n2598 VGND.n2597 9.3005
R3174 VGND.n2595 VGND.n2594 9.3005
R3175 VGND.n2592 VGND.n2591 9.3005
R3176 VGND.n2590 VGND.n845 9.3005
R3177 VGND.n2589 VGND.n2588 9.3005
R3178 VGND.n2587 VGND.n847 9.3005
R3179 VGND.n2586 VGND.n2585 9.3005
R3180 VGND.n850 VGND.n848 9.3005
R3181 VGND.n921 VGND.n920 9.3005
R3182 VGND.n919 VGND.n852 9.3005
R3183 VGND.n917 VGND.n855 9.3005
R3184 VGND.n916 VGND.n856 9.3005
R3185 VGND.n915 VGND.n914 9.3005
R3186 VGND.n913 VGND.n857 9.3005
R3187 VGND.n912 VGND.n911 9.3005
R3188 VGND.n910 VGND.n858 9.3005
R3189 VGND.n908 VGND.n907 9.3005
R3190 VGND.n906 VGND.n905 9.3005
R3191 VGND.n904 VGND.n862 9.3005
R3192 VGND.n903 VGND.n902 9.3005
R3193 VGND.n865 VGND.n863 9.3005
R3194 VGND.n876 VGND.n872 9.3005
R3195 VGND.n892 VGND.n891 9.3005
R3196 VGND.n889 VGND.n873 9.3005
R3197 VGND.n887 VGND.n881 9.3005
R3198 VGND.n1838 VGND.n1294 9.3005
R3199 VGND.n1838 VGND.n1293 9.3005
R3200 VGND.n1840 VGND.n1839 9.3005
R3201 VGND.n1842 VGND.n1841 9.3005
R3202 VGND.n1847 VGND.n1846 9.3005
R3203 VGND.n1848 VGND.n1289 9.3005
R3204 VGND.n1851 VGND.n1849 9.3005
R3205 VGND.n1852 VGND.n1287 9.3005
R3206 VGND.n1855 VGND.n1854 9.3005
R3207 VGND.n1856 VGND.n1286 9.3005
R3208 VGND.n1858 VGND.n1857 9.3005
R3209 VGND.n1860 VGND.n1859 9.3005
R3210 VGND.n1861 VGND.n1285 9.3005
R3211 VGND.n1863 VGND.n1862 9.3005
R3212 VGND.n1865 VGND.n1282 9.3005
R3213 VGND.n1868 VGND.n1867 9.3005
R3214 VGND.n1866 VGND.n1274 9.3005
R3215 VGND.n1880 VGND.n1273 9.3005
R3216 VGND.n1882 VGND.n1881 9.3005
R3217 VGND.n1884 VGND.n1883 9.3005
R3218 VGND.n1885 VGND.n1272 9.3005
R3219 VGND.n1887 VGND.n1886 9.3005
R3220 VGND.n1888 VGND.n1269 9.3005
R3221 VGND.n1893 VGND.n1892 9.3005
R3222 VGND.n1894 VGND.n1268 9.3005
R3223 VGND.n1915 VGND.n1895 9.3005
R3224 VGND.n1913 VGND.n1912 9.3005
R3225 VGND.n1911 VGND.n1896 9.3005
R3226 VGND.n1904 VGND.n1897 9.3005
R3227 VGND.n1906 VGND.n1905 9.3005
R3228 VGND.n1241 VGND.n1238 9.3005
R3229 VGND.n1980 VGND.n1979 9.3005
R3230 VGND.n1978 VGND.n1239 9.3005
R3231 VGND.n1976 VGND.n1975 9.3005
R3232 VGND.n1974 VGND.n1242 9.3005
R3233 VGND.n1973 VGND.n1972 9.3005
R3234 VGND.n1246 VGND.n1243 9.3005
R3235 VGND.n1967 VGND.n1966 9.3005
R3236 VGND.n1965 VGND.n1245 9.3005
R3237 VGND.n1964 VGND.n1963 9.3005
R3238 VGND.n1962 VGND.n1247 9.3005
R3239 VGND.n1961 VGND.n1960 9.3005
R3240 VGND.n1959 VGND.n1958 9.3005
R3241 VGND.n1957 VGND.n1956 9.3005
R3242 VGND.n1264 VGND.n1253 9.3005
R3243 VGND.n1948 VGND.n1947 9.3005
R3244 VGND.n1946 VGND.n1261 9.3005
R3245 VGND.n1944 VGND.n1943 9.3005
R3246 VGND.n1942 VGND.n1265 9.3005
R3247 VGND.n1941 VGND.n1940 9.3005
R3248 VGND.n1936 VGND.n1266 9.3005
R3249 VGND.n1935 VGND.n1934 9.3005
R3250 VGND.n1933 VGND.n1267 9.3005
R3251 VGND.n1932 VGND.n1931 9.3005
R3252 VGND.n1930 VGND.n1929 9.3005
R3253 VGND.n1928 VGND.n1927 9.3005
R3254 VGND.n1924 VGND.n1923 9.3005
R3255 VGND.n1922 VGND.n929 9.3005
R3256 VGND.n1920 VGND.n930 9.3005
R3257 VGND.n2561 VGND.n2560 9.3005
R3258 VGND.n2559 VGND.n935 9.3005
R3259 VGND.n2558 VGND.n2557 9.3005
R3260 VGND.n2556 VGND.n2555 9.3005
R3261 VGND.n2554 VGND.n938 9.3005
R3262 VGND.n2553 VGND.n2552 9.3005
R3263 VGND.n2551 VGND.n940 9.3005
R3264 VGND.n2550 VGND.n2549 9.3005
R3265 VGND.n2548 VGND.n941 9.3005
R3266 VGND.n2547 VGND.n2546 9.3005
R3267 VGND.n2545 VGND.n2544 9.3005
R3268 VGND.n2540 VGND.n945 9.3005
R3269 VGND.n2538 VGND.n2537 9.3005
R3270 VGND.n961 VGND.n950 9.3005
R3271 VGND.n962 VGND.n958 9.3005
R3272 VGND.n978 VGND.n977 9.3005
R3273 VGND.n976 VGND.n959 9.3005
R3274 VGND.n975 VGND.n974 9.3005
R3275 VGND.n973 VGND.n972 9.3005
R3276 VGND.n970 VGND.n965 9.3005
R3277 VGND.n2440 VGND.n2439 9.3005
R3278 VGND.n2442 VGND.n2441 9.3005
R3279 VGND.n1744 VGND.n1742 9.3005
R3280 VGND.n1757 VGND.n1756 9.3005
R3281 VGND.n1825 VGND.n1824 9.3005
R3282 VGND.n1823 VGND.n1759 9.3005
R3283 VGND.n1822 VGND.n1821 9.3005
R3284 VGND.n1820 VGND.n1760 9.3005
R3285 VGND.n1819 VGND.n1818 9.3005
R3286 VGND.n1817 VGND.n1761 9.3005
R3287 VGND.n1816 VGND.n1815 9.3005
R3288 VGND.n1814 VGND.n1813 9.3005
R3289 VGND.n1812 VGND.n1764 9.3005
R3290 VGND.n1809 VGND.n1808 9.3005
R3291 VGND.n1807 VGND.n1765 9.3005
R3292 VGND.n1806 VGND.n1805 9.3005
R3293 VGND.n1804 VGND.n1803 9.3005
R3294 VGND.n1775 VGND.n1768 9.3005
R3295 VGND.n1779 VGND.n1777 9.3005
R3296 VGND.n1793 VGND.n1792 9.3005
R3297 VGND.n1791 VGND.n1778 9.3005
R3298 VGND.n1788 VGND.n1787 9.3005
R3299 VGND.n1786 VGND.n1784 9.3005
R3300 VGND.n1785 VGND.n1223 9.3005
R3301 VGND.n2029 VGND.n1224 9.3005
R3302 VGND.n2028 VGND.n2027 9.3005
R3303 VGND.n2026 VGND.n2025 9.3005
R3304 VGND.n2024 VGND.n2023 9.3005
R3305 VGND.n2012 VGND.n1229 9.3005
R3306 VGND.n2012 VGND.n1990 9.3005
R3307 VGND.n2013 VGND.n2012 9.3005
R3308 VGND.n2011 VGND.n2010 9.3005
R3309 VGND.n2009 VGND.n1992 9.3005
R3310 VGND.n2008 VGND.n2007 9.3005
R3311 VGND.n2006 VGND.n2005 9.3005
R3312 VGND.n2004 VGND.n1993 9.3005
R3313 VGND.n2003 VGND.n2002 9.3005
R3314 VGND.n2001 VGND.n1994 9.3005
R3315 VGND.n1997 VGND.n989 9.3005
R3316 VGND.n2520 VGND.n2519 9.3005
R3317 VGND.n2518 VGND.n2517 9.3005
R3318 VGND.n2512 VGND.n991 9.3005
R3319 VGND.n2511 VGND.n2510 9.3005
R3320 VGND.n2508 VGND.n995 9.3005
R3321 VGND.n2507 VGND.n2506 9.3005
R3322 VGND.n2505 VGND.n2504 9.3005
R3323 VGND.n2503 VGND.n2502 9.3005
R3324 VGND.n2501 VGND.n999 9.3005
R3325 VGND.n2500 VGND.n2499 9.3005
R3326 VGND.n2498 VGND.n2396 9.3005
R3327 VGND.n2497 VGND.n2496 9.3005
R3328 VGND.n2495 VGND.n2494 9.3005
R3329 VGND.n2493 VGND.n2398 9.3005
R3330 VGND.n2492 VGND.n2491 9.3005
R3331 VGND.n2407 VGND.n2399 9.3005
R3332 VGND.n2475 VGND.n2409 9.3005
R3333 VGND.n2481 VGND.n2480 9.3005
R3334 VGND.n2473 VGND.n2410 9.3005
R3335 VGND.n2472 VGND.n2471 9.3005
R3336 VGND.n2470 VGND.n2413 9.3005
R3337 VGND.n2469 VGND.n2468 9.3005
R3338 VGND.n2467 VGND.n2466 9.3005
R3339 VGND.n2465 VGND.n2414 9.3005
R3340 VGND.n2464 VGND.n2463 9.3005
R3341 VGND.n2462 VGND.n2415 9.3005
R3342 VGND.n2460 VGND.n2418 9.3005
R3343 VGND.n2459 VGND.n2458 9.3005
R3344 VGND.n2431 VGND.n2421 9.3005
R3345 VGND.n2450 VGND.n2449 9.3005
R3346 VGND.n2448 VGND.n2447 9.3005
R3347 VGND.n2446 VGND.n2432 9.3005
R3348 VGND.n2445 VGND.n2444 9.3005
R3349 VGND.n2443 VGND.n2433 9.3005
R3350 VGND.n244 VGND.n241 9.3005
R3351 VGND.n255 VGND.n254 9.3005
R3352 VGND.n3041 VGND.n3040 9.3005
R3353 VGND.n3038 VGND.n239 9.3005
R3354 VGND.n3035 VGND.n3034 9.3005
R3355 VGND.n3033 VGND.n256 9.3005
R3356 VGND.n3032 VGND.n3031 9.3005
R3357 VGND.n3030 VGND.n257 9.3005
R3358 VGND.n3029 VGND.n3028 9.3005
R3359 VGND.n3027 VGND.n259 9.3005
R3360 VGND.n3026 VGND.n3025 9.3005
R3361 VGND.n262 VGND.n260 9.3005
R3362 VGND.n3020 VGND.n3019 9.3005
R3363 VGND.n3018 VGND.n264 9.3005
R3364 VGND.n272 VGND.n265 9.3005
R3365 VGND.n3010 VGND.n3009 9.3005
R3366 VGND.n3008 VGND.n3007 9.3005
R3367 VGND.n3001 VGND.n273 9.3005
R3368 VGND.n3000 VGND.n2999 9.3005
R3369 VGND.n2998 VGND.n274 9.3005
R3370 VGND.n2997 VGND.n2996 9.3005
R3371 VGND.n2995 VGND.n2994 9.3005
R3372 VGND.n2993 VGND.n276 9.3005
R3373 VGND.n2992 VGND.n2991 9.3005
R3374 VGND.n2990 VGND.n2989 9.3005
R3375 VGND.n2988 VGND.n279 9.3005
R3376 VGND.n1058 VGND.n278 9.3005
R3377 VGND.n1063 VGND.n1062 9.3005
R3378 VGND.n1065 VGND.n1055 9.3005
R3379 VGND.n1074 VGND.n1073 9.3005
R3380 VGND.n1076 VGND.n1053 9.3005
R3381 VGND.n1113 VGND.n1112 9.3005
R3382 VGND.n1111 VGND.n1054 9.3005
R3383 VGND.n1110 VGND.n1109 9.3005
R3384 VGND.n1108 VGND.n1077 9.3005
R3385 VGND.n1107 VGND.n1106 9.3005
R3386 VGND.n1105 VGND.n1078 9.3005
R3387 VGND.n1103 VGND.n1102 9.3005
R3388 VGND.n1101 VGND.n1079 9.3005
R3389 VGND.n1100 VGND.n1099 9.3005
R3390 VGND.n1097 VGND 9.3005
R3391 VGND.n1096 VGND.n1095 9.3005
R3392 VGND.n1094 VGND.n1093 9.3005
R3393 VGND.n1092 VGND.n1091 9.3005
R3394 VGND.n1084 VGND.n1082 9.3005
R3395 VGND.n2972 VGND.n499 9.3005
R3396 VGND.n2974 VGND.n2973 9.3005
R3397 VGND.n2975 VGND.n498 9.3005
R3398 VGND.n2977 VGND.n2976 9.3005
R3399 VGND.n2979 VGND.n2978 9.3005
R3400 VGND.n2980 VGND.n496 9.3005
R3401 VGND.n2982 VGND.n2981 9.3005
R3402 VGND.n2984 VGND.n2983 9.3005
R3403 VGND.n2985 VGND.n494 9.3005
R3404 VGND.n1040 VGND.n493 9.3005
R3405 VGND.n1042 VGND.n1041 9.3005
R3406 VGND.n1044 VGND.n1043 9.3005
R3407 VGND.n2314 VGND.n2313 9.3005
R3408 VGND.n2316 VGND.n2315 9.3005
R3409 VGND.n1036 VGND.n1035 9.3005
R3410 VGND.n2322 VGND.n2321 9.3005
R3411 VGND.n2323 VGND.n1033 9.3005
R3412 VGND.n2329 VGND.n2328 9.3005
R3413 VGND.n2331 VGND.n2330 9.3005
R3414 VGND.n2333 VGND.n2332 9.3005
R3415 VGND.n2334 VGND.n1031 9.3005
R3416 VGND.n2336 VGND.n2335 9.3005
R3417 VGND.n2337 VGND.n1029 9.3005
R3418 VGND.n2340 VGND.n2339 9.3005
R3419 VGND.n2341 VGND.n1028 9.3005
R3420 VGND.n2343 VGND.n2342 9.3005
R3421 VGND.n2344 VGND.n1025 9.3005
R3422 VGND.n2371 VGND.n2370 9.3005
R3423 VGND.n2369 VGND.n2368 9.3005
R3424 VGND.n2366 VGND.n2345 9.3005
R3425 VGND.n2365 VGND.n2364 9.3005
R3426 VGND.n2363 VGND.n2348 9.3005
R3427 VGND.n2362 VGND.n2361 9.3005
R3428 VGND.n2360 VGND.n2359 9.3005
R3429 VGND.n2358 VGND.n2357 9.3005
R3430 VGND.n2356 VGND.n2355 9.3005
R3431 VGND.n1446 VGND.n1415 9.12791
R3432 VGND.n1477 VGND.n1476 9.03579
R3433 VGND.n1393 VGND.n1392 9.03579
R3434 VGND.n1674 VGND.n1575 9.03579
R3435 VGND.n2626 VGND.n2624 8.9684
R3436 VGND.n328 VGND.n327 8.44328
R3437 VGND.n350 VGND.n349 8.44328
R3438 VGND.n3220 VGND.n3219 8.44328
R3439 VGND.n3274 VGND.n3273 8.44328
R3440 VGND.t594 VGND.t94 8.42962
R3441 VGND.t552 VGND.t474 8.42962
R3442 VGND.t196 VGND.t1082 8.42962
R3443 VGND VGND.n3406 8.3721
R3444 VGND.n331 VGND.n330 8.33966
R3445 VGND.n3384 VGND.n3383 8.33966
R3446 VGND.n200 VGND.n181 8.31061
R3447 VGND.n3054 VGND.n227 8.30267
R3448 VGND.n918 VGND.n917 8.28285
R3449 VGND.n2223 VGND.n1153 8.23546
R3450 VGND.n2934 VGND.n2933 8.23546
R3451 VGND.n2933 VGND.n2932 8.23546
R3452 VGND.n2932 VGND.n526 8.23546
R3453 VGND.n562 VGND.n545 8.23546
R3454 VGND.n2830 VGND.n678 8.23546
R3455 VGND.n2834 VGND.n678 8.23546
R3456 VGND.n2803 VGND.n684 8.23546
R3457 VGND.n2813 VGND.n684 8.23546
R3458 VGND.n2821 VGND.n682 8.23546
R3459 VGND.n2824 VGND.n2821 8.23546
R3460 VGND.n2726 VGND.n2725 8.23546
R3461 VGND.n2619 VGND.n2618 8.23546
R3462 VGND.n2618 VGND.n785 8.23546
R3463 VGND.n802 VGND.n801 8.23546
R3464 VGND.n1424 VGND.n1423 8.23546
R3465 VGND.n2641 VGND.n2640 8.23546
R3466 VGND.n2637 VGND.n2636 8.23546
R3467 VGND.n2633 VGND.n777 8.23546
R3468 VGND.n1352 VGND.n1351 8.23546
R3469 VGND.n1354 VGND.n1352 8.23546
R3470 VGND.n1358 VGND.n1308 8.23546
R3471 VGND.n1514 VGND.n1363 8.23546
R3472 VGND.n1510 VGND.n1363 8.23546
R3473 VGND.n1508 VGND.n1507 8.23546
R3474 VGND.n1507 VGND.n1366 8.23546
R3475 VGND.n1503 VGND.n1366 8.23546
R3476 VGND.n1501 VGND.n1500 8.23546
R3477 VGND.n1500 VGND.n1369 8.23546
R3478 VGND.n1967 VGND.n1245 8.23546
R3479 VGND.n1963 VGND.n1245 8.23546
R3480 VGND.n1963 VGND.n1962 8.23546
R3481 VGND.n1962 VGND.n1961 8.23546
R3482 VGND.n1958 VGND.n1957 8.23546
R3483 VGND.n1947 VGND.n1264 8.23546
R3484 VGND.n1947 VGND.n1946 8.23546
R3485 VGND.n2339 VGND.n1028 8.23546
R3486 VGND.n2343 VGND.n1028 8.23546
R3487 VGND.n2344 VGND.n2343 8.23546
R3488 VGND.n2370 VGND.n2344 8.23546
R3489 VGND.n2370 VGND.n2369 8.23546
R3490 VGND.n2369 VGND.n2345 8.23546
R3491 VGND.n2364 VGND.n2363 8.23546
R3492 VGND.n2363 VGND.n2362 8.23546
R3493 VGND.n1093 VGND.n1092 8.23546
R3494 VGND.n1092 VGND.n1082 8.23546
R3495 VGND.n1082 VGND.n499 8.23546
R3496 VGND.n2974 VGND.n499 8.23546
R3497 VGND.n2975 VGND.n2974 8.23546
R3498 VGND.n2976 VGND.n2975 8.23546
R3499 VGND.n2980 VGND.n2979 8.23546
R3500 VGND.n2981 VGND.n2980 8.23546
R3501 VGND.n1112 VGND.n1076 8.23546
R3502 VGND.n1112 VGND.n1111 8.23546
R3503 VGND.n1111 VGND.n1110 8.23546
R3504 VGND.n1110 VGND.n1077 8.23546
R3505 VGND.n1106 VGND.n1077 8.23546
R3506 VGND.n1106 VGND.n1105 8.23546
R3507 VGND.n1103 VGND.n1079 8.23546
R3508 VGND.n1099 VGND.n1079 8.23546
R3509 VGND.n3009 VGND.n272 8.23546
R3510 VGND.n3009 VGND.n3008 8.23546
R3511 VGND.n3008 VGND.n273 8.23546
R3512 VGND.n2999 VGND.n273 8.23546
R3513 VGND.n2999 VGND.n2998 8.23546
R3514 VGND.n2998 VGND.n2997 8.23546
R3515 VGND.n2994 VGND.n2993 8.23546
R3516 VGND.n2993 VGND.n2992 8.23546
R3517 VGND.n2815 VGND.n2814 8.14595
R3518 VGND.n537 VGND.n536 8.05644
R3519 VGND.n329 VGND.n287 7.97888
R3520 VGND.n374 VGND.n228 7.97888
R3521 VGND.n3240 VGND.n78 7.97888
R3522 VGND.n3201 VGND.n3200 7.97888
R3523 VGND.n328 VGND.n288 7.97601
R3524 VGND.n351 VGND.n350 7.97601
R3525 VGND.n3273 VGND.n3272 7.97601
R3526 VGND.n3221 VGND.n3220 7.97601
R3527 VGND.n1470 VGND.n1469 7.90638
R3528 VGND.n1628 VGND.n1612 7.90638
R3529 VGND.n2549 VGND.n943 7.90638
R3530 VGND.n1360 VGND.n1359 7.78791
R3531 VGND.n1970 VGND.n1969 7.72113
R3532 VGND.n2236 VGND.n2226 7.6984
R3533 VGND.n2934 VGND.n525 7.6984
R3534 VGND.n2830 VGND.n2829 7.6984
R3535 VGND.n2818 VGND.n2816 7.6984
R3536 VGND.n2621 VGND.n781 7.6984
R3537 VGND.n1429 VGND.n1428 7.6984
R3538 VGND.n1428 VGND.n1425 7.6984
R3539 VGND.n2629 VGND.n2628 7.6984
R3540 VGND.n1361 VGND.n1360 7.6984
R3541 VGND.n1370 VGND.n1369 7.6984
R3542 VGND.n1968 VGND.n1967 7.6984
R3543 VGND.n1946 VGND.n1945 7.6984
R3544 VGND.n2339 VGND.n2338 7.6984
R3545 VGND.n2362 VGND.n2350 7.6984
R3546 VGND.n1093 VGND.n1080 7.6984
R3547 VGND.n2981 VGND.n495 7.6984
R3548 VGND.n1076 VGND.n1075 7.6984
R3549 VGND.n1099 VGND.n1098 7.6984
R3550 VGND.n272 VGND.n271 7.6984
R3551 VGND.n2992 VGND.n277 7.6984
R3552 VGND.n3144 VGND.n212 7.64725
R3553 VGND.n3169 VGND.n3167 7.64725
R3554 VGND.n3089 VGND.n221 7.64725
R3555 VGND.n3108 VGND.n3107 7.64725
R3556 VGND.n948 VGND.n947 7.6005
R3557 VGND.n1509 VGND.n1508 7.51938
R3558 VGND.n2824 VGND.n2823 7.34036
R3559 VGND.n1958 VGND.n1249 7.34036
R3560 VGND.n793 VGND.n785 7.25085
R3561 VGND.n1516 VGND.n1515 7.25085
R3562 VGND.n390 VGND.n227 7.16724
R3563 VGND.n3241 VGND.n3240 7.16724
R3564 VGND.n3272 VGND.n3271 7.16724
R3565 VGND.n3223 VGND.n3221 7.16724
R3566 VGND.n3219 VGND.n3218 7.16724
R3567 VGND.n3200 VGND.n3199 7.16724
R3568 VGND.n3385 VGND.n3384 7.16724
R3569 VGND.n3275 VGND.n3274 7.16724
R3570 VGND.n2620 VGND.n2619 7.16134
R3571 VGND.n3461 VGND.n3460 7.15344
R3572 VGND.n3329 VGND.n113 7.15344
R3573 VGND.n2237 VGND.n2236 7.11268
R3574 VGND.n2790 VGND.n694 7.11268
R3575 VGND.n537 VGND.n533 6.98232
R3576 VGND.n2835 VGND.n2834 6.88949
R3577 VGND.n1351 VGND.n1311 6.88949
R3578 VGND.n1423 VGND.n772 6.62428
R3579 VGND.n2286 VGND.n1125 6.61527
R3580 VGND.n2739 VGND.n718 6.61527
R3581 VGND.n2382 VGND.t395 6.6005
R3582 VGND.n2382 VGND.t391 6.6005
R3583 VGND.n2384 VGND.t563 6.6005
R3584 VGND.n2384 VGND.t760 6.6005
R3585 VGND.n1017 VGND.t393 6.6005
R3586 VGND.n1017 VGND.t473 6.6005
R3587 VGND.n2219 VGND.n1125 6.57117
R3588 VGND.n2729 VGND.n718 6.57117
R3589 VGND.n1714 VGND.n1549 6.57117
R3590 VGND.n1716 VGND.n1714 6.57117
R3591 VGND.n803 VGND.n802 6.53477
R3592 VGND.n3449 VGND.n3448 6.50373
R3593 VGND.n3104 VGND.n209 6.50373
R3594 VGND.n3357 VGND.n3355 6.50373
R3595 VGND.n49 VGND.n48 6.4005
R3596 VGND.n3311 VGND.n3310 6.4005
R3597 VGND.n1939 VGND.n1936 6.4005
R3598 VGND.n1922 VGND.n1921 6.4005
R3599 VGND.n56 VGND.n55 6.26433
R3600 VGND.n3441 VGND.n3440 6.26433
R3601 VGND.n3304 VGND.n3303 6.26433
R3602 VGND.n103 VGND.n102 6.26433
R3603 VGND.n1442 VGND.n1441 6.26433
R3604 VGND.n1711 VGND.n1710 6.26433
R3605 VGND.n1846 VGND.n1842 6.26433
R3606 VGND.n1813 VGND.n1812 6.26433
R3607 VGND.n1792 VGND.n1791 6.26433
R3608 VGND.n2025 VGND.n2024 6.26433
R3609 VGND.n2002 VGND.n2001 6.26433
R3610 VGND.n2508 VGND.n2507 6.26433
R3611 VGND.n2494 VGND.n2493 6.26433
R3612 VGND.n2493 VGND.n2492 6.26433
R3613 VGND.n2463 VGND.n2462 6.26433
R3614 VGND.n2315 VGND.n2314 6.26433
R3615 VGND.n2315 VGND.n1035 6.26433
R3616 VGND.n3031 VGND.n3030 6.26433
R3617 VGND.n3030 VGND.n3029 6.26433
R3618 VGND.n890 VGND.n889 6.12816
R3619 VGND.n622 VGND.n621 6.06007
R3620 VGND.n315 VGND.n295 6.05269
R3621 VGND.n305 VGND.n301 6.05269
R3622 VGND.n326 VGND.n325 6.05269
R3623 VGND.n336 VGND.n332 6.05269
R3624 VGND.n380 VGND.n375 6.05269
R3625 VGND.n357 VGND.n352 6.05269
R3626 VGND.n364 VGND.n345 6.05269
R3627 VGND.n202 VGND.n201 6.05269
R3628 VGND.n2202 VGND.n2201 6.02861
R3629 VGND.n2118 VGND.n1217 6.02861
R3630 VGND.n2068 VGND.n2067 6.02861
R3631 VGND.n2904 VGND.n2903 6.02861
R3632 VGND.n2709 VGND.n2708 6.02861
R3633 VGND.n1476 VGND.n1474 6.02403
R3634 VGND.n1484 VGND.n1483 6.02403
R3635 VGND.n1666 VGND.n1578 5.98311
R3636 VGND.n1927 VGND.n1918 5.98311
R3637 VGND.n2544 VGND.n944 5.98311
R3638 VGND.n1744 VGND.n1741 5.98311
R3639 VGND.n2439 VGND.n2435 5.98311
R3640 VGND.n2355 VGND.n2351 5.98311
R3641 VGND.n1062 VGND.n1059 5.98311
R3642 VGND.n3039 VGND.n3038 5.98311
R3643 VGND.n244 VGND.n240 5.98311
R3644 VGND.n55 VGND.n42 5.85582
R3645 VGND.n3441 VGND.n40 5.85582
R3646 VGND.n32 VGND.n31 5.85582
R3647 VGND.n6 VGND.n3 5.85582
R3648 VGND.n10 VGND.n7 5.85582
R3649 VGND.n3305 VGND.n3304 5.85582
R3650 VGND.n103 VGND.n97 5.85582
R3651 VGND.n3319 VGND.n115 5.85582
R3652 VGND.n3321 VGND.n3320 5.85582
R3653 VGND.n3349 VGND.n3341 5.85582
R3654 VGND.n622 VGND.n610 5.85582
R3655 VGND.n1442 VGND.n1418 5.85582
R3656 VGND.n1717 VGND.n1541 5.85582
R3657 VGND.n891 VGND.n877 5.85582
R3658 VGND.n1842 VGND.n1290 5.85582
R3659 VGND.n961 VGND.n960 5.85582
R3660 VGND.n1813 VGND.n1763 5.85582
R3661 VGND.n1792 VGND.n1780 5.85582
R3662 VGND.n2025 VGND.n1225 5.85582
R3663 VGND.n2002 VGND.n1995 5.85582
R3664 VGND.n2509 VGND.n2508 5.85582
R3665 VGND.n2494 VGND.n2397 5.85582
R3666 VGND.n2463 VGND.n2416 5.85582
R3667 VGND.n2314 VGND.n1039 5.85582
R3668 VGND.n3031 VGND.n258 5.85582
R3669 VGND.n2492 VGND.n2399 5.65809
R3670 VGND.n2322 VGND.n1035 5.65809
R3671 VGND.n3029 VGND.n259 5.65809
R3672 VGND.n2217 VGND.n1153 5.63966
R3673 VGND.n2803 VGND.n2802 5.63966
R3674 VGND.n2791 VGND.n2790 5.63966
R3675 VGND.n2726 VGND.n730 5.63966
R3676 VGND.n2890 VGND.n581 5.5878
R3677 VGND.n2640 VGND.n774 5.55015
R3678 VGND.n2104 VGND.n2038 5.48621
R3679 VGND.n2081 VGND.n2058 5.48128
R3680 VGND.n962 VGND.n961 5.37524
R3681 VGND.n2594 VGND.n2593 5.27109
R3682 VGND.n1709 VGND.n1708 5.24958
R3683 VGND.n1174 VGND.n1172 5.13108
R3684 VGND.n1174 VGND.n1173 5.13108
R3685 VGND.n2172 VGND.n1175 5.13108
R3686 VGND.n2172 VGND.n2171 5.13108
R3687 VGND.n550 VGND.n548 5.13108
R3688 VGND.n550 VGND.n549 5.13108
R3689 VGND.n2143 VGND.n1185 5.13108
R3690 VGND.n2143 VGND.n1187 5.13108
R3691 VGND.n2142 VGND.n1188 5.13108
R3692 VGND.n2142 VGND.n1197 5.13108
R3693 VGND.n614 VGND.n612 5.13108
R3694 VGND.n614 VGND.n613 5.13108
R3695 VGND.n2845 VGND.n2842 5.13108
R3696 VGND.n2845 VGND.n2844 5.13108
R3697 VGND.n753 VGND.n751 5.13108
R3698 VGND.n753 VGND.n752 5.13108
R3699 VGND.n2679 VGND.n754 5.13108
R3700 VGND.n2679 VGND.n2678 5.13108
R3701 VGND.n1328 VGND.n1320 5.13108
R3702 VGND.n1328 VGND.n1321 5.13108
R3703 VGND.n808 VGND.n806 5.13108
R3704 VGND.n808 VGND.n807 5.13108
R3705 VGND.n1721 VGND.n1538 5.13108
R3706 VGND.n1721 VGND.n1540 5.13108
R3707 VGND.n886 VGND.n883 5.13108
R3708 VGND.n886 VGND.n884 5.13108
R3709 VGND.n1838 VGND.n1292 5.13108
R3710 VGND.n1838 VGND.n1837 5.13108
R3711 VGND.n969 VGND.n966 5.13108
R3712 VGND.n969 VGND.n967 5.13108
R3713 VGND.n2629 VGND.n780 4.92358
R3714 VGND.n2987 VGND.n492 4.89029
R3715 VGND.n2084 VGND.n2057 4.85762
R3716 VGND.n1702 VGND.n1555 4.85762
R3717 VGND.n2478 VGND.n2477 4.85762
R3718 VGND.n3023 VGND.n263 4.85762
R3719 VGND.n2326 VGND.n2325 4.85762
R3720 VGND.n1927 VGND.n1926 4.8005
R3721 VGND.n1745 VGND.n1744 4.8005
R3722 VGND.n2439 VGND.n2438 4.8005
R3723 VGND.n2355 VGND.n2354 4.8005
R3724 VGND.n1062 VGND.n1061 4.8005
R3725 VGND.n3038 VGND.n3037 4.8005
R3726 VGND.n245 VGND.n244 4.8005
R3727 VGND.n3448 VGND.n36 4.788
R3728 VGND.n209 VGND.n194 4.788
R3729 VGND.n3358 VGND.n3357 4.788
R3730 VGND.n2261 VGND.n2260 4.72533
R3731 VGND.n2760 VGND.n2759 4.72533
R3732 VGND.n2187 VGND.n2186 4.67352
R3733 VGND.n2206 VGND.n2205 4.67352
R3734 VGND.n2208 VGND.n2206 4.67352
R3735 VGND.n2212 VGND.n1155 4.67352
R3736 VGND.n2213 VGND.n2212 4.67352
R3737 VGND.n2276 VGND.n2275 4.67352
R3738 VGND.n2275 VGND.n1128 4.67352
R3739 VGND.n2271 VGND.n1128 4.67352
R3740 VGND.n2271 VGND.n2270 4.67352
R3741 VGND.n2268 VGND.n1130 4.67352
R3742 VGND.n2249 VGND.n1147 4.67352
R3743 VGND.n2249 VGND.n2248 4.67352
R3744 VGND.n2248 VGND.n2247 4.67352
R3745 VGND.n2247 VGND.n1148 4.67352
R3746 VGND.n2243 VGND.n2242 4.67352
R3747 VGND.n2229 VGND.n2228 4.67352
R3748 VGND.n2228 VGND.n517 4.67352
R3749 VGND.n2951 VGND.n517 4.67352
R3750 VGND.n2951 VGND.n2950 4.67352
R3751 VGND.n2950 VGND.n518 4.67352
R3752 VGND.n2946 VGND.n518 4.67352
R3753 VGND.n2944 VGND.n2943 4.67352
R3754 VGND.n2943 VGND.n520 4.67352
R3755 VGND.n2130 VGND.n1205 4.67352
R3756 VGND.n2116 VGND.n2115 4.67352
R3757 VGND.n2115 VGND.n1218 4.67352
R3758 VGND.n2111 VGND.n2110 4.67352
R3759 VGND.n2110 VGND.n2109 4.67352
R3760 VGND.n2077 VGND.n2076 4.67352
R3761 VGND.n2074 VGND.n2061 4.67352
R3762 VGND.n2070 VGND.n2061 4.67352
R3763 VGND.n2915 VGND.n575 4.67352
R3764 VGND.n2915 VGND.n2914 4.67352
R3765 VGND.n2900 VGND.n2899 4.67352
R3766 VGND.n2897 VGND.n579 4.67352
R3767 VGND.n2893 VGND.n579 4.67352
R3768 VGND.n2694 VGND.n2693 4.67352
R3769 VGND.n2713 VGND.n2712 4.67352
R3770 VGND.n2715 VGND.n2713 4.67352
R3771 VGND.n2719 VGND.n734 4.67352
R3772 VGND.n2720 VGND.n2719 4.67352
R3773 VGND.n2743 VGND.n714 4.67352
R3774 VGND.n2747 VGND.n714 4.67352
R3775 VGND.n2748 VGND.n2747 4.67352
R3776 VGND.n2749 VGND.n2748 4.67352
R3777 VGND.n2753 VGND.n2752 4.67352
R3778 VGND.n2763 VGND.n698 4.67352
R3779 VGND.n2777 VGND.n698 4.67352
R3780 VGND.n2778 VGND.n2777 4.67352
R3781 VGND.n2779 VGND.n2778 4.67352
R3782 VGND.n2783 VGND.n2782 4.67352
R3783 VGND.n2286 VGND.n1123 4.63943
R3784 VGND.n2260 VGND.n1133 4.63943
R3785 VGND.n2740 VGND.n2739 4.63943
R3786 VGND.n2761 VGND.n2760 4.63943
R3787 VGND.n887 VGND.n880 4.62124
R3788 VGND.n2460 VGND.n2419 4.62124
R3789 VGND.n2260 VGND.n2259 4.62124
R3790 VGND.n2801 VGND.n2794 4.62124
R3791 VGND.n2760 VGND.n709 4.62124
R3792 VGND.n1714 VGND.n1713 4.62124
R3793 VGND.n2219 VGND.n2217 4.6085
R3794 VGND.n2729 VGND.n730 4.6085
R3795 VGND.n2262 VGND.n2261 4.60638
R3796 VGND.n2759 VGND.n2758 4.60638
R3797 VGND.n473 VGND.n472 4.5578
R3798 VGND.n2278 VGND.n1123 4.55559
R3799 VGND.n1142 VGND.n1133 4.55559
R3800 VGND.n2741 VGND.n2740 4.55559
R3801 VGND.n2765 VGND.n2761 4.55559
R3802 VGND.n1460 VGND.n1459 4.51815
R3803 VGND.n1469 VGND.n1394 4.51815
R3804 VGND.n1680 VGND.n1679 4.51815
R3805 VGND.n1656 VGND.n1655 4.51815
R3806 VGND.n1915 VGND.n1914 4.51815
R3807 VGND.n1046 VGND.n1045 4.51401
R3808 VGND.n2320 VGND.n2319 4.51401
R3809 VGND.n247 VGND.n243 4.51401
R3810 VGND.n3043 VGND.n3042 4.51401
R3811 VGND.n2570 VGND.n927 4.51401
R3812 VGND.n932 VGND.n931 4.51401
R3813 VGND.n1064 VGND.n1057 4.51401
R3814 VGND.n1115 VGND.n1114 4.51401
R3815 VGND.n2578 VGND.n846 4.51401
R3816 VGND.n2582 VGND.n922 4.51401
R3817 VGND.n1085 VGND.n1081 4.51401
R3818 VGND.n2971 VGND.n2970 4.51401
R3819 VGND.n2961 VGND.n511 4.51401
R3820 VGND.n516 VGND.n515 4.51401
R3821 VGND.n2290 VGND.n1120 4.51401
R3822 VGND VGND.n2284 4.51401
R3823 VGND.n2194 VGND.n1165 4.51401
R3824 VGND.n2199 VGND.n2198 4.51401
R3825 VGND.n2163 VGND.n2153 4.51401
R3826 VGND.n2169 VGND.n2168 4.51401
R3827 VGND.n2930 VGND.n2929 4.51401
R3828 VGND.n565 VGND.n564 4.51401
R3829 VGND.n2258 VGND.n2257 4.51401
R3830 VGND.n2252 VGND.n2251 4.51401
R3831 VGND.n1207 VGND.n1203 4.51401
R3832 VGND.n2121 VGND.n2120 4.51401
R3833 VGND.n2147 VGND.n1182 4.51401
R3834 VGND.n1195 VGND.n1194 4.51401
R3835 VGND.n646 VGND.n645 4.51401
R3836 VGND.n640 VGND.n639 4.51401
R3837 VGND.n587 VGND.n586 4.51401
R3838 VGND.n667 VGND.n666 4.51401
R3839 VGND.n2045 VGND.n2041 4.51401
R3840 VGND.n2089 VGND.n2088 4.51401
R3841 VGND.n2919 VGND.n572 4.51401
R3842 VGND.n2910 VGND.n2906 4.51401
R3843 VGND.n2701 VGND.n744 4.51401
R3844 VGND.n2706 VGND.n2705 4.51401
R3845 VGND.n2671 VGND.n2661 4.51401
R3846 VGND.n2676 VGND.n2675 4.51401
R3847 VGND.n2867 VGND.n674 4.51401
R3848 VGND.n2860 VGND.n2859 4.51401
R3849 VGND.n2797 VGND.n2795 4.51401
R3850 VGND.n2811 VGND.n2810 4.51401
R3851 VGND.n2733 VGND.n725 4.51401
R3852 VGND VGND.n2737 4.51401
R3853 VGND.n2769 VGND.n704 4.51401
R3854 VGND.n2774 VGND.n2773 4.51401
R3855 VGND.n1327 VGND.n1326 4.51401
R3856 VGND.n1336 VGND.n1335 4.51401
R3857 VGND.n2616 VGND.n2615 4.51401
R3858 VGND.n823 VGND.n822 4.51401
R3859 VGND.n2651 VGND.n765 4.51401
R3860 VGND.n770 VGND.n769 4.51401
R3861 VGND.n1383 VGND.n1381 4.51401
R3862 VGND.n1487 VGND 4.51401
R3863 VGND.n1527 VGND.n1301 4.51401
R3864 VGND.n1306 VGND.n1305 4.51401
R3865 VGND.n1407 VGND.n1399 4.51401
R3866 VGND.n1452 VGND.n1451 4.51401
R3867 VGND.n1257 VGND.n1250 4.51401
R3868 VGND.n1950 VGND.n1949 4.51401
R3869 VGND.n2523 VGND.n986 4.51401
R3870 VGND.n2514 VGND.n2513 4.51401
R3871 VGND.n1616 VGND.n1613 4.51401
R3872 VGND.n2605 VGND.n2604 4.51401
R3873 VGND.n1562 VGND.n1557 4.51401
R3874 VGND.n1684 VGND.n1683 4.51401
R3875 VGND.n1725 VGND.n1535 4.51401
R3876 VGND.n1548 VGND.n1547 4.51401
R3877 VGND.n866 VGND.n864 4.51401
R3878 VGND.n894 VGND.n893 4.51401
R3879 VGND.n1590 VGND.n1588 4.51401
R3880 VGND.n1645 VGND.n1644 4.51401
R3881 VGND.n1230 VGND.n1226 4.51401
R3882 VGND.n2015 VGND.n2014 4.51401
R3883 VGND.n1910 VGND.n1909 4.51401
R3884 VGND.n1982 VGND.n1981 4.51401
R3885 VGND.n1836 VGND.n1835 4.51401
R3886 VGND.n1735 VGND.n1291 4.51401
R3887 VGND.n951 VGND.n949 4.51401
R3888 VGND.n980 VGND.n979 4.51401
R3889 VGND.n1874 VGND.n1280 4.51401
R3890 VGND.n1879 VGND.n1878 4.51401
R3891 VGND.n1769 VGND.n1766 4.51401
R3892 VGND.n1795 VGND.n1794 4.51401
R3893 VGND.n1747 VGND.n1743 4.51401
R3894 VGND.n1827 VGND.n1826 4.51401
R3895 VGND.n2427 VGND.n2424 4.51401
R3896 VGND.n2452 VGND.n2451 4.51401
R3897 VGND.n2402 VGND.n2400 4.51401
R3898 VGND.n2483 VGND.n2482 4.51401
R3899 VGND.n2374 VGND.n1024 4.51401
R3900 VGND.n2367 VGND.n1022 4.51401
R3901 VGND.n3017 VGND.n3016 4.51401
R3902 VGND.n3006 VGND.n3005 4.51401
R3903 VGND.n3448 VGND.n3447 4.50726
R3904 VGND.n3174 VGND.n209 4.50726
R3905 VGND.n3357 VGND.n3356 4.50726
R3906 VGND.n534 VGND.n528 4.5005
R3907 VGND.n542 VGND.n541 4.5005
R3908 VGND.n543 VGND.n532 4.5005
R3909 VGND.n2162 VGND.n2161 4.5005
R3910 VGND.n2159 VGND.n2158 4.5005
R3911 VGND.n2155 VGND.n1176 4.5005
R3912 VGND.n2193 VGND.n2192 4.5005
R3913 VGND.n2191 VGND.n2190 4.5005
R3914 VGND.n1160 VGND.n1159 4.5005
R3915 VGND.n2289 VGND.n2288 4.5005
R3916 VGND.n2280 VGND.n1122 4.5005
R3917 VGND.n2283 VGND.n1126 4.5005
R3918 VGND.n2960 VGND.n2959 4.5005
R3919 VGND.n2958 VGND.n2957 4.5005
R3920 VGND.n2954 VGND.n2953 4.5005
R3921 VGND.n1141 VGND.n1134 4.5005
R3922 VGND.n1145 VGND.n1144 4.5005
R3923 VGND.n1138 VGND.n1137 4.5005
R3924 VGND.n2051 VGND.n2049 4.5005
R3925 VGND.n2879 VGND.n2878 4.5005
R3926 VGND.n592 VGND.n588 4.5005
R3927 VGND.n594 VGND.n591 4.5005
R3928 VGND.n630 VGND.n606 4.5005
R3929 VGND.n633 VGND.n632 4.5005
R3930 VGND.n634 VGND.n609 4.5005
R3931 VGND.n2146 VGND.n2145 4.5005
R3932 VGND.n1189 VGND.n1184 4.5005
R3933 VGND.n1193 VGND.n1192 4.5005
R3934 VGND.n2128 VGND.n2127 4.5005
R3935 VGND.n1208 VGND.n1206 4.5005
R3936 VGND.n1213 VGND.n1211 4.5005
R3937 VGND.n2096 VGND.n2095 4.5005
R3938 VGND.n2050 VGND.n2046 4.5005
R3939 VGND.n2918 VGND.n2917 4.5005
R3940 VGND.n2907 VGND.n574 4.5005
R3941 VGND.n2912 VGND.n2911 4.5005
R3942 VGND.n720 VGND.n719 4.5005
R3943 VGND.n2799 VGND.n2798 4.5005
R3944 VGND.n2806 VGND.n2805 4.5005
R3945 VGND.n689 VGND.n686 4.5005
R3946 VGND.n2866 VGND.n2865 4.5005
R3947 VGND.n2855 VGND.n677 4.5005
R3948 VGND.n2858 VGND.n2838 4.5005
R3949 VGND.n2670 VGND.n2669 4.5005
R3950 VGND.n2667 VGND.n2666 4.5005
R3951 VGND.n2663 VGND.n755 4.5005
R3952 VGND.n2700 VGND.n2699 4.5005
R3953 VGND.n2698 VGND.n2697 4.5005
R3954 VGND.n739 VGND.n738 4.5005
R3955 VGND.n2732 VGND.n2731 4.5005
R3956 VGND.n728 VGND.n727 4.5005
R3957 VGND.n2768 VGND.n2767 4.5005
R3958 VGND.n708 VGND.n707 4.5005
R3959 VGND.n700 VGND.n699 4.5005
R3960 VGND.n1382 VGND.n1375 4.5005
R3961 VGND.n1492 VGND.n1491 4.5005
R3962 VGND.n1378 VGND.n1376 4.5005
R3963 VGND.n2650 VGND.n2649 4.5005
R3964 VGND.n2648 VGND.n2647 4.5005
R3965 VGND.n2644 VGND.n2643 4.5005
R3966 VGND.n794 VGND.n787 4.5005
R3967 VGND.n799 VGND.n798 4.5005
R3968 VGND.n795 VGND.n790 4.5005
R3969 VGND.n1323 VGND.n1322 4.5005
R3970 VGND.n1331 VGND.n1330 4.5005
R3971 VGND.n1319 VGND.n1315 4.5005
R3972 VGND.n1526 VGND.n1525 4.5005
R3973 VGND.n1524 VGND.n1523 4.5005
R3974 VGND.n1520 VGND.n1519 4.5005
R3975 VGND.n1406 VGND.n1402 4.5005
R3976 VGND.n1457 VGND.n1456 4.5005
R3977 VGND.n1410 VGND.n1405 4.5005
R3978 VGND.n871 VGND.n869 4.5005
R3979 VGND.n1724 VGND.n1723 4.5005
R3980 VGND.n1542 VGND.n1537 4.5005
R3981 VGND.n1546 VGND.n1545 4.5005
R3982 VGND.n1691 VGND.n1690 4.5005
R3983 VGND.n1563 VGND.n1561 4.5005
R3984 VGND.n1568 VGND.n1565 4.5005
R3985 VGND.n1617 VGND.n1614 4.5005
R3986 VGND.n1622 VGND.n1621 4.5005
R3987 VGND.n833 VGND.n832 4.5005
R3988 VGND.n2577 VGND.n2576 4.5005
R3989 VGND.n2574 VGND.n849 4.5005
R3990 VGND.n2584 VGND.n2583 4.5005
R3991 VGND.n901 VGND.n900 4.5005
R3992 VGND.n870 VGND.n867 4.5005
R3993 VGND.n1652 VGND.n1651 4.5005
R3994 VGND.n1594 VGND.n1591 4.5005
R3995 VGND.n1595 VGND.n1593 4.5005
R3996 VGND.n957 VGND.n955 4.5005
R3997 VGND.n1296 VGND.n1295 4.5005
R3998 VGND.n1731 VGND.n1730 4.5005
R3999 VGND.n1734 VGND.n1733 4.5005
R4000 VGND.n1908 VGND.n1907 4.5005
R4001 VGND.n1903 VGND.n1902 4.5005
R4002 VGND.n1900 VGND.n1237 4.5005
R4003 VGND.n1256 VGND.n1252 4.5005
R4004 VGND.n1955 VGND.n1954 4.5005
R4005 VGND.n1260 VGND.n1255 4.5005
R4006 VGND.n2569 VGND.n2568 4.5005
R4007 VGND.n2567 VGND.n2566 4.5005
R4008 VGND.n2563 VGND.n2562 4.5005
R4009 VGND.n2536 VGND.n2535 4.5005
R4010 VGND.n956 VGND.n952 4.5005
R4011 VGND.n1873 VGND.n1872 4.5005
R4012 VGND.n1871 VGND.n1870 4.5005
R4013 VGND.n1283 VGND.n1275 4.5005
R4014 VGND.n2430 VGND.n2423 4.5005
R4015 VGND.n1749 VGND.n1748 4.5005
R4016 VGND.n1754 VGND.n1753 4.5005
R4017 VGND.n1755 VGND.n1740 4.5005
R4018 VGND.n1802 VGND.n1801 4.5005
R4019 VGND.n1774 VGND.n1770 4.5005
R4020 VGND.n1776 VGND.n1773 4.5005
R4021 VGND.n2022 VGND.n2021 4.5005
R4022 VGND.n1988 VGND.n1231 4.5005
R4023 VGND.n1989 VGND.n1987 4.5005
R4024 VGND.n2522 VGND.n2521 4.5005
R4025 VGND.n992 VGND.n988 4.5005
R4026 VGND.n2516 VGND.n2515 4.5005
R4027 VGND.n2426 VGND.n2425 4.5005
R4028 VGND.n2457 VGND.n2456 4.5005
R4029 VGND.n2490 VGND.n2489 4.5005
R4030 VGND.n2403 VGND.n2401 4.5005
R4031 VGND.n2408 VGND.n2406 4.5005
R4032 VGND.n2347 VGND.n2346 4.5005
R4033 VGND.n249 VGND.n248 4.5005
R4034 VGND.n252 VGND.n251 4.5005
R4035 VGND.n253 VGND.n238 4.5005
R4036 VGND.n1067 VGND.n1066 4.5005
R4037 VGND.n1072 VGND.n1071 4.5005
R4038 VGND.n1056 VGND.n1052 4.5005
R4039 VGND.n1086 VGND.n1083 4.5005
R4040 VGND.n1090 VGND.n1089 4.5005
R4041 VGND.n501 VGND.n500 4.5005
R4042 VGND.n2312 VGND.n2311 4.5005
R4043 VGND.n1047 VGND.n1038 4.5005
R4044 VGND.n2318 VGND.n2317 4.5005
R4045 VGND.n2373 VGND.n2372 4.5005
R4046 VGND.n1027 VGND.n1026 4.5005
R4047 VGND.n269 VGND.n266 4.5005
R4048 VGND.n3012 VGND.n3011 4.5005
R4049 VGND.n3002 VGND.n270 4.5005
R4050 VGND.n2389 VGND.n2388 4.4805
R4051 VGND.n2543 VGND.n2542 4.38311
R4052 VGND.n2186 VGND.n2185 4.36875
R4053 VGND.n2187 VGND.n1158 4.36875
R4054 VGND.n2205 VGND.n1157 4.36875
R4055 VGND.n2214 VGND.n2213 4.36875
R4056 VGND.n2277 VGND.n2276 4.36875
R4057 VGND.n2264 VGND.n2263 4.36875
R4058 VGND.n1147 VGND.n1140 4.36875
R4059 VGND.n2240 VGND.n1151 4.36875
R4060 VGND.n2229 VGND.n2227 4.36875
R4061 VGND.n521 VGND.n520 4.36875
R4062 VGND.n2131 VGND.n2130 4.36875
R4063 VGND.n1216 VGND.n1205 4.36875
R4064 VGND.n2117 VGND.n2116 4.36875
R4065 VGND.n2109 VGND.n1221 4.36875
R4066 VGND.n2077 VGND.n2060 4.36875
R4067 VGND.n2070 VGND.n2069 4.36875
R4068 VGND.n2914 VGND.n576 4.36875
R4069 VGND.n2900 VGND.n577 4.36875
R4070 VGND.n2893 VGND.n2892 4.36875
R4071 VGND.n2693 VGND.n2692 4.36875
R4072 VGND.n2694 VGND.n737 4.36875
R4073 VGND.n2712 VGND.n736 4.36875
R4074 VGND.n2721 VGND.n2720 4.36875
R4075 VGND.n2743 VGND.n2742 4.36875
R4076 VGND.n2755 VGND.n710 4.36875
R4077 VGND.n2764 VGND.n2763 4.36875
R4078 VGND.n2786 VGND.n2785 4.36875
R4079 VGND.n1717 VGND.n1716 4.28986
R4080 VGND.n1711 VGND.n1549 4.28986
R4081 VGND.n889 VGND.n888 4.28986
R4082 VGND.n1791 VGND.n1790 4.28986
R4083 VGND.n2024 VGND.n1228 4.28986
R4084 VGND.n2001 VGND.n2000 4.28986
R4085 VGND.n2462 VGND.n2461 4.28986
R4086 VGND.n1693 VGND.n1560 4.14168
R4087 VGND.n2818 VGND.n2817 4.11798
R4088 VGND.n2817 VGND.n682 4.11798
R4089 VGND.n2636 VGND.n2635 4.11798
R4090 VGND.n1354 VGND.n1353 4.11798
R4091 VGND.n1353 VGND.n1308 4.11798
R4092 VGND.n1503 VGND.n1502 4.11798
R4093 VGND.n1502 VGND.n1501 4.11798
R4094 VGND.n1957 VGND.n1251 4.11798
R4095 VGND.n2349 VGND.n2345 4.11798
R4096 VGND.n2364 VGND.n2349 4.11798
R4097 VGND.n2976 VGND.n497 4.11798
R4098 VGND.n2979 VGND.n497 4.11798
R4099 VGND.n1105 VGND.n1104 4.11798
R4100 VGND.n1104 VGND.n1103 4.11798
R4101 VGND.n2997 VGND.n275 4.11798
R4102 VGND.n2994 VGND.n275 4.11798
R4103 VGND.n2801 VGND.n691 4.09013
R4104 VGND.n888 VGND.n887 4.07323
R4105 VGND.n1790 VGND.n1789 4.07323
R4106 VGND.n2012 VGND.n1228 4.07323
R4107 VGND.n2000 VGND.n1999 4.07323
R4108 VGND.n2461 VGND.n2460 4.07323
R4109 VGND.n562 VGND.n561 4.03876
R4110 VGND.n820 VGND.n819 4.03876
R4111 VGND.n3053 VGND 4.02175
R4112 VGND.n230 VGND 4.02175
R4113 VGND.n3382 VGND 4.02175
R4114 VGND.n231 VGND 4.02175
R4115 VGND.n2223 VGND.n1152 3.97459
R4116 VGND.n2725 VGND.n732 3.97459
R4117 VGND.n2177 VGND.n2176 3.96548
R4118 VGND.n2180 VGND.n2177 3.96548
R4119 VGND.n557 VGND.n556 3.96548
R4120 VGND.n2138 VGND.n2137 3.96548
R4121 VGND.n2137 VGND.n2136 3.96548
R4122 VGND.n2885 VGND.n2884 3.96548
R4123 VGND.n2863 VGND.n2862 3.96548
R4124 VGND.n2862 VGND.n2837 3.96548
R4125 VGND.n2852 VGND.n2851 3.96548
R4126 VGND.n2684 VGND.n2683 3.96548
R4127 VGND.n2687 VGND.n2684 3.96548
R4128 VGND.n815 VGND.n814 3.96548
R4129 VGND.n1345 VGND.n1344 3.96548
R4130 VGND.n1347 VGND.n1345 3.96548
R4131 VGND.n841 VGND.n839 3.90948
R4132 VGND.n841 VGND.n840 3.90948
R4133 VGND.n390 VGND.n389 3.78485
R4134 VGND.n3241 VGND.n3239 3.78485
R4135 VGND.n3271 VGND.n3260 3.78485
R4136 VGND.n3223 VGND.n3222 3.78485
R4137 VGND.n3218 VGND.n3217 3.78485
R4138 VGND.n3199 VGND.n182 3.78485
R4139 VGND.n3385 VGND.n77 3.78485
R4140 VGND.n3275 VGND.n3255 3.78485
R4141 VGND.n2634 VGND.n2633 3.75994
R4142 VGND.n412 VGND.n409 3.75517
R4143 VGND.n2176 VGND.n1171 3.7069
R4144 VGND.n557 VGND.n546 3.7069
R4145 VGND.n2138 VGND.n1198 3.7069
R4146 VGND.n2885 VGND.n582 3.7069
R4147 VGND.n2100 VGND.n2039 3.7069
R4148 VGND.n2100 VGND.n2099 3.7069
R4149 VGND.n2863 VGND.n2836 3.7069
R4150 VGND.n2849 VGND.n2841 3.7069
R4151 VGND.n2683 VGND.n750 3.7069
R4152 VGND.n815 VGND.n804 3.7069
R4153 VGND.n1344 VGND.n1313 3.7069
R4154 VGND.n1347 VGND.n1346 3.7069
R4155 VGND.n1705 VGND.n1552 3.50735
R4156 VGND.n2476 VGND.n2475 3.50735
R4157 VGND.n2324 VGND.n2323 3.50735
R4158 VGND.n3025 VGND.n261 3.50735
R4159 VGND.n490 VGND.n401 3.46461
R4160 VGND.n422 VGND.n401 3.46461
R4161 VGND.t551 VGND.t371 3.46461
R4162 VGND.t551 VGND.t457 3.46461
R4163 VGND.n424 VGND.n420 3.46461
R4164 VGND.n469 VGND.n424 3.46461
R4165 VGND.n977 VGND.n976 3.44377
R4166 VGND.n976 VGND.n975 3.44377
R4167 VGND.n931 VGND.n924 3.43925
R4168 VGND.n2571 VGND.n2570 3.43925
R4169 VGND.n2582 VGND.n2581 3.43925
R4170 VGND.n2579 VGND.n2578 3.43925
R4171 VGND.n515 VGND.n508 3.43925
R4172 VGND.n2962 VGND.n2961 3.43925
R4173 VGND.n2284 VGND.n1117 3.43925
R4174 VGND.n2291 VGND.n2290 3.43925
R4175 VGND.n2198 VGND.n2197 3.43925
R4176 VGND.n2195 VGND.n2194 3.43925
R4177 VGND.n566 VGND.n565 3.43925
R4178 VGND.n2929 VGND.n2928 3.43925
R4179 VGND.n2253 VGND.n2252 3.43925
R4180 VGND.n2257 VGND.n2256 3.43925
R4181 VGND.n2122 VGND.n2121 3.43925
R4182 VGND.n2124 VGND.n1207 3.43925
R4183 VGND.n1194 VGND.n1180 3.43925
R4184 VGND.n2148 VGND.n2147 3.43925
R4185 VGND.n641 VGND.n640 3.43925
R4186 VGND.n645 VGND.n644 3.43925
R4187 VGND.n668 VGND.n667 3.43925
R4188 VGND.n2875 VGND.n587 3.43925
R4189 VGND.n2090 VGND.n2089 3.43925
R4190 VGND.n2092 VGND.n2045 3.43925
R4191 VGND.n2910 VGND.n569 3.43925
R4192 VGND.n2920 VGND.n2919 3.43925
R4193 VGND.n2705 VGND.n2704 3.43925
R4194 VGND.n2702 VGND.n2701 3.43925
R4195 VGND.n2675 VGND.n2674 3.43925
R4196 VGND.n2672 VGND.n2671 3.43925
R4197 VGND.n2859 VGND.n671 3.43925
R4198 VGND.n2868 VGND.n2867 3.43925
R4199 VGND.n2810 VGND.n2809 3.43925
R4200 VGND.n2797 VGND.n2796 3.43925
R4201 VGND.n2737 VGND.n2736 3.43925
R4202 VGND.n2734 VGND.n2733 3.43925
R4203 VGND.n2773 VGND.n2772 3.43925
R4204 VGND.n2770 VGND.n2769 3.43925
R4205 VGND.n824 VGND.n823 3.43925
R4206 VGND.n2615 VGND.n2614 3.43925
R4207 VGND.n769 VGND.n762 3.43925
R4208 VGND.n2652 VGND.n2651 3.43925
R4209 VGND.n1488 VGND.n1487 3.43925
R4210 VGND.n1384 VGND.n1383 3.43925
R4211 VGND.n1305 VGND.n1299 3.43925
R4212 VGND.n1528 VGND.n1527 3.43925
R4213 VGND.n1453 VGND.n1452 3.43925
R4214 VGND.n1408 VGND.n1407 3.43925
R4215 VGND.n1951 VGND.n1950 3.43925
R4216 VGND.n1258 VGND.n1257 3.43925
R4217 VGND.n2514 VGND.n984 3.43925
R4218 VGND.n2524 VGND.n2523 3.43925
R4219 VGND.n1685 VGND.n1684 3.43925
R4220 VGND.n1687 VGND.n1562 3.43925
R4221 VGND.n1547 VGND.n1533 3.43925
R4222 VGND.n1726 VGND.n1725 3.43925
R4223 VGND.n895 VGND.n894 3.43925
R4224 VGND.n897 VGND.n866 3.43925
R4225 VGND.n1646 VGND.n1645 3.43925
R4226 VGND.n1648 VGND.n1590 3.43925
R4227 VGND.n2016 VGND.n2015 3.43925
R4228 VGND.n2018 VGND.n1230 3.43925
R4229 VGND.n981 VGND.n980 3.43925
R4230 VGND.n2532 VGND.n951 3.43925
R4231 VGND.n1878 VGND.n1877 3.43925
R4232 VGND.n1875 VGND.n1874 3.43925
R4233 VGND.n1796 VGND.n1795 3.43925
R4234 VGND.n1798 VGND.n1769 3.43925
R4235 VGND.n2453 VGND.n2452 3.43925
R4236 VGND.n2428 VGND.n2427 3.43925
R4237 VGND.n2484 VGND.n2483 3.43925
R4238 VGND.n2486 VGND.n2402 3.43925
R4239 VGND.n3044 VGND.n3043 3.41839
R4240 VGND.n243 VGND.n242 3.41839
R4241 VGND.n3005 VGND.n3004 3.41636
R4242 VGND.n3016 VGND.n3015 3.41636
R4243 VGND.n1116 VGND.n1115 3.41624
R4244 VGND.n1057 VGND.n1050 3.41624
R4245 VGND.n2970 VGND.n2969 3.41605
R4246 VGND.n1085 VGND.n503 3.41605
R4247 VGND.n2168 VGND.n2167 3.41514
R4248 VGND.n1335 VGND.n1334 3.41514
R4249 VGND.n1736 VGND.n1735 3.41514
R4250 VGND.n250 VGND.n235 3.4105
R4251 VGND.n3045 VGND.n236 3.4105
R4252 VGND.n928 VGND.n926 3.4105
R4253 VGND.n2565 VGND.n2564 3.4105
R4254 VGND.n1069 VGND.n1068 3.4105
R4255 VGND.n1070 VGND.n1051 3.4105
R4256 VGND.n2575 VGND.n2573 3.4105
R4257 VGND.n923 VGND.n851 3.4105
R4258 VGND.n1087 VGND.n1048 3.4105
R4259 VGND.n1088 VGND.n502 3.4105
R4260 VGND.n512 VGND.n510 3.4105
R4261 VGND.n2956 VGND.n2955 3.4105
R4262 VGND.n1121 VGND.n1119 3.4105
R4263 VGND.n2282 VGND.n2281 3.4105
R4264 VGND.n1166 VGND.n1164 3.4105
R4265 VGND.n2189 VGND.n1161 3.4105
R4266 VGND.n2164 VGND.n2163 3.4105
R4267 VGND.n2154 VGND.n2152 3.4105
R4268 VGND.n2157 VGND.n1177 3.4105
R4269 VGND.n539 VGND.n529 3.4105
R4270 VGND.n540 VGND.n531 3.4105
R4271 VGND.n2255 VGND.n1135 3.4105
R4272 VGND.n2254 VGND.n1136 3.4105
R4273 VGND.n2126 VGND.n2125 3.4105
R4274 VGND.n1210 VGND.n1209 3.4105
R4275 VGND.n1183 VGND.n1181 3.4105
R4276 VGND.n1191 VGND.n1190 3.4105
R4277 VGND.n643 VGND.n607 3.4105
R4278 VGND.n642 VGND.n608 3.4105
R4279 VGND.n2877 VGND.n2876 3.4105
R4280 VGND.n590 VGND.n589 3.4105
R4281 VGND.n2094 VGND.n2093 3.4105
R4282 VGND.n2048 VGND.n2047 3.4105
R4283 VGND.n573 VGND.n571 3.4105
R4284 VGND.n2909 VGND.n2908 3.4105
R4285 VGND.n745 VGND.n743 3.4105
R4286 VGND.n2696 VGND.n740 3.4105
R4287 VGND.n2662 VGND.n2660 3.4105
R4288 VGND.n2665 VGND.n756 3.4105
R4289 VGND.n675 VGND.n673 3.4105
R4290 VGND.n2857 VGND.n2856 3.4105
R4291 VGND.n688 VGND.n687 3.4105
R4292 VGND.n2808 VGND.n2807 3.4105
R4293 VGND.n729 VGND.n724 3.4105
R4294 VGND.n726 VGND.n721 3.4105
R4295 VGND.n705 VGND.n703 3.4105
R4296 VGND.n706 VGND.n701 3.4105
R4297 VGND.n1326 VGND.n1325 3.4105
R4298 VGND.n1317 VGND.n1316 3.4105
R4299 VGND.n1333 VGND.n1332 3.4105
R4300 VGND.n796 VGND.n788 3.4105
R4301 VGND.n797 VGND.n789 3.4105
R4302 VGND.n766 VGND.n764 3.4105
R4303 VGND.n2646 VGND.n2645 3.4105
R4304 VGND.n1379 VGND.n1377 3.4105
R4305 VGND.n1490 VGND.n1489 3.4105
R4306 VGND.n1302 VGND.n1300 3.4105
R4307 VGND.n1522 VGND.n1521 3.4105
R4308 VGND.n1409 VGND.n1404 3.4105
R4309 VGND.n1455 VGND.n1454 3.4105
R4310 VGND.n1259 VGND.n1254 3.4105
R4311 VGND.n1953 VGND.n1952 3.4105
R4312 VGND.n987 VGND.n985 3.4105
R4313 VGND.n994 VGND.n993 3.4105
R4314 VGND.n2607 VGND.n2606 3.4105
R4315 VGND.n2607 VGND.n829 3.4105
R4316 VGND.n2606 VGND.n2605 3.4105
R4317 VGND.n1616 VGND.n829 3.4105
R4318 VGND.n1619 VGND.n1618 3.4105
R4319 VGND.n1620 VGND.n831 3.4105
R4320 VGND.n1689 VGND.n1688 3.4105
R4321 VGND.n1686 VGND.n1564 3.4105
R4322 VGND.n1536 VGND.n1534 3.4105
R4323 VGND.n1544 VGND.n1543 3.4105
R4324 VGND.n899 VGND.n898 3.4105
R4325 VGND.n896 VGND.n868 3.4105
R4326 VGND.n1650 VGND.n1649 3.4105
R4327 VGND.n1647 VGND.n1592 3.4105
R4328 VGND.n2020 VGND.n2019 3.4105
R4329 VGND.n1986 VGND.n1232 3.4105
R4330 VGND.n1984 VGND.n1983 3.4105
R4331 VGND.n1984 VGND.n1235 3.4105
R4332 VGND.n1983 VGND.n1982 3.4105
R4333 VGND.n1909 VGND.n1235 3.4105
R4334 VGND.n1899 VGND.n1898 3.4105
R4335 VGND.n1901 VGND.n1236 3.4105
R4336 VGND.n1835 VGND.n1834 3.4105
R4337 VGND.n1729 VGND.n1298 3.4105
R4338 VGND.n1732 VGND.n1728 3.4105
R4339 VGND.n2534 VGND.n2533 3.4105
R4340 VGND.n954 VGND.n953 3.4105
R4341 VGND.n1281 VGND.n1279 3.4105
R4342 VGND.n1869 VGND.n1276 3.4105
R4343 VGND.n1800 VGND.n1799 3.4105
R4344 VGND.n1772 VGND.n1771 3.4105
R4345 VGND.n1829 VGND.n1828 3.4105
R4346 VGND.n1829 VGND.n1738 3.4105
R4347 VGND.n1828 VGND.n1827 3.4105
R4348 VGND.n1743 VGND.n1738 3.4105
R4349 VGND.n1751 VGND.n1750 3.4105
R4350 VGND.n1752 VGND.n1739 3.4105
R4351 VGND.n2429 VGND.n2422 3.4105
R4352 VGND.n2455 VGND.n2454 3.4105
R4353 VGND.n2488 VGND.n2487 3.4105
R4354 VGND.n2405 VGND.n2404 3.4105
R4355 VGND.n2375 VGND.n2374 3.4105
R4356 VGND.n3014 VGND.n3013 3.4105
R4357 VGND.n3003 VGND.n268 3.4105
R4358 VGND.n2319 VGND.n1019 3.4105
R4359 VGND.n2305 VGND.n1046 3.4105
R4360 VGND.n2310 VGND.n2309 3.4105
R4361 VGND.n2308 VGND.n1037 3.4105
R4362 VGND.n2375 VGND.n1022 3.4105
R4363 VGND.n2375 VGND.n1021 3.4105
R4364 VGND.n2375 VGND.n1020 3.4105
R4365 VGND.n30 VGND.n29 3.40476
R4366 VGND.n3348 VGND.n3347 3.40476
R4367 VGND.n780 VGND.n777 3.31239
R4368 VGND.n1263 VGND.n1251 3.22288
R4369 VGND.n977 VGND.n963 3.21921
R4370 VGND.n972 VGND.n971 3.21921
R4371 VGND.n1703 VGND.n1554 3.2005
R4372 VGND.n2480 VGND.n2411 3.2005
R4373 VGND.n2328 VGND.n1034 3.2005
R4374 VGND.n3024 VGND.n262 3.2005
R4375 VGND.n57 VGND.n56 3.13241
R4376 VGND.n3440 VGND.n3436 3.13241
R4377 VGND.n29 VGND.n25 3.13241
R4378 VGND.n10 VGND.n9 3.13241
R4379 VGND.n3303 VGND.n3302 3.13241
R4380 VGND.n102 VGND.n98 3.13241
R4381 VGND.n3322 VGND.n3321 3.13241
R4382 VGND.n3347 VGND.n3346 3.13241
R4383 VGND.n620 VGND.n619 3.13241
R4384 VGND.n1441 VGND.n1440 3.13241
R4385 VGND.n1812 VGND.n1811 3.13241
R4386 VGND.n2507 VGND.n996 3.13241
R4387 VGND.n1016 VGND.n1015 3.1005
R4388 VGND.n2043 VGND.n2042 3.09945
R4389 VGND.n2215 VGND.n1152 3.05276
R4390 VGND.n2722 VGND.n732 3.05276
R4391 VGND.n551 VGND.n550 3.04861
R4392 VGND.n2172 VGND.n2170 3.04861
R4393 VGND.n615 VGND.n614 3.04861
R4394 VGND.n2142 VGND.n1196 3.04861
R4395 VGND.n2845 VGND.n2843 3.04861
R4396 VGND.n2679 VGND.n2677 3.04861
R4397 VGND.n809 VGND.n808 3.04861
R4398 VGND.n886 VGND.n885 3.04861
R4399 VGND.n969 VGND.n968 3.04861
R4400 VGND.n1789 VGND.n1782 3.04861
R4401 VGND.n1999 VGND.n1998 3.04861
R4402 VGND.n1892 VGND.n1889 3.01226
R4403 VGND.n1666 VGND.n1665 2.92224
R4404 VGND.n2802 VGND.n2801 2.92166
R4405 VGND.n3468 VGND.n3467 2.90519
R4406 VGND.n3071 VGND.t298 2.89674
R4407 VGND.n2180 VGND.n2179 2.88804
R4408 VGND.n2136 VGND.n1201 2.88804
R4409 VGND.n2687 VGND.n2686 2.88804
R4410 VGND.n3134 VGND.n3133 2.88636
R4411 VGND.n31 VGND.n30 2.86007
R4412 VGND.n3349 VGND.n3348 2.86007
R4413 VGND.n2179 VGND.n2178 2.79323
R4414 VGND.n1201 VGND.n1200 2.79323
R4415 VGND.n2686 VGND.n2685 2.79323
R4416 VGND.n561 VGND.n560 2.77203
R4417 VGND.n819 VGND.n818 2.77203
R4418 VGND.n58 VGND.n57 2.7239
R4419 VGND.n3437 VGND.n3436 2.7239
R4420 VGND.n26 VGND.n25 2.7239
R4421 VGND.n9 VGND.n8 2.7239
R4422 VGND.n3302 VGND.n81 2.7239
R4423 VGND.n99 VGND.n98 2.7239
R4424 VGND.n3323 VGND.n3322 2.7239
R4425 VGND.n3346 VGND.n3345 2.7239
R4426 VGND.n619 VGND.n618 2.7239
R4427 VGND.n1440 VGND.n1439 2.7239
R4428 VGND.n1844 VGND.n1843 2.7239
R4429 VGND.n1811 VGND.n1810 2.7239
R4430 VGND.n997 VGND.n996 2.7239
R4431 VGND.n2637 VGND.n774 2.68581
R4432 VGND.n3467 VGND.n3466 2.63717
R4433 VGND.n3298 VGND.n3297 2.63717
R4434 VGND.n1701 VGND.n1700 2.63064
R4435 VGND.n2479 VGND.n2474 2.63064
R4436 VGND.n2327 VGND.n1032 2.63064
R4437 VGND.n3022 VGND.n3021 2.63064
R4438 VGND.n3408 VGND.n3407 2.59858
R4439 VGND VGND.n229 2.56738
R4440 VGND.n2086 VGND.n2055 2.55412
R4441 VGND.n2938 VGND.n2937 2.50679
R4442 VGND.n1432 VGND.n1421 2.50679
R4443 VGND.n1971 VGND.n1243 2.50679
R4444 VGND.n692 VGND.n691 2.38348
R4445 VGND.n2208 VGND.n2207 2.33701
R4446 VGND.n2207 VGND.n1155 2.33701
R4447 VGND.n2270 VGND.n2269 2.33701
R4448 VGND.n2269 VGND.n2268 2.33701
R4449 VGND.n1132 VGND.n1130 2.33701
R4450 VGND.n2264 VGND.n1132 2.33701
R4451 VGND.n1150 VGND.n1148 2.33701
R4452 VGND.n2243 VGND.n1150 2.33701
R4453 VGND.n2242 VGND.n2241 2.33701
R4454 VGND.n2241 VGND.n2240 2.33701
R4455 VGND.n2946 VGND.n2945 2.33701
R4456 VGND.n2945 VGND.n2944 2.33701
R4457 VGND.n1220 VGND.n1218 2.33701
R4458 VGND.n2111 VGND.n1220 2.33701
R4459 VGND.n2076 VGND.n2075 2.33701
R4460 VGND.n2075 VGND.n2074 2.33701
R4461 VGND.n2063 VGND.n575 2.33701
R4462 VGND.n2899 VGND.n2898 2.33701
R4463 VGND.n2898 VGND.n2897 2.33701
R4464 VGND.n2715 VGND.n2714 2.33701
R4465 VGND.n2714 VGND.n734 2.33701
R4466 VGND.n2749 VGND.n712 2.33701
R4467 VGND.n2752 VGND.n712 2.33701
R4468 VGND.n2754 VGND.n2753 2.33701
R4469 VGND.n2755 VGND.n2754 2.33701
R4470 VGND.n2779 VGND.n696 2.33701
R4471 VGND.n2782 VGND.n696 2.33701
R4472 VGND.n2784 VGND.n2783 2.33701
R4473 VGND.n2786 VGND.n2784 2.33701
R4474 VGND.n2085 VGND.n2056 2.33067
R4475 VGND.n295 VGND.n288 2.3255
R4476 VGND.n301 VGND.n287 2.3255
R4477 VGND.n327 VGND.n326 2.3255
R4478 VGND.n332 VGND.n331 2.3255
R4479 VGND.n375 VGND.n374 2.3255
R4480 VGND.n352 VGND.n351 2.3255
R4481 VGND.n349 VGND.n345 2.3255
R4482 VGND.n201 VGND.n200 2.3255
R4483 VGND.n3088 VGND.n3087 2.25932
R4484 VGND.n3128 VGND.n3098 2.25932
R4485 VGND.n629 VGND.n628 2.25932
R4486 VGND.n1478 VGND.n1393 2.25932
R4487 VGND.n1679 VGND.n1678 2.25932
R4488 VGND.n1657 VGND.n1656 2.25932
R4489 VGND.n1598 VGND.n1587 2.25932
R4490 VGND.n1599 VGND.n1598 2.25932
R4491 VGND.n919 VGND.n918 2.25932
R4492 VGND.n1853 VGND.n1852 2.25932
R4493 VGND.n1892 VGND.n1891 2.25932
R4494 VGND.n1920 VGND.n934 2.25932
R4495 VGND.n2182 VGND.n1169 2.25312
R4496 VGND.n2134 VGND.n1202 2.25312
R4497 VGND.n2689 VGND.n748 2.25312
R4498 VGND.n2596 VGND.n841 2.25293
R4499 VGND.n3050 VGND.n3049 2.23999
R4500 VGND.n1169 VGND.n1168 2.2228
R4501 VGND.n1204 VGND.n1202 2.2228
R4502 VGND.n748 VGND.n747 2.2228
R4503 VGND.n1845 VGND.n1844 2.17922
R4504 VGND.n3295 VGND.n3294 2.14347
R4505 VGND.n1716 VGND.n1715 2.13383
R4506 VGND.n1125 VGND.n1124 2.11085
R4507 VGND.n718 VGND.n717 2.11085
R4508 VGND.n2851 VGND.n2850 2.06919
R4509 VGND.n3067 VGND.n3066 2.03479
R4510 VGND.n2064 VGND.n2063 2.03225
R4511 VGND.n556 VGND.n555 1.98299
R4512 VGND.n2884 VGND.n2883 1.98299
R4513 VGND.n2840 VGND.n2837 1.98299
R4514 VGND.n2852 VGND.n2840 1.98299
R4515 VGND.n814 VGND.n813 1.98299
R4516 VGND.n2539 VGND.n2538 1.97497
R4517 VGND.n2083 VGND.n2082 1.91571
R4518 VGND.n2850 VGND.n2849 1.8968
R4519 VGND.n875 VGND.n874 1.88285
R4520 VGND.n1665 VGND.n1664 1.87876
R4521 VGND.n975 VGND.n964 1.79699
R4522 VGND.n3068 VGND.n3067 1.77326
R4523 VGND.n2627 VGND.n2626 1.75824
R4524 VGND.n3435 VGND.n3434 1.753
R4525 VGND.n3433 VGND.n3432 1.753
R4526 VGND.n3166 VGND.n3165 1.753
R4527 VGND.n3164 VGND.n3163 1.753
R4528 VGND.n96 VGND.n79 1.753
R4529 VGND.n3380 VGND.n3379 1.753
R4530 VGND.n1671 VGND.n1669 1.7528
R4531 VGND.n555 VGND.n554 1.72441
R4532 VGND.n2883 VGND.n2882 1.72441
R4533 VGND.n813 VGND.n812 1.72441
R4534 VGND.n2307 VGND.n507 1.70468
R4535 VGND.n2306 VGND.n507 1.70468
R4536 VGND.n1832 VGND.n1736 1.70393
R4537 VGND.n1833 VGND.n1832 1.70393
R4538 VGND.n1334 VGND.n760 1.70393
R4539 VGND.n1324 VGND.n760 1.70393
R4540 VGND.n2167 VGND.n2166 1.70393
R4541 VGND.n2166 VGND.n2165 1.70393
R4542 VGND.n2969 VGND.n2968 1.70348
R4543 VGND.n2968 VGND.n503 1.70348
R4544 VGND.n2294 VGND.n1116 1.70338
R4545 VGND.n2294 VGND.n1050 1.70338
R4546 VGND.n3004 VGND.n267 1.70332
R4547 VGND.n3015 VGND.n267 1.70332
R4548 VGND.n3044 VGND.n237 1.70231
R4549 VGND.n242 VGND.n237 1.70231
R4550 VGND.n820 VGND.n803 1.7012
R4551 VGND.n2525 VGND.n984 1.69188
R4552 VGND.n2525 VGND.n2524 1.69188
R4553 VGND.n1951 VGND.n830 1.69188
R4554 VGND.n1258 VGND.n830 1.69188
R4555 VGND.n1453 VGND.n827 1.69188
R4556 VGND.n1408 VGND.n827 1.69188
R4557 VGND.n2772 VGND.n2771 1.69188
R4558 VGND.n2771 VGND.n2770 1.69188
R4559 VGND.n2921 VGND.n569 1.69188
R4560 VGND.n2921 VGND.n2920 1.69188
R4561 VGND.n2253 VGND.n504 1.69188
R4562 VGND.n2256 VGND.n504 1.69188
R4563 VGND.n2607 VGND.n828 1.69188
R4564 VGND.n2017 VGND.n2016 1.69188
R4565 VGND.n2018 VGND.n2017 1.69188
R4566 VGND.n1646 VGND.n1233 1.69188
R4567 VGND.n1648 VGND.n1233 1.69188
R4568 VGND.n1488 VGND.n1385 1.69188
R4569 VGND.n1385 VGND.n1384 1.69188
R4570 VGND.n2736 VGND.n2735 1.69188
R4571 VGND.n2735 VGND.n2734 1.69188
R4572 VGND.n2091 VGND.n2090 1.69188
R4573 VGND.n2092 VGND.n2091 1.69188
R4574 VGND.n2292 VGND.n1117 1.69188
R4575 VGND.n2292 VGND.n2291 1.69188
R4576 VGND.n1984 VGND.n1234 1.69188
R4577 VGND.n1797 VGND.n1796 1.69188
R4578 VGND.n1798 VGND.n1797 1.69188
R4579 VGND.n1877 VGND.n1876 1.69188
R4580 VGND.n1876 VGND.n1875 1.69188
R4581 VGND.n1685 VGND.n1277 1.69188
R4582 VGND.n1687 VGND.n1277 1.69188
R4583 VGND.n1529 VGND.n1299 1.69188
R4584 VGND.n1529 VGND.n1528 1.69188
R4585 VGND.n2704 VGND.n2703 1.69188
R4586 VGND.n2703 VGND.n2702 1.69188
R4587 VGND.n2123 VGND.n2122 1.69188
R4588 VGND.n2124 VGND.n2123 1.69188
R4589 VGND.n2197 VGND.n2196 1.69188
R4590 VGND.n2196 VGND.n2195 1.69188
R4591 VGND.n1727 VGND.n1533 1.69188
R4592 VGND.n1727 VGND.n1726 1.69188
R4593 VGND.n2674 VGND.n2673 1.69188
R4594 VGND.n2673 VGND.n2672 1.69188
R4595 VGND.n2149 VGND.n1180 1.69188
R4596 VGND.n2149 VGND.n2148 1.69188
R4597 VGND.n1829 VGND.n1737 1.69188
R4598 VGND.n2485 VGND.n2484 1.69188
R4599 VGND.n2486 VGND.n2485 1.69188
R4600 VGND.n2572 VGND.n924 1.69188
R4601 VGND.n2572 VGND.n2571 1.69188
R4602 VGND.n2581 VGND.n2580 1.69188
R4603 VGND.n2580 VGND.n2579 1.69188
R4604 VGND.n2653 VGND.n762 1.69188
R4605 VGND.n2653 VGND.n2652 1.69188
R4606 VGND.n2809 VGND.n669 1.69188
R4607 VGND.n2796 VGND.n669 1.69188
R4608 VGND.n2874 VGND.n668 1.69188
R4609 VGND.n2875 VGND.n2874 1.69188
R4610 VGND.n2963 VGND.n508 1.69188
R4611 VGND.n2963 VGND.n2962 1.69188
R4612 VGND.n2453 VGND.n982 1.69188
R4613 VGND.n2428 VGND.n982 1.69188
R4614 VGND.n2531 VGND.n981 1.69188
R4615 VGND.n2532 VGND.n2531 1.69188
R4616 VGND.n895 VGND.n825 1.69188
R4617 VGND.n897 VGND.n825 1.69188
R4618 VGND.n2613 VGND.n824 1.69188
R4619 VGND.n2614 VGND.n2613 1.69188
R4620 VGND.n2869 VGND.n671 1.69188
R4621 VGND.n2869 VGND.n2868 1.69188
R4622 VGND.n641 VGND.n567 1.69188
R4623 VGND.n644 VGND.n567 1.69188
R4624 VGND.n2927 VGND.n566 1.69188
R4625 VGND.n2928 VGND.n2927 1.69188
R4626 VGND.n972 VGND.n964 1.64728
R4627 VGND.n2641 VGND.n772 1.61169
R4628 VGND.n3401 VGND 1.54822
R4629 VGND.n3160 VGND.n3146 1.50638
R4630 VGND.n3154 VGND.n3148 1.50638
R4631 VGND.n191 VGND.n189 1.50638
R4632 VGND.n3182 VGND.n192 1.50638
R4633 VGND.n3096 VGND.n3095 1.50638
R4634 VGND.n3097 VGND.n3096 1.50638
R4635 VGND.n3125 VGND.n3124 1.50638
R4636 VGND.n3118 VGND.n3101 1.50638
R4637 VGND.n3118 VGND.n3117 1.50638
R4638 VGND.n3109 VGND.n3108 1.50638
R4639 VGND.n2891 VGND.n2890 1.47352
R4640 VGND.n3067 VGND.n3054 1.44312
R4641 VGND.n2106 VGND.n2105 1.34658
R4642 VGND.n3052 VGND.n229 1.3415
R4643 VGND.n691 VGND.n690 1.3283
R4644 VGND.n3051 VGND.n3050 1.31337
R4645 VGND.n2184 VGND.n1168 1.29527
R4646 VGND.n2132 VGND.n1204 1.29527
R4647 VGND.n2691 VGND.n747 1.29527
R4648 VGND.n545 VGND.n533 1.25365
R4649 VGND.n2104 VGND.n2103 1.25033
R4650 VGND.n17 VGND.n1 1.21169
R4651 VGND.n3133 VGND.n3132 1.21169
R4652 VGND.n3296 VGND.n111 1.21169
R4653 VGND.n1341 VGND.n1340 1.20723
R4654 VGND.n1664 VGND.n1663 1.18311
R4655 VGND.n1926 VGND.n1925 1.18311
R4656 VGND.n2542 VGND.n2541 1.18311
R4657 VGND.n1746 VGND.n1745 1.18311
R4658 VGND.n2438 VGND.n2437 1.18311
R4659 VGND.n2354 VGND.n2353 1.18311
R4660 VGND.n1061 VGND.n1060 1.18311
R4661 VGND.n3037 VGND.n3036 1.18311
R4662 VGND.n246 VGND.n245 1.18311
R4663 VGND.n450 VGND.n409 1.15795
R4664 VGND.n1701 VGND.n1554 1.14023
R4665 VGND.n2480 VGND.n2479 1.14023
R4666 VGND.n2328 VGND.n2327 1.14023
R4667 VGND.n3022 VGND.n262 1.14023
R4668 VGND.n1604 VGND.n1601 1.12991
R4669 VGND.n2889 VGND.n2888 1.12954
R4670 VGND.n2296 VGND 1.12383
R4671 VGND.n2295 VGND 1.11689
R4672 VGND.n2300 VGND 1.11689
R4673 VGND.n3050 VGND.n232 1.11056
R4674 VGND.n2299 VGND 1.07702
R4675 VGND.n2621 VGND.n2620 1.07463
R4676 VGND.n3469 VGND 1.06996
R4677 VGND.n3052 VGND.n3051 1.05425
R4678 VGND.n3433 VGND 1.00137
R4679 VGND.n2381 VGND.n2380 0.993972
R4680 VGND.n801 VGND.n793 0.985115
R4681 VGND.n1846 VGND.n1845 0.953691
R4682 VGND.n888 VGND.n879 0.952566
R4683 VGND.n1790 VGND.n1781 0.952566
R4684 VGND.n1228 VGND.n1227 0.952566
R4685 VGND.n2000 VGND.n1996 0.952566
R4686 VGND.n2461 VGND.n2417 0.952566
R4687 VGND.n472 VGND.n0 0.927421
R4688 VGND.n887 VGND.n882 0.899674
R4689 VGND.n1961 VGND.n1249 0.895605
R4690 VGND.n1264 VGND.n1263 0.895605
R4691 VGND.n2179 VGND.n1169 0.892621
R4692 VGND.n1202 VGND.n1201 0.892621
R4693 VGND.n2686 VGND.n748 0.892621
R4694 VGND.n2375 VGND.n1023 0.853
R4695 VGND.n2379 VGND.n2378 0.842928
R4696 VGND.n2475 VGND.n2411 0.833377
R4697 VGND.n2323 VGND.n1034 0.833377
R4698 VGND.n3025 VGND.n3024 0.833377
R4699 VGND.n2083 VGND.n2056 0.830425
R4700 VGND.n2054 VGND.n2042 0.798505
R4701 VGND.n2388 VGND.n2387 0.777453
R4702 VGND.n3434 VGND.n3433 0.761313
R4703 VGND.n3165 VGND.n3164 0.761313
R4704 VGND.n3380 VGND.n79 0.761313
R4705 VGND.n3156 VGND.n3155 0.753441
R4706 VGND.n3150 VGND.n188 0.753441
R4707 VGND.n3184 VGND.n3183 0.753441
R4708 VGND.n3178 VGND.n3177 0.753441
R4709 VGND.n3129 VGND.n3128 0.753441
R4710 VGND.n3122 VGND.n3121 0.753441
R4711 VGND.n3115 VGND.n3114 0.753441
R4712 VGND.n1483 VGND.n1482 0.753441
R4713 VGND.n1674 VGND.n1673 0.753441
R4714 VGND.n908 VGND.n861 0.753441
R4715 VGND.n1510 VGND.n1509 0.716584
R4716 VGND.n2086 VGND.n2085 0.606984
R4717 VGND.n468 VGND.n426 0.577852
R4718 VGND.t643 VGND.t467 0.577852
R4719 VGND.n460 VGND.n438 0.577852
R4720 VGND.n2233 VGND.n2226 0.537563
R4721 VGND.n2829 VGND.n2828 0.537563
R4722 VGND.n2816 VGND.n2815 0.537563
R4723 VGND.n2827 VGND.n680 0.537563
R4724 VGND.n2624 VGND.n781 0.537563
R4725 VGND.n1425 VGND.n1424 0.537563
R4726 VGND.n2628 VGND.n2627 0.537563
R4727 VGND.n1362 VGND.n1361 0.537563
R4728 VGND.n1517 VGND.n1516 0.537563
R4729 VGND.n1496 VGND.n1370 0.537563
R4730 VGND.n1945 VGND.n1944 0.537563
R4731 VGND.n2338 VGND.n2337 0.537563
R4732 VGND.n2359 VGND.n2350 0.537563
R4733 VGND.n1096 VGND.n1080 0.537563
R4734 VGND.n2984 VGND.n495 0.537563
R4735 VGND.n1075 VGND.n1074 0.537563
R4736 VGND.n1098 VGND.n1097 0.537563
R4737 VGND.n271 VGND.n264 0.537563
R4738 VGND.n2989 VGND.n277 0.537563
R4739 VGND.n1 VGND 0.531208
R4740 VGND.n3133 VGND 0.531208
R4741 VGND.n1708 VGND.n1552 0.526527
R4742 VGND.n1705 VGND.n1704 0.526527
R4743 VGND.n2476 VGND.n2399 0.526527
R4744 VGND.n2324 VGND.n2322 0.526527
R4745 VGND.n261 VGND.n259 0.526527
R4746 VGND.n1532 VGND.n1531 0.500125
R4747 VGND.n1831 VGND.n1830 0.500125
R4748 VGND.n1179 VGND.n1178 0.500125
R4749 VGND.n2151 VGND.n2150 0.500125
R4750 VGND.n759 VGND.n758 0.500125
R4751 VGND.n2659 VGND.n2658 0.500125
R4752 VGND.n3382 VGND.n3381 0.482665
R4753 VGND.n3049 VGND.n0 0.473674
R4754 VGND.n329 VGND.n328 0.467019
R4755 VGND.n350 VGND.n228 0.467019
R4756 VGND.n3220 VGND.n3201 0.467019
R4757 VGND.n3273 VGND.n78 0.467019
R4758 VGND.n3294 VGND 0.448179
R4759 VGND.n525 VGND.n523 0.448052
R4760 VGND.n1359 VGND.n1358 0.448052
R4761 VGND.n1515 VGND.n1514 0.448052
R4762 VGND.n232 VGND.n210 0.426643
R4763 VGND.n1669 VGND.n1578 0.417891
R4764 VGND.n1663 VGND.n1662 0.417891
R4765 VGND.n1930 VGND.n1918 0.417891
R4766 VGND.n1925 VGND.n1924 0.417891
R4767 VGND.n2547 VGND.n944 0.417891
R4768 VGND.n2544 VGND.n2543 0.417891
R4769 VGND.n2541 VGND.n2540 0.417891
R4770 VGND.n1757 VGND.n1741 0.417891
R4771 VGND.n2442 VGND.n2435 0.417891
R4772 VGND.n2358 VGND.n2351 0.417891
R4773 VGND.n1059 VGND.n278 0.417891
R4774 VGND.n1060 VGND.n1055 0.417891
R4775 VGND.n3040 VGND.n3039 0.417891
R4776 VGND.n3036 VGND.n3035 0.417891
R4777 VGND.n255 VGND.n240 0.417891
R4778 VGND.n2387 VGND.n1016 0.410656
R4779 VGND.n3430 VGND.n58 0.409011
R4780 VGND.n3444 VGND.n40 0.409011
R4781 VGND.n33 VGND.n32 0.409011
R4782 VGND.n3464 VGND.n3 0.409011
R4783 VGND.n7 VGND.n6 0.409011
R4784 VGND.n8 VGND.n4 0.409011
R4785 VGND.n3377 VGND.n81 0.409011
R4786 VGND.n97 VGND.n92 0.409011
R4787 VGND.n3316 VGND.n115 0.409011
R4788 VGND.n3320 VGND.n3319 0.409011
R4789 VGND.n3324 VGND.n3323 0.409011
R4790 VGND.n3352 VGND.n3341 0.409011
R4791 VGND.n625 VGND.n610 0.409011
R4792 VGND.n618 VGND.n617 0.409011
R4793 VGND.n1418 VGND.n1415 0.409011
R4794 VGND.n1720 VGND.n1541 0.409011
R4795 VGND.n1710 VGND.n1709 0.409011
R4796 VGND.n877 VGND.n876 0.409011
R4797 VGND.n1839 VGND.n1290 0.409011
R4798 VGND.n1843 VGND.n1289 0.409011
R4799 VGND.n1816 VGND.n1763 0.409011
R4800 VGND.n1810 VGND.n1809 0.409011
R4801 VGND.n1780 VGND.n1779 0.409011
R4802 VGND.n2028 VGND.n1225 0.409011
R4803 VGND.n1995 VGND.n1993 0.409011
R4804 VGND.n2510 VGND.n2509 0.409011
R4805 VGND.n2504 VGND.n997 0.409011
R4806 VGND.n2497 VGND.n2397 0.409011
R4807 VGND.n2416 VGND.n2414 0.409011
R4808 VGND.n1043 VGND.n1039 0.409011
R4809 VGND.n258 VGND.n256 0.409011
R4810 VGND.n2055 VGND.n2054 0.383542
R4811 VGND.n1834 VGND.n1297 0.381255
R4812 VGND.n2656 VGND.n702 0.3805
R4813 VGND.n670 VGND.n570 0.3805
R4814 VGND.n2923 VGND.n2922 0.3805
R4815 VGND.n2967 VGND.n2966 0.3805
R4816 VGND.n2527 VGND.n2526 0.3805
R4817 VGND.n2609 VGND.n2608 0.3805
R4818 VGND.n2293 VGND.n505 0.3805
R4819 VGND.n1118 VGND.n568 0.3805
R4820 VGND.n757 VGND.n722 0.3805
R4821 VGND.n2657 VGND.n723 0.3805
R4822 VGND.n1380 VGND.n826 0.3805
R4823 VGND.n1985 VGND.n983 0.3805
R4824 VGND.n1178 VGND.n1162 0.3805
R4825 VGND.n2150 VGND.n1163 0.3805
R4826 VGND.n758 VGND.n741 0.3805
R4827 VGND.n2658 VGND.n742 0.3805
R4828 VGND.n1531 VGND.n1530 0.3805
R4829 VGND.n1830 VGND.n1278 0.3805
R4830 VGND.n2965 VGND.n2964 0.3805
R4831 VGND.n2924 VGND.n509 0.3805
R4832 VGND.n2873 VGND.n2872 0.3805
R4833 VGND.n2655 VGND.n2654 0.3805
R4834 VGND.n2610 VGND.n763 0.3805
R4835 VGND.n2528 VGND.n925 0.3805
R4836 VGND.n761 VGND.n672 0.3805
R4837 VGND.n2871 VGND.n2870 0.3805
R4838 VGND.n2926 VGND.n2925 0.3805
R4839 VGND.n530 VGND.n506 0.3805
R4840 VGND.n2530 VGND.n2529 0.3805
R4841 VGND.n2612 VGND.n2611 0.3805
R4842 VGND.n874 VGND.n863 0.376971
R4843 uio_oe[7] VGND.n3491 0.371345
R4844 VGND VGND.n3295 0.366908
R4845 VGND.n3049 VGND.n3048 0.364419
R4846 VGND.n3297 VGND.n116 0.358995
R4847 VGND.n2823 VGND.n680 0.358542
R4848 VGND.n1430 VGND.n1429 0.358542
R4849 VGND.n2635 VGND.n2634 0.358542
R4850 VGND.n1969 VGND.n1243 0.358542
R4851 VGND.n1438 VGND.n1437 0.340926
R4852 VGND.n3048 VGND.n3047 0.335802
R4853 VGND.n3469 uo_out[0] 0.3295
R4854 VGND.n3470 uo_out[1] 0.3295
R4855 VGND.n3471 uo_out[2] 0.3295
R4856 VGND.n3472 uo_out[3] 0.3295
R4857 VGND.n3473 uo_out[4] 0.3295
R4858 VGND.n3474 uo_out[5] 0.3295
R4859 VGND.n3475 uo_out[6] 0.3295
R4860 VGND.n3476 uo_out[7] 0.3295
R4861 VGND.n3477 uio_out[0] 0.3295
R4862 VGND.n3478 uio_out[1] 0.3295
R4863 VGND.n3479 uio_out[2] 0.3295
R4864 VGND.n3480 uio_out[3] 0.3295
R4865 VGND.n3481 uio_out[4] 0.3295
R4866 VGND.n3482 uio_out[5] 0.3295
R4867 VGND.n3483 uio_out[6] 0.3295
R4868 VGND.n3484 uio_out[7] 0.3295
R4869 VGND.n3485 uio_oe[0] 0.3295
R4870 VGND.n3486 uio_oe[1] 0.3295
R4871 VGND.n3487 uio_oe[2] 0.3295
R4872 VGND.n3488 uio_oe[3] 0.3295
R4873 VGND.n3489 uio_oe[4] 0.3295
R4874 VGND.n3490 uio_oe[5] 0.3295
R4875 VGND.n3491 uio_oe[6] 0.3295
R4876 VGND.n1704 VGND.n1703 0.307349
R4877 VGND.n2185 VGND.n2184 0.305262
R4878 VGND.n2201 VGND.n1158 0.305262
R4879 VGND.n2202 VGND.n1157 0.305262
R4880 VGND.n2215 VGND.n2214 0.305262
R4881 VGND.n2278 VGND.n2277 0.305262
R4882 VGND.n2263 VGND.n2262 0.305262
R4883 VGND.n1142 VGND.n1140 0.305262
R4884 VGND.n2237 VGND.n1151 0.305262
R4885 VGND.n2232 VGND.n2227 0.305262
R4886 VGND.n2939 VGND.n521 0.305262
R4887 VGND.n2132 VGND.n2131 0.305262
R4888 VGND.n1217 VGND.n1216 0.305262
R4889 VGND.n2118 VGND.n2117 0.305262
R4890 VGND.n2106 VGND.n1221 0.305262
R4891 VGND.n2060 VGND.n2058 0.305262
R4892 VGND.n2069 VGND.n2068 0.305262
R4893 VGND.n2067 VGND.n2064 0.305262
R4894 VGND.n2904 VGND.n576 0.305262
R4895 VGND.n2903 VGND.n577 0.305262
R4896 VGND.n2892 VGND.n2891 0.305262
R4897 VGND.n2692 VGND.n2691 0.305262
R4898 VGND.n2708 VGND.n737 0.305262
R4899 VGND.n2709 VGND.n736 0.305262
R4900 VGND.n2722 VGND.n2721 0.305262
R4901 VGND.n2742 VGND.n2741 0.305262
R4902 VGND.n2758 VGND.n710 0.305262
R4903 VGND.n2765 VGND.n2764 0.305262
R4904 VGND.n2785 VGND.n694 0.305262
R4905 VGND.n2380 VGND.n2379 0.298799
R4906 VGND.n2182 VGND.n2181 0.298074
R4907 VGND.n2135 VGND.n2134 0.298074
R4908 VGND.n2689 VGND.n2688 0.298074
R4909 VGND.n471 VGND 0.286698
R4910 VGND.n1325 VGND.n1297 0.281546
R4911 VGND.n2164 VGND.n233 0.281132
R4912 VGND.n2302 VGND.n2301 0.278782
R4913 VGND VGND.n3468 0.268171
R4914 VGND.n1700 VGND.n1699 0.263514
R4915 VGND.n2474 VGND.n2473 0.263514
R4916 VGND.n2331 VGND.n1032 0.263514
R4917 VGND.n3021 VGND.n3020 0.263514
R4918 VGND.n3296 VGND 0.260439
R4919 VGND.n2173 VGND.n1171 0.259086
R4920 VGND.n560 VGND.n546 0.259086
R4921 VGND.n554 VGND.n553 0.259086
R4922 VGND.n2141 VGND.n1198 0.259086
R4923 VGND.n2888 VGND.n582 0.259086
R4924 VGND.n2882 VGND.n2881 0.259086
R4925 VGND.n2103 VGND.n2039 0.259086
R4926 VGND.n2099 VGND.n2098 0.259086
R4927 VGND.n2836 VGND.n2835 0.259086
R4928 VGND.n2846 VGND.n2841 0.259086
R4929 VGND.n2680 VGND.n750 0.259086
R4930 VGND.n818 VGND.n804 0.259086
R4931 VGND.n812 VGND.n811 0.259086
R4932 VGND.n1341 VGND.n1313 0.259086
R4933 VGND.n1346 VGND.n1311 0.259086
R4934 VGND.n1015 VGND.n1005 0.2565
R4935 VGND.n3467 VGND.n1 0.249698
R4936 VGND.n1782 VGND.n1778 0.239381
R4937 VGND.n1998 VGND.n1994 0.239381
R4938 VGND VGND.n2596 0.237784
R4939 VGND.n2379 VGND.n116 0.23574
R4940 VGND.n963 VGND.n962 0.225061
R4941 VGND.n971 VGND.n970 0.225061
R4942 VGND.n2380 VGND.n2376 0.224703
R4943 VGND.n2297 VGND.n237 0.218753
R4944 VGND.n621 VGND.n620 0.204755
R4945 VGND.n2538 VGND.n948 0.204755
R4946 VGND.n960 VGND.n948 0.204755
R4947 VGND.n2596 VGND 0.200023
R4948 VGND VGND.n2182 0.199635
R4949 VGND.n2134 VGND 0.199635
R4950 VGND VGND.n2689 0.199635
R4951 VGND.n231 VGND.n181 0.198729
R4952 VGND.n2298 VGND.n2297 0.196532
R4953 VGND.n1049 VGND.n234 0.196532
R4954 VGND.n2301 VGND.n2300 0.195539
R4955 VGND.n3054 VGND.n3053 0.194976
R4956 VGND.n2082 VGND.n2081 0.192021
R4957 VGND.n3047 VGND.n234 0.18942
R4958 VGND.n2376 VGND.n1019 0.184476
R4959 VGND.n330 VGND.n230 0.1838
R4960 VGND.n3383 VGND.n3382 0.1838
R4961 VGND.n2419 VGND.n2415 0.180304
R4962 VGND.n885 VGND 0.17983
R4963 VGND.n968 VGND 0.17983
R4964 VGND.n536 VGND.n526 0.179521
R4965 VGND.n1430 VGND.n1421 0.179521
R4966 VGND.n1969 VGND.n1968 0.179521
R4967 VGND VGND.n551 0.179485
R4968 VGND VGND.n615 0.179485
R4969 VGND.n2843 VGND 0.179485
R4970 VGND VGND.n809 0.179485
R4971 VGND.n2305 VGND.n2304 0.175416
R4972 VGND.n2387 VGND.n2386 0.173577
R4973 VGND.n2607 VGND.n830 0.1603
R4974 VGND.n1984 VGND.n1233 0.1603
R4975 VGND.n1876 VGND.n1277 0.1603
R4976 VGND.n1832 VGND.n1727 0.1603
R4977 VGND.n2580 VGND.n2572 0.1603
R4978 VGND.n2531 VGND.n825 0.1603
R4979 VGND.n2608 VGND.n827 0.159712
R4980 VGND.n1385 VGND.n1380 0.159712
R4981 VGND.n1530 VGND.n1529 0.159712
R4982 VGND.n1532 VGND.n760 0.159712
R4983 VGND.n2653 VGND.n763 0.159712
R4984 VGND.n2613 VGND.n2612 0.159712
R4985 VGND.n2259 VGND 0.158169
R4986 VGND VGND.n709 0.158169
R4987 VGND.n2794 VGND 0.158169
R4988 VGND VGND.n880 0.156867
R4989 VGND.n2424 VGND.n2419 0.151658
R4990 VGND.n2170 VGND.n2169 0.143027
R4991 VGND.n1196 VGND.n1195 0.143027
R4992 VGND.n2677 VGND.n2676 0.143027
R4993 VGND.n2170 VGND 0.14207
R4994 VGND.n551 VGND 0.14207
R4995 VGND VGND.n1196 0.14207
R4996 VGND.n615 VGND 0.14207
R4997 VGND.n2677 VGND 0.14207
R4998 VGND.n2843 VGND 0.14207
R4999 VGND.n809 VGND 0.14207
R5000 VGND VGND.n1782 0.14207
R5001 VGND.n1998 VGND 0.14207
R5002 VGND.n885 VGND 0.141725
R5003 VGND.n968 VGND 0.141725
R5004 VGND.n1297 VGND.n233 0.141676
R5005 VGND.n3111 VGND.n3105 0.141672
R5006 VGND.n3143 VGND.n211 0.141672
R5007 VGND.n2967 VGND.n504 0.137387
R5008 VGND.n2293 VGND.n2292 0.137387
R5009 VGND.n2196 VGND.n1162 0.137387
R5010 VGND.n2166 VGND.n1179 0.137387
R5011 VGND.n2964 VGND.n2963 0.137387
R5012 VGND.n2927 VGND.n530 0.137387
R5013 VGND.n891 VGND.n890 0.13667
R5014 VGND.n2526 VGND.n2525 0.126812
R5015 VGND.n2017 VGND.n1985 0.126812
R5016 VGND.n1797 VGND.n1278 0.126812
R5017 VGND.n1831 VGND.n1829 0.126812
R5018 VGND.n2485 VGND.n925 0.126812
R5019 VGND.n2530 VGND.n982 0.126812
R5020 VGND.n2105 VGND.n2104 0.126617
R5021 VGND.n2771 VGND.n702 0.125637
R5022 VGND.n2735 VGND.n723 0.125637
R5023 VGND.n2703 VGND.n742 0.125637
R5024 VGND.n2673 VGND.n2659 0.125637
R5025 VGND.n2654 VGND.n669 0.125637
R5026 VGND.n2869 VGND.n672 0.125637
R5027 VGND.n3447 VGND.n37 0.1255
R5028 VGND.n3174 VGND.n3173 0.1255
R5029 VGND.n3356 VGND.n106 0.1255
R5030 VGND.n3297 VGND.n3296 0.122556
R5031 VGND.n3105 VGND 0.121778
R5032 VGND.n3168 VGND 0.121778
R5033 VGND.n2890 VGND.n2889 0.120632
R5034 VGND.n1713 VGND 0.120408
R5035 VGND.n54 VGND.n53 0.120292
R5036 VGND.n54 VGND.n41 0.120292
R5037 VGND.n3427 VGND.n59 0.120292
R5038 VGND.n3427 VGND.n3426 0.120292
R5039 VGND.n3425 VGND.n61 0.120292
R5040 VGND.n62 VGND.n61 0.120292
R5041 VGND.n3418 VGND.n3410 0.120292
R5042 VGND.n3418 VGND.n3417 0.120292
R5043 VGND.n3416 VGND.n3413 0.120292
R5044 VGND.n3413 VGND.n3412 0.120292
R5045 VGND.n3443 VGND.n3442 0.120292
R5046 VGND.n3439 VGND.n3438 0.120292
R5047 VGND.n51 VGND.n43 0.120292
R5048 VGND.n46 VGND.n43 0.120292
R5049 VGND.n46 VGND.n45 0.120292
R5050 VGND.n12 VGND.n11 0.120292
R5051 VGND.n3456 VGND.n18 0.120292
R5052 VGND.n19 VGND.n18 0.120292
R5053 VGND.n3450 VGND.n20 0.120292
R5054 VGND.n34 VGND.n23 0.120292
R5055 VGND.n28 VGND.n23 0.120292
R5056 VGND.n28 VGND.n27 0.120292
R5057 VGND.n3141 VGND.n213 0.120292
R5058 VGND.n3136 VGND.n213 0.120292
R5059 VGND.n3136 VGND.n3135 0.120292
R5060 VGND.n3092 VGND.n3091 0.120292
R5061 VGND.n3126 VGND.n3099 0.120292
R5062 VGND.n3120 VGND.n3099 0.120292
R5063 VGND.n3119 VGND.n3102 0.120292
R5064 VGND.n3112 VGND.n3111 0.120292
R5065 VGND.n3159 VGND.n3158 0.120292
R5066 VGND.n3158 VGND.n3147 0.120292
R5067 VGND.n3153 VGND.n3152 0.120292
R5068 VGND.n3152 VGND.n3149 0.120292
R5069 VGND.n3187 VGND.n3186 0.120292
R5070 VGND.n3186 VGND.n190 0.120292
R5071 VGND.n3181 VGND.n3180 0.120292
R5072 VGND.n3180 VGND.n193 0.120292
R5073 VGND.n3172 VGND.n3171 0.120292
R5074 VGND.n3306 VGND.n3301 0.120292
R5075 VGND.n3301 VGND.n80 0.120292
R5076 VGND.n3374 VGND.n82 0.120292
R5077 VGND.n3374 VGND.n3373 0.120292
R5078 VGND.n3372 VGND.n84 0.120292
R5079 VGND.n85 VGND.n84 0.120292
R5080 VGND.n3365 VGND.n88 0.120292
R5081 VGND.n3365 VGND.n3364 0.120292
R5082 VGND.n3363 VGND.n90 0.120292
R5083 VGND.n91 VGND.n90 0.120292
R5084 VGND.n105 VGND.n104 0.120292
R5085 VGND.n101 VGND.n100 0.120292
R5086 VGND.n3312 VGND.n3300 0.120292
R5087 VGND.n3313 VGND.n3312 0.120292
R5088 VGND.n3314 VGND.n3313 0.120292
R5089 VGND.n3325 VGND.n114 0.120292
R5090 VGND.n3333 VGND.n109 0.120292
R5091 VGND.n3337 VGND.n109 0.120292
R5092 VGND.n3339 VGND.n3338 0.120292
R5093 VGND.n3351 VGND.n3350 0.120292
R5094 VGND.n3350 VGND.n3342 0.120292
R5095 VGND.n3344 VGND.n3342 0.120292
R5096 VGND.n2175 VGND.n2174 0.120292
R5097 VGND.n2175 VGND.n1170 0.120292
R5098 VGND.n2181 VGND.n1170 0.120292
R5099 VGND.n2204 VGND.n2203 0.120292
R5100 VGND.n2204 VGND.n1156 0.120292
R5101 VGND.n2209 VGND.n1156 0.120292
R5102 VGND.n2210 VGND.n2209 0.120292
R5103 VGND.n2211 VGND.n2210 0.120292
R5104 VGND.n2211 VGND.n1154 0.120292
R5105 VGND.n2216 VGND.n1154 0.120292
R5106 VGND.n2279 VGND.n1127 0.120292
R5107 VGND.n2274 VGND.n1127 0.120292
R5108 VGND.n2274 VGND.n2273 0.120292
R5109 VGND.n2273 VGND.n2272 0.120292
R5110 VGND.n2272 VGND.n1129 0.120292
R5111 VGND.n2267 VGND.n1129 0.120292
R5112 VGND.n2267 VGND.n2266 0.120292
R5113 VGND.n2266 VGND.n2265 0.120292
R5114 VGND.n2265 VGND.n1131 0.120292
R5115 VGND.n2250 VGND.n1139 0.120292
R5116 VGND.n2246 VGND.n1139 0.120292
R5117 VGND.n2246 VGND.n2245 0.120292
R5118 VGND.n2245 VGND.n2244 0.120292
R5119 VGND.n2244 VGND.n1149 0.120292
R5120 VGND.n2239 VGND.n1149 0.120292
R5121 VGND.n2239 VGND.n2238 0.120292
R5122 VGND.n2231 VGND.n2230 0.120292
R5123 VGND.n2949 VGND.n2948 0.120292
R5124 VGND.n2948 VGND.n2947 0.120292
R5125 VGND.n2947 VGND.n519 0.120292
R5126 VGND.n2942 VGND.n519 0.120292
R5127 VGND.n2942 VGND.n2941 0.120292
R5128 VGND.n2941 VGND.n2940 0.120292
R5129 VGND.n2936 VGND.n2935 0.120292
R5130 VGND.n2935 VGND.n524 0.120292
R5131 VGND.n2931 VGND.n524 0.120292
R5132 VGND.n559 VGND.n558 0.120292
R5133 VGND.n558 VGND.n547 0.120292
R5134 VGND.n552 VGND.n547 0.120292
R5135 VGND.n2140 VGND.n2139 0.120292
R5136 VGND.n2139 VGND.n1199 0.120292
R5137 VGND.n2135 VGND.n1199 0.120292
R5138 VGND.n2119 VGND.n1215 0.120292
R5139 VGND.n2114 VGND.n1215 0.120292
R5140 VGND.n2114 VGND.n2113 0.120292
R5141 VGND.n2113 VGND.n2112 0.120292
R5142 VGND.n2112 VGND.n1219 0.120292
R5143 VGND.n2108 VGND.n1219 0.120292
R5144 VGND.n2108 VGND.n2107 0.120292
R5145 VGND.n2102 VGND.n2101 0.120292
R5146 VGND.n2087 VGND.n2053 0.120292
R5147 VGND.n2080 VGND.n2053 0.120292
R5148 VGND.n2079 VGND.n2078 0.120292
R5149 VGND.n2078 VGND.n2059 0.120292
R5150 VGND.n2073 VGND.n2059 0.120292
R5151 VGND.n2073 VGND.n2072 0.120292
R5152 VGND.n2072 VGND.n2071 0.120292
R5153 VGND.n2071 VGND.n2062 0.120292
R5154 VGND.n2066 VGND.n2065 0.120292
R5155 VGND.n2902 VGND.n2901 0.120292
R5156 VGND.n2901 VGND.n578 0.120292
R5157 VGND.n2896 VGND.n578 0.120292
R5158 VGND.n2896 VGND.n2895 0.120292
R5159 VGND.n2895 VGND.n2894 0.120292
R5160 VGND.n2894 VGND.n580 0.120292
R5161 VGND.n2887 VGND.n2886 0.120292
R5162 VGND.n2886 VGND.n584 0.120292
R5163 VGND.n665 VGND.n596 0.120292
R5164 VGND.n661 VGND.n596 0.120292
R5165 VGND.n661 VGND.n660 0.120292
R5166 VGND.n660 VGND.n659 0.120292
R5167 VGND.n659 VGND.n601 0.120292
R5168 VGND.n653 VGND.n601 0.120292
R5169 VGND.n653 VGND.n652 0.120292
R5170 VGND.n652 VGND.n651 0.120292
R5171 VGND.n651 VGND.n603 0.120292
R5172 VGND.n647 VGND.n603 0.120292
R5173 VGND.n624 VGND.n623 0.120292
R5174 VGND.n623 VGND.n611 0.120292
R5175 VGND.n2682 VGND.n2681 0.120292
R5176 VGND.n2682 VGND.n749 0.120292
R5177 VGND.n2688 VGND.n749 0.120292
R5178 VGND.n2711 VGND.n2710 0.120292
R5179 VGND.n2711 VGND.n735 0.120292
R5180 VGND.n2716 VGND.n735 0.120292
R5181 VGND.n2717 VGND.n2716 0.120292
R5182 VGND.n2718 VGND.n2717 0.120292
R5183 VGND.n2718 VGND.n733 0.120292
R5184 VGND.n2723 VGND.n733 0.120292
R5185 VGND.n2744 VGND.n715 0.120292
R5186 VGND.n2745 VGND.n2744 0.120292
R5187 VGND.n2746 VGND.n2745 0.120292
R5188 VGND.n2746 VGND.n713 0.120292
R5189 VGND.n2750 VGND.n713 0.120292
R5190 VGND.n2751 VGND.n2750 0.120292
R5191 VGND.n2751 VGND.n711 0.120292
R5192 VGND.n2756 VGND.n711 0.120292
R5193 VGND.n2757 VGND.n2756 0.120292
R5194 VGND.n2776 VGND.n2775 0.120292
R5195 VGND.n2776 VGND.n697 0.120292
R5196 VGND.n2780 VGND.n697 0.120292
R5197 VGND.n2781 VGND.n2780 0.120292
R5198 VGND.n2781 VGND.n695 0.120292
R5199 VGND.n2787 VGND.n695 0.120292
R5200 VGND.n2788 VGND.n2787 0.120292
R5201 VGND.n2819 VGND.n683 0.120292
R5202 VGND.n2820 VGND.n2819 0.120292
R5203 VGND VGND.n2820 0.120292
R5204 VGND.n2826 VGND.n2825 0.120292
R5205 VGND.n2831 VGND.n679 0.120292
R5206 VGND.n2832 VGND.n2831 0.120292
R5207 VGND.n2854 VGND.n2853 0.120292
R5208 VGND.n2853 VGND.n2839 0.120292
R5209 VGND.n2848 VGND.n2839 0.120292
R5210 VGND.n2848 VGND.n2847 0.120292
R5211 VGND.n1343 VGND.n1342 0.120292
R5212 VGND.n1343 VGND.n1312 0.120292
R5213 VGND.n1348 VGND.n1312 0.120292
R5214 VGND.n1349 VGND.n1348 0.120292
R5215 VGND.n1355 VGND.n1309 0.120292
R5216 VGND.n1357 VGND.n1356 0.120292
R5217 VGND.n1512 VGND.n1511 0.120292
R5218 VGND.n1511 VGND.n1364 0.120292
R5219 VGND.n1506 VGND.n1364 0.120292
R5220 VGND.n1506 VGND.n1505 0.120292
R5221 VGND.n1505 VGND.n1504 0.120292
R5222 VGND.n1504 VGND.n1367 0.120292
R5223 VGND.n1498 VGND.n1497 0.120292
R5224 VGND.n1481 VGND.n1480 0.120292
R5225 VGND.n1480 VGND.n1479 0.120292
R5226 VGND.n1479 VGND.n1390 0.120292
R5227 VGND.n1473 VGND.n1390 0.120292
R5228 VGND.n1473 VGND.n1472 0.120292
R5229 VGND.n1472 VGND.n1471 0.120292
R5230 VGND.n1471 VGND.n1395 0.120292
R5231 VGND.n1464 VGND.n1395 0.120292
R5232 VGND.n1464 VGND.n1463 0.120292
R5233 VGND.n1463 VGND.n1462 0.120292
R5234 VGND.n1450 VGND.n1411 0.120292
R5235 VGND.n1444 VGND.n1443 0.120292
R5236 VGND.n1443 VGND.n1417 0.120292
R5237 VGND.n1436 VGND.n1417 0.120292
R5238 VGND.n2639 VGND.n2638 0.120292
R5239 VGND.n2638 VGND.n775 0.120292
R5240 VGND.n2632 VGND.n775 0.120292
R5241 VGND.n2632 VGND.n2631 0.120292
R5242 VGND.n2631 VGND.n2630 0.120292
R5243 VGND.n2630 VGND.n778 0.120292
R5244 VGND.n2623 VGND.n2622 0.120292
R5245 VGND.n2622 VGND.n782 0.120292
R5246 VGND.n2617 VGND.n782 0.120292
R5247 VGND.n817 VGND.n816 0.120292
R5248 VGND.n816 VGND.n805 0.120292
R5249 VGND.n810 VGND.n805 0.120292
R5250 VGND.n1719 VGND.n1718 0.120292
R5251 VGND.n1712 VGND.n1550 0.120292
R5252 VGND.n1707 VGND.n1550 0.120292
R5253 VGND.n1707 VGND.n1706 0.120292
R5254 VGND.n1706 VGND.n1553 0.120292
R5255 VGND.n1698 VGND.n1553 0.120292
R5256 VGND.n1697 VGND.n1696 0.120292
R5257 VGND.n1682 VGND.n1567 0.120292
R5258 VGND.n1676 VGND.n1567 0.120292
R5259 VGND.n1676 VGND.n1675 0.120292
R5260 VGND.n1675 VGND.n1576 0.120292
R5261 VGND.n1668 VGND.n1667 0.120292
R5262 VGND.n1667 VGND.n1579 0.120292
R5263 VGND.n1659 VGND.n1584 0.120292
R5264 VGND.n1639 VGND.n1638 0.120292
R5265 VGND.n1638 VGND.n1602 0.120292
R5266 VGND.n1634 VGND.n1602 0.120292
R5267 VGND.n1634 VGND.n1633 0.120292
R5268 VGND.n1633 VGND.n1632 0.120292
R5269 VGND.n1632 VGND.n1607 0.120292
R5270 VGND.n2603 VGND.n834 0.120292
R5271 VGND.n837 VGND.n834 0.120292
R5272 VGND.n2591 VGND.n2590 0.120292
R5273 VGND.n2590 VGND.n2589 0.120292
R5274 VGND.n921 VGND.n852 0.120292
R5275 VGND.n855 VGND.n852 0.120292
R5276 VGND.n856 VGND.n855 0.120292
R5277 VGND.n914 VGND.n856 0.120292
R5278 VGND.n914 VGND.n913 0.120292
R5279 VGND.n913 VGND.n912 0.120292
R5280 VGND.n912 VGND.n858 0.120292
R5281 VGND.n907 VGND.n858 0.120292
R5282 VGND.n907 VGND.n906 0.120292
R5283 VGND.n892 VGND.n873 0.120292
R5284 VGND.n1841 VGND.n1840 0.120292
R5285 VGND.n1849 VGND.n1287 0.120292
R5286 VGND.n1855 VGND.n1287 0.120292
R5287 VGND.n1856 VGND.n1855 0.120292
R5288 VGND.n1857 VGND.n1856 0.120292
R5289 VGND.n1862 VGND.n1861 0.120292
R5290 VGND.n1885 VGND.n1884 0.120292
R5291 VGND.n1886 VGND.n1885 0.120292
R5292 VGND.n1893 VGND.n1269 0.120292
R5293 VGND.n1894 VGND.n1893 0.120292
R5294 VGND.n1980 VGND.n1239 0.120292
R5295 VGND.n1975 VGND.n1239 0.120292
R5296 VGND.n1974 VGND.n1973 0.120292
R5297 VGND.n1966 VGND.n1246 0.120292
R5298 VGND.n1964 VGND.n1247 0.120292
R5299 VGND.n1960 VGND.n1247 0.120292
R5300 VGND.n1960 VGND.n1959 0.120292
R5301 VGND.n1948 VGND.n1261 0.120292
R5302 VGND.n1943 VGND.n1261 0.120292
R5303 VGND.n1942 VGND.n1941 0.120292
R5304 VGND.n1941 VGND.n1266 0.120292
R5305 VGND.n1934 VGND.n1266 0.120292
R5306 VGND.n1934 VGND.n1933 0.120292
R5307 VGND.n2557 VGND.n935 0.120292
R5308 VGND.n2557 VGND.n2556 0.120292
R5309 VGND.n2556 VGND.n938 0.120292
R5310 VGND.n2552 VGND.n938 0.120292
R5311 VGND.n2552 VGND.n2551 0.120292
R5312 VGND.n2551 VGND.n2550 0.120292
R5313 VGND.n2550 VGND.n941 0.120292
R5314 VGND.n2546 VGND.n2545 0.120292
R5315 VGND.n2545 VGND.n945 0.120292
R5316 VGND.n978 VGND.n959 0.120292
R5317 VGND.n974 VGND.n959 0.120292
R5318 VGND.n974 VGND.n973 0.120292
R5319 VGND.n973 VGND.n965 0.120292
R5320 VGND.n1821 VGND.n1759 0.120292
R5321 VGND.n1820 VGND.n1819 0.120292
R5322 VGND.n1819 VGND.n1761 0.120292
R5323 VGND.n1815 VGND.n1814 0.120292
R5324 VGND.n1814 VGND.n1764 0.120292
R5325 VGND.n1808 VGND.n1764 0.120292
R5326 VGND.n1793 VGND.n1778 0.120292
R5327 VGND.n1786 VGND.n1785 0.120292
R5328 VGND.n2027 VGND.n2026 0.120292
R5329 VGND.n2009 VGND.n2008 0.120292
R5330 VGND.n2004 VGND.n2003 0.120292
R5331 VGND.n2003 VGND.n1994 0.120292
R5332 VGND.n2511 VGND.n995 0.120292
R5333 VGND.n2506 VGND.n995 0.120292
R5334 VGND.n2506 VGND.n2505 0.120292
R5335 VGND.n2501 VGND.n2500 0.120292
R5336 VGND.n2496 VGND.n2495 0.120292
R5337 VGND.n2495 VGND.n2398 0.120292
R5338 VGND.n2481 VGND.n2410 0.120292
R5339 VGND.n2470 VGND.n2469 0.120292
R5340 VGND.n2465 VGND.n2464 0.120292
R5341 VGND.n2464 VGND.n2415 0.120292
R5342 VGND.n2445 VGND.n2433 0.120292
R5343 VGND.n2441 VGND.n2440 0.120292
R5344 VGND.n2440 VGND.n2436 0.120292
R5345 VGND.n3041 VGND.n239 0.120292
R5346 VGND.n3034 VGND.n239 0.120292
R5347 VGND.n3033 VGND.n3032 0.120292
R5348 VGND.n3032 VGND.n257 0.120292
R5349 VGND.n3028 VGND.n257 0.120292
R5350 VGND.n3028 VGND.n3027 0.120292
R5351 VGND.n3027 VGND.n3026 0.120292
R5352 VGND.n3026 VGND.n260 0.120292
R5353 VGND.n3019 VGND.n260 0.120292
R5354 VGND.n3001 VGND.n3000 0.120292
R5355 VGND.n3000 VGND.n274 0.120292
R5356 VGND.n2996 VGND.n274 0.120292
R5357 VGND.n2996 VGND.n2995 0.120292
R5358 VGND.n2995 VGND.n276 0.120292
R5359 VGND.n2991 VGND.n276 0.120292
R5360 VGND.n2991 VGND.n2990 0.120292
R5361 VGND.n1063 VGND.n1058 0.120292
R5362 VGND.n1113 VGND.n1054 0.120292
R5363 VGND.n1109 VGND.n1054 0.120292
R5364 VGND.n1109 VGND.n1108 0.120292
R5365 VGND.n1108 VGND.n1107 0.120292
R5366 VGND.n1107 VGND.n1078 0.120292
R5367 VGND.n1102 VGND.n1078 0.120292
R5368 VGND.n1102 VGND.n1101 0.120292
R5369 VGND.n1101 VGND.n1100 0.120292
R5370 VGND.n1100 VGND 0.120292
R5371 VGND.n1095 VGND.n1094 0.120292
R5372 VGND.n2973 VGND.n2972 0.120292
R5373 VGND.n2973 VGND.n498 0.120292
R5374 VGND.n2977 VGND.n498 0.120292
R5375 VGND.n2978 VGND.n2977 0.120292
R5376 VGND.n2978 VGND.n496 0.120292
R5377 VGND.n2982 VGND.n496 0.120292
R5378 VGND.n2983 VGND.n2982 0.120292
R5379 VGND.n1041 VGND.n1040 0.120292
R5380 VGND.n2321 VGND.n1033 0.120292
R5381 VGND.n2329 VGND.n1033 0.120292
R5382 VGND.n2330 VGND.n2329 0.120292
R5383 VGND.n2335 VGND.n2334 0.120292
R5384 VGND.n2340 VGND.n1029 0.120292
R5385 VGND.n2341 VGND.n2340 0.120292
R5386 VGND.n2342 VGND.n2341 0.120292
R5387 VGND.n2366 VGND.n2365 0.120292
R5388 VGND.n2365 VGND.n2348 0.120292
R5389 VGND.n2361 VGND.n2348 0.120292
R5390 VGND.n2361 VGND.n2360 0.120292
R5391 VGND.n2357 VGND.n2356 0.120292
R5392 VGND.n2356 VGND.n2352 0.120292
R5393 VGND.n1531 VGND.n826 0.120125
R5394 VGND.n2609 VGND.n826 0.120125
R5395 VGND.n2610 VGND.n2609 0.120125
R5396 VGND.n2611 VGND.n2610 0.120125
R5397 VGND.n1830 VGND.n983 0.120125
R5398 VGND.n2527 VGND.n983 0.120125
R5399 VGND.n2528 VGND.n2527 0.120125
R5400 VGND.n2529 VGND.n2528 0.120125
R5401 VGND.n1178 VGND.n505 0.120125
R5402 VGND.n2966 VGND.n505 0.120125
R5403 VGND.n2966 VGND.n2965 0.120125
R5404 VGND.n2965 VGND.n506 0.120125
R5405 VGND.n2150 VGND.n568 0.120125
R5406 VGND.n2923 VGND.n568 0.120125
R5407 VGND.n2924 VGND.n2923 0.120125
R5408 VGND.n2925 VGND.n2924 0.120125
R5409 VGND.n758 VGND.n757 0.120125
R5410 VGND.n757 VGND.n670 0.120125
R5411 VGND.n2872 VGND.n670 0.120125
R5412 VGND.n2872 VGND.n2871 0.120125
R5413 VGND.n2658 VGND.n2657 0.120125
R5414 VGND.n2657 VGND.n2656 0.120125
R5415 VGND.n2656 VGND.n2655 0.120125
R5416 VGND.n2655 VGND.n761 0.120125
R5417 VGND.n116 VGND 0.114397
R5418 VGND.n330 VGND.n329 0.113648
R5419 VGND.n3383 VGND.n78 0.113648
R5420 VGND.n229 VGND 0.11275
R5421 VGND.n130 VGND.n129 0.111077
R5422 VGND.n135 VGND.n134 0.111077
R5423 VGND.n140 VGND.n139 0.111077
R5424 VGND.n145 VGND.n144 0.111077
R5425 VGND.n150 VGND.n149 0.111077
R5426 VGND.n155 VGND.n154 0.111077
R5427 VGND.n160 VGND.n159 0.111077
R5428 VGND.n165 VGND.n164 0.111077
R5429 VGND.n170 VGND.n169 0.111077
R5430 VGND.n2795 VGND.n2794 0.109992
R5431 VGND.n2304 VGND.n2303 0.10744
R5432 VGND.n2922 VGND.n2921 0.103312
R5433 VGND.n2091 VGND.n1118 0.103312
R5434 VGND.n2123 VGND.n1163 0.103312
R5435 VGND.n2151 VGND.n2149 0.103312
R5436 VGND.n2874 VGND.n509 0.103312
R5437 VGND.n2926 VGND.n567 0.103312
R5438 VGND.n1513 VGND.n1306 0.102062
R5439 VGND.n1683 VGND.n1682 0.102062
R5440 VGND.n1880 VGND.n1879 0.102062
R5441 VGND.n1794 VGND.n1793 0.102062
R5442 VGND.n3006 VGND.n3001 0.102062
R5443 VGND.n11 VGND 0.0981562
R5444 VGND.n3091 VGND 0.0981562
R5445 VGND VGND.n114 0.0981562
R5446 VGND.n2203 VGND 0.0981562
R5447 VGND.n2222 VGND 0.0981562
R5448 VGND.n2235 VGND 0.0981562
R5449 VGND.n2936 VGND 0.0981562
R5450 VGND VGND.n2119 0.0981562
R5451 VGND.n2040 VGND 0.0981562
R5452 VGND.n2066 VGND 0.0981562
R5453 VGND.n2902 VGND 0.0981562
R5454 VGND.n583 VGND 0.0981562
R5455 VGND.n2710 VGND 0.0981562
R5456 VGND.n2724 VGND 0.0981562
R5457 VGND.n2789 VGND 0.0981562
R5458 VGND VGND.n679 0.0981562
R5459 VGND VGND.n1309 0.0981562
R5460 VGND.n1481 VGND 0.0981562
R5461 VGND.n1427 VGND 0.0981562
R5462 VGND.n2623 VGND 0.0981562
R5463 VGND.n1627 VGND 0.0981562
R5464 VGND.n1848 VGND 0.0981562
R5465 VGND.n1884 VGND 0.0981562
R5466 VGND VGND.n1964 0.0981562
R5467 VGND.n1923 VGND 0.0981562
R5468 VGND.n279 VGND 0.0981562
R5469 VGND.n1095 VGND 0.0981562
R5470 VGND VGND.n494 0.0981562
R5471 VGND.n2357 VGND 0.0981562
R5472 VGND.n2949 VGND.n516 0.0968542
R5473 VGND.n666 VGND.n665 0.0968542
R5474 VGND.n2812 VGND.n2811 0.0968542
R5475 VGND.n2639 VGND.n770 0.0968542
R5476 VGND VGND.n1639 0.0968542
R5477 VGND.n1861 VGND 0.0968542
R5478 VGND.n2482 VGND.n2481 0.0968542
R5479 VGND.n2321 VGND.n2320 0.0968542
R5480 VGND.n1759 VGND 0.0955521
R5481 VGND VGND.n1806 0.0955521
R5482 VGND VGND.n1786 0.0955521
R5483 VGND VGND.n2009 0.0955521
R5484 VGND VGND.n2501 0.0955521
R5485 VGND VGND.n2470 0.0955521
R5486 VGND VGND.n2445 0.0955521
R5487 VGND.n2334 VGND 0.0955521
R5488 VGND.n2311 VGND.n1046 0.0950946
R5489 VGND.n2319 VGND.n2318 0.0950946
R5490 VGND.n249 VGND.n243 0.0950946
R5491 VGND.n3043 VGND.n238 0.0950946
R5492 VGND.n2570 VGND.n2569 0.0950946
R5493 VGND.n2563 VGND.n931 0.0950946
R5494 VGND.n1067 VGND.n1057 0.0950946
R5495 VGND.n1115 VGND.n1052 0.0950946
R5496 VGND.n2578 VGND.n2577 0.0950946
R5497 VGND.n2583 VGND.n2582 0.0950946
R5498 VGND.n1086 VGND.n1085 0.0950946
R5499 VGND.n2970 VGND.n501 0.0950946
R5500 VGND.n2961 VGND.n2960 0.0950946
R5501 VGND.n2954 VGND.n515 0.0950946
R5502 VGND.n2290 VGND.n2289 0.0950946
R5503 VGND.n2284 VGND.n2283 0.0950946
R5504 VGND.n2194 VGND.n2193 0.0950946
R5505 VGND.n2198 VGND.n1160 0.0950946
R5506 VGND.n2163 VGND.n2162 0.0950946
R5507 VGND.n2168 VGND.n1176 0.0950946
R5508 VGND.n2929 VGND.n528 0.0950946
R5509 VGND.n565 VGND.n532 0.0950946
R5510 VGND.n2257 VGND.n1134 0.0950946
R5511 VGND.n2252 VGND.n1137 0.0950946
R5512 VGND.n2127 VGND.n1207 0.0950946
R5513 VGND.n2121 VGND.n1211 0.0950946
R5514 VGND.n2147 VGND.n2146 0.0950946
R5515 VGND.n1194 VGND.n1193 0.0950946
R5516 VGND.n645 VGND.n606 0.0950946
R5517 VGND.n640 VGND.n609 0.0950946
R5518 VGND.n2878 VGND.n587 0.0950946
R5519 VGND.n667 VGND.n591 0.0950946
R5520 VGND.n2095 VGND.n2045 0.0950946
R5521 VGND.n2089 VGND.n2049 0.0950946
R5522 VGND.n2919 VGND.n2918 0.0950946
R5523 VGND.n2911 VGND.n2910 0.0950946
R5524 VGND.n2701 VGND.n2700 0.0950946
R5525 VGND.n2705 VGND.n739 0.0950946
R5526 VGND.n2671 VGND.n2670 0.0950946
R5527 VGND.n2675 VGND.n755 0.0950946
R5528 VGND.n2867 VGND.n2866 0.0950946
R5529 VGND.n2859 VGND.n2858 0.0950946
R5530 VGND.n2798 VGND.n2797 0.0950946
R5531 VGND.n2810 VGND.n686 0.0950946
R5532 VGND.n2733 VGND.n2732 0.0950946
R5533 VGND.n2737 VGND.n720 0.0950946
R5534 VGND.n2769 VGND.n2768 0.0950946
R5535 VGND.n2773 VGND.n700 0.0950946
R5536 VGND.n1326 VGND.n1323 0.0950946
R5537 VGND.n1335 VGND.n1315 0.0950946
R5538 VGND.n2615 VGND.n787 0.0950946
R5539 VGND.n823 VGND.n790 0.0950946
R5540 VGND.n2651 VGND.n2650 0.0950946
R5541 VGND.n2644 VGND.n769 0.0950946
R5542 VGND.n1383 VGND.n1382 0.0950946
R5543 VGND.n1487 VGND.n1378 0.0950946
R5544 VGND.n1527 VGND.n1526 0.0950946
R5545 VGND.n1520 VGND.n1305 0.0950946
R5546 VGND.n1407 VGND.n1406 0.0950946
R5547 VGND.n1452 VGND.n1405 0.0950946
R5548 VGND.n1257 VGND.n1256 0.0950946
R5549 VGND.n1950 VGND.n1255 0.0950946
R5550 VGND.n2523 VGND.n2522 0.0950946
R5551 VGND.n2515 VGND.n2514 0.0950946
R5552 VGND.n1617 VGND.n1616 0.0950946
R5553 VGND.n2605 VGND.n832 0.0950946
R5554 VGND.n1690 VGND.n1562 0.0950946
R5555 VGND.n1684 VGND.n1565 0.0950946
R5556 VGND.n1725 VGND.n1724 0.0950946
R5557 VGND.n1547 VGND.n1546 0.0950946
R5558 VGND.n900 VGND.n866 0.0950946
R5559 VGND.n894 VGND.n869 0.0950946
R5560 VGND.n1651 VGND.n1590 0.0950946
R5561 VGND.n1645 VGND.n1593 0.0950946
R5562 VGND.n2021 VGND.n1230 0.0950946
R5563 VGND.n2015 VGND.n1987 0.0950946
R5564 VGND.n1909 VGND.n1908 0.0950946
R5565 VGND.n1982 VGND.n1237 0.0950946
R5566 VGND.n1835 VGND.n1296 0.0950946
R5567 VGND.n1735 VGND.n1734 0.0950946
R5568 VGND.n2535 VGND.n951 0.0950946
R5569 VGND.n980 VGND.n955 0.0950946
R5570 VGND.n1874 VGND.n1873 0.0950946
R5571 VGND.n1878 VGND.n1275 0.0950946
R5572 VGND.n1801 VGND.n1769 0.0950946
R5573 VGND.n1795 VGND.n1773 0.0950946
R5574 VGND.n1749 VGND.n1743 0.0950946
R5575 VGND.n1827 VGND.n1740 0.0950946
R5576 VGND.n2427 VGND.n2426 0.0950946
R5577 VGND.n2452 VGND.n2423 0.0950946
R5578 VGND.n2489 VGND.n2402 0.0950946
R5579 VGND.n2483 VGND.n2406 0.0950946
R5580 VGND.n2374 VGND.n2373 0.0950946
R5581 VGND.n2346 VGND.n1022 0.0950946
R5582 VGND.n3016 VGND.n266 0.0950946
R5583 VGND.n3005 VGND.n3002 0.0950946
R5584 VGND.n52 VGND 0.09425
R5585 VGND.n3142 VGND 0.09425
R5586 VGND VGND.n3307 0.09425
R5587 VGND.n3168 VGND.n3166 0.0934947
R5588 VGND.n2931 VGND.n2930 0.0916458
R5589 VGND.n647 VGND.n646 0.0916458
R5590 VGND.n2617 VGND.n2616 0.0916458
R5591 VGND.n864 VGND.n862 0.0916458
R5592 VGND.n2342 VGND.n1024 0.0916458
R5593 VGND.n2921 VGND.n570 0.0915625
R5594 VGND.n2091 VGND.n722 0.0915625
R5595 VGND.n2123 VGND.n741 0.0915625
R5596 VGND.n2149 VGND.n759 0.0915625
R5597 VGND.n2874 VGND.n2873 0.0915625
R5598 VGND.n2870 VGND.n567 0.0915625
R5599 VGND.n2378 VGND 0.0907344
R5600 VGND.n129 VGND 0.0906442
R5601 VGND.n134 VGND 0.0906442
R5602 VGND.n139 VGND 0.0906442
R5603 VGND.n144 VGND 0.0906442
R5604 VGND.n149 VGND 0.0906442
R5605 VGND.n154 VGND 0.0906442
R5606 VGND.n159 VGND 0.0906442
R5607 VGND.n164 VGND 0.0906442
R5608 VGND.n169 VGND 0.0906442
R5609 VGND.n2937 VGND.n523 0.0900105
R5610 VGND.n2814 VGND.n2813 0.0900105
R5611 VGND.n2302 VGND.n2298 0.0898892
R5612 VGND.n2303 VGND.n1049 0.0898892
R5613 VGND.n3434 VGND 0.0881354
R5614 VGND.n3165 VGND 0.0881354
R5615 VGND.n79 VGND 0.0881354
R5616 VGND.n2220 VGND.n1120 0.0864375
R5617 VGND.n2101 VGND.n2041 0.0864375
R5618 VGND.n2728 VGND.n725 0.0864375
R5619 VGND.n1588 VGND.n1584 0.0864375
R5620 VGND.n2026 VGND.n1226 0.0864375
R5621 VGND.n1064 VGND.n1063 0.0864375
R5622 VGND.n3468 VGND.n0 0.0853293
R5623 VGND.n2192 VGND.n2191 0.0838333
R5624 VGND.n1126 VGND.n1122 0.0838333
R5625 VGND.n2251 VGND.n1138 0.0838333
R5626 VGND.n2959 VGND.n2958 0.0838333
R5627 VGND.n543 VGND.n542 0.0838333
R5628 VGND.n2128 VGND.n1206 0.0838333
R5629 VGND.n2051 VGND.n2050 0.0838333
R5630 VGND.n2917 VGND.n572 0.0838333
R5631 VGND.n2912 VGND.n2906 0.0838333
R5632 VGND.n634 VGND.n633 0.0838333
R5633 VGND.n2699 VGND.n2698 0.0838333
R5634 VGND.n727 VGND.n719 0.0838333
R5635 VGND.n2774 VGND.n699 0.0838333
R5636 VGND.n2838 VGND.n677 0.0838333
R5637 VGND.n1525 VGND.n1524 0.0838333
R5638 VGND.n1492 VGND.n1376 0.0838333
R5639 VGND.n1402 VGND.n1399 0.0838333
R5640 VGND.n1451 VGND.n1410 0.0838333
R5641 VGND.n2649 VGND.n2648 0.0838333
R5642 VGND.n799 VGND.n795 0.0838333
R5643 VGND.n1691 VGND.n1561 0.0838333
R5644 VGND.n1595 VGND.n1594 0.0838333
R5645 VGND.n1614 VGND.n1613 0.0838333
R5646 VGND.n2604 VGND.n833 0.0838333
R5647 VGND.n2576 VGND.n849 0.0838333
R5648 VGND.n1872 VGND.n1871 0.0838333
R5649 VGND.n1903 VGND.n1900 0.0838333
R5650 VGND.n1949 VGND.n1260 0.0838333
R5651 VGND.n2568 VGND.n2567 0.0838333
R5652 VGND.n1989 VGND.n1988 0.0838333
R5653 VGND.n2490 VGND.n2401 0.0838333
R5654 VGND.n3011 VGND.n269 0.0838333
R5655 VGND.n1072 VGND.n1056 0.0838333
R5656 VGND.n1083 VGND.n1081 0.0838333
R5657 VGND.n2971 VGND.n500 0.0838333
R5658 VGND.n2312 VGND.n1038 0.0838333
R5659 VGND.n2347 VGND.n1027 0.0838333
R5660 VGND.n2611 VGND 0.0827875
R5661 VGND.n2529 VGND 0.0827875
R5662 VGND.n506 VGND 0.0827875
R5663 VGND.n2925 VGND 0.0827875
R5664 VGND.n2871 VGND 0.0827875
R5665 VGND.n761 VGND 0.0827875
R5666 VGND VGND.n880 0.082648
R5667 VGND.n1713 VGND 0.082648
R5668 VGND.n2430 VGND 0.0773229
R5669 VGND.n3054 VGND.n228 0.0766574
R5670 VGND.n3201 VGND.n181 0.0766574
R5671 VGND.n1167 VGND.n1165 0.0760208
R5672 VGND.n2129 VGND.n1203 0.0760208
R5673 VGND.n746 VGND.n744 0.0760208
R5674 VGND.n1303 VGND.n1301 0.0760208
R5675 VGND.n1692 VGND.n1557 0.0760208
R5676 VGND.n1282 VGND.n1280 0.0760208
R5677 VGND.n1803 VGND.n1766 0.0760208
R5678 VGND.n3017 VGND.n265 0.0760208
R5679 VGND.n2377 VGND.n1016 0.0747188
R5680 VGND.n3439 VGND.n3435 0.0721146
R5681 VGND.n101 VGND.n96 0.0721146
R5682 VGND.n3164 VGND.n210 0.0708554
R5683 VGND.n3458 VGND.n17 0.0708125
R5684 VGND.n3132 VGND.n3131 0.0708125
R5685 VGND.n3331 VGND.n111 0.0708125
R5686 VGND.n2159 VGND.n2156 0.0708125
R5687 VGND.n2288 VGND.n2287 0.0708125
R5688 VGND.n513 VGND.n511 0.0708125
R5689 VGND.n1186 VGND.n1184 0.0708125
R5690 VGND.n2096 VGND.n2044 0.0708125
R5691 VGND.n2880 VGND.n586 0.0708125
R5692 VGND.n2667 VGND.n2664 0.0708125
R5693 VGND.n2731 VGND.n716 0.0708125
R5694 VGND.n2800 VGND.n2795 0.0708125
R5695 VGND.n1330 VGND.n1329 0.0708125
R5696 VGND.n1493 VGND.n1375 0.0708125
R5697 VGND.n767 VGND.n765 0.0708125
R5698 VGND.n1539 VGND.n1537 0.0708125
R5699 VGND.n1652 VGND.n1589 0.0708125
R5700 VGND.n847 VGND.n846 0.0708125
R5701 VGND.n1730 VGND.n1293 0.0708125
R5702 VGND.n1907 VGND.n1906 0.0708125
R5703 VGND.n1756 VGND.n1754 0.0708125
R5704 VGND.n2022 VGND.n1229 0.0708125
R5705 VGND.n2491 VGND.n2400 0.0708125
R5706 VGND.n254 VGND.n252 0.0708125
R5707 VGND.n2313 VGND.n1045 0.0708125
R5708 VGND.n1141 VGND 0.0695104
R5709 VGND.n2767 VGND 0.0695104
R5710 VGND.n2771 VGND.n570 0.0692375
R5711 VGND.n2735 VGND.n722 0.0692375
R5712 VGND.n2703 VGND.n741 0.0692375
R5713 VGND.n2673 VGND.n759 0.0692375
R5714 VGND.n2873 VGND.n669 0.0692375
R5715 VGND.n2870 VGND.n2869 0.0692375
R5716 VGND.n1439 VGND.n1438 0.0685851
R5717 VGND.n2259 VGND.n2258 0.068325
R5718 VGND.n709 VGND.n704 0.068325
R5719 VGND.n2310 VGND.n1047 0.0680676
R5720 VGND.n1047 VGND.n1037 0.0680676
R5721 VGND.n251 VGND.n250 0.0680676
R5722 VGND.n251 VGND.n236 0.0680676
R5723 VGND.n2566 VGND.n928 0.0680676
R5724 VGND.n2566 VGND.n2565 0.0680676
R5725 VGND.n1071 VGND.n1069 0.0680676
R5726 VGND.n1071 VGND.n1070 0.0680676
R5727 VGND.n2575 VGND.n2574 0.0680676
R5728 VGND.n2574 VGND.n851 0.0680676
R5729 VGND.n1089 VGND.n1087 0.0680676
R5730 VGND.n1089 VGND.n1088 0.0680676
R5731 VGND.n2957 VGND.n512 0.0680676
R5732 VGND.n2957 VGND.n2956 0.0680676
R5733 VGND.n2280 VGND.n1121 0.0680676
R5734 VGND.n2282 VGND.n2280 0.0680676
R5735 VGND.n2190 VGND.n1166 0.0680676
R5736 VGND.n2190 VGND.n2189 0.0680676
R5737 VGND.n2158 VGND.n2154 0.0680676
R5738 VGND.n2158 VGND.n2157 0.0680676
R5739 VGND.n541 VGND.n539 0.0680676
R5740 VGND.n541 VGND.n540 0.0680676
R5741 VGND.n1144 VGND.n1135 0.0680676
R5742 VGND.n1144 VGND.n1136 0.0680676
R5743 VGND.n2126 VGND.n1208 0.0680676
R5744 VGND.n1210 VGND.n1208 0.0680676
R5745 VGND.n1189 VGND.n1183 0.0680676
R5746 VGND.n1191 VGND.n1189 0.0680676
R5747 VGND.n632 VGND.n607 0.0680676
R5748 VGND.n632 VGND.n608 0.0680676
R5749 VGND.n2877 VGND.n588 0.0680676
R5750 VGND.n590 VGND.n588 0.0680676
R5751 VGND.n2094 VGND.n2046 0.0680676
R5752 VGND.n2048 VGND.n2046 0.0680676
R5753 VGND.n2907 VGND.n573 0.0680676
R5754 VGND.n2909 VGND.n2907 0.0680676
R5755 VGND.n2697 VGND.n745 0.0680676
R5756 VGND.n2697 VGND.n2696 0.0680676
R5757 VGND.n2666 VGND.n2662 0.0680676
R5758 VGND.n2666 VGND.n2665 0.0680676
R5759 VGND.n2855 VGND.n675 0.0680676
R5760 VGND.n2857 VGND.n2855 0.0680676
R5761 VGND.n2806 VGND.n688 0.0680676
R5762 VGND.n2807 VGND.n2806 0.0680676
R5763 VGND.n729 VGND.n728 0.0680676
R5764 VGND.n728 VGND.n726 0.0680676
R5765 VGND.n707 VGND.n705 0.0680676
R5766 VGND.n707 VGND.n706 0.0680676
R5767 VGND.n1331 VGND.n1317 0.0680676
R5768 VGND.n1332 VGND.n1331 0.0680676
R5769 VGND.n798 VGND.n796 0.0680676
R5770 VGND.n798 VGND.n797 0.0680676
R5771 VGND.n2647 VGND.n766 0.0680676
R5772 VGND.n2647 VGND.n2646 0.0680676
R5773 VGND.n1491 VGND.n1377 0.0680676
R5774 VGND.n1491 VGND.n1490 0.0680676
R5775 VGND.n1523 VGND.n1302 0.0680676
R5776 VGND.n1523 VGND.n1522 0.0680676
R5777 VGND.n1456 VGND.n1404 0.0680676
R5778 VGND.n1456 VGND.n1455 0.0680676
R5779 VGND.n1954 VGND.n1254 0.0680676
R5780 VGND.n1954 VGND.n1953 0.0680676
R5781 VGND.n992 VGND.n987 0.0680676
R5782 VGND.n994 VGND.n992 0.0680676
R5783 VGND.n1621 VGND.n1619 0.0680676
R5784 VGND.n1621 VGND.n1620 0.0680676
R5785 VGND.n1689 VGND.n1563 0.0680676
R5786 VGND.n1564 VGND.n1563 0.0680676
R5787 VGND.n1542 VGND.n1536 0.0680676
R5788 VGND.n1544 VGND.n1542 0.0680676
R5789 VGND.n899 VGND.n867 0.0680676
R5790 VGND.n868 VGND.n867 0.0680676
R5791 VGND.n1650 VGND.n1591 0.0680676
R5792 VGND.n1592 VGND.n1591 0.0680676
R5793 VGND.n2020 VGND.n1231 0.0680676
R5794 VGND.n1986 VGND.n1231 0.0680676
R5795 VGND.n1902 VGND.n1899 0.0680676
R5796 VGND.n1902 VGND.n1901 0.0680676
R5797 VGND.n1731 VGND.n1729 0.0680676
R5798 VGND.n1732 VGND.n1731 0.0680676
R5799 VGND.n2534 VGND.n952 0.0680676
R5800 VGND.n954 VGND.n952 0.0680676
R5801 VGND.n1870 VGND.n1281 0.0680676
R5802 VGND.n1870 VGND.n1869 0.0680676
R5803 VGND.n1800 VGND.n1770 0.0680676
R5804 VGND.n1772 VGND.n1770 0.0680676
R5805 VGND.n1753 VGND.n1751 0.0680676
R5806 VGND.n1753 VGND.n1752 0.0680676
R5807 VGND.n2456 VGND.n2422 0.0680676
R5808 VGND.n2456 VGND.n2455 0.0680676
R5809 VGND.n2488 VGND.n2403 0.0680676
R5810 VGND.n2405 VGND.n2403 0.0680676
R5811 VGND.n1026 VGND.n1021 0.0680676
R5812 VGND.n1026 VGND.n1020 0.0680676
R5813 VGND.n3013 VGND.n3012 0.0680676
R5814 VGND.n3012 VGND.n268 0.0680676
R5815 VGND.n2521 VGND 0.0669062
R5816 VGND.n2200 VGND.n1159 0.0656042
R5817 VGND.n1146 VGND.n1145 0.0656042
R5818 VGND.n538 VGND.n534 0.0656042
R5819 VGND.n1214 VGND.n1213 0.0656042
R5820 VGND.n2913 VGND.n574 0.0656042
R5821 VGND.n631 VGND.n630 0.0656042
R5822 VGND.n2707 VGND.n738 0.0656042
R5823 VGND.n2762 VGND.n708 0.0656042
R5824 VGND.n2865 VGND.n2864 0.0656042
R5825 VGND.n2861 VGND.n2860 0.0656042
R5826 VGND.n1519 VGND.n1518 0.0656042
R5827 VGND.n1457 VGND.n1403 0.0656042
R5828 VGND.n800 VGND.n794 0.0656042
R5829 VGND.n822 VGND.n791 0.0656042
R5830 VGND.n1568 VGND.n1566 0.0656042
R5831 VGND.n1622 VGND.n1615 0.0656042
R5832 VGND.n901 VGND.n865 0.0656042
R5833 VGND.n893 VGND.n872 0.0656042
R5834 VGND.n1283 VGND.n1274 0.0656042
R5835 VGND.n1955 VGND.n1253 0.0656042
R5836 VGND.n2536 VGND.n950 0.0656042
R5837 VGND.n979 VGND.n958 0.0656042
R5838 VGND.n2517 VGND.n988 0.0656042
R5839 VGND.n2451 VGND.n2431 0.0656042
R5840 VGND.n3007 VGND.n270 0.0656042
R5841 VGND.n1090 VGND.n1084 0.0656042
R5842 VGND.n2372 VGND.n2371 0.0656042
R5843 VGND.n2368 VGND.n2367 0.0656042
R5844 VGND.n227 VGND 0.064875
R5845 VGND.n288 VGND 0.064875
R5846 VGND.n287 VGND 0.064875
R5847 VGND.n327 VGND 0.064875
R5848 VGND.n331 VGND 0.064875
R5849 VGND.n374 VGND 0.064875
R5850 VGND.n351 VGND 0.064875
R5851 VGND.n349 VGND 0.064875
R5852 VGND.n3240 VGND 0.064875
R5853 VGND.n3272 VGND 0.064875
R5854 VGND.n3221 VGND 0.064875
R5855 VGND.n3219 VGND 0.064875
R5856 VGND.n200 VGND 0.064875
R5857 VGND.n3200 VGND 0.064875
R5858 VGND.n3384 VGND 0.064875
R5859 VGND.n3274 VGND 0.064875
R5860 VGND.n2161 VGND 0.0643021
R5861 VGND.n2145 VGND 0.0643021
R5862 VGND.n2669 VGND 0.0643021
R5863 VGND.n1322 VGND 0.0643021
R5864 VGND.n1723 VGND 0.0643021
R5865 VGND.n1295 VGND 0.0643021
R5866 VGND VGND.n1910 0.0643021
R5867 VGND.n1748 VGND 0.0643021
R5868 VGND.n248 VGND 0.0643021
R5869 VGND.n3053 VGND.n3052 0.063797
R5870 VGND.n3068 VGND 0.063625
R5871 VGND.n3048 VGND.n233 0.0635047
R5872 VGND.n3066 VGND 0.063
R5873 VGND.n3432 VGND.n41 0.0616979
R5874 VGND.n3163 VGND.n211 0.0616979
R5875 VGND.n3379 VGND.n80 0.0616979
R5876 VGND.n59 VGND 0.0603958
R5877 VGND VGND.n3425 0.0603958
R5878 VGND.n3409 VGND 0.0603958
R5879 VGND.n3410 VGND 0.0603958
R5880 VGND VGND.n3416 0.0603958
R5881 VGND VGND.n36 0.0603958
R5882 VGND.n3443 VGND 0.0603958
R5883 VGND.n45 VGND 0.0603958
R5884 VGND.n5 VGND 0.0603958
R5885 VGND.n13 VGND 0.0603958
R5886 VGND.n14 VGND 0.0603958
R5887 VGND.n3458 VGND 0.0603958
R5888 VGND VGND.n3457 0.0603958
R5889 VGND VGND.n3456 0.0603958
R5890 VGND.n20 VGND 0.0603958
R5891 VGND.n3450 VGND 0.0603958
R5892 VGND VGND.n34 0.0603958
R5893 VGND.n3135 VGND 0.0603958
R5894 VGND.n3086 VGND 0.0603958
R5895 VGND.n3093 VGND 0.0603958
R5896 VGND VGND.n217 0.0603958
R5897 VGND.n3131 VGND 0.0603958
R5898 VGND.n3127 VGND 0.0603958
R5899 VGND VGND.n3126 0.0603958
R5900 VGND VGND.n3119 0.0603958
R5901 VGND VGND.n3102 0.0603958
R5902 VGND VGND.n3112 0.0603958
R5903 VGND.n3159 VGND 0.0603958
R5904 VGND.n3153 VGND 0.0603958
R5905 VGND.n3188 VGND 0.0603958
R5906 VGND VGND.n3187 0.0603958
R5907 VGND.n3181 VGND 0.0603958
R5908 VGND.n194 VGND 0.0603958
R5909 VGND VGND.n3172 0.0603958
R5910 VGND.n82 VGND 0.0603958
R5911 VGND VGND.n3372 0.0603958
R5912 VGND.n87 VGND 0.0603958
R5913 VGND.n88 VGND 0.0603958
R5914 VGND VGND.n3363 0.0603958
R5915 VGND.n3358 VGND 0.0603958
R5916 VGND VGND.n105 0.0603958
R5917 VGND.n3314 VGND 0.0603958
R5918 VGND.n3318 VGND 0.0603958
R5919 VGND.n3326 VGND 0.0603958
R5920 VGND.n3327 VGND 0.0603958
R5921 VGND VGND.n3331 0.0603958
R5922 VGND.n3332 VGND 0.0603958
R5923 VGND.n3333 VGND 0.0603958
R5924 VGND.n3338 VGND 0.0603958
R5925 VGND.n3339 VGND 0.0603958
R5926 VGND.n3351 VGND 0.0603958
R5927 VGND.n2174 VGND 0.0603958
R5928 VGND.n2183 VGND 0.0603958
R5929 VGND VGND.n2221 0.0603958
R5930 VGND VGND.n2220 0.0603958
R5931 VGND VGND.n2279 0.0603958
R5932 VGND VGND.n2234 0.0603958
R5933 VGND.n2231 VGND 0.0603958
R5934 VGND.n2953 VGND.n514 0.0603958
R5935 VGND.n2953 VGND.n2952 0.0603958
R5936 VGND.n559 VGND 0.0603958
R5937 VGND.n2140 VGND 0.0603958
R5938 VGND VGND.n2133 0.0603958
R5939 VGND.n2102 VGND 0.0603958
R5940 VGND.n2088 VGND.n2052 0.0603958
R5941 VGND.n2088 VGND.n2087 0.0603958
R5942 VGND VGND.n2079 0.0603958
R5943 VGND.n2887 VGND 0.0603958
R5944 VGND.n595 VGND.n594 0.0603958
R5945 VGND.n635 VGND 0.0603958
R5946 VGND.n624 VGND 0.0603958
R5947 VGND VGND.n611 0.0603958
R5948 VGND.n616 VGND 0.0603958
R5949 VGND.n2681 VGND 0.0603958
R5950 VGND.n2690 VGND 0.0603958
R5951 VGND.n2727 VGND 0.0603958
R5952 VGND.n2728 VGND 0.0603958
R5953 VGND VGND.n715 0.0603958
R5954 VGND.n2793 VGND 0.0603958
R5955 VGND.n2804 VGND.n689 0.0603958
R5956 VGND.n689 VGND.n685 0.0603958
R5957 VGND VGND.n683 0.0603958
R5958 VGND.n2825 VGND 0.0603958
R5959 VGND.n2833 VGND 0.0603958
R5960 VGND.n1338 VGND 0.0603958
R5961 VGND.n1342 VGND 0.0603958
R5962 VGND.n1350 VGND 0.0603958
R5963 VGND VGND.n1355 0.0603958
R5964 VGND.n1356 VGND 0.0603958
R5965 VGND VGND.n1512 0.0603958
R5966 VGND.n1499 VGND 0.0603958
R5967 VGND VGND.n1498 0.0603958
R5968 VGND VGND.n1386 0.0603958
R5969 VGND VGND.n1486 0.0603958
R5970 VGND VGND.n1411 0.0603958
R5971 VGND.n1414 VGND 0.0603958
R5972 VGND VGND.n1414 0.0603958
R5973 VGND.n1445 VGND 0.0603958
R5974 VGND VGND.n1444 0.0603958
R5975 VGND VGND.n1435 0.0603958
R5976 VGND VGND.n1434 0.0603958
R5977 VGND.n1426 VGND 0.0603958
R5978 VGND.n2643 VGND.n768 0.0603958
R5979 VGND.n2643 VGND.n2642 0.0603958
R5980 VGND.n821 VGND 0.0603958
R5981 VGND.n817 VGND 0.0603958
R5982 VGND VGND.n1712 0.0603958
R5983 VGND VGND.n1697 0.0603958
R5984 VGND.n1668 VGND 0.0603958
R5985 VGND.n1660 VGND 0.0603958
R5986 VGND VGND.n1659 0.0603958
R5987 VGND.n1644 VGND.n1596 0.0603958
R5988 VGND.n1644 VGND.n1643 0.0603958
R5989 VGND.n1640 VGND 0.0603958
R5990 VGND VGND.n1607 0.0603958
R5991 VGND.n1609 VGND 0.0603958
R5992 VGND VGND.n1626 0.0603958
R5993 VGND VGND.n837 0.0603958
R5994 VGND.n2597 VGND 0.0603958
R5995 VGND VGND.n2595 0.0603958
R5996 VGND.n2591 VGND 0.0603958
R5997 VGND.n2585 VGND.n2584 0.0603958
R5998 VGND.n2584 VGND.n850 0.0603958
R5999 VGND VGND.n921 0.0603958
R6000 VGND.n862 VGND 0.0603958
R6001 VGND.n881 VGND 0.0603958
R6002 VGND.n1847 VGND 0.0603958
R6003 VGND.n1849 VGND 0.0603958
R6004 VGND.n1857 VGND 0.0603958
R6005 VGND.n1860 VGND 0.0603958
R6006 VGND VGND.n1880 0.0603958
R6007 VGND.n1881 VGND 0.0603958
R6008 VGND VGND.n1269 0.0603958
R6009 VGND VGND.n1894 0.0603958
R6010 VGND.n1895 VGND 0.0603958
R6011 VGND.n1912 VGND 0.0603958
R6012 VGND VGND.n1911 0.0603958
R6013 VGND.n1981 VGND.n1238 0.0603958
R6014 VGND.n1981 VGND.n1980 0.0603958
R6015 VGND.n1975 VGND 0.0603958
R6016 VGND VGND.n1974 0.0603958
R6017 VGND.n1246 VGND 0.0603958
R6018 VGND VGND.n1965 0.0603958
R6019 VGND VGND.n1942 0.0603958
R6020 VGND VGND.n1932 0.0603958
R6021 VGND.n1929 VGND 0.0603958
R6022 VGND VGND.n1928 0.0603958
R6023 VGND.n929 VGND 0.0603958
R6024 VGND.n2562 VGND.n930 0.0603958
R6025 VGND.n2562 VGND.n2561 0.0603958
R6026 VGND.n935 VGND 0.0603958
R6027 VGND.n2546 VGND 0.0603958
R6028 VGND.n1821 VGND 0.0603958
R6029 VGND VGND.n1820 0.0603958
R6030 VGND.n1815 VGND 0.0603958
R6031 VGND VGND.n1807 0.0603958
R6032 VGND.n1777 VGND 0.0603958
R6033 VGND.n1787 VGND 0.0603958
R6034 VGND.n1785 VGND 0.0603958
R6035 VGND VGND.n1224 0.0603958
R6036 VGND.n2027 VGND 0.0603958
R6037 VGND.n2014 VGND.n1990 0.0603958
R6038 VGND.n2014 VGND.n2013 0.0603958
R6039 VGND.n2010 VGND 0.0603958
R6040 VGND.n2008 VGND 0.0603958
R6041 VGND.n2005 VGND 0.0603958
R6042 VGND VGND.n2004 0.0603958
R6043 VGND VGND.n1997 0.0603958
R6044 VGND VGND.n2511 0.0603958
R6045 VGND.n2502 VGND 0.0603958
R6046 VGND.n2500 VGND 0.0603958
R6047 VGND.n2396 VGND 0.0603958
R6048 VGND.n2496 VGND 0.0603958
R6049 VGND.n2408 VGND.n2407 0.0603958
R6050 VGND.n2409 VGND.n2408 0.0603958
R6051 VGND.n2471 VGND 0.0603958
R6052 VGND.n2469 VGND 0.0603958
R6053 VGND.n2466 VGND 0.0603958
R6054 VGND VGND.n2465 0.0603958
R6055 VGND.n2458 VGND 0.0603958
R6056 VGND.n2450 VGND 0.0603958
R6057 VGND.n2447 VGND 0.0603958
R6058 VGND VGND.n2446 0.0603958
R6059 VGND VGND.n2433 0.0603958
R6060 VGND.n2441 VGND 0.0603958
R6061 VGND VGND.n3033 0.0603958
R6062 VGND VGND.n3018 0.0603958
R6063 VGND.n1058 VGND 0.0603958
R6064 VGND.n1073 VGND 0.0603958
R6065 VGND.n1114 VGND.n1053 0.0603958
R6066 VGND.n1114 VGND.n1113 0.0603958
R6067 VGND.n1040 VGND 0.0603958
R6068 VGND.n1044 VGND 0.0603958
R6069 VGND.n2317 VGND.n2316 0.0603958
R6070 VGND.n2317 VGND.n1036 0.0603958
R6071 VGND.n2333 VGND 0.0603958
R6072 VGND.n2335 VGND 0.0603958
R6073 VGND VGND.n1029 0.0603958
R6074 VGND.n3432 VGND.n3431 0.0590938
R6075 VGND VGND.n3449 0.0590938
R6076 VGND.n3104 VGND 0.0590938
R6077 VGND.n3163 VGND.n3162 0.0590938
R6078 VGND.n3379 VGND.n3378 0.0590938
R6079 VGND.n3355 VGND 0.0590938
R6080 VGND.n2922 VGND.n504 0.0574875
R6081 VGND.n2292 VGND.n1118 0.0574875
R6082 VGND.n2196 VGND.n1163 0.0574875
R6083 VGND.n2166 VGND.n2151 0.0574875
R6084 VGND.n2963 VGND.n509 0.0574875
R6085 VGND.n2927 VGND.n2926 0.0574875
R6086 VGND.n2564 VGND.n926 0.0574697
R6087 VGND.n2573 VGND.n923 0.0574697
R6088 VGND.n2955 VGND.n510 0.0574697
R6089 VGND.n2281 VGND.n1119 0.0574697
R6090 VGND.n1164 VGND.n1161 0.0574697
R6091 VGND.n531 VGND.n529 0.0574697
R6092 VGND.n2255 VGND.n2254 0.0574697
R6093 VGND.n2125 VGND.n1209 0.0574697
R6094 VGND.n1190 VGND.n1181 0.0574697
R6095 VGND.n643 VGND.n642 0.0574697
R6096 VGND.n2876 VGND.n589 0.0574697
R6097 VGND.n2093 VGND.n2047 0.0574697
R6098 VGND.n2908 VGND.n571 0.0574697
R6099 VGND.n743 VGND.n740 0.0574697
R6100 VGND.n2660 VGND.n756 0.0574697
R6101 VGND.n2856 VGND.n673 0.0574697
R6102 VGND.n2808 VGND.n687 0.0574697
R6103 VGND.n724 VGND.n721 0.0574697
R6104 VGND.n703 VGND.n701 0.0574697
R6105 VGND.n789 VGND.n788 0.0574697
R6106 VGND.n2645 VGND.n764 0.0574697
R6107 VGND.n1489 VGND.n1379 0.0574697
R6108 VGND.n1521 VGND.n1300 0.0574697
R6109 VGND.n1454 VGND.n1409 0.0574697
R6110 VGND.n1952 VGND.n1259 0.0574697
R6111 VGND.n993 VGND.n985 0.0574697
R6112 VGND.n1618 VGND.n829 0.0574697
R6113 VGND.n2606 VGND.n831 0.0574697
R6114 VGND.n1688 VGND.n1686 0.0574697
R6115 VGND.n1543 VGND.n1534 0.0574697
R6116 VGND.n898 VGND.n896 0.0574697
R6117 VGND.n1649 VGND.n1647 0.0574697
R6118 VGND.n2019 VGND.n1232 0.0574697
R6119 VGND.n1898 VGND.n1235 0.0574697
R6120 VGND.n1983 VGND.n1236 0.0574697
R6121 VGND.n2533 VGND.n953 0.0574697
R6122 VGND.n1279 VGND.n1276 0.0574697
R6123 VGND.n1799 VGND.n1771 0.0574697
R6124 VGND.n1750 VGND.n1738 0.0574697
R6125 VGND.n1828 VGND.n1739 0.0574697
R6126 VGND.n2454 VGND.n2429 0.0574697
R6127 VGND.n2487 VGND.n2404 0.0574697
R6128 VGND.n232 VGND.n231 0.0574529
R6129 VGND VGND.n3399 0.0557885
R6130 VGND VGND.n3398 0.0557885
R6131 VGND VGND.n3397 0.0557885
R6132 VGND.n126 VGND 0.0557885
R6133 VGND.n128 VGND 0.0557885
R6134 VGND.n133 VGND 0.0557885
R6135 VGND.n138 VGND 0.0557885
R6136 VGND.n143 VGND 0.0557885
R6137 VGND.n148 VGND 0.0557885
R6138 VGND.n153 VGND 0.0557885
R6139 VGND.n158 VGND 0.0557885
R6140 VGND.n163 VGND 0.0557885
R6141 VGND.n168 VGND 0.0557885
R6142 VGND.n3293 VGND 0.0557885
R6143 VGND.n2188 VGND.n1159 0.0551875
R6144 VGND.n1145 VGND.n1143 0.0551875
R6145 VGND.n534 VGND.n527 0.0551875
R6146 VGND.n564 VGND.n563 0.0551875
R6147 VGND.n1213 VGND.n1212 0.0551875
R6148 VGND.n2916 VGND.n574 0.0551875
R6149 VGND.n630 VGND.n605 0.0551875
R6150 VGND.n639 VGND.n638 0.0551875
R6151 VGND.n2695 VGND.n738 0.0551875
R6152 VGND.n2766 VGND.n708 0.0551875
R6153 VGND.n2865 VGND.n676 0.0551875
R6154 VGND.n2860 VGND.n2854 0.0551875
R6155 VGND.n1458 VGND.n1457 0.0551875
R6156 VGND.n794 VGND.n786 0.0551875
R6157 VGND.n822 VGND.n821 0.0551875
R6158 VGND.n1569 VGND.n1568 0.0551875
R6159 VGND.n1623 VGND.n1622 0.0551875
R6160 VGND.n902 VGND.n901 0.0551875
R6161 VGND.n893 VGND.n892 0.0551875
R6162 VGND.n1868 VGND.n1283 0.0551875
R6163 VGND.n1956 VGND.n1955 0.0551875
R6164 VGND.n2537 VGND.n2536 0.0551875
R6165 VGND.n979 VGND.n978 0.0551875
R6166 VGND.n2520 VGND.n988 0.0551875
R6167 VGND.n2451 VGND.n2450 0.0551875
R6168 VGND.n3010 VGND.n270 0.0551875
R6169 VGND.n1091 VGND.n1090 0.0551875
R6170 VGND.n2372 VGND.n1025 0.0551875
R6171 VGND.n2367 VGND.n2366 0.0551875
R6172 VGND.n3381 VGND 0.0527529
R6173 VGND VGND.n1250 0.0525833
R6174 VGND.n1802 VGND 0.0525833
R6175 VGND.n3381 VGND.n3380 0.0519696
R6176 VGND.n3295 VGND 0.0518289
R6177 VGND.n17 VGND.n14 0.0499792
R6178 VGND.n3132 VGND.n217 0.0499792
R6179 VGND.n3327 VGND.n111 0.0499792
R6180 VGND.n2160 VGND.n2159 0.0499792
R6181 VGND.n2230 VGND.n511 0.0499792
R6182 VGND.n2144 VGND.n1184 0.0499792
R6183 VGND.n586 VGND.n584 0.0499792
R6184 VGND.n2668 VGND.n2667 0.0499792
R6185 VGND.n1330 VGND.n1318 0.0499792
R6186 VGND.n1427 VGND.n765 0.0499792
R6187 VGND.n1722 VGND.n1537 0.0499792
R6188 VGND.n1653 VGND.n1652 0.0499792
R6189 VGND.n2589 VGND.n846 0.0499792
R6190 VGND.n1730 VGND.n1294 0.0499792
R6191 VGND.n1907 VGND.n1897 0.0499792
R6192 VGND.n1754 VGND.n1742 0.0499792
R6193 VGND.n2023 VGND.n2022 0.0499792
R6194 VGND.n2400 VGND.n2398 0.0499792
R6195 VGND.n252 VGND.n241 0.0499792
R6196 VGND.n1045 VGND.n1044 0.0499792
R6197 VGND.n3442 VGND.n3435 0.0486771
R6198 VGND.n3171 VGND.n3166 0.0486771
R6199 VGND.n104 VGND.n96 0.0486771
R6200 VGND.n2155 VGND 0.047375
R6201 VGND.n1192 VGND 0.047375
R6202 VGND.n2663 VGND 0.047375
R6203 VGND.n1319 VGND 0.047375
R6204 VGND.n1545 VGND 0.047375
R6205 VGND.n1733 VGND 0.047375
R6206 VGND.n1755 VGND 0.047375
R6207 VGND.n253 VGND 0.047375
R6208 VGND.n3466 VGND 0.0460729
R6209 VGND VGND.n3134 0.0460729
R6210 VGND VGND.n3298 0.0460729
R6211 VGND.n2183 VGND.n1165 0.0447708
R6212 VGND.n2133 VGND.n1203 0.0447708
R6213 VGND.n2690 VGND.n744 0.0447708
R6214 VGND.n1357 VGND.n1301 0.0447708
R6215 VGND.n1696 VGND.n1557 0.0447708
R6216 VGND.n1862 VGND.n1280 0.0447708
R6217 VGND.n1806 VGND.n1766 0.0447708
R6218 VGND.n3018 VGND.n3017 0.0447708
R6219 VGND.n3470 VGND.n3469 0.0423452
R6220 VGND.n3471 VGND.n3470 0.0423452
R6221 VGND.n3472 VGND.n3471 0.0423452
R6222 VGND.n3473 VGND.n3472 0.0423452
R6223 VGND.n3474 VGND.n3473 0.0423452
R6224 VGND.n3475 VGND.n3474 0.0423452
R6225 VGND.n3476 VGND.n3475 0.0423452
R6226 VGND.n3477 VGND.n3476 0.0423452
R6227 VGND.n3478 VGND.n3477 0.0423452
R6228 VGND.n3479 VGND.n3478 0.0423452
R6229 VGND.n3480 VGND.n3479 0.0423452
R6230 VGND.n3481 VGND.n3480 0.0423452
R6231 VGND.n3482 VGND.n3481 0.0423452
R6232 VGND.n3483 VGND.n3482 0.0423452
R6233 VGND.n3484 VGND.n3483 0.0423452
R6234 VGND.n3485 VGND.n3484 0.0423452
R6235 VGND.n3486 VGND.n3485 0.0423452
R6236 VGND.n3487 VGND.n3486 0.0423452
R6237 VGND.n3488 VGND.n3487 0.0423452
R6238 VGND.n3489 VGND.n3488 0.0423452
R6239 VGND.n3490 VGND.n3489 0.0423452
R6240 VGND.n3491 VGND.n3490 0.0423452
R6241 VGND.n871 VGND 0.0421667
R6242 VGND.n957 VGND 0.0421667
R6243 VGND.n2516 VGND 0.0421667
R6244 VGND.n2513 VGND 0.0421667
R6245 VGND.n3051 VGND.n230 0.0416941
R6246 VGND.n2385 VGND.n2383 0.0414836
R6247 VGND.n2311 VGND.n2310 0.0410405
R6248 VGND.n2318 VGND.n1037 0.0410405
R6249 VGND.n250 VGND.n249 0.0410405
R6250 VGND.n238 VGND.n236 0.0410405
R6251 VGND.n2569 VGND.n928 0.0410405
R6252 VGND.n2565 VGND.n2563 0.0410405
R6253 VGND.n1069 VGND.n1067 0.0410405
R6254 VGND.n1070 VGND.n1052 0.0410405
R6255 VGND.n2577 VGND.n2575 0.0410405
R6256 VGND.n2583 VGND.n851 0.0410405
R6257 VGND.n1087 VGND.n1086 0.0410405
R6258 VGND.n1088 VGND.n501 0.0410405
R6259 VGND.n2960 VGND.n512 0.0410405
R6260 VGND.n2956 VGND.n2954 0.0410405
R6261 VGND.n2289 VGND.n1121 0.0410405
R6262 VGND.n2283 VGND.n2282 0.0410405
R6263 VGND.n2193 VGND.n1166 0.0410405
R6264 VGND.n2189 VGND.n1160 0.0410405
R6265 VGND.n2162 VGND.n2154 0.0410405
R6266 VGND.n2157 VGND.n1176 0.0410405
R6267 VGND.n539 VGND.n528 0.0410405
R6268 VGND.n540 VGND.n532 0.0410405
R6269 VGND.n1135 VGND.n1134 0.0410405
R6270 VGND.n1137 VGND.n1136 0.0410405
R6271 VGND.n2127 VGND.n2126 0.0410405
R6272 VGND.n1211 VGND.n1210 0.0410405
R6273 VGND.n2146 VGND.n1183 0.0410405
R6274 VGND.n1193 VGND.n1191 0.0410405
R6275 VGND.n607 VGND.n606 0.0410405
R6276 VGND.n609 VGND.n608 0.0410405
R6277 VGND.n2878 VGND.n2877 0.0410405
R6278 VGND.n591 VGND.n590 0.0410405
R6279 VGND.n2095 VGND.n2094 0.0410405
R6280 VGND.n2049 VGND.n2048 0.0410405
R6281 VGND.n2918 VGND.n573 0.0410405
R6282 VGND.n2911 VGND.n2909 0.0410405
R6283 VGND.n2700 VGND.n745 0.0410405
R6284 VGND.n2696 VGND.n739 0.0410405
R6285 VGND.n2670 VGND.n2662 0.0410405
R6286 VGND.n2665 VGND.n755 0.0410405
R6287 VGND.n2866 VGND.n675 0.0410405
R6288 VGND.n2858 VGND.n2857 0.0410405
R6289 VGND.n2798 VGND.n688 0.0410405
R6290 VGND.n2807 VGND.n686 0.0410405
R6291 VGND.n2732 VGND.n729 0.0410405
R6292 VGND.n726 VGND.n720 0.0410405
R6293 VGND.n2768 VGND.n705 0.0410405
R6294 VGND.n706 VGND.n700 0.0410405
R6295 VGND.n1323 VGND.n1317 0.0410405
R6296 VGND.n1332 VGND.n1315 0.0410405
R6297 VGND.n796 VGND.n787 0.0410405
R6298 VGND.n797 VGND.n790 0.0410405
R6299 VGND.n2650 VGND.n766 0.0410405
R6300 VGND.n2646 VGND.n2644 0.0410405
R6301 VGND.n1382 VGND.n1377 0.0410405
R6302 VGND.n1490 VGND.n1378 0.0410405
R6303 VGND.n1526 VGND.n1302 0.0410405
R6304 VGND.n1522 VGND.n1520 0.0410405
R6305 VGND.n1406 VGND.n1404 0.0410405
R6306 VGND.n1455 VGND.n1405 0.0410405
R6307 VGND.n1256 VGND.n1254 0.0410405
R6308 VGND.n1953 VGND.n1255 0.0410405
R6309 VGND.n2522 VGND.n987 0.0410405
R6310 VGND.n2515 VGND.n994 0.0410405
R6311 VGND.n1619 VGND.n1617 0.0410405
R6312 VGND.n1620 VGND.n832 0.0410405
R6313 VGND.n1690 VGND.n1689 0.0410405
R6314 VGND.n1565 VGND.n1564 0.0410405
R6315 VGND.n1724 VGND.n1536 0.0410405
R6316 VGND.n1546 VGND.n1544 0.0410405
R6317 VGND.n900 VGND.n899 0.0410405
R6318 VGND.n869 VGND.n868 0.0410405
R6319 VGND.n1651 VGND.n1650 0.0410405
R6320 VGND.n1593 VGND.n1592 0.0410405
R6321 VGND.n2021 VGND.n2020 0.0410405
R6322 VGND.n1987 VGND.n1986 0.0410405
R6323 VGND.n1908 VGND.n1899 0.0410405
R6324 VGND.n1901 VGND.n1237 0.0410405
R6325 VGND.n1729 VGND.n1296 0.0410405
R6326 VGND.n1734 VGND.n1732 0.0410405
R6327 VGND.n2535 VGND.n2534 0.0410405
R6328 VGND.n955 VGND.n954 0.0410405
R6329 VGND.n1873 VGND.n1281 0.0410405
R6330 VGND.n1869 VGND.n1275 0.0410405
R6331 VGND.n1801 VGND.n1800 0.0410405
R6332 VGND.n1773 VGND.n1772 0.0410405
R6333 VGND.n1751 VGND.n1749 0.0410405
R6334 VGND.n1752 VGND.n1740 0.0410405
R6335 VGND.n2426 VGND.n2422 0.0410405
R6336 VGND.n2455 VGND.n2423 0.0410405
R6337 VGND.n2489 VGND.n2488 0.0410405
R6338 VGND.n2406 VGND.n2405 0.0410405
R6339 VGND.n2373 VGND.n1021 0.0410405
R6340 VGND.n2346 VGND.n1020 0.0410405
R6341 VGND.n3013 VGND.n266 0.0410405
R6342 VGND.n3002 VGND.n268 0.0410405
R6343 VGND.n2301 VGND.n2299 0.0393869
R6344 VGND.n594 VGND 0.0382604
R6345 VGND.n2169 VGND 0.0369583
R6346 VGND.n1195 VGND 0.0369583
R6347 VGND.n592 VGND 0.0369583
R6348 VGND.n2676 VGND 0.0369583
R6349 VGND.n2805 VGND 0.0369583
R6350 VGND.n1336 VGND 0.0369583
R6351 VGND.n1548 VGND 0.0369583
R6352 VGND.n922 VGND 0.0369583
R6353 VGND VGND.n1291 0.0369583
R6354 VGND VGND.n932 0.0369583
R6355 VGND.n1826 VGND 0.0369583
R6356 VGND.n3042 VGND 0.0369583
R6357 VGND.n2378 VGND.n2377 0.0352656
R6358 VGND.n827 VGND.n702 0.0351625
R6359 VGND.n1385 VGND.n723 0.0351625
R6360 VGND.n1529 VGND.n742 0.0351625
R6361 VGND.n2659 VGND.n760 0.0351625
R6362 VGND.n2654 VGND.n2653 0.0351625
R6363 VGND.n2613 VGND.n672 0.0351625
R6364 VGND.n210 VGND 0.0346243
R6365 VGND.n3465 VGND 0.0343542
R6366 VGND VGND.n216 0.0343542
R6367 VGND VGND.n3317 0.0343542
R6368 VGND.n2161 VGND.n2160 0.0343542
R6369 VGND.n2218 VGND.n1120 0.0343542
R6370 VGND.n2145 VGND.n2144 0.0343542
R6371 VGND.n2097 VGND.n2041 0.0343542
R6372 VGND.n2669 VGND.n2668 0.0343542
R6373 VGND.n2730 VGND.n725 0.0343542
R6374 VGND.n1322 VGND.n1318 0.0343542
R6375 VGND.n1338 VGND 0.0343542
R6376 VGND.n1381 VGND.n1371 0.0343542
R6377 VGND.n1723 VGND.n1722 0.0343542
R6378 VGND.n1718 VGND 0.0343542
R6379 VGND.n1653 VGND.n1588 0.0343542
R6380 VGND.n1295 VGND.n1294 0.0343542
R6381 VGND.n1841 VGND 0.0343542
R6382 VGND.n1910 VGND.n1897 0.0343542
R6383 VGND.n1973 VGND 0.0343542
R6384 VGND.n1929 VGND 0.0343542
R6385 VGND.n1748 VGND.n1742 0.0343542
R6386 VGND.n2023 VGND.n1226 0.0343542
R6387 VGND.n248 VGND.n241 0.0343542
R6388 VGND.n1065 VGND.n1064 0.0343542
R6389 VGND.n1041 VGND 0.0343542
R6390 VGND.n2526 VGND.n830 0.0339875
R6391 VGND.n1985 VGND.n1984 0.0339875
R6392 VGND.n1876 VGND.n1278 0.0339875
R6393 VGND.n1832 VGND.n1831 0.0339875
R6394 VGND.n2572 VGND.n925 0.0339875
R6395 VGND.n2531 VGND.n2530 0.0339875
R6396 VGND VGND.n3409 0.0330521
R6397 VGND VGND.n13 0.0330521
R6398 VGND.n3093 VGND 0.0330521
R6399 VGND.n3188 VGND 0.0330521
R6400 VGND VGND.n87 0.0330521
R6401 VGND VGND.n3326 0.0330521
R6402 VGND.n2222 VGND 0.0330521
R6403 VGND.n2235 VGND 0.0330521
R6404 VGND VGND.n2040 0.0330521
R6405 VGND VGND.n583 0.0330521
R6406 VGND.n2724 VGND 0.0330521
R6407 VGND.n2789 VGND 0.0330521
R6408 VGND.n1519 VGND 0.0330521
R6409 VGND.n1499 VGND 0.0330521
R6410 VGND.n1435 VGND 0.0330521
R6411 VGND.n1660 VGND 0.0330521
R6412 VGND VGND.n1895 0.0330521
R6413 VGND.n1932 VGND 0.0330521
R6414 VGND VGND.n1224 0.0330521
R6415 VGND VGND.n2396 0.0330521
R6416 VGND.n2425 VGND 0.0330521
R6417 VGND VGND.n279 0.0330521
R6418 VGND VGND.n494 0.0330521
R6419 VGND VGND.n37 0.03175
R6420 VGND.n3173 VGND 0.03175
R6421 VGND.n106 VGND 0.03175
R6422 VGND.n2221 VGND 0.03175
R6423 VGND.n563 VGND 0.03175
R6424 VGND VGND.n2727 0.03175
R6425 VGND.n2833 VGND 0.03175
R6426 VGND VGND.n674 0.03175
R6427 VGND VGND.n1337 0.03175
R6428 VGND.n1445 VGND 0.03175
R6429 VGND.n1434 VGND 0.03175
R6430 VGND.n1912 VGND 0.03175
R6431 VGND.n1252 VGND 0.03175
R6432 VGND.n949 VGND 0.03175
R6433 VGND.n1774 VGND 0.03175
R6434 VGND VGND.n1775 0.03175
R6435 VGND.n2005 VGND 0.03175
R6436 VGND.n2512 VGND 0.03175
R6437 VGND.n2466 VGND 0.03175
R6438 VGND.n2447 VGND 0.03175
R6439 VGND.n2381 VGND.n1018 0.0308279
R6440 VGND.n3399 VGND 0.0305481
R6441 VGND.n3398 VGND 0.0305481
R6442 VGND.n3397 VGND 0.0305481
R6443 VGND VGND.n126 0.0305481
R6444 VGND VGND.n3293 0.0305481
R6445 VGND.n2524 VGND.n985 0.0292489
R6446 VGND.n993 VGND.n984 0.0292489
R6447 VGND.n1259 VGND.n1258 0.0292489
R6448 VGND.n1952 VGND.n1951 0.0292489
R6449 VGND.n1409 VGND.n1408 0.0292489
R6450 VGND.n1454 VGND.n1453 0.0292489
R6451 VGND.n2770 VGND.n703 0.0292489
R6452 VGND.n2772 VGND.n701 0.0292489
R6453 VGND.n2920 VGND.n571 0.0292489
R6454 VGND.n2908 VGND.n569 0.0292489
R6455 VGND.n2256 VGND.n2255 0.0292489
R6456 VGND.n2254 VGND.n2253 0.0292489
R6457 VGND.n831 VGND.n828 0.0292489
R6458 VGND.n1618 VGND.n828 0.0292489
R6459 VGND.n2019 VGND.n2018 0.0292489
R6460 VGND.n2016 VGND.n1232 0.0292489
R6461 VGND.n1649 VGND.n1648 0.0292489
R6462 VGND.n1647 VGND.n1646 0.0292489
R6463 VGND.n1384 VGND.n1379 0.0292489
R6464 VGND.n1489 VGND.n1488 0.0292489
R6465 VGND.n2734 VGND.n724 0.0292489
R6466 VGND.n2736 VGND.n721 0.0292489
R6467 VGND.n2093 VGND.n2092 0.0292489
R6468 VGND.n2090 VGND.n2047 0.0292489
R6469 VGND.n2291 VGND.n1119 0.0292489
R6470 VGND.n2281 VGND.n1117 0.0292489
R6471 VGND.n1236 VGND.n1234 0.0292489
R6472 VGND.n1898 VGND.n1234 0.0292489
R6473 VGND.n1799 VGND.n1798 0.0292489
R6474 VGND.n1796 VGND.n1771 0.0292489
R6475 VGND.n1875 VGND.n1279 0.0292489
R6476 VGND.n1877 VGND.n1276 0.0292489
R6477 VGND.n1688 VGND.n1687 0.0292489
R6478 VGND.n1686 VGND.n1685 0.0292489
R6479 VGND.n1528 VGND.n1300 0.0292489
R6480 VGND.n1521 VGND.n1299 0.0292489
R6481 VGND.n2702 VGND.n743 0.0292489
R6482 VGND.n2704 VGND.n740 0.0292489
R6483 VGND.n2125 VGND.n2124 0.0292489
R6484 VGND.n2122 VGND.n1209 0.0292489
R6485 VGND.n2195 VGND.n1164 0.0292489
R6486 VGND.n2197 VGND.n1161 0.0292489
R6487 VGND.n1726 VGND.n1534 0.0292489
R6488 VGND.n1543 VGND.n1533 0.0292489
R6489 VGND.n2672 VGND.n2660 0.0292489
R6490 VGND.n2674 VGND.n756 0.0292489
R6491 VGND.n2148 VGND.n1181 0.0292489
R6492 VGND.n1190 VGND.n1180 0.0292489
R6493 VGND.n1739 VGND.n1737 0.0292489
R6494 VGND.n1750 VGND.n1737 0.0292489
R6495 VGND.n2487 VGND.n2486 0.0292489
R6496 VGND.n2484 VGND.n2404 0.0292489
R6497 VGND.n2571 VGND.n926 0.0292489
R6498 VGND.n2564 VGND.n924 0.0292489
R6499 VGND.n2579 VGND.n2573 0.0292489
R6500 VGND.n2581 VGND.n923 0.0292489
R6501 VGND.n2652 VGND.n764 0.0292489
R6502 VGND.n2645 VGND.n762 0.0292489
R6503 VGND.n2796 VGND.n687 0.0292489
R6504 VGND.n2809 VGND.n2808 0.0292489
R6505 VGND.n2876 VGND.n2875 0.0292489
R6506 VGND.n668 VGND.n589 0.0292489
R6507 VGND.n2962 VGND.n510 0.0292489
R6508 VGND.n2955 VGND.n508 0.0292489
R6509 VGND.n2429 VGND.n2428 0.0292489
R6510 VGND.n2454 VGND.n2453 0.0292489
R6511 VGND.n2533 VGND.n2532 0.0292489
R6512 VGND.n981 VGND.n953 0.0292489
R6513 VGND.n898 VGND.n897 0.0292489
R6514 VGND.n896 VGND.n895 0.0292489
R6515 VGND.n2614 VGND.n788 0.0292489
R6516 VGND.n824 VGND.n789 0.0292489
R6517 VGND.n2868 VGND.n673 0.0292489
R6518 VGND.n2856 VGND.n671 0.0292489
R6519 VGND.n644 VGND.n643 0.0292489
R6520 VGND.n642 VGND.n641 0.0292489
R6521 VGND.n2928 VGND.n529 0.0292489
R6522 VGND.n566 VGND.n531 0.0292489
R6523 VGND.n2191 VGND.n2188 0.0291458
R6524 VGND.n1143 VGND.n1141 0.0291458
R6525 VGND.n2930 VGND.n527 0.0291458
R6526 VGND.n1212 VGND.n1206 0.0291458
R6527 VGND.n2917 VGND.n2916 0.0291458
R6528 VGND.n646 VGND.n605 0.0291458
R6529 VGND.n2698 VGND.n2695 0.0291458
R6530 VGND.n2767 VGND.n2766 0.0291458
R6531 VGND.n676 VGND.n674 0.0291458
R6532 VGND.n1524 VGND.n1304 0.0291458
R6533 VGND.n1458 VGND.n1402 0.0291458
R6534 VGND.n2616 VGND.n786 0.0291458
R6535 VGND.n1569 VGND.n1561 0.0291458
R6536 VGND.n1623 VGND.n1614 0.0291458
R6537 VGND.n902 VGND.n864 0.0291458
R6538 VGND.n1871 VGND.n1868 0.0291458
R6539 VGND.n1956 VGND.n1252 0.0291458
R6540 VGND.n2537 VGND.n949 0.0291458
R6541 VGND.n1775 VGND.n1774 0.0291458
R6542 VGND.n2521 VGND.n2520 0.0291458
R6543 VGND.n2424 VGND.n2418 0.0291458
R6544 VGND.n3011 VGND.n3010 0.0291458
R6545 VGND.n1091 VGND.n1083 0.0291458
R6546 VGND.n1025 VGND.n1024 0.0291458
R6547 VGND.n2288 VGND 0.0278438
R6548 VGND VGND.n2096 0.0278438
R6549 VGND.n2731 VGND 0.0278438
R6550 VGND.n1375 VGND 0.0278438
R6551 VGND VGND.n927 0.0278438
R6552 VGND.n1066 VGND 0.0278438
R6553 VGND.n1381 VGND 0.0265417
R6554 VGND.n1825 VGND 0.0252396
R6555 VGND.n1807 VGND 0.0252396
R6556 VGND.n1787 VGND 0.0252396
R6557 VGND.n2010 VGND 0.0252396
R6558 VGND.n2502 VGND 0.0252396
R6559 VGND.n2471 VGND 0.0252396
R6560 VGND.n2446 VGND 0.0252396
R6561 VGND VGND.n2333 0.0252396
R6562 VGND.n2376 VGND.n2375 0.024993
R6563 VGND.n2285 VGND.n1126 0.0239375
R6564 VGND.n2958 VGND.n514 0.0239375
R6565 VGND.n2952 VGND.n516 0.0239375
R6566 VGND.n2052 VGND.n2051 0.0239375
R6567 VGND.n593 VGND.n592 0.0239375
R6568 VGND.n666 VGND.n595 0.0239375
R6569 VGND.n2738 VGND.n719 0.0239375
R6570 VGND.n2805 VGND.n2804 0.0239375
R6571 VGND.n2811 VGND.n685 0.0239375
R6572 VGND.n1337 VGND.n1336 0.0239375
R6573 VGND.n1386 VGND.n1376 0.0239375
R6574 VGND.n2648 VGND.n768 0.0239375
R6575 VGND.n2642 VGND.n770 0.0239375
R6576 VGND.n1719 VGND.n1548 0.0239375
R6577 VGND.n1596 VGND.n1595 0.0239375
R6578 VGND.n1640 VGND 0.0239375
R6579 VGND.n2585 VGND.n849 0.0239375
R6580 VGND.n922 VGND.n850 0.0239375
R6581 VGND.n881 VGND 0.0239375
R6582 VGND.n1840 VGND.n1291 0.0239375
R6583 VGND VGND.n1860 0.0239375
R6584 VGND.n1900 VGND.n1238 0.0239375
R6585 VGND.n2567 VGND.n930 0.0239375
R6586 VGND.n2561 VGND.n932 0.0239375
R6587 VGND.n1826 VGND.n1825 0.0239375
R6588 VGND.n1776 VGND 0.0239375
R6589 VGND.n1990 VGND.n1989 0.0239375
R6590 VGND.n2407 VGND.n2401 0.0239375
R6591 VGND.n2482 VGND.n2409 0.0239375
R6592 VGND.n3042 VGND.n3041 0.0239375
R6593 VGND.n1056 VGND.n1053 0.0239375
R6594 VGND.n2316 VGND.n1038 0.0239375
R6595 VGND.n2320 VGND.n1036 0.0239375
R6596 VGND.n2968 VGND.n2967 0.0234125
R6597 VGND.n2294 VGND.n2293 0.0234125
R6598 VGND.n1162 VGND.n267 0.0234125
R6599 VGND.n1179 VGND.n237 0.0234125
R6600 VGND.n2964 VGND.n507 0.0234125
R6601 VGND.n1023 VGND.n530 0.0234125
R6602 VGND.n3431 VGND 0.0226354
R6603 VGND.n3426 VGND 0.0226354
R6604 VGND VGND.n62 0.0226354
R6605 VGND.n3417 VGND 0.0226354
R6606 VGND.n3412 VGND 0.0226354
R6607 VGND.n3438 VGND 0.0226354
R6608 VGND.n5 VGND 0.0226354
R6609 VGND VGND.n12 0.0226354
R6610 VGND.n3457 VGND 0.0226354
R6611 VGND VGND.n19 0.0226354
R6612 VGND.n35 VGND 0.0226354
R6613 VGND.n27 VGND 0.0226354
R6614 VGND.n3086 VGND 0.0226354
R6615 VGND VGND.n3092 0.0226354
R6616 VGND.n3127 VGND 0.0226354
R6617 VGND.n3120 VGND 0.0226354
R6618 VGND.n3113 VGND 0.0226354
R6619 VGND.n3162 VGND 0.0226354
R6620 VGND VGND.n3147 0.0226354
R6621 VGND.n3149 VGND 0.0226354
R6622 VGND VGND.n190 0.0226354
R6623 VGND VGND.n193 0.0226354
R6624 VGND.n3378 VGND 0.0226354
R6625 VGND.n3373 VGND 0.0226354
R6626 VGND VGND.n85 0.0226354
R6627 VGND.n3364 VGND 0.0226354
R6628 VGND VGND.n91 0.0226354
R6629 VGND.n100 VGND 0.0226354
R6630 VGND.n3318 VGND 0.0226354
R6631 VGND VGND.n3325 0.0226354
R6632 VGND VGND.n3332 0.0226354
R6633 VGND VGND.n3337 0.0226354
R6634 VGND.n3354 VGND 0.0226354
R6635 VGND.n3344 VGND 0.0226354
R6636 VGND VGND.n2216 0.0226354
R6637 VGND.n2218 VGND 0.0226354
R6638 VGND.n2285 VGND 0.0226354
R6639 VGND VGND.n1131 0.0226354
R6640 VGND.n2238 VGND 0.0226354
R6641 VGND.n2234 VGND 0.0226354
R6642 VGND.n2940 VGND 0.0226354
R6643 VGND.n544 VGND 0.0226354
R6644 VGND.n552 VGND 0.0226354
R6645 VGND.n2107 VGND 0.0226354
R6646 VGND.n2097 VGND 0.0226354
R6647 VGND.n2080 VGND 0.0226354
R6648 VGND VGND.n2062 0.0226354
R6649 VGND.n2905 VGND 0.0226354
R6650 VGND VGND.n580 0.0226354
R6651 VGND VGND.n593 0.0226354
R6652 VGND.n638 VGND 0.0226354
R6653 VGND.n616 VGND 0.0226354
R6654 VGND VGND.n2723 0.0226354
R6655 VGND VGND.n2730 0.0226354
R6656 VGND.n2738 VGND 0.0226354
R6657 VGND.n2757 VGND 0.0226354
R6658 VGND VGND.n2788 0.0226354
R6659 VGND VGND.n2793 0.0226354
R6660 VGND.n2826 VGND 0.0226354
R6661 VGND VGND.n2832 0.0226354
R6662 VGND.n2847 VGND 0.0226354
R6663 VGND VGND.n1349 0.0226354
R6664 VGND.n1350 VGND 0.0226354
R6665 VGND VGND.n1304 0.0226354
R6666 VGND.n1513 VGND 0.0226354
R6667 VGND VGND.n1367 0.0226354
R6668 VGND.n1497 VGND 0.0226354
R6669 VGND VGND.n1371 0.0226354
R6670 VGND.n1486 VGND 0.0226354
R6671 VGND.n1436 VGND 0.0226354
R6672 VGND VGND.n1426 0.0226354
R6673 VGND VGND.n778 0.0226354
R6674 VGND.n810 VGND 0.0226354
R6675 VGND.n1698 VGND 0.0226354
R6676 VGND VGND.n1576 0.0226354
R6677 VGND VGND.n1579 0.0226354
R6678 VGND.n1643 VGND 0.0226354
R6679 VGND VGND.n1609 0.0226354
R6680 VGND.n1627 VGND 0.0226354
R6681 VGND.n2595 VGND 0.0226354
R6682 VGND.n906 VGND 0.0226354
R6683 VGND VGND.n873 0.0226354
R6684 VGND VGND.n1847 0.0226354
R6685 VGND VGND.n1848 0.0226354
R6686 VGND.n1881 VGND 0.0226354
R6687 VGND.n1886 VGND 0.0226354
R6688 VGND.n1911 VGND 0.0226354
R6689 VGND.n1966 VGND 0.0226354
R6690 VGND.n1965 VGND 0.0226354
R6691 VGND.n1943 VGND 0.0226354
R6692 VGND.n1933 VGND 0.0226354
R6693 VGND.n1928 VGND 0.0226354
R6694 VGND.n1923 VGND 0.0226354
R6695 VGND VGND.n941 0.0226354
R6696 VGND VGND.n945 0.0226354
R6697 VGND VGND.n965 0.0226354
R6698 VGND.n1808 VGND 0.0226354
R6699 VGND.n2013 VGND 0.0226354
R6700 VGND.n2505 VGND 0.0226354
R6701 VGND VGND.n2410 0.0226354
R6702 VGND VGND.n2418 0.0226354
R6703 VGND.n2436 VGND 0.0226354
R6704 VGND.n3034 VGND 0.0226354
R6705 VGND.n3019 VGND 0.0226354
R6706 VGND.n2990 VGND 0.0226354
R6707 VGND VGND.n1065 0.0226354
R6708 VGND.n2983 VGND 0.0226354
R6709 VGND.n2330 VGND 0.0226354
R6710 VGND.n2360 VGND 0.0226354
R6711 VGND.n2352 VGND 0.0226354
R6712 VGND.n3294 VGND 0.0219286
R6713 VGND.n2303 VGND.n2302 0.0218125
R6714 VGND.n2812 VGND 0.0213333
R6715 VGND.n2597 VGND 0.0213333
R6716 VGND VGND.n128 0.0209327
R6717 VGND.n130 VGND 0.0209327
R6718 VGND VGND.n133 0.0209327
R6719 VGND.n135 VGND 0.0209327
R6720 VGND VGND.n138 0.0209327
R6721 VGND.n140 VGND 0.0209327
R6722 VGND VGND.n143 0.0209327
R6723 VGND.n145 VGND 0.0209327
R6724 VGND VGND.n148 0.0209327
R6725 VGND.n150 VGND 0.0209327
R6726 VGND VGND.n153 0.0209327
R6727 VGND.n155 VGND 0.0209327
R6728 VGND VGND.n158 0.0209327
R6729 VGND.n160 VGND 0.0209327
R6730 VGND VGND.n163 0.0209327
R6731 VGND.n165 VGND 0.0209327
R6732 VGND VGND.n168 0.0209327
R6733 VGND.n170 VGND 0.0209327
R6734 VGND VGND.n2153 0.0200312
R6735 VGND VGND.n1182 0.0200312
R6736 VGND VGND.n2661 0.0200312
R6737 VGND.n1327 VGND 0.0200312
R6738 VGND VGND.n1535 0.0200312
R6739 VGND.n1836 VGND 0.0200312
R6740 VGND VGND.n1747 0.0200312
R6741 VGND VGND.n1761 0.0200312
R6742 VGND VGND.n247 0.0200312
R6743 VGND.n2200 VGND.n2199 0.0187292
R6744 VGND.n1146 VGND.n1138 0.0187292
R6745 VGND.n2251 VGND.n2250 0.0187292
R6746 VGND.n542 VGND.n538 0.0187292
R6747 VGND.n544 VGND.n543 0.0187292
R6748 VGND.n2120 VGND.n1214 0.0187292
R6749 VGND.n2913 VGND.n2912 0.0187292
R6750 VGND.n2906 VGND.n2905 0.0187292
R6751 VGND.n633 VGND.n631 0.0187292
R6752 VGND.n635 VGND.n634 0.0187292
R6753 VGND.n2707 VGND.n2706 0.0187292
R6754 VGND.n2762 VGND.n699 0.0187292
R6755 VGND.n2775 VGND.n2774 0.0187292
R6756 VGND.n2864 VGND.n677 0.0187292
R6757 VGND.n2861 VGND.n2838 0.0187292
R6758 VGND.n1518 VGND.n1306 0.0187292
R6759 VGND.n1410 VGND.n1403 0.0187292
R6760 VGND.n1451 VGND.n1450 0.0187292
R6761 VGND.n800 VGND.n799 0.0187292
R6762 VGND.n795 VGND.n791 0.0187292
R6763 VGND.n1683 VGND.n1566 0.0187292
R6764 VGND.n1615 VGND.n833 0.0187292
R6765 VGND.n2604 VGND.n2603 0.0187292
R6766 VGND.n870 VGND.n865 0.0187292
R6767 VGND.n872 VGND.n871 0.0187292
R6768 VGND.n1879 VGND.n1274 0.0187292
R6769 VGND.n1260 VGND.n1253 0.0187292
R6770 VGND.n1949 VGND.n1948 0.0187292
R6771 VGND.n956 VGND.n950 0.0187292
R6772 VGND.n958 VGND.n957 0.0187292
R6773 VGND.n1794 VGND.n1777 0.0187292
R6774 VGND.n2517 VGND.n2516 0.0187292
R6775 VGND.n2513 VGND.n2512 0.0187292
R6776 VGND.n2458 VGND.n2457 0.0187292
R6777 VGND.n2431 VGND.n2430 0.0187292
R6778 VGND.n3007 VGND.n3006 0.0187292
R6779 VGND.n1084 VGND.n500 0.0187292
R6780 VGND.n2972 VGND.n2971 0.0187292
R6781 VGND.n2371 VGND.n1027 0.0187292
R6782 VGND.n2368 VGND.n2347 0.0187292
R6783 VGND.n2297 VGND.n2296 0.0183038
R6784 VGND.n2298 VGND.n2295 0.0182893
R6785 VGND VGND.n986 0.0174271
R6786 VGND.n472 VGND.n471 0.0158654
R6787 VGND.n3466 VGND.n3465 0.0148229
R6788 VGND.n3134 VGND.n216 0.0148229
R6789 VGND.n3317 VGND.n3298 0.0148229
R6790 VGND.n2258 VGND 0.0148229
R6791 VGND VGND.n704 0.0148229
R6792 VGND.n3047 VGND 0.0140546
R6793 VGND.n2156 VGND.n2155 0.0135208
R6794 VGND.n2287 VGND.n1122 0.0135208
R6795 VGND.n2959 VGND.n513 0.0135208
R6796 VGND.n1192 VGND.n1186 0.0135208
R6797 VGND.n2050 VGND.n2044 0.0135208
R6798 VGND.n2880 VGND.n2879 0.0135208
R6799 VGND.n2664 VGND.n2663 0.0135208
R6800 VGND.n727 VGND.n716 0.0135208
R6801 VGND.n2800 VGND.n2799 0.0135208
R6802 VGND.n1329 VGND.n1319 0.0135208
R6803 VGND.n1493 VGND.n1492 0.0135208
R6804 VGND.n2649 VGND.n767 0.0135208
R6805 VGND.n1545 VGND.n1539 0.0135208
R6806 VGND.n1594 VGND.n1589 0.0135208
R6807 VGND.n2576 VGND.n847 0.0135208
R6808 VGND.n1733 VGND.n1293 0.0135208
R6809 VGND.n1906 VGND.n1903 0.0135208
R6810 VGND.n2568 VGND.n929 0.0135208
R6811 VGND.n1756 VGND.n1755 0.0135208
R6812 VGND.n1988 VGND.n1229 0.0135208
R6813 VGND.n2491 VGND.n2490 0.0135208
R6814 VGND.n254 VGND.n253 0.0135208
R6815 VGND.n1073 VGND.n1072 0.0135208
R6816 VGND.n2313 VGND.n2312 0.0135208
R6817 VGND VGND.n927 0.0109167
R6818 VGND.n1066 VGND 0.0109167
R6819 VGND.n2879 VGND 0.00961458
R6820 VGND.n2799 VGND 0.00961458
R6821 VGND.n2152 VGND.n1177 0.00878194
R6822 VGND.n1333 VGND.n1316 0.00878194
R6823 VGND.n1728 VGND.n1298 0.00878194
R6824 VGND.n242 VGND.n235 0.00838554
R6825 VGND.n3045 VGND.n3044 0.00838554
R6826 VGND.n2192 VGND.n1167 0.0083125
R6827 VGND.n2129 VGND.n2128 0.0083125
R6828 VGND.n2065 VGND.n572 0.0083125
R6829 VGND.n2699 VGND.n746 0.0083125
R6830 VGND.n1525 VGND.n1303 0.0083125
R6831 VGND.n1462 VGND.n1399 0.0083125
R6832 VGND.n1692 VGND.n1691 0.0083125
R6833 VGND.n1626 VGND.n1613 0.0083125
R6834 VGND.n1872 VGND.n1282 0.0083125
R6835 VGND.n1959 VGND.n1250 0.0083125
R6836 VGND.n1803 VGND.n1802 0.0083125
R6837 VGND.n1997 VGND.n986 0.0083125
R6838 VGND.n269 VGND.n265 0.0083125
R6839 VGND.n1094 VGND.n1081 0.0083125
R6840 VGND.n2386 VGND.n2381 0.00808197
R6841 VGND.n3046 VGND.n235 0.00790157
R6842 VGND.n3046 VGND.n3045 0.00790157
R6843 VGND.n2525 VGND 0.00755
R6844 VGND.n2017 VGND 0.00755
R6845 VGND.n1797 VGND 0.00755
R6846 VGND.n1829 VGND 0.00755
R6847 VGND.n2485 VGND 0.00755
R6848 VGND.n982 VGND 0.00755
R6849 VGND.n3047 VGND.n3046 0.0070355
R6850 VGND.n2457 VGND 0.00701042
R6851 VGND.n1051 VGND.n1049 0.00653911
R6852 VGND.n3003 VGND.n234 0.00640857
R6853 VGND.n3015 VGND.n3014 0.00636298
R6854 VGND.n3004 VGND.n3003 0.00636298
R6855 VGND.n2304 VGND.n502 0.00631183
R6856 VGND.n1068 VGND.n1050 0.00624332
R6857 VGND.n1116 VGND.n1051 0.00624332
R6858 VGND.n1048 VGND.n503 0.00604629
R6859 VGND.n2969 VGND.n502 0.00604629
R6860 VGND.n2309 VGND.n2308 0.00579577
R6861 VGND.n564 VGND 0.00570833
R6862 VGND.n639 VGND 0.00570833
R6863 VGND VGND.n1776 0.00570833
R6864 VGND.n2425 VGND 0.00570833
R6865 VGND.n3014 VGND.n234 0.00533429
R6866 VGND.n2295 VGND.n2294 0.0052
R6867 VGND.n2296 VGND.n267 0.0052
R6868 VGND.n2299 VGND.n507 0.0052
R6869 VGND.n2300 VGND.n1023 0.0052
R6870 VGND.n2165 VGND.n2164 0.00513595
R6871 VGND.n1325 VGND.n1324 0.00513595
R6872 VGND.n1834 VGND.n1833 0.00513595
R6873 VGND.n1833 VGND.n1298 0.00513595
R6874 VGND.n1736 VGND.n1728 0.00513595
R6875 VGND.n1324 VGND.n1316 0.00513595
R6876 VGND.n1334 VGND.n1333 0.00513595
R6877 VGND.n2165 VGND.n2152 0.00513595
R6878 VGND.n2167 VGND.n1177 0.00513595
R6879 VGND.n1068 VGND.n1049 0.00496369
R6880 VGND.n2304 VGND.n1048 0.0047957
R6881 VGND.n52 VGND.n51 0.00440625
R6882 VGND.n3142 VGND.n3141 0.00440625
R6883 VGND.n3307 VGND.n3300 0.00440625
R6884 VGND.n2199 VGND 0.00440625
R6885 VGND.n2120 VGND 0.00440625
R6886 VGND.n2706 VGND 0.00440625
R6887 VGND VGND.n956 0.00440625
R6888 VGND.n2309 VGND.n2306 0.00364583
R6889 VGND.n2307 VGND.n1019 0.00364583
R6890 VGND.n2308 VGND.n2307 0.00364583
R6891 VGND.n2306 VGND.n2305 0.00364583
R6892 VGND VGND.n870 0.00310417
R6893 VGND.n37 VGND.n36 0.00180208
R6894 VGND.n3449 VGND.n35 0.00180208
R6895 VGND.n3113 VGND.n3104 0.00180208
R6896 VGND.n3173 VGND.n194 0.00180208
R6897 VGND.n3358 VGND.n106 0.00180208
R6898 VGND.n3355 VGND.n3354 0.00180208
R6899 VGND.n2386 VGND.n2385 0.00152459
R6900 VGND.n2608 VGND.n2607 0.0010875
R6901 VGND.n1380 VGND.n1233 0.0010875
R6902 VGND.n1530 VGND.n1277 0.0010875
R6903 VGND.n1727 VGND.n1532 0.0010875
R6904 VGND.n2580 VGND.n763 0.0010875
R6905 VGND.n2612 VGND.n825 0.0010875
R6906 VDPWR.n711 VDPWR.n707 8629.41
R6907 VDPWR.n711 VDPWR.n708 8629.41
R6908 VDPWR.n713 VDPWR.n707 8629.41
R6909 VDPWR.n713 VDPWR.n708 8629.41
R6910 VDPWR.n696 VDPWR.n692 8629.41
R6911 VDPWR.n696 VDPWR.n693 8629.41
R6912 VDPWR.n698 VDPWR.n692 8629.41
R6913 VDPWR.n698 VDPWR.n693 8629.41
R6914 VDPWR.n680 VDPWR.n676 8629.41
R6915 VDPWR.n680 VDPWR.n677 8629.41
R6916 VDPWR.n682 VDPWR.n676 8629.41
R6917 VDPWR.n682 VDPWR.n677 8629.41
R6918 VDPWR.n666 VDPWR.n660 8629.41
R6919 VDPWR.n664 VDPWR.n660 8629.41
R6920 VDPWR.n666 VDPWR.n662 8629.41
R6921 VDPWR.n664 VDPWR.n662 8629.41
R6922 VDPWR.n522 VDPWR.n518 8629.41
R6923 VDPWR.n522 VDPWR.n519 8629.41
R6924 VDPWR.n524 VDPWR.n518 8629.41
R6925 VDPWR.n524 VDPWR.n519 8629.41
R6926 VDPWR.n507 VDPWR.n503 8629.41
R6927 VDPWR.n507 VDPWR.n504 8629.41
R6928 VDPWR.n509 VDPWR.n503 8629.41
R6929 VDPWR.n509 VDPWR.n504 8629.41
R6930 VDPWR.n491 VDPWR.n487 8629.41
R6931 VDPWR.n491 VDPWR.n488 8629.41
R6932 VDPWR.n493 VDPWR.n487 8629.41
R6933 VDPWR.n493 VDPWR.n488 8629.41
R6934 VDPWR.n474 VDPWR.n470 8629.41
R6935 VDPWR.n474 VDPWR.n471 8629.41
R6936 VDPWR.n476 VDPWR.n470 8629.41
R6937 VDPWR.n476 VDPWR.n471 8629.41
R6938 VDPWR.n412 VDPWR.n406 8629.41
R6939 VDPWR.n412 VDPWR.n407 8629.41
R6940 VDPWR.n410 VDPWR.n407 8629.41
R6941 VDPWR.n410 VDPWR.n406 8629.41
R6942 VDPWR.n385 VDPWR.n379 8629.41
R6943 VDPWR.n382 VDPWR.n381 8629.41
R6944 VDPWR.n397 VDPWR.n391 8629.41
R6945 VDPWR.n394 VDPWR.n393 8629.41
R6946 VDPWR.n453 VDPWR.n449 8629.41
R6947 VDPWR.n453 VDPWR.n450 8629.41
R6948 VDPWR.n455 VDPWR.n449 8629.41
R6949 VDPWR.n455 VDPWR.n450 8629.41
R6950 VDPWR.n437 VDPWR.n433 8629.41
R6951 VDPWR.n437 VDPWR.n434 8629.41
R6952 VDPWR.n439 VDPWR.n433 8629.41
R6953 VDPWR.n439 VDPWR.n434 8629.41
R6954 VDPWR.n423 VDPWR.n417 8629.41
R6955 VDPWR.n421 VDPWR.n417 8629.41
R6956 VDPWR.n423 VDPWR.n419 8629.41
R6957 VDPWR.n421 VDPWR.n419 8629.41
R6958 VDPWR.n766 VDPWR.n762 8629.41
R6959 VDPWR.n766 VDPWR.n763 8629.41
R6960 VDPWR.n768 VDPWR.n762 8629.41
R6961 VDPWR.n768 VDPWR.n763 8629.41
R6962 VDPWR.n3160 VDPWR.n3154 8629.41
R6963 VDPWR.n3160 VDPWR.n3155 8629.41
R6964 VDPWR.n3158 VDPWR.n3155 8629.41
R6965 VDPWR.n3158 VDPWR.n3154 8629.41
R6966 VDPWR.n3144 VDPWR.n3138 8629.41
R6967 VDPWR.n3144 VDPWR.n3139 8629.41
R6968 VDPWR.n3142 VDPWR.n3139 8629.41
R6969 VDPWR.n3142 VDPWR.n3138 8629.41
R6970 VDPWR.n3125 VDPWR.n3121 8629.41
R6971 VDPWR.n3125 VDPWR.n3122 8629.41
R6972 VDPWR.n3127 VDPWR.n3121 8629.41
R6973 VDPWR.n3127 VDPWR.n3122 8629.41
R6974 VDPWR.n734 VDPWR.n731 5460
R6975 VDPWR.n736 VDPWR.n731 5460
R6976 VDPWR.n734 VDPWR.n732 5460
R6977 VDPWR.n736 VDPWR.n732 5460
R6978 VDPWR.n748 VDPWR.n742 4260
R6979 VDPWR.n746 VDPWR.n745 4260
R6980 VDPWR.t315 VDPWR.n711 2459.29
R6981 VDPWR.n713 VDPWR.t314 2459.29
R6982 VDPWR.t760 VDPWR.n696 2459.29
R6983 VDPWR.n698 VDPWR.t761 2459.29
R6984 VDPWR.t281 VDPWR.n680 2459.29
R6985 VDPWR.n682 VDPWR.t282 2459.29
R6986 VDPWR.t763 VDPWR.n660 2459.29
R6987 VDPWR.t762 VDPWR.n662 2459.29
R6988 VDPWR.t1036 VDPWR.n522 2459.29
R6989 VDPWR.n524 VDPWR.t1035 2459.29
R6990 VDPWR.t67 VDPWR.n507 2459.29
R6991 VDPWR.n509 VDPWR.t13 2459.29
R6992 VDPWR.t122 VDPWR.n491 2459.29
R6993 VDPWR.n493 VDPWR.t121 2459.29
R6994 VDPWR.t956 VDPWR.n474 2459.29
R6995 VDPWR.n476 VDPWR.t957 2459.29
R6996 VDPWR.t345 VDPWR.n410 2459.29
R6997 VDPWR.n412 VDPWR.t1037 2459.29
R6998 VDPWR.t68 VDPWR.n453 2459.29
R6999 VDPWR.n455 VDPWR.t69 2459.29
R7000 VDPWR.t120 VDPWR.n437 2459.29
R7001 VDPWR.n439 VDPWR.t123 2459.29
R7002 VDPWR.t958 VDPWR.n417 2459.29
R7003 VDPWR.t959 VDPWR.n419 2459.29
R7004 VDPWR.t1012 VDPWR.n766 2459.29
R7005 VDPWR.n768 VDPWR.t118 2459.29
R7006 VDPWR.t239 VDPWR.n3158 2459.29
R7007 VDPWR.n3160 VDPWR.t1093 2459.29
R7008 VDPWR.t49 VDPWR.n3142 2459.29
R7009 VDPWR.n3144 VDPWR.t50 2459.29
R7010 VDPWR.t1094 VDPWR.n3125 2459.29
R7011 VDPWR.n3127 VDPWR.t1095 2459.29
R7012 VDPWR.n712 VDPWR.t315 2298.92
R7013 VDPWR.t314 VDPWR.n712 2298.92
R7014 VDPWR.n697 VDPWR.t760 2298.92
R7015 VDPWR.t761 VDPWR.n697 2298.92
R7016 VDPWR.n681 VDPWR.t281 2298.92
R7017 VDPWR.t282 VDPWR.n681 2298.92
R7018 VDPWR.n665 VDPWR.t763 2298.92
R7019 VDPWR.n665 VDPWR.t762 2298.92
R7020 VDPWR.n523 VDPWR.t1036 2298.92
R7021 VDPWR.t1035 VDPWR.n523 2298.92
R7022 VDPWR.n508 VDPWR.t67 2298.92
R7023 VDPWR.t13 VDPWR.n508 2298.92
R7024 VDPWR.n492 VDPWR.t122 2298.92
R7025 VDPWR.t121 VDPWR.n492 2298.92
R7026 VDPWR.n475 VDPWR.t956 2298.92
R7027 VDPWR.t957 VDPWR.n475 2298.92
R7028 VDPWR.n411 VDPWR.t345 2298.92
R7029 VDPWR.t1037 VDPWR.n411 2298.92
R7030 VDPWR.n454 VDPWR.t68 2298.92
R7031 VDPWR.t69 VDPWR.n454 2298.92
R7032 VDPWR.n438 VDPWR.t120 2298.92
R7033 VDPWR.t123 VDPWR.n438 2298.92
R7034 VDPWR.n422 VDPWR.t958 2298.92
R7035 VDPWR.n422 VDPWR.t959 2298.92
R7036 VDPWR.n767 VDPWR.t1012 2298.92
R7037 VDPWR.t118 VDPWR.n767 2298.92
R7038 VDPWR.n3159 VDPWR.t239 2298.92
R7039 VDPWR.t1093 VDPWR.n3159 2298.92
R7040 VDPWR.n3143 VDPWR.t49 2298.92
R7041 VDPWR.t50 VDPWR.n3143 2298.92
R7042 VDPWR.n3126 VDPWR.t1094 2298.92
R7043 VDPWR.t1095 VDPWR.n3126 2298.92
R7044 VDPWR.n1367 VDPWR.n1349 2296.22
R7045 VDPWR.n1700 VDPWR.n1682 2296.22
R7046 VDPWR.n1623 VDPWR.n1622 2296.22
R7047 VDPWR.n2453 VDPWR.n2452 2291.62
R7048 VDPWR.n2452 VDPWR.n2442 1418.92
R7049 VDPWR.n1367 VDPWR.n1366 1408
R7050 VDPWR.n1700 VDPWR.n1699 1408
R7051 VDPWR.n1622 VDPWR.n1621 1408
R7052 VDPWR VDPWR.t565 975.178
R7053 VDPWR VDPWR.t465 975.178
R7054 VDPWR VDPWR.t459 975.178
R7055 VDPWR.n710 VDPWR.n709 920.471
R7056 VDPWR.n695 VDPWR.n694 920.471
R7057 VDPWR.n679 VDPWR.n678 920.471
R7058 VDPWR.n663 VDPWR.n659 920.471
R7059 VDPWR.n521 VDPWR.n520 920.471
R7060 VDPWR.n506 VDPWR.n505 920.471
R7061 VDPWR.n490 VDPWR.n489 920.471
R7062 VDPWR.n473 VDPWR.n472 920.471
R7063 VDPWR.n409 VDPWR.n408 920.471
R7064 VDPWR.n386 VDPWR.n380 920.471
R7065 VDPWR.n398 VDPWR.n392 920.471
R7066 VDPWR.n452 VDPWR.n451 920.471
R7067 VDPWR.n436 VDPWR.n435 920.471
R7068 VDPWR.n420 VDPWR.n416 920.471
R7069 VDPWR.n765 VDPWR.n764 920.471
R7070 VDPWR.n3157 VDPWR.n3156 920.471
R7071 VDPWR.n3141 VDPWR.n3140 920.471
R7072 VDPWR.n3124 VDPWR.n3123 920.471
R7073 VDPWR.n387 VDPWR.n386 917.46
R7074 VDPWR.n399 VDPWR.n398 917.46
R7075 VDPWR.n709 VDPWR.n705 914.447
R7076 VDPWR.n694 VDPWR.n689 914.447
R7077 VDPWR.n678 VDPWR.n673 914.447
R7078 VDPWR.n663 VDPWR.n658 914.447
R7079 VDPWR.n520 VDPWR.n516 914.447
R7080 VDPWR.n505 VDPWR.n500 914.447
R7081 VDPWR.n489 VDPWR.n484 914.447
R7082 VDPWR.n472 VDPWR.n468 914.447
R7083 VDPWR.n408 VDPWR.n404 914.447
R7084 VDPWR.n451 VDPWR.n446 914.447
R7085 VDPWR.n435 VDPWR.n430 914.447
R7086 VDPWR.n420 VDPWR.n415 914.447
R7087 VDPWR.n764 VDPWR.n760 914.447
R7088 VDPWR.n3156 VDPWR.n3151 914.447
R7089 VDPWR.n3140 VDPWR.n3135 914.447
R7090 VDPWR.n3123 VDPWR.n3119 914.447
R7091 VDPWR.t565 VDPWR 877.827
R7092 VDPWR.t465 VDPWR 877.827
R7093 VDPWR.t459 VDPWR 877.827
R7094 VDPWR.n2359 VDPWR.t389 843.261
R7095 VDPWR.n1871 VDPWR.t43 842.073
R7096 VDPWR.n3051 VDPWR.t1151 842.073
R7097 VDPWR.n1184 VDPWR.t349 832.876
R7098 VDPWR.n1826 VDPWR.t576 812.014
R7099 VDPWR.n2107 VDPWR.t493 811.918
R7100 VDPWR.n2172 VDPWR.t706 811.793
R7101 VDPWR.n2865 VDPWR.t309 808.141
R7102 VDPWR.n1239 VDPWR.t612 807.567
R7103 VDPWR.n2459 VDPWR.t512 807.548
R7104 VDPWR.n1796 VDPWR.t651 807.481
R7105 VDPWR.n1767 VDPWR.t753 807.481
R7106 VDPWR.n1761 VDPWR.t552 807.462
R7107 VDPWR.n1834 VDPWR.t454 806.484
R7108 VDPWR.n1327 VDPWR.t675 806.423
R7109 VDPWR.n1127 VDPWR.t547 806.423
R7110 VDPWR.n807 VDPWR.t266 804.845
R7111 VDPWR.n1528 VDPWR.t609 804.731
R7112 VDPWR.n1521 VDPWR.t608 804.731
R7113 VDPWR.n1528 VDPWR.t461 804.731
R7114 VDPWR.n1521 VDPWR.t460 804.731
R7115 VDPWR.n1520 VDPWR.t655 804.731
R7116 VDPWR.n1296 VDPWR.t654 804.731
R7117 VDPWR.n1482 VDPWR.t623 804.731
R7118 VDPWR.n1311 VDPWR.t622 804.731
R7119 VDPWR.n1482 VDPWR.t467 804.731
R7120 VDPWR.n1311 VDPWR.t466 804.731
R7121 VDPWR.n1312 VDPWR.t710 804.731
R7122 VDPWR.n1323 VDPWR.t709 804.731
R7123 VDPWR.n1312 VDPWR.t567 804.731
R7124 VDPWR.n1323 VDPWR.t566 804.731
R7125 VDPWR.n1326 VDPWR.t488 804.731
R7126 VDPWR.n1328 VDPWR.t621 804.731
R7127 VDPWR.n1405 VDPWR.t674 804.731
R7128 VDPWR.n1397 VDPWR.t620 804.731
R7129 VDPWR.n1339 VDPWR.t524 804.731
R7130 VDPWR.n1350 VDPWR.t523 804.731
R7131 VDPWR.n1353 VDPWR.t458 804.731
R7132 VDPWR.n1356 VDPWR.t647 804.731
R7133 VDPWR.n1360 VDPWR.t431 804.731
R7134 VDPWR.n1365 VDPWR.t634 804.731
R7135 VDPWR.n1540 VDPWR.t452 804.731
R7136 VDPWR.n1543 VDPWR.t649 804.731
R7137 VDPWR.n1213 VDPWR.t455 804.731
R7138 VDPWR.n1829 VDPWR.t745 804.731
R7139 VDPWR.n1798 VDPWR.t575 804.731
R7140 VDPWR.n1810 VDPWR.t652 804.731
R7141 VDPWR.n1769 VDPWR.t611 804.731
R7142 VDPWR.n1791 VDPWR.t754 804.731
R7143 VDPWR.n1260 VDPWR.t725 804.731
R7144 VDPWR.n1743 VDPWR.t470 804.731
R7145 VDPWR.n1735 VDPWR.t551 804.731
R7146 VDPWR.n1727 VDPWR.t469 804.731
R7147 VDPWR.n1275 VDPWR.t582 804.731
R7148 VDPWR.n1683 VDPWR.t581 804.731
R7149 VDPWR.n1686 VDPWR.t691 804.731
R7150 VDPWR.n1689 VDPWR.t538 804.731
R7151 VDPWR.n1693 VDPWR.t521 804.731
R7152 VDPWR.n1698 VDPWR.t703 804.731
R7153 VDPWR.n1201 VDPWR.t748 804.731
R7154 VDPWR.n1204 VDPWR.t615 804.731
R7155 VDPWR.n1208 VDPWR.t743 804.731
R7156 VDPWR.n1895 VDPWR.t604 804.731
R7157 VDPWR.n1602 VDPWR.t578 804.731
R7158 VDPWR.n1628 VDPWR.t560 804.731
R7159 VDPWR.n1644 VDPWR.t579 804.731
R7160 VDPWR.n2059 VDPWR.t561 804.731
R7161 VDPWR.n1639 VDPWR.t546 804.731
R7162 VDPWR.t448 VDPWR.n2048 804.731
R7163 VDPWR.n2047 VDPWR.t750 804.731
R7164 VDPWR.n1134 VDPWR.t665 804.731
R7165 VDPWR.n2027 VDPWR.t751 804.731
R7166 VDPWR.n1155 VDPWR.t666 804.731
R7167 VDPWR.n1153 VDPWR.t644 804.731
R7168 VDPWR.n1156 VDPWR.t659 804.731
R7169 VDPWR.n1177 VDPWR.t645 804.731
R7170 VDPWR.n1995 VDPWR.t660 804.731
R7171 VDPWR.n1606 VDPWR.t618 804.731
R7172 VDPWR.n1612 VDPWR.t695 804.731
R7173 VDPWR.n1615 VDPWR.t443 804.731
R7174 VDPWR.n1619 VDPWR.t535 804.731
R7175 VDPWR.t606 VDPWR.n1924 804.731
R7176 VDPWR.n1939 VDPWR.t515 804.731
R7177 VDPWR.n1942 VDPWR.t593 804.731
R7178 VDPWR.n2098 VDPWR.t527 804.731
R7179 VDPWR.n2101 VDPWR.t636 804.731
R7180 VDPWR.n2265 VDPWR.t591 804.731
R7181 VDPWR.n2284 VDPWR.t590 804.731
R7182 VDPWR.n1051 VDPWR.t632 804.731
R7183 VDPWR.n1029 VDPWR.t631 804.731
R7184 VDPWR.n2316 VDPWR.t738 804.731
R7185 VDPWR.n2207 VDPWR.t737 804.731
R7186 VDPWR.n2203 VDPWR.t434 804.731
R7187 VDPWR.n2185 VDPWR.t433 804.731
R7188 VDPWR.n1108 VDPWR.t563 804.731
R7189 VDPWR.n2166 VDPWR.t642 804.731
R7190 VDPWR.n2141 VDPWR.t705 804.731
R7191 VDPWR.n2136 VDPWR.t641 804.731
R7192 VDPWR.n2080 VDPWR.t494 804.731
R7193 VDPWR.n2094 VDPWR.t679 804.731
R7194 VDPWR.n1071 VDPWR.t585 804.731
R7195 VDPWR.n1074 VDPWR.t693 804.731
R7196 VDPWR.n2731 VDPWR.t626 804.731
R7197 VDPWR.n2734 VDPWR.t723 804.731
R7198 VDPWR.n2959 VDPWR.t689 804.731
R7199 VDPWR.n2940 VDPWR.t688 804.731
R7200 VDPWR.n939 VDPWR.t716 804.731
R7201 VDPWR.n2903 VDPWR.t715 804.731
R7202 VDPWR.t588 VDPWR.n2726 804.731
R7203 VDPWR.n2728 VDPWR.t572 804.731
R7204 VDPWR.n2743 VDPWR.t587 804.731
R7205 VDPWR.n932 VDPWR.t677 804.731
R7206 VDPWR.n2972 VDPWR.t446 804.731
R7207 VDPWR.n2552 VDPWR.t708 804.731
R7208 VDPWR.n2555 VDPWR.t491 804.731
R7209 VDPWR.n2559 VDPWR.t721 804.731
R7210 VDPWR.n2564 VDPWR.t500 804.731
R7211 VDPWR.n2597 VDPWR.t497 804.731
R7212 VDPWR.n891 VDPWR.t732 804.731
R7213 VDPWR.n2991 VDPWR.t428 804.731
R7214 VDPWR.n2999 VDPWR.t549 804.731
R7215 VDPWR.n819 VDPWR.t509 804.731
R7216 VDPWR.n2373 VDPWR.t476 804.731
R7217 VDPWR.n2376 VDPWR.t595 804.731
R7218 VDPWR.n2474 VDPWR.t734 804.731
R7219 VDPWR.n2450 VDPWR.t511 804.731
R7220 VDPWR.n834 VDPWR.t533 804.731
R7221 VDPWR.n838 VDPWR.t657 804.731
R7222 VDPWR.n1003 VDPWR.t1119 783.403
R7223 VDPWR.n2210 VDPWR.t419 779.372
R7224 VDPWR.n1065 VDPWR.t1082 779.372
R7225 VDPWR.t664 VDPWR.t749 772.086
R7226 VDPWR.t658 VDPWR.t643 772.086
R7227 VDPWR.t745 VDPWR.n1828 751.692
R7228 VDPWR.t725 VDPWR.n1259 751.692
R7229 VDPWR.t748 VDPWR.n1200 751.692
R7230 VDPWR.t615 VDPWR.n1203 751.692
R7231 VDPWR.n2049 VDPWR.t448 751.692
R7232 VDPWR.n1925 VDPWR.t606 751.692
R7233 VDPWR.t563 VDPWR.n1107 751.692
R7234 VDPWR.n2740 VDPWR.t588 751.692
R7235 VDPWR.t572 VDPWR.n2727 751.692
R7236 VDPWR.t587 VDPWR.n2742 751.692
R7237 VDPWR.t721 VDPWR.n2558 751.692
R7238 VDPWR.t500 VDPWR.n2563 751.692
R7239 VDPWR.t734 VDPWR.n2473 751.692
R7240 VDPWR.t488 VDPWR.n1325 725.173
R7241 VDPWR.t458 VDPWR.n1352 725.173
R7242 VDPWR.t647 VDPWR.n1355 725.173
R7243 VDPWR.t431 VDPWR.n1359 725.173
R7244 VDPWR.t634 VDPWR.n1364 725.173
R7245 VDPWR.t452 VDPWR.n1539 725.173
R7246 VDPWR.t649 VDPWR.n1542 725.173
R7247 VDPWR.t691 VDPWR.n1685 725.173
R7248 VDPWR.t538 VDPWR.n1688 725.173
R7249 VDPWR.t521 VDPWR.n1692 725.173
R7250 VDPWR.t703 VDPWR.n1697 725.173
R7251 VDPWR.t743 VDPWR.n1207 725.173
R7252 VDPWR.t604 VDPWR.n1894 725.173
R7253 VDPWR.t618 VDPWR.n1605 725.173
R7254 VDPWR.t695 VDPWR.n1611 725.173
R7255 VDPWR.t443 VDPWR.n1614 725.173
R7256 VDPWR.t535 VDPWR.n1618 725.173
R7257 VDPWR.t515 VDPWR.n1938 725.173
R7258 VDPWR.t593 VDPWR.n1941 725.173
R7259 VDPWR.t527 VDPWR.n2097 725.173
R7260 VDPWR.t636 VDPWR.n2100 725.173
R7261 VDPWR.t679 VDPWR.n2093 725.173
R7262 VDPWR.t585 VDPWR.n1070 725.173
R7263 VDPWR.t693 VDPWR.n1073 725.173
R7264 VDPWR.t626 VDPWR.n2730 725.173
R7265 VDPWR.t723 VDPWR.n2733 725.173
R7266 VDPWR.t677 VDPWR.n931 725.173
R7267 VDPWR.t446 VDPWR.n2971 725.173
R7268 VDPWR.t708 VDPWR.n2551 725.173
R7269 VDPWR.t491 VDPWR.n2554 725.173
R7270 VDPWR.t497 VDPWR.n2596 725.173
R7271 VDPWR.t732 VDPWR.n890 725.173
R7272 VDPWR.t428 VDPWR.n2990 725.173
R7273 VDPWR.t549 VDPWR.n2998 725.173
R7274 VDPWR.t509 VDPWR.n818 725.173
R7275 VDPWR.t476 VDPWR.n2372 725.173
R7276 VDPWR.t595 VDPWR.n2375 725.173
R7277 VDPWR.t533 VDPWR.n833 725.173
R7278 VDPWR.t657 VDPWR.n837 725.173
R7279 VDPWR.n2637 VDPWR.n2636 717.729
R7280 VDPWR.n2643 VDPWR.n2642 717.729
R7281 VDPWR.n1919 VDPWR.n1916 713.462
R7282 VDPWR.n571 VDPWR.t1024 675.542
R7283 VDPWR.n291 VDPWR.t107 675.542
R7284 VDPWR.n33 VDPWR.t927 675.542
R7285 VDPWR.n879 VDPWR.t915 671.408
R7286 VDPWR.n789 VDPWR.t871 671.408
R7287 VDPWR.n3091 VDPWR.t869 671.408
R7288 VDPWR.n560 VDPWR.t146 671.376
R7289 VDPWR.n280 VDPWR.t765 671.376
R7290 VDPWR.n22 VDPWR.t988 671.376
R7291 VDPWR.n2852 VDPWR.t365 669.655
R7292 VDPWR.n1872 VDPWR.t3 667.734
R7293 VDPWR.n1966 VDPWR.t997 667.734
R7294 VDPWR.n965 VDPWR.t380 667.734
R7295 VDPWR.n2714 VDPWR.t830 667.734
R7296 VDPWR.n2714 VDPWR.t1145 667.734
R7297 VDPWR.n3045 VDPWR.t205 667.734
R7298 VDPWR.n3040 VDPWR.t213 667.734
R7299 VDPWR.n2834 VDPWR.t1135 666.677
R7300 VDPWR.n2668 VDPWR.t1161 666.677
R7301 VDPWR.n2700 VDPWR.t12 666.677
R7302 VDPWR.n2700 VDPWR.t264 666.677
R7303 VDPWR.n3024 VDPWR.t251 666.677
R7304 VDPWR.n3019 VDPWR.t10 666.677
R7305 VDPWR.t504 VDPWR 666.343
R7306 VDPWR.t717 VDPWR 666.343
R7307 VDPWR VDPWR.t752 666.343
R7308 VDPWR VDPWR.t650 666.343
R7309 VDPWR.t477 VDPWR 666.343
R7310 VDPWR.t556 VDPWR 666.343
R7311 VDPWR VDPWR.t684 664.664
R7312 VDPWR.n2657 VDPWR.t35 664.37
R7313 VDPWR.n2909 VDPWR.t813 664.279
R7314 VDPWR.n2677 VDPWR.t382 664.279
R7315 VDPWR.n2684 VDPWR.t317 664.279
R7316 VDPWR.n2938 VDPWR.t978 663.024
R7317 VDPWR.n1841 VDPWR.t175 662.571
R7318 VDPWR.n1987 VDPWR.t919 662.571
R7319 VDPWR.n2793 VDPWR.t162 659.593
R7320 VDPWR.n2417 VDPWR.t834 659.593
R7321 VDPWR.n2434 VDPWR.t325 659.593
R7322 VDPWR.n980 VDPWR.n979 642.188
R7323 VDPWR.n251 VDPWR.t892 633.369
R7324 VDPWR VDPWR.t516 630.375
R7325 VDPWR VDPWR.t435 630.375
R7326 VDPWR VDPWR.t568 630.375
R7327 VDPWR.t673 VDPWR.t619 617.668
R7328 VDPWR.t550 VDPWR.t468 617.668
R7329 VDPWR.t545 VDPWR.t559 617.668
R7330 VDPWR.n814 VDPWR.n813 614.562
R7331 VDPWR.n2860 VDPWR.n2859 613.71
R7332 VDPWR.n1968 VDPWR.n1967 611.178
R7333 VDPWR.n2633 VDPWR.n2625 611.178
R7334 VDPWR.n2657 VDPWR.n2647 611.178
R7335 VDPWR.n2782 VDPWR.n2781 610.861
R7336 VDPWR.n2773 VDPWR.n2772 609.847
R7337 VDPWR.n1001 VDPWR.n1000 609.717
R7338 VDPWR.n1057 VDPWR.n1050 609.303
R7339 VDPWR.n2202 VDPWR.n2201 606.42
R7340 VDPWR.n2231 VDPWR.n2199 606.42
R7341 VDPWR.n2205 VDPWR.n2204 606.42
R7342 VDPWR.n1062 VDPWR.n1061 606.42
R7343 VDPWR.n2282 VDPWR.n1058 606.42
R7344 VDPWR.n998 VDPWR.n997 606.42
R7345 VDPWR.n2221 VDPWR.n2208 605.581
R7346 VDPWR.n2276 VDPWR.n1064 605.581
R7347 VDPWR.n2196 VDPWR.n2195 605.186
R7348 VDPWR.n2194 VDPWR.n1098 605.186
R7349 VDPWR.n1100 VDPWR.n1099 605.186
R7350 VDPWR.n1041 VDPWR.n1040 605.186
R7351 VDPWR.n1039 VDPWR.n1038 605.186
R7352 VDPWR.n2303 VDPWR.n1035 605.186
R7353 VDPWR.n2790 VDPWR.n996 605.186
R7354 VDPWR.n2794 VDPWR.n2792 605.186
R7355 VDPWR.n2814 VDPWR.n983 605.186
R7356 VDPWR.n1990 VDPWR.n1989 604.394
R7357 VDPWR.n2830 VDPWR.n2829 604.394
R7358 VDPWR.n2620 VDPWR.n2619 604.394
R7359 VDPWR.n2649 VDPWR.n2648 604.394
R7360 VDPWR.n2587 VDPWR.n2585 604.394
R7361 VDPWR.n2587 VDPWR.n2586 604.394
R7362 VDPWR.n916 VDPWR.n915 604.394
R7363 VDPWR.n2635 VDPWR.n2634 603.231
R7364 VDPWR.n2353 VDPWR.n2352 603.231
R7365 VDPWR.n1960 VDPWR.n1927 603.052
R7366 VDPWR.n630 VDPWR.n565 602.456
R7367 VDPWR.n651 VDPWR.n540 602.456
R7368 VDPWR.n350 VDPWR.n285 602.456
R7369 VDPWR.n371 VDPWR.n260 602.456
R7370 VDPWR.n2777 VDPWR.n2776 602.456
R7371 VDPWR.n92 VDPWR.n27 602.456
R7372 VDPWR.n113 VDPWR.n2 602.456
R7373 VDPWR.n1221 VDPWR.n1220 601.097
R7374 VDPWR.n937 VDPWR.n936 601.097
R7375 VDPWR.n3014 VDPWR.n919 601.097
R7376 VDPWR.n2890 VDPWR.n2887 599.159
R7377 VDPWR.n2791 VDPWR.n995 596.442
R7378 VDPWR.n2421 VDPWR.n2419 596.442
R7379 VDPWR.n2519 VDPWR.n2436 596.442
R7380 VDPWR.n2771 VDPWR.n2770 589.481
R7381 VDPWR.n2872 VDPWR.n961 588.318
R7382 VDPWR.n546 VDPWR.n545 585
R7383 VDPWR.n544 VDPWR.n543 585
R7384 VDPWR.n266 VDPWR.n265 585
R7385 VDPWR.n264 VDPWR.n263 585
R7386 VDPWR.n2836 VDPWR.n2835 585
R7387 VDPWR.n2874 VDPWR.n2873 585
R7388 VDPWR.n2769 VDPWR.n2768 585
R7389 VDPWR.n8 VDPWR.n7 585
R7390 VDPWR.n6 VDPWR.n5 585
R7391 VDPWR.n737 VDPWR.n730 582.4
R7392 VDPWR.n733 VDPWR.n730 582.4
R7393 VDPWR.t610 VDPWR 568.994
R7394 VDPWR.t574 VDPWR 568.994
R7395 VDPWR VDPWR.t447 568.994
R7396 VDPWR.t498 VDPWR.t489 540.46
R7397 VDPWR VDPWR.n250 535.705
R7398 VDPWR.n733 VDPWR.n729 531.923
R7399 VDPWR.n738 VDPWR.n737 531.427
R7400 VDPWR.t640 VDPWR 511.926
R7401 VDPWR VDPWR.t670 510.248
R7402 VDPWR.t1081 VDPWR.t696 496.82
R7403 VDPWR VDPWR.n1166 491.784
R7404 VDPWR.n409 VDPWR.n405 480.764
R7405 VDPWR.n3157 VDPWR.n3152 480.764
R7406 VDPWR.n3141 VDPWR.n3136 480.764
R7407 VDPWR.n710 VDPWR.n706 480.764
R7408 VDPWR.n695 VDPWR.n690 480.764
R7409 VDPWR.n679 VDPWR.n674 480.764
R7410 VDPWR.n667 VDPWR.n659 480.764
R7411 VDPWR.n521 VDPWR.n517 480.764
R7412 VDPWR.n506 VDPWR.n501 480.764
R7413 VDPWR.n490 VDPWR.n485 480.764
R7414 VDPWR.n473 VDPWR.n469 480.764
R7415 VDPWR.n380 VDPWR.n378 480.764
R7416 VDPWR.n392 VDPWR.n390 480.764
R7417 VDPWR.n452 VDPWR.n447 480.764
R7418 VDPWR.n436 VDPWR.n431 480.764
R7419 VDPWR.n424 VDPWR.n416 480.764
R7420 VDPWR.n765 VDPWR.n761 480.764
R7421 VDPWR.n3124 VDPWR.n3120 480.764
R7422 VDPWR VDPWR.t370 470.562
R7423 VDPWR VDPWR.t76 470.562
R7424 VDPWR VDPWR.t246 470.562
R7425 VDPWR VDPWR.t84 470.562
R7426 VDPWR VDPWR.t90 470.562
R7427 VDPWR VDPWR.t310 470.562
R7428 VDPWR VDPWR.t273 470.562
R7429 VDPWR VDPWR.t279 470.562
R7430 VDPWR.t429 VDPWR.t456 463.252
R7431 VDPWR.t519 VDPWR.t536 463.252
R7432 VDPWR.t616 VDPWR.t441 463.252
R7433 VDPWR.t678 VDPWR.t525 463.252
R7434 VDPWR.t704 VDPWR.t640 463.252
R7435 VDPWR.t687 VDPWR.t462 463.252
R7436 VDPWR VDPWR.t699 458.724
R7437 VDPWR.t516 VDPWR 458.724
R7438 VDPWR VDPWR.t596 458.724
R7439 VDPWR.t435 VDPWR 458.724
R7440 VDPWR VDPWR.t711 458.724
R7441 VDPWR.t568 VDPWR 458.724
R7442 VDPWR.t998 VDPWR.t128 458.216
R7443 VDPWR.n749 VDPWR.n741 454.401
R7444 VDPWR.n743 VDPWR.n741 454.401
R7445 VDPWR.n743 VDPWR.n740 448.736
R7446 VDPWR.n750 VDPWR.n749 448.288
R7447 VDPWR.n178 VDPWR 435.082
R7448 VDPWR.n621 VDPWR.t943 420.25
R7449 VDPWR.n341 VDPWR.t1096 420.25
R7450 VDPWR.t904 VDPWR.n176 420.25
R7451 VDPWR.n83 VDPWR.t949 420.25
R7452 VDPWR.t653 VDPWR 414.577
R7453 VDPWR VDPWR.t492 414.577
R7454 VDPWR VDPWR.t704 414.577
R7455 VDPWR.t462 VDPWR 414.577
R7456 VDPWR.t670 VDPWR 414.577
R7457 VDPWR.n857 VDPWR.t473 390.875
R7458 VDPWR.n1257 VDPWR.t726 389.526
R7459 VDPWR.n2471 VDPWR.t735 389.361
R7460 VDPWR.n1222 VDPWR.t746 388.721
R7461 VDPWR.n320 VDPWR.t437 388.656
R7462 VDPWR.n1350 VDPWR.t505 388.656
R7463 VDPWR.n1391 VDPWR.t506 388.656
R7464 VDPWR.n1503 VDPWR.t685 388.656
R7465 VDPWR.n1292 VDPWR.t686 388.656
R7466 VDPWR.n1683 VDPWR.t718 388.656
R7467 VDPWR.n1721 VDPWR.t719 388.656
R7468 VDPWR.n1133 VDPWR.t449 388.656
R7469 VDPWR.n1602 VDPWR.t478 388.656
R7470 VDPWR.n1627 VDPWR.t479 388.656
R7471 VDPWR.n2090 VDPWR.t557 388.656
R7472 VDPWR.n2082 VDPWR.t558 388.656
R7473 VDPWR.n2179 VDPWR.t564 388.656
R7474 VDPWR.n2628 VDPWR.t484 388.656
R7475 VDPWR.n884 VDPWR.t485 388.656
R7476 VDPWR.n830 VDPWR.t544 388.656
R7477 VDPWR.n596 VDPWR.t517 388.656
R7478 VDPWR.n600 VDPWR.t518 388.656
R7479 VDPWR.n588 VDPWR.t700 388.656
R7480 VDPWR.n624 VDPWR.t701 388.656
R7481 VDPWR.n574 VDPWR.t668 388.656
R7482 VDPWR.n583 VDPWR.t669 388.656
R7483 VDPWR.n548 VDPWR.t682 388.656
R7484 VDPWR.n553 VDPWR.t683 388.656
R7485 VDPWR.n316 VDPWR.t436 388.656
R7486 VDPWR.n308 VDPWR.t597 388.656
R7487 VDPWR.n344 VDPWR.t598 388.656
R7488 VDPWR.n294 VDPWR.t600 388.656
R7489 VDPWR.n303 VDPWR.t601 388.656
R7490 VDPWR.n268 VDPWR.t540 388.656
R7491 VDPWR.n273 VDPWR.t541 388.656
R7492 VDPWR.n1179 VDPWR.t740 388.656
R7493 VDPWR.n1995 VDPWR.t741 388.656
R7494 VDPWR.n1928 VDPWR.t607 388.656
R7495 VDPWR.n2211 VDPWR.t728 388.656
R7496 VDPWR.n1019 VDPWR.t729 388.656
R7497 VDPWR.n1066 VDPWR.t697 388.656
R7498 VDPWR.n2265 VDPWR.t698 388.656
R7499 VDPWR.n2884 VDPWR.t502 388.656
R7500 VDPWR.n2889 VDPWR.t503 388.656
R7501 VDPWR.n2762 VDPWR.t573 388.656
R7502 VDPWR.n2952 VDPWR.t463 388.656
R7503 VDPWR.n2959 VDPWR.t464 388.656
R7504 VDPWR.n917 VDPWR.t554 388.656
R7505 VDPWR.n2987 VDPWR.t555 388.656
R7506 VDPWR.n2411 VDPWR.t638 388.656
R7507 VDPWR.n2420 VDPWR.t639 388.656
R7508 VDPWR.n2398 VDPWR.t439 388.656
R7509 VDPWR.n2357 VDPWR.t440 388.656
R7510 VDPWR.n2525 VDPWR.t481 388.656
R7511 VDPWR.n2437 VDPWR.t482 388.656
R7512 VDPWR.n2450 VDPWR.t671 388.656
R7513 VDPWR.n2485 VDPWR.t672 388.656
R7514 VDPWR.n792 VDPWR.t628 388.656
R7515 VDPWR.n798 VDPWR.t629 388.656
R7516 VDPWR.n864 VDPWR.t472 388.656
R7517 VDPWR.n58 VDPWR.t569 388.656
R7518 VDPWR.n62 VDPWR.t570 388.656
R7519 VDPWR.n50 VDPWR.t712 388.656
R7520 VDPWR.n86 VDPWR.t713 388.656
R7521 VDPWR.n36 VDPWR.t529 388.656
R7522 VDPWR.n45 VDPWR.t530 388.656
R7523 VDPWR.n10 VDPWR.t662 388.656
R7524 VDPWR.n15 VDPWR.t663 388.656
R7525 VDPWR.n1199 VDPWR.t747 387.682
R7526 VDPWR.n1202 VDPWR.t614 387.682
R7527 VDPWR.n2557 VDPWR.t720 387.682
R7528 VDPWR.n2562 VDPWR.t499 387.682
R7529 VDPWR.n1167 VDPWR.t739 386.043
R7530 VDPWR.n820 VDPWR.t543 385.026
R7531 VDPWR.n2091 VDPWR.t680 383.42
R7532 VDPWR VDPWR.t837 381.007
R7533 VDPWR.n1324 VDPWR.t487 380.193
R7534 VDPWR.n1351 VDPWR.t457 380.193
R7535 VDPWR.n1354 VDPWR.t646 380.193
R7536 VDPWR.n1358 VDPWR.t430 380.193
R7537 VDPWR.n1363 VDPWR.t633 380.193
R7538 VDPWR.n1538 VDPWR.t451 380.193
R7539 VDPWR.n1541 VDPWR.t648 380.193
R7540 VDPWR.n1684 VDPWR.t690 380.193
R7541 VDPWR.n1687 VDPWR.t537 380.193
R7542 VDPWR.n1691 VDPWR.t520 380.193
R7543 VDPWR.n1696 VDPWR.t702 380.193
R7544 VDPWR.n1206 VDPWR.t742 380.193
R7545 VDPWR.n1893 VDPWR.t603 380.193
R7546 VDPWR.n1604 VDPWR.t617 380.193
R7547 VDPWR.n1610 VDPWR.t694 380.193
R7548 VDPWR.n1613 VDPWR.t442 380.193
R7549 VDPWR.n1617 VDPWR.t534 380.193
R7550 VDPWR.n1937 VDPWR.t514 380.193
R7551 VDPWR.n1940 VDPWR.t592 380.193
R7552 VDPWR.n2096 VDPWR.t526 380.193
R7553 VDPWR.n2099 VDPWR.t635 380.193
R7554 VDPWR.n1069 VDPWR.t584 380.193
R7555 VDPWR.n1072 VDPWR.t692 380.193
R7556 VDPWR.n2729 VDPWR.t625 380.193
R7557 VDPWR.n2732 VDPWR.t722 380.193
R7558 VDPWR.n930 VDPWR.t676 380.193
R7559 VDPWR.n2970 VDPWR.t445 380.193
R7560 VDPWR.n2550 VDPWR.t707 380.193
R7561 VDPWR.n2553 VDPWR.t490 380.193
R7562 VDPWR.n2595 VDPWR.t496 380.193
R7563 VDPWR.n889 VDPWR.t731 380.193
R7564 VDPWR.n2989 VDPWR.t427 380.193
R7565 VDPWR.n2997 VDPWR.t548 380.193
R7566 VDPWR.n817 VDPWR.t508 380.193
R7567 VDPWR.n2371 VDPWR.t475 380.193
R7568 VDPWR.n2374 VDPWR.t594 380.193
R7569 VDPWR.n832 VDPWR.t532 380.193
R7570 VDPWR.n836 VDPWR.t656 380.193
R7571 VDPWR.n716 VDPWR.n706 379.2
R7572 VDPWR.n700 VDPWR.n690 379.2
R7573 VDPWR.n684 VDPWR.n674 379.2
R7574 VDPWR.n668 VDPWR.n667 379.2
R7575 VDPWR.n527 VDPWR.n517 379.2
R7576 VDPWR.n511 VDPWR.n501 379.2
R7577 VDPWR.n495 VDPWR.n485 379.2
R7578 VDPWR.n479 VDPWR.n469 379.2
R7579 VDPWR.n463 VDPWR.n405 379.2
R7580 VDPWR.n388 VDPWR.n378 379.2
R7581 VDPWR.n400 VDPWR.n390 379.2
R7582 VDPWR.n457 VDPWR.n447 379.2
R7583 VDPWR.n441 VDPWR.n431 379.2
R7584 VDPWR.n425 VDPWR.n424 379.2
R7585 VDPWR.n3168 VDPWR.n761 379.2
R7586 VDPWR.n3162 VDPWR.n3152 379.2
R7587 VDPWR.n3146 VDPWR.n3136 379.2
R7588 VDPWR.n3130 VDPWR.n3120 379.2
R7589 VDPWR VDPWR.t116 369.938
R7590 VDPWR VDPWR.t853 369.938
R7591 VDPWR VDPWR.t1045 369.938
R7592 VDPWR VDPWR.t237 369.938
R7593 VDPWR.t172 VDPWR 369.938
R7594 VDPWR.t182 VDPWR 369.938
R7595 VDPWR.t888 VDPWR 369.938
R7596 VDPWR.t884 VDPWR 369.938
R7597 VDPWR.t291 VDPWR 369.938
R7598 VDPWR.t842 VDPWR 369.938
R7599 VDPWR.t840 VDPWR 369.938
R7600 VDPWR.t898 VDPWR 369.938
R7601 VDPWR VDPWR.t1021 369.938
R7602 VDPWR VDPWR.t59 369.938
R7603 VDPWR VDPWR.t613 360.866
R7604 VDPWR.t619 VDPWR 357.51
R7605 VDPWR.t468 VDPWR 357.51
R7606 VDPWR.t559 VDPWR 357.51
R7607 VDPWR.t586 VDPWR 355.83
R7608 VDPWR.t157 VDPWR.t812 352.474
R7609 VDPWR.t829 VDPWR.t320 352.474
R7610 VDPWR.n141 VDPWR.t859 348.849
R7611 VDPWR.n2828 VDPWR.t774 340.212
R7612 VDPWR VDPWR.t474 337.368
R7613 VDPWR.n2177 VDPWR.t255 336.524
R7614 VDPWR.n1028 VDPWR.t1157 336.524
R7615 VDPWR.n2687 VDPWR.n2603 334.247
R7616 VDPWR VDPWR.t624 334.012
R7617 VDPWR.n1922 VDPWR.n1921 333.99
R7618 VDPWR.n1875 VDPWR.n1874 333.348
R7619 VDPWR.n953 VDPWR.n952 333.348
R7620 VDPWR.n2547 VDPWR.n2546 333.348
R7621 VDPWR.n894 VDPWR.n893 333.348
R7622 VDPWR.n2866 VDPWR.n964 333.346
R7623 VDPWR.n2608 VDPWR.n2607 333.346
R7624 VDPWR.n2547 VDPWR.n2545 333.346
R7625 VDPWR.n897 VDPWR.n896 333.346
R7626 VDPWR.n2386 VDPWR.n2366 328.036
R7627 VDPWR.n1403 VDPWR.t1192 328.005
R7628 VDPWR.n1733 VDPWR.t1286 328.005
R7629 VDPWR.n1630 VDPWR.t1208 328.005
R7630 VDPWR.n2470 VDPWR.n2461 326.202
R7631 VDPWR.n3052 VDPWR.n887 325.639
R7632 VDPWR.n1876 VDPWR.n1873 324.74
R7633 VDPWR.n577 VDPWR.n570 322.329
R7634 VDPWR.n555 VDPWR.n551 322.329
R7635 VDPWR.n297 VDPWR.n290 322.329
R7636 VDPWR.n275 VDPWR.n271 322.329
R7637 VDPWR.n2627 VDPWR.n2626 322.329
R7638 VDPWR.n796 VDPWR.n795 322.329
R7639 VDPWR.n39 VDPWR.n32 322.329
R7640 VDPWR.n17 VDPWR.n13 322.329
R7641 VDPWR.t269 VDPWR.t214 322.262
R7642 VDPWR.n1031 VDPWR.t1216 321.911
R7643 VDPWR.n140 VDPWR.n139 320.976
R7644 VDPWR.n1848 VDPWR.n1847 320.976
R7645 VDPWR.n2916 VDPWR.n2915 320.976
R7646 VDPWR.n2676 VDPWR.n2609 320.976
R7647 VDPWR.n2707 VDPWR.n2582 320.976
R7648 VDPWR.n900 VDPWR.n899 320.976
R7649 VDPWR.n1918 VDPWR.n1917 320.976
R7650 VDPWR.n2853 VDPWR.n2851 320.976
R7651 VDPWR.n2669 VDPWR.n2612 320.976
R7652 VDPWR.n2707 VDPWR.n2581 320.976
R7653 VDPWR.n3026 VDPWR.n913 320.976
R7654 VDPWR.t147 VDPWR.t11 315.548
R7655 VDPWR.t167 VDPWR.t388 315.548
R7656 VDPWR.n2816 VDPWR.n2815 315.089
R7657 VDPWR.n2824 VDPWR.n2823 314.447
R7658 VDPWR.t379 VDPWR.t308 313.87
R7659 VDPWR.n1982 VDPWR.n1981 312.829
R7660 VDPWR.n2406 VDPWR.n2355 312.053
R7661 VDPWR.n2386 VDPWR.n2368 312.053
R7662 VDPWR.n2381 VDPWR.n2370 312.053
R7663 VDPWR.n2513 VDPWR.n2441 312.053
R7664 VDPWR.n2824 VDPWR.n2822 312.051
R7665 VDPWR.n2179 VDPWR.n2178 311.151
R7666 VDPWR.n2310 VDPWR.n1030 311.151
R7667 VDPWR.n2186 VDPWR.n1102 310.904
R7668 VDPWR.n1034 VDPWR.n1033 310.904
R7669 VDPWR.n2514 VDPWR.n2438 310.5
R7670 VDPWR.t522 VDPWR.t504 308.834
R7671 VDPWR.n1430 VDPWR.t486 308.834
R7672 VDPWR.t580 VDPWR.t717 308.834
R7673 VDPWR.t752 VDPWR.t610 308.834
R7674 VDPWR.t650 VDPWR.t574 308.834
R7675 VDPWR.t577 VDPWR.t477 308.834
R7676 VDPWR.t736 VDPWR.t727 308.834
R7677 VDPWR.t571 VDPWR.t586 308.834
R7678 VDPWR.n826 VDPWR.n825 308.755
R7679 VDPWR.n800 VDPWR.n799 308.755
R7680 VDPWR.n2463 VDPWR.n2462 308.755
R7681 VDPWR.n2480 VDPWR.n2458 308.755
R7682 VDPWR.n2531 VDPWR.n2347 308.755
R7683 VDPWR VDPWR.n821 308.755
R7684 VDPWR.n1519 VDPWR.n1291 308.755
R7685 VDPWR.n2761 VDPWR.n1005 308.755
R7686 VDPWR.n2784 VDPWR.n2783 307.204
R7687 VDPWR.n2431 VDPWR.n2348 307.204
R7688 VDPWR.n1440 VDPWR.t1252 306.735
R7689 VDPWR.n1440 VDPWR.t1281 306.735
R7690 VDPWR.n1309 VDPWR.t1168 306.735
R7691 VDPWR.n1309 VDPWR.t1191 306.735
R7692 VDPWR.n1343 VDPWR.t1272 306.735
R7693 VDPWR.n1411 VDPWR.t1213 306.735
R7694 VDPWR.n1506 VDPWR.t1222 306.735
R7695 VDPWR.n1524 VDPWR.t1170 306.735
R7696 VDPWR.n1524 VDPWR.t1195 306.735
R7697 VDPWR.n1279 VDPWR.t1246 306.735
R7698 VDPWR.n1741 VDPWR.t1260 306.735
R7699 VDPWR.n1776 VDPWR.t1235 306.735
R7700 VDPWR.n1770 VDPWR.t1175 306.735
R7701 VDPWR.n1804 VDPWR.t1177 306.735
R7702 VDPWR.n1237 VDPWR.t1223 306.735
R7703 VDPWR.n1835 VDPWR.t1219 306.735
R7704 VDPWR.n1158 VDPWR.t1174 306.735
R7705 VDPWR.n1154 VDPWR.t1184 306.735
R7706 VDPWR.n1150 VDPWR.t1172 306.735
R7707 VDPWR.n1132 VDPWR.t1271 306.735
R7708 VDPWR.n1633 VDPWR.t1224 306.735
R7709 VDPWR.n1625 VDPWR.t1210 306.735
R7710 VDPWR.n2117 VDPWR.t1238 306.735
R7711 VDPWR.n2079 VDPWR.t1209 306.735
R7712 VDPWR.n2077 VDPWR.t1279 306.735
R7713 VDPWR.n2192 VDPWR.t1283 306.735
R7714 VDPWR.n2209 VDPWR.t1173 306.735
R7715 VDPWR.n1063 VDPWR.t1230 306.735
R7716 VDPWR.n950 VDPWR.t1178 306.735
R7717 VDPWR.n2945 VDPWR.t1187 306.735
R7718 VDPWR.n2456 VDPWR.t1264 306.735
R7719 VDPWR.t418 VDPWR 290.372
R7720 VDPWR VDPWR.t450 280.3
R7721 VDPWR VDPWR.t602 280.3
R7722 VDPWR.t994 VDPWR 280.3
R7723 VDPWR VDPWR.t513 280.3
R7724 VDPWR VDPWR.t583 280.3
R7725 VDPWR VDPWR.t444 280.3
R7726 VDPWR VDPWR.t426 280.3
R7727 VDPWR VDPWR.t531 280.3
R7728 VDPWR.t790 VDPWR.t220 278.623
R7729 VDPWR.n147 VDPWR.n146 272.274
R7730 VDPWR.n147 VDPWR.n134 272.274
R7731 VDPWR.n176 VDPWR.n134 272.274
R7732 VDPWR.t47 VDPWR 261.837
R7733 VDPWR VDPWR.t522 260.159
R7734 VDPWR VDPWR.t673 260.159
R7735 VDPWR VDPWR.t580 260.159
R7736 VDPWR VDPWR.t550 260.159
R7737 VDPWR.t724 VDPWR 260.159
R7738 VDPWR.t744 VDPWR 260.159
R7739 VDPWR.t613 VDPWR 260.159
R7740 VDPWR VDPWR.t577 260.159
R7741 VDPWR VDPWR.t545 260.159
R7742 VDPWR.t739 VDPWR 260.159
R7743 VDPWR.t727 VDPWR 260.159
R7744 VDPWR.t696 VDPWR 260.159
R7745 VDPWR VDPWR.t498 260.159
R7746 VDPWR VDPWR.t438 260.159
R7747 VDPWR.t922 VDPWR 260.159
R7748 VDPWR.t63 VDPWR 260.159
R7749 VDPWR.t38 VDPWR 260.159
R7750 VDPWR.n634 VDPWR.n632 259.697
R7751 VDPWR.n354 VDPWR.n352 259.697
R7752 VDPWR.n96 VDPWR.n94 259.697
R7753 VDPWR.n610 VDPWR.t854 255.905
R7754 VDPWR.n615 VDPWR.t117 255.905
R7755 VDPWR.n591 VDPWR.t944 255.905
R7756 VDPWR.n631 VDPWR.t970 255.905
R7757 VDPWR.n539 VDPWR.t187 255.905
R7758 VDPWR.n330 VDPWR.t238 255.905
R7759 VDPWR.n335 VDPWR.t1046 255.905
R7760 VDPWR.n311 VDPWR.t1097 255.905
R7761 VDPWR.n351 VDPWR.t850 255.905
R7762 VDPWR.n259 VDPWR.t177 255.905
R7763 VDPWR.n183 VDPWR.t899 255.905
R7764 VDPWR.n188 VDPWR.t841 255.905
R7765 VDPWR.n193 VDPWR.t843 255.905
R7766 VDPWR.n198 VDPWR.t292 255.905
R7767 VDPWR.n129 VDPWR.t885 255.905
R7768 VDPWR.n159 VDPWR.t889 255.905
R7769 VDPWR.n164 VDPWR.t183 255.905
R7770 VDPWR.n169 VDPWR.t173 255.905
R7771 VDPWR.n135 VDPWR.t905 255.905
R7772 VDPWR.n72 VDPWR.t60 255.905
R7773 VDPWR.n77 VDPWR.t1022 255.905
R7774 VDPWR.n53 VDPWR.t950 255.905
R7775 VDPWR.n93 VDPWR.t1138 255.905
R7776 VDPWR.n1 VDPWR.t881 255.905
R7777 VDPWR.n246 VDPWR.t371 255.904
R7778 VDPWR.n123 VDPWR.t77 255.904
R7779 VDPWR.n124 VDPWR.t247 255.904
R7780 VDPWR.n125 VDPWR.t85 255.904
R7781 VDPWR.n126 VDPWR.t91 255.904
R7782 VDPWR.n204 VDPWR.t311 255.904
R7783 VDPWR.n205 VDPWR.t274 255.904
R7784 VDPWR.n206 VDPWR.t280 255.904
R7785 VDPWR.n119 VDPWR.t893 255.904
R7786 VDPWR.n581 VDPWR.t982 254.475
R7787 VDPWR.n301 VDPWR.t1009 254.475
R7788 VDPWR.n43 VDPWR.t211 254.475
R7789 VDPWR.n606 VDPWR.t58 252.95
R7790 VDPWR.n611 VDPWR.t115 252.95
R7791 VDPWR.n616 VDPWR.t953 252.95
R7792 VDPWR.n650 VDPWR.t185 252.95
R7793 VDPWR.n645 VDPWR.t1163 252.95
R7794 VDPWR.n326 VDPWR.t234 252.95
R7795 VDPWR.n331 VDPWR.t815 252.95
R7796 VDPWR.n336 VDPWR.t1099 252.95
R7797 VDPWR.n370 VDPWR.t179 252.95
R7798 VDPWR.n365 VDPWR.t73 252.95
R7799 VDPWR.n179 VDPWR.t897 252.95
R7800 VDPWR.n184 VDPWR.t839 252.95
R7801 VDPWR.n189 VDPWR.t845 252.95
R7802 VDPWR.n194 VDPWR.t290 252.95
R7803 VDPWR.n199 VDPWR.t883 252.95
R7804 VDPWR.n155 VDPWR.t887 252.95
R7805 VDPWR.n160 VDPWR.t181 252.95
R7806 VDPWR.n165 VDPWR.t171 252.95
R7807 VDPWR.n170 VDPWR.t903 252.95
R7808 VDPWR.n68 VDPWR.t1032 252.95
R7809 VDPWR.n73 VDPWR.t929 252.95
R7810 VDPWR.n78 VDPWR.t947 252.95
R7811 VDPWR.n112 VDPWR.t879 252.95
R7812 VDPWR.n107 VDPWR.t305 252.95
R7813 VDPWR.n120 VDPWR.t369 252.948
R7814 VDPWR.n245 VDPWR.t75 252.948
R7815 VDPWR.n240 VDPWR.t245 252.948
R7816 VDPWR.n235 VDPWR.t87 252.948
R7817 VDPWR.n230 VDPWR.t89 252.948
R7818 VDPWR.n225 VDPWR.t313 252.948
R7819 VDPWR.n220 VDPWR.t276 252.948
R7820 VDPWR.n215 VDPWR.t278 252.948
R7821 VDPWR.n210 VDPWR.t895 252.948
R7822 VDPWR.n630 VDPWR.t980 251.516
R7823 VDPWR.n350 VDPWR.t1011 251.516
R7824 VDPWR.n92 VDPWR.t209 251.516
R7825 VDPWR.n541 VDPWR.t1165 250.724
R7826 VDPWR.n261 VDPWR.t71 250.724
R7827 VDPWR.n3 VDPWR.t307 250.724
R7828 VDPWR.n144 VDPWR.t241 249.363
R7829 VDPWR.t943 VDPWR.t952 248.599
R7830 VDPWR.t116 VDPWR.t114 248.599
R7831 VDPWR.t853 VDPWR.t57 248.599
R7832 VDPWR.t1096 VDPWR.t1098 248.599
R7833 VDPWR.t1045 VDPWR.t814 248.599
R7834 VDPWR.t237 VDPWR.t233 248.599
R7835 VDPWR.t370 VDPWR.t368 248.599
R7836 VDPWR.t76 VDPWR.t74 248.599
R7837 VDPWR.t246 VDPWR.t244 248.599
R7838 VDPWR.t84 VDPWR.t86 248.599
R7839 VDPWR.t90 VDPWR.t88 248.599
R7840 VDPWR.t310 VDPWR.t312 248.599
R7841 VDPWR.t273 VDPWR.t275 248.599
R7842 VDPWR.t279 VDPWR.t277 248.599
R7843 VDPWR.t892 VDPWR.t894 248.599
R7844 VDPWR.t860 VDPWR.t858 248.599
R7845 VDPWR.t242 VDPWR.t860 248.599
R7846 VDPWR.t240 VDPWR.t242 248.599
R7847 VDPWR.t902 VDPWR.t904 248.599
R7848 VDPWR.t170 VDPWR.t172 248.599
R7849 VDPWR.t180 VDPWR.t182 248.599
R7850 VDPWR.t886 VDPWR.t888 248.599
R7851 VDPWR.t882 VDPWR.t884 248.599
R7852 VDPWR.t289 VDPWR.t291 248.599
R7853 VDPWR.t844 VDPWR.t842 248.599
R7854 VDPWR.t838 VDPWR.t840 248.599
R7855 VDPWR.t896 VDPWR.t898 248.599
R7856 VDPWR.t949 VDPWR.t946 248.599
R7857 VDPWR.t1021 VDPWR.t928 248.599
R7858 VDPWR.t59 VDPWR.t1031 248.599
R7859 VDPWR.n633 VDPWR.t972 248.219
R7860 VDPWR.n353 VDPWR.t852 248.219
R7861 VDPWR.n95 VDPWR.t1137 248.219
R7862 VDPWR.n2093 VDPWR.t1188 246.71
R7863 VDPWR.n1325 VDPWR.t1244 245.667
R7864 VDPWR.n1352 VDPWR.t1258 245.667
R7865 VDPWR.n1355 VDPWR.t1225 245.667
R7866 VDPWR.n1359 VDPWR.t1262 245.667
R7867 VDPWR.n1364 VDPWR.t1233 245.667
R7868 VDPWR.n1539 VDPWR.t1257 245.667
R7869 VDPWR.n1542 VDPWR.t1226 245.667
R7870 VDPWR.n1685 VDPWR.t1221 245.667
R7871 VDPWR.n1688 VDPWR.t1266 245.667
R7872 VDPWR.n1692 VDPWR.t1227 245.667
R7873 VDPWR.n1697 VDPWR.t1197 245.667
R7874 VDPWR.n1207 VDPWR.t1220 245.667
R7875 VDPWR.n1894 VDPWR.t1242 245.667
R7876 VDPWR.n1605 VDPWR.t1186 245.667
R7877 VDPWR.n1611 VDPWR.t1169 245.667
R7878 VDPWR.n1614 VDPWR.t1251 245.667
R7879 VDPWR.n1618 VDPWR.t1229 245.667
R7880 VDPWR.n1938 VDPWR.t1232 245.667
R7881 VDPWR.n1941 VDPWR.t1203 245.667
R7882 VDPWR.n2097 VDPWR.t1254 245.667
R7883 VDPWR.n2100 VDPWR.t1183 245.667
R7884 VDPWR.n1070 VDPWR.t1234 245.667
R7885 VDPWR.n1073 VDPWR.t1167 245.667
R7886 VDPWR.n2730 VDPWR.t1218 245.667
R7887 VDPWR.n2733 VDPWR.t1277 245.667
R7888 VDPWR.n931 VDPWR.t1190 245.667
R7889 VDPWR.n2971 VDPWR.t1253 245.667
R7890 VDPWR.n2551 VDPWR.t1179 245.667
R7891 VDPWR.n2554 VDPWR.t1278 245.667
R7892 VDPWR.n2596 VDPWR.t1267 245.667
R7893 VDPWR.n890 VDPWR.t1180 245.667
R7894 VDPWR.n2990 VDPWR.t1285 245.667
R7895 VDPWR.n2998 VDPWR.t1256 245.667
R7896 VDPWR.n818 VDPWR.t1265 245.667
R7897 VDPWR.n2372 VDPWR.t1274 245.667
R7898 VDPWR.n2375 VDPWR.t1211 245.667
R7899 VDPWR.n833 VDPWR.t1248 245.667
R7900 VDPWR.n837 VDPWR.t1185 245.667
R7901 VDPWR.n962 VDPWR.t796 245.064
R7902 VDPWR.n1182 VDPWR.t103 243.512
R7903 VDPWR.n797 VDPWR.t129 241.767
R7904 VDPWR.n2946 VDPWR.t873 240.215
R7905 VDPWR.n2987 VDPWR.t877 240.214
R7906 VDPWR.n1828 VDPWR.t1181 235.319
R7907 VDPWR.n2432 VDPWR.t7 234.982
R7908 VDPWR VDPWR.t872 233.304
R7909 VDPWR.t733 VDPWR.t846 231.625
R7910 VDPWR.t795 VDPWR.t14 229.947
R7911 VDPWR.n146 VDPWR 224.923
R7912 VDPWR.n2405 VDPWR.n2356 223.868
R7913 VDPWR.t831 VDPWR 223.233
R7914 VDPWR.t318 VDPWR 223.233
R7915 VDPWR.n621 VDPWR 221.964
R7916 VDPWR.n341 VDPWR 221.964
R7917 VDPWR.n83 VDPWR 221.964
R7918 VDPWR.t168 VDPWR.t26 221.555
R7919 VDPWR.t920 VDPWR.t1053 221.555
R7920 VDPWR.t200 VDPWR.t198 221.555
R7921 VDPWR.n2633 VDPWR.n2623 221.314
R7922 VDPWR.n1259 VDPWR.t1189 215.827
R7923 VDPWR.n2473 VDPWR.t1280 215.827
R7924 VDPWR VDPWR.t153 213.163
R7925 VDPWR VDPWR.t974 213.163
R7926 VDPWR.n1200 VDPWR.t1166 213.148
R7927 VDPWR.n1203 VDPWR.t1237 213.148
R7928 VDPWR.n2558 VDPWR.t1176 213.148
R7929 VDPWR.n2563 VDPWR.t1276 213.148
R7930 VDPWR.n581 VDPWR.n578 213.119
R7931 VDPWR.n301 VDPWR.n298 213.119
R7932 VDPWR.n43 VDPWR.n40 213.119
R7933 VDPWR.n622 VDPWR.n621 213.119
R7934 VDPWR.n641 VDPWR.n640 213.119
R7935 VDPWR.n342 VDPWR.n341 213.119
R7936 VDPWR.n361 VDPWR.n360 213.119
R7937 VDPWR.n176 VDPWR.n175 213.119
R7938 VDPWR.n136 VDPWR.n134 213.119
R7939 VDPWR.n148 VDPWR.n147 213.119
R7940 VDPWR.n146 VDPWR.n145 213.119
R7941 VDPWR.n2811 VDPWR.n954 213.119
R7942 VDPWR.n3053 VDPWR.n886 213.119
R7943 VDPWR.n3096 VDPWR.n791 213.119
R7944 VDPWR.n84 VDPWR.n83 213.119
R7945 VDPWR.n103 VDPWR.n102 213.119
R7946 VDPWR.n533 VDPWR.t942 212.081
R7947 VDPWR.n534 VDPWR.t951 212.081
R7948 VDPWR.n3173 VDPWR.t948 212.081
R7949 VDPWR.n3174 VDPWR.t945 212.081
R7950 VDPWR.n1106 VDPWR.t1240 211.263
R7951 VDPWR.n598 VDPWR.t1205 210.964
R7952 VDPWR.n589 VDPWR.t1261 210.964
R7953 VDPWR.n575 VDPWR.t1214 210.964
R7954 VDPWR.n550 VDPWR.t1207 210.964
R7955 VDPWR.n318 VDPWR.t1263 210.964
R7956 VDPWR.n309 VDPWR.t1201 210.964
R7957 VDPWR.n295 VDPWR.t1200 210.964
R7958 VDPWR.n270 VDPWR.t1228 210.964
R7959 VDPWR.n1181 VDPWR.t1275 210.964
R7960 VDPWR.n1018 VDPWR.t1273 210.964
R7961 VDPWR.n1068 VDPWR.t1284 210.964
R7962 VDPWR.n2885 VDPWR.t1236 210.964
R7963 VDPWR.n878 VDPWR.t1270 210.964
R7964 VDPWR.n2399 VDPWR.t1269 210.964
R7965 VDPWR.n60 VDPWR.t1215 210.964
R7966 VDPWR.n51 VDPWR.t1282 210.964
R7967 VDPWR.n37 VDPWR.t1268 210.964
R7968 VDPWR.n12 VDPWR.t1217 210.964
R7969 VDPWR.n1431 VDPWR.n1430 209.368
R7970 VDPWR.n1825 VDPWR.n1223 209.368
R7971 VDPWR.n1760 VDPWR.n1262 209.368
R7972 VDPWR.n2001 VDPWR.n1167 209.368
R7973 VDPWR.n1166 VDPWR.n1126 209.368
R7974 VDPWR.n2317 VDPWR.n1024 209.368
R7975 VDPWR.n1110 VDPWR.n1109 209.368
R7976 VDPWR.n2813 VDPWR.n2812 209.368
R7977 VDPWR.n2686 VDPWR.n2685 209.368
R7978 VDPWR.t267 VDPWR 206.45
R7979 VDPWR VDPWR.t744 203.093
R7980 VDPWR.t447 VDPWR 203.093
R7981 VDPWR.t749 VDPWR 203.093
R7982 VDPWR.t643 VDPWR 203.093
R7983 VDPWR VDPWR.t471 203.093
R7984 VDPWR VDPWR.t918 201.413
R7985 VDPWR VDPWR.t992 199.736
R7986 VDPWR VDPWR.t194 199.736
R7987 VDPWR.t952 VDPWR 198.287
R7988 VDPWR.t114 VDPWR 198.287
R7989 VDPWR.t57 VDPWR 198.287
R7990 VDPWR.t1098 VDPWR 198.287
R7991 VDPWR.t814 VDPWR 198.287
R7992 VDPWR.t233 VDPWR 198.287
R7993 VDPWR VDPWR.t902 198.287
R7994 VDPWR VDPWR.t170 198.287
R7995 VDPWR VDPWR.t180 198.287
R7996 VDPWR VDPWR.t886 198.287
R7997 VDPWR VDPWR.t882 198.287
R7998 VDPWR VDPWR.t289 198.287
R7999 VDPWR VDPWR.t844 198.287
R8000 VDPWR VDPWR.t838 198.287
R8001 VDPWR VDPWR.t896 198.287
R8002 VDPWR.t946 VDPWR 198.287
R8003 VDPWR.t928 VDPWR 198.287
R8004 VDPWR.t1031 VDPWR 198.287
R8005 VDPWR.t1150 VDPWR.t202 198.058
R8006 VDPWR.n2051 VDPWR.n2050 197.508
R8007 VDPWR.t25 VDPWR.t2 191.344
R8008 VDPWR.t812 VDPWR.t803 191.344
R8009 VDPWR.t152 VDPWR.t829 191.344
R8010 VDPWR.t1146 VDPWR.t248 189.665
R8011 VDPWR VDPWR.t240 189.409
R8012 VDPWR.n2811 VDPWR 184.63
R8013 VDPWR.n791 VDPWR 184.63
R8014 VDPWR.n643 VDPWR.n642 183.673
R8015 VDPWR.n363 VDPWR.n362 183.673
R8016 VDPWR.n105 VDPWR.n104 183.673
R8017 VDPWR.n535 VDPWR.n534 183.441
R8018 VDPWR.n3175 VDPWR.n3174 183.441
R8019 VDPWR VDPWR.t4 182.952
R8020 VDPWR VDPWR.n641 182.952
R8021 VDPWR.t287 VDPWR 182.952
R8022 VDPWR VDPWR.t302 182.952
R8023 VDPWR VDPWR.n361 182.952
R8024 VDPWR.t285 VDPWR 182.952
R8025 VDPWR VDPWR.t429 182.952
R8026 VDPWR.t486 VDPWR 182.952
R8027 VDPWR.t450 VDPWR 182.952
R8028 VDPWR VDPWR.t519 182.952
R8029 VDPWR.n1223 VDPWR 182.952
R8030 VDPWR.t602 VDPWR 182.952
R8031 VDPWR VDPWR.t616 182.952
R8032 VDPWR.t513 VDPWR 182.952
R8033 VDPWR.t583 VDPWR 182.952
R8034 VDPWR.t444 VDPWR 182.952
R8035 VDPWR.t426 VDPWR 182.952
R8036 VDPWR.t507 VDPWR 182.952
R8037 VDPWR.t531 VDPWR 182.952
R8038 VDPWR VDPWR.t206 182.952
R8039 VDPWR VDPWR.n103 182.952
R8040 VDPWR.t260 VDPWR 182.952
R8041 VDPWR.t1132 VDPWR.t354 181.273
R8042 VDPWR.n1429 VDPWR 179.595
R8043 VDPWR.n1262 VDPWR 179.595
R8044 VDPWR.n1109 VDPWR 179.595
R8045 VDPWR.n1024 VDPWR 179.595
R8046 VDPWR.n2432 VDPWR 179.595
R8047 VDPWR.t356 VDPWR.t1040 174.559
R8048 VDPWR.t227 VDPWR.t799 174.559
R8049 VDPWR.t165 VDPWR.t168 172.881
R8050 VDPWR.t1053 VDPWR.t155 172.881
R8051 VDPWR.t149 VDPWR.t200 172.881
R8052 VDPWR.t1000 VDPWR.t80 172.881
R8053 VDPWR.t914 VDPWR 169.524
R8054 VDPWR.t1040 VDPWR.t833 167.845
R8055 VDPWR.t163 VDPWR.t453 164.488
R8056 VDPWR.t366 VDPWR.t1148 162.81
R8057 VDPWR.t862 VDPWR.t293 162.81
R8058 VDPWR.t250 VDPWR.t973 161.131
R8059 VDPWR.t912 VDPWR.t352 161.131
R8060 VDPWR.n545 VDPWR.n544 159.476
R8061 VDPWR.n265 VDPWR.n264 159.476
R8062 VDPWR.n2873 VDPWR.n2872 159.476
R8063 VDPWR.n2770 VDPWR.n2769 159.476
R8064 VDPWR.n7 VDPWR.n6 159.476
R8065 VDPWR.t24 VDPWR.t165 159.452
R8066 VDPWR.t827 VDPWR.t983 159.452
R8067 VDPWR.t190 VDPWR.t986 159.452
R8068 VDPWR.t155 VDPWR.t804 159.452
R8069 VDPWR.t198 VDPWR.t150 159.452
R8070 VDPWR.t151 VDPWR.t149 159.452
R8071 VDPWR.t142 VDPWR.t283 159.452
R8072 VDPWR.t962 VDPWR.t542 157.774
R8073 VDPWR.n632 VDPWR.t925 157.014
R8074 VDPWR.n352 VDPWR.t105 157.014
R8075 VDPWR.n94 VDPWR.t931 157.014
R8076 VDPWR.t1164 VDPWR.t910 154.417
R8077 VDPWR.t70 VDPWR.t1089 154.417
R8078 VDPWR.t684 VDPWR.t653 154.417
R8079 VDPWR.t346 VDPWR.t134 154.417
R8080 VDPWR.t492 VDPWR.t556 154.417
R8081 VDPWR.t973 VDPWR.t334 154.417
R8082 VDPWR.t306 VDPWR.t55 154.417
R8083 VDPWR VDPWR.t126 152.739
R8084 VDPWR.t453 VDPWR.t174 151.06
R8085 VDPWR.t501 VDPWR.t1141 151.06
R8086 VDPWR.t324 VDPWR.t480 151.06
R8087 VDPWR.t1002 VDPWR.t94 149.382
R8088 VDPWR.t932 VDPWR.t47 149.382
R8089 VDPWR.t30 VDPWR.t924 147.703
R8090 VDPWR.t848 VDPWR.t104 147.703
R8091 VDPWR.t1087 VDPWR.t40 147.703
R8092 VDPWR.t954 VDPWR.t900 147.703
R8093 VDPWR.t194 VDPWR.t22 147.703
R8094 VDPWR.t7 VDPWR.t801 147.703
R8095 VDPWR.t223 VDPWR.t922 147.703
R8096 VDPWR.t159 VDPWR.t63 147.703
R8097 VDPWR.t757 VDPWR.t962 147.703
R8098 VDPWR.t938 VDPWR.t78 147.703
R8099 VDPWR.t960 VDPWR.t930 147.703
R8100 VDPWR.t759 VDPWR.t932 144.346
R8101 VDPWR.t254 VDPWR.t1019 144.346
R8102 VDPWR.t258 VDPWR.t256 144.346
R8103 VDPWR.t256 VDPWR.t416 144.346
R8104 VDPWR.t416 VDPWR.t410 144.346
R8105 VDPWR.t410 VDPWR.t420 144.346
R8106 VDPWR.t420 VDPWR.t424 144.346
R8107 VDPWR.t424 VDPWR.t396 144.346
R8108 VDPWR.t400 VDPWR.t422 144.346
R8109 VDPWR.t422 VDPWR.t394 144.346
R8110 VDPWR.t398 VDPWR.t402 144.346
R8111 VDPWR.t402 VDPWR.t412 144.346
R8112 VDPWR.t406 VDPWR.t408 144.346
R8113 VDPWR.t408 VDPWR.t404 144.346
R8114 VDPWR.t404 VDPWR.t414 144.346
R8115 VDPWR.t414 VDPWR.t418 144.346
R8116 VDPWR.t1156 VDPWR.t1152 144.346
R8117 VDPWR.t1152 VDPWR.t779 144.346
R8118 VDPWR.t779 VDPWR.t1154 144.346
R8119 VDPWR.t1154 VDPWR.t1061 144.346
R8120 VDPWR.t1061 VDPWR.t1067 144.346
R8121 VDPWR.t1071 VDPWR.t1075 144.346
R8122 VDPWR.t1075 VDPWR.t1065 144.346
R8123 VDPWR.t1065 VDPWR.t1069 144.346
R8124 VDPWR.t1069 VDPWR.t1073 144.346
R8125 VDPWR.t1073 VDPWR.t1063 144.346
R8126 VDPWR.t1079 VDPWR.t1085 144.346
R8127 VDPWR.t1085 VDPWR.t1057 144.346
R8128 VDPWR.t1057 VDPWR.t1059 144.346
R8129 VDPWR.t1059 VDPWR.t1083 144.346
R8130 VDPWR.t1083 VDPWR.t1055 144.346
R8131 VDPWR.t1055 VDPWR.t1077 144.346
R8132 VDPWR.t1112 VDPWR.t1118 144.346
R8133 VDPWR.t1122 VDPWR.t1130 144.346
R8134 VDPWR.t1116 VDPWR.t1126 144.346
R8135 VDPWR.t1106 VDPWR.t1108 144.346
R8136 VDPWR.t775 VDPWR.t773 144.346
R8137 VDPWR.t799 VDPWR.t297 144.346
R8138 VDPWR.t174 VDPWR.t24 142.668
R8139 VDPWR.t394 VDPWR.t398 142.668
R8140 VDPWR.t1124 VDPWR.t1120 142.668
R8141 VDPWR.t804 VDPWR.t977 142.668
R8142 VDPWR.t11 VDPWR.t151 142.668
R8143 VDPWR.t1160 VDPWR.t1000 142.668
R8144 VDPWR.t1033 VDPWR.t1023 140.989
R8145 VDPWR.t924 VDPWR.t971 140.989
R8146 VDPWR.t184 VDPWR.t186 140.989
R8147 VDPWR.t1162 VDPWR.t1164 140.989
R8148 VDPWR.t145 VDPWR.t328 140.989
R8149 VDPWR.t1091 VDPWR.t106 140.989
R8150 VDPWR.t104 VDPWR.t851 140.989
R8151 VDPWR.t178 VDPWR.t176 140.989
R8152 VDPWR.t72 VDPWR.t70 140.989
R8153 VDPWR.t764 VDPWR.t61 140.989
R8154 VDPWR.t825 VDPWR.t163 140.989
R8155 VDPWR.t42 VDPWR.t936 140.989
R8156 VDPWR.t992 VDPWR.t994 140.989
R8157 VDPWR.t810 VDPWR.t157 140.989
R8158 VDPWR.t803 VDPWR.t156 140.989
R8159 VDPWR.t153 VDPWR.t390 140.989
R8160 VDPWR.t320 VDPWR.t831 140.989
R8161 VDPWR.t150 VDPWR.t152 140.989
R8162 VDPWR.t783 VDPWR.t147 140.989
R8163 VDPWR.t80 VDPWR.t322 140.989
R8164 VDPWR.t1029 VDPWR.t221 140.989
R8165 VDPWR.t771 VDPWR.t326 140.989
R8166 VDPWR.t337 VDPWR.t336 140.989
R8167 VDPWR.t974 VDPWR.t392 140.989
R8168 VDPWR.t96 VDPWR.t387 140.989
R8169 VDPWR.t805 VDPWR.t96 140.989
R8170 VDPWR.t868 VDPWR.t916 140.989
R8171 VDPWR.t908 VDPWR.t926 140.989
R8172 VDPWR.t930 VDPWR.t1136 140.989
R8173 VDPWR.t878 VDPWR.t880 140.989
R8174 VDPWR.t304 VDPWR.t306 140.989
R8175 VDPWR.t987 VDPWR.t792 140.989
R8176 VDPWR.n533 VDPWR.t1193 139.78
R8177 VDPWR.n534 VDPWR.t1202 139.78
R8178 VDPWR.n3173 VDPWR.t1206 139.78
R8179 VDPWR.n3174 VDPWR.t1212 139.78
R8180 VDPWR.t1148 VDPWR.t1134 139.311
R8181 VDPWR.t936 VDPWR.t906 137.633
R8182 VDPWR.t940 VDPWR.t0 137.633
R8183 VDPWR.n632 VDPWR.t29 137.079
R8184 VDPWR.n352 VDPWR.t111 137.079
R8185 VDPWR.n94 VDPWR.t1039 137.079
R8186 VDPWR.t348 VDPWR.t133 135.954
R8187 VDPWR.t781 VDPWR.t331 135.954
R8188 VDPWR.t92 VDPWR.t231 135.954
R8189 VDPWR.t81 VDPWR.t797 135.954
R8190 VDPWR.t294 VDPWR.t1015 135.954
R8191 VDPWR.t876 VDPWR 135.954
R8192 VDPWR.n2835 VDPWR.t93 135.268
R8193 VDPWR.t300 VDPWR.t1049 134.276
R8194 VDPWR.t336 VDPWR.t212 130.919
R8195 VDPWR.t338 VDPWR.t890 130.919
R8196 VDPWR.n934 VDPWR.t1247 129.344
R8197 VDPWR.n3015 VDPWR.t1250 129.344
R8198 VDPWR.n863 VDPWR.t1259 129.344
R8199 VDPWR.n2524 VDPWR.t1255 129.344
R8200 VDPWR.n2351 VDPWR.t1194 129.344
R8201 VDPWR VDPWR.t166 129.24
R8202 VDPWR.n2453 VDPWR.t1182 127.695
R8203 VDPWR.t866 VDPWR.t1114 127.562
R8204 VDPWR.n2685 VDPWR.t316 127.562
R8205 VDPWR.t350 VDPWR.t358 127.562
R8206 VDPWR VDPWR.t1132 127.562
R8207 VDPWR.n578 VDPWR 125.883
R8208 VDPWR.n642 VDPWR 125.883
R8209 VDPWR.n298 VDPWR 125.883
R8210 VDPWR.n362 VDPWR 125.883
R8211 VDPWR.t456 VDPWR 125.883
R8212 VDPWR.n1430 VDPWR 125.883
R8213 VDPWR VDPWR.n1429 125.883
R8214 VDPWR.t536 VDPWR 125.883
R8215 VDPWR.n1262 VDPWR 125.883
R8216 VDPWR VDPWR.n1223 125.883
R8217 VDPWR.t441 VDPWR 125.883
R8218 VDPWR.n1166 VDPWR 125.883
R8219 VDPWR.n1167 VDPWR 125.883
R8220 VDPWR.t525 VDPWR 125.883
R8221 VDPWR.n1109 VDPWR 125.883
R8222 VDPWR VDPWR.n1024 125.883
R8223 VDPWR.t624 VDPWR 125.883
R8224 VDPWR.t828 VDPWR.t362 125.883
R8225 VDPWR VDPWR.n2811 125.883
R8226 VDPWR.t489 VDPWR 125.883
R8227 VDPWR.n2685 VDPWR 125.883
R8228 VDPWR.t283 VDPWR.t381 125.883
R8229 VDPWR.t755 VDPWR.t98 125.883
R8230 VDPWR VDPWR.n886 125.883
R8231 VDPWR.t474 VDPWR 125.883
R8232 VDPWR VDPWR.n791 125.883
R8233 VDPWR.n40 VDPWR 125.883
R8234 VDPWR.n104 VDPWR 125.883
R8235 VDPWR.n2741 VDPWR.t1231 124.953
R8236 VDPWR.t968 VDPWR.t1112 124.206
R8237 VDPWR.t316 VDPWR.t383 124.206
R8238 VDPWR.t32 VDPWR.t1025 124.206
R8239 VDPWR.t46 VDPWR 122.526
R8240 VDPWR.t1128 VDPWR.t360 122.526
R8241 VDPWR.t1102 VDPWR.t1042 122.526
R8242 VDPWR.n2812 VDPWR.t1106 122.526
R8243 VDPWR.t53 VDPWR.t1143 122.526
R8244 VDPWR.t589 VDPWR.t1081 120.849
R8245 VDPWR.t299 VDPWR.t364 120.849
R8246 VDPWR.t872 VDPWR.t1044 120.849
R8247 VDPWR.t967 VDPWR.t876 120.849
R8248 VDPWR.n823 VDPWR.t1245 120.76
R8249 VDPWR.n2727 VDPWR.t1204 119.007
R8250 VDPWR.n1925 VDPWR.t1196 118.853
R8251 VDPWR.n2835 VDPWR.t1048 118.549
R8252 VDPWR.t202 VDPWR.t991 117.492
R8253 VDPWR.n2783 VDPWR.t361 117.451
R8254 VDPWR.n2348 VDPWR.t1052 117.451
R8255 VDPWR.n2438 VDPWR.t298 117.451
R8256 VDPWR.n1505 VDPWR.t1171 117.294
R8257 VDPWR.n2116 VDPWR.t1243 117.294
R8258 VDPWR.n3090 VDPWR.t1198 117.294
R8259 VDPWR.n2461 VDPWR.t127 116.343
R8260 VDPWR.n570 VDPWR.t1034 116.341
R8261 VDPWR.n551 VDPWR.t329 116.341
R8262 VDPWR.n290 VDPWR.t1092 116.341
R8263 VDPWR.n271 VDPWR.t62 116.341
R8264 VDPWR.n2626 VDPWR.t355 116.341
R8265 VDPWR.n795 VDPWR.t917 116.341
R8266 VDPWR.n32 VDPWR.t909 116.341
R8267 VDPWR.n13 VDPWR.t793 116.341
R8268 VDPWR.t1027 VDPWR 115.814
R8269 VDPWR.n2859 VDPWR.t363 114.918
R8270 VDPWR.n813 VDPWR.t1147 114.918
R8271 VDPWR.n1349 VDPWR.t1239 114.546
R8272 VDPWR.n1682 VDPWR.t1199 114.546
R8273 VDPWR.n1623 VDPWR.t1241 114.546
R8274 VDPWR.t102 VDPWR.t136 114.135
R8275 VDPWR.t1120 VDPWR.t262 114.135
R8276 VDPWR.n1847 VDPWR.t169 113.98
R8277 VDPWR.n1917 VDPWR.t1003 113.98
R8278 VDPWR.n2851 VDPWR.t232 113.98
R8279 VDPWR.n2915 VDPWR.t1054 113.98
R8280 VDPWR.n2612 VDPWR.t1001 113.98
R8281 VDPWR.n2609 VDPWR.t376 113.98
R8282 VDPWR.n2582 VDPWR.t201 113.98
R8283 VDPWR.n2581 VDPWR.t794 113.98
R8284 VDPWR.n913 VDPWR.t891 113.98
R8285 VDPWR.n899 VDPWR.t865 113.98
R8286 VDPWR.t1023 VDPWR 112.457
R8287 VDPWR.t971 VDPWR 112.457
R8288 VDPWR VDPWR.t145 112.457
R8289 VDPWR.t106 VDPWR 112.457
R8290 VDPWR.t851 VDPWR 112.457
R8291 VDPWR VDPWR.t764 112.457
R8292 VDPWR VDPWR.t868 112.457
R8293 VDPWR.t926 VDPWR 112.457
R8294 VDPWR.t1136 VDPWR 112.457
R8295 VDPWR VDPWR.t987 112.457
R8296 VDPWR.t1004 VDPWR 110.778
R8297 VDPWR.t1019 VDPWR 110.778
R8298 VDPWR.t204 VDPWR.t36 110.778
R8299 VDPWR VDPWR.t964 109.1
R8300 VDPWR VDPWR.t188 109.1
R8301 VDPWR.t40 VDPWR 109.1
R8302 VDPWR VDPWR.t954 109.1
R8303 VDPWR VDPWR.t385 109.1
R8304 VDPWR.t1141 VDPWR 109.1
R8305 VDPWR.t100 VDPWR 109.1
R8306 VDPWR.t192 VDPWR 109.1
R8307 VDPWR VDPWR.t140 109.1
R8308 VDPWR VDPWR.t807 109.1
R8309 VDPWR.t51 VDPWR 109.1
R8310 VDPWR.t248 VDPWR 109.1
R8311 VDPWR.t78 VDPWR 109.1
R8312 VDPWR VDPWR.t216 109.1
R8313 VDPWR.t6 VDPWR 107.421
R8314 VDPWR.t934 VDPWR.t996 107.421
R8315 VDPWR.t1044 VDPWR 107.421
R8316 VDPWR.t553 VDPWR 107.421
R8317 VDPWR.n1429 VDPWR.n1297 106.561
R8318 VDPWR.n2433 VDPWR.n2432 106.559
R8319 VDPWR.n717 VDPWR.n705 105.788
R8320 VDPWR.n701 VDPWR.n689 105.788
R8321 VDPWR.n685 VDPWR.n673 105.788
R8322 VDPWR.n669 VDPWR.n658 105.788
R8323 VDPWR.n528 VDPWR.n516 105.788
R8324 VDPWR.n512 VDPWR.n500 105.788
R8325 VDPWR.n496 VDPWR.n484 105.788
R8326 VDPWR.n480 VDPWR.n468 105.788
R8327 VDPWR.n464 VDPWR.n404 105.788
R8328 VDPWR.n458 VDPWR.n446 105.788
R8329 VDPWR.n442 VDPWR.n430 105.788
R8330 VDPWR.n426 VDPWR.n415 105.788
R8331 VDPWR.n3169 VDPWR.n760 105.788
R8332 VDPWR.n3163 VDPWR.n3151 105.788
R8333 VDPWR.n3147 VDPWR.n3135 105.788
R8334 VDPWR.n3131 VDPWR.n3119 105.788
R8335 VDPWR VDPWR.t664 105.743
R8336 VDPWR VDPWR.t658 105.743
R8337 VDPWR VDPWR.t571 105.743
R8338 VDPWR.t510 VDPWR 105.743
R8339 VDPWR.t265 VDPWR.t38 105.743
R8340 VDPWR.t667 VDPWR.t1033 104.064
R8341 VDPWR.t328 VDPWR.t681 104.064
R8342 VDPWR.t599 VDPWR.t1091 104.064
R8343 VDPWR.t61 VDPWR.t539 104.064
R8344 VDPWR.t1104 VDPWR 104.064
R8345 VDPWR.t1158 VDPWR 104.064
R8346 VDPWR VDPWR.t835 104.064
R8347 VDPWR.t916 VDPWR.t627 104.064
R8348 VDPWR.t528 VDPWR.t908 104.064
R8349 VDPWR.t792 VDPWR.t661 104.064
R8350 VDPWR.t855 VDPWR 102.385
R8351 VDPWR.t235 VDPWR 102.385
R8352 VDPWR.t377 VDPWR.t795 102.385
R8353 VDPWR.t977 VDPWR 102.385
R8354 VDPWR.t34 VDPWR 102.385
R8355 VDPWR.t542 VDPWR 102.385
R8356 VDPWR.t130 VDPWR 102.385
R8357 VDPWR.n2050 VDPWR.n2049 101.591
R8358 VDPWR VDPWR.t20 100.707
R8359 VDPWR.t981 VDPWR 99.0288
R8360 VDPWR.t1008 VDPWR 99.0288
R8361 VDPWR.t630 VDPWR.t1071 99.0288
R8362 VDPWR.t14 VDPWR 99.0288
R8363 VDPWR VDPWR.t768 99.0288
R8364 VDPWR.t210 VDPWR 99.0288
R8365 VDPWR.t368 VDPWR 97.6641
R8366 VDPWR.t74 VDPWR 97.6641
R8367 VDPWR.t244 VDPWR 97.6641
R8368 VDPWR.t86 VDPWR 97.6641
R8369 VDPWR.t88 VDPWR 97.6641
R8370 VDPWR.t312 VDPWR 97.6641
R8371 VDPWR.t275 VDPWR 97.6641
R8372 VDPWR.t277 VDPWR 97.6641
R8373 VDPWR.t894 VDPWR 97.6641
R8374 VDPWR.t1047 VDPWR.t827 97.3503
R8375 VDPWR.n565 VDPWR.t31 96.1553
R8376 VDPWR.n540 VDPWR.t19 96.1553
R8377 VDPWR.n285 VDPWR.t849 96.1553
R8378 VDPWR.n260 VDPWR.t990 96.1553
R8379 VDPWR.n979 VDPWR.t1149 96.1553
R8380 VDPWR.n2887 VDPWR.t23 96.1553
R8381 VDPWR.n2776 VDPWR.t867 96.1553
R8382 VDPWR.n27 VDPWR.t961 96.1553
R8383 VDPWR.n2 VDPWR.t197 96.1553
R8384 VDPWR.t381 VDPWR.t375 95.6719
R8385 VDPWR.t375 VDPWR.t817 95.6719
R8386 VDPWR.t83 VDPWR.t766 95.6719
R8387 VDPWR.n1916 VDPWR.t45 93.81
R8388 VDPWR.n2636 VDPWR.t756 93.81
R8389 VDPWR.n2642 VDPWR.t798 93.81
R8390 VDPWR.n746 VDPWR.n741 92.5005
R8391 VDPWR.n742 VDPWR.n740 92.5005
R8392 VDPWR VDPWR.t18 92.315
R8393 VDPWR VDPWR.t989 92.315
R8394 VDPWR.t1100 VDPWR.t225 92.315
R8395 VDPWR VDPWR.t196 92.315
R8396 VDPWR.t166 VDPWR.t857 90.6365
R8397 VDPWR.t483 VDPWR.t914 90.6365
R8398 VDPWR.t976 VDPWR.t333 90.6365
R8399 VDPWR.t271 VDPWR.t338 90.6365
R8400 VDPWR.n744 VDPWR.n742 89.0328
R8401 VDPWR.n747 VDPWR.n746 89.0328
R8402 VDPWR.t412 VDPWR 88.9581
R8403 VDPWR.t65 VDPWR.t44 87.2797
R8404 VDPWR.t124 VDPWR.t870 87.2797
R8405 VDPWR VDPWR.t966 87.2797
R8406 VDPWR.n544 VDPWR.t911 86.7743
R8407 VDPWR.n264 VDPWR.t1090 86.7743
R8408 VDPWR.n2872 VDPWR.t195 86.7743
R8409 VDPWR.n2770 VDPWR.t969 86.7743
R8410 VDPWR.n995 VDPWR.t1043 86.7743
R8411 VDPWR.n995 VDPWR.t226 86.7743
R8412 VDPWR.n2419 VDPWR.t1041 86.7743
R8413 VDPWR.n2419 VDPWR.t357 86.7743
R8414 VDPWR.n2436 VDPWR.t228 86.7743
R8415 VDPWR.n2436 VDPWR.t800 86.7743
R8416 VDPWR.n6 VDPWR.t56 86.7743
R8417 VDPWR VDPWR.t1079 85.6012
R8418 VDPWR.t837 VDPWR 85.6012
R8419 VDPWR.n578 VDPWR.t981 83.9228
R8420 VDPWR.n298 VDPWR.t1008 83.9228
R8421 VDPWR.t135 VDPWR.t1017 83.9228
R8422 VDPWR.t132 VDPWR.t934 83.9228
R8423 VDPWR.t768 VDPWR.t495 83.9228
R8424 VDPWR.n40 VDPWR.t210 83.9228
R8425 VDPWR.t773 VDPWR 82.2443
R8426 VDPWR.t864 VDPWR.t976 82.2443
R8427 VDPWR.n641 VDPWR.t28 80.5659
R8428 VDPWR.n361 VDPWR.t110 80.5659
R8429 VDPWR.t777 VDPWR 80.5659
R8430 VDPWR.t156 VDPWR.t714 80.5659
R8431 VDPWR.t390 VDPWR 80.5659
R8432 VDPWR VDPWR.t783 80.5659
R8433 VDPWR.t785 VDPWR 80.5659
R8434 VDPWR.t36 VDPWR.t337 80.5659
R8435 VDPWR.t392 VDPWR 80.5659
R8436 VDPWR.n103 VDPWR.t1038 80.5659
R8437 VDPWR.t364 VDPWR.t190 78.8874
R8438 VDPWR.t714 VDPWR.t920 78.8874
R8439 VDPWR.t138 VDPWR.t1160 78.8874
R8440 VDPWR VDPWR.t1051 78.8874
R8441 VDPWR.t297 VDPWR 78.8874
R8442 VDPWR.t4 VDPWR.t667 77.209
R8443 VDPWR.t681 VDPWR.t287 77.209
R8444 VDPWR.t302 VDPWR.t599 77.209
R8445 VDPWR.t539 VDPWR.t285 77.209
R8446 VDPWR.t817 VDPWR.t143 77.209
R8447 VDPWR.t627 VDPWR.t998 77.209
R8448 VDPWR.t471 VDPWR.t507 77.209
R8449 VDPWR.t206 VDPWR.t528 77.209
R8450 VDPWR.t661 VDPWR.t260 77.209
R8451 VDPWR.t396 VDPWR.t432 75.5305
R8452 VDPWR.t161 VDPWR.t1100 75.5305
R8453 VDPWR VDPWR.t912 75.5305
R8454 VDPWR.t1051 VDPWR 75.5305
R8455 VDPWR.t339 VDPWR.n734 75.1466
R8456 VDPWR.n736 VDPWR.t343 75.1466
R8457 VDPWR.t2 VDPWR.t42 73.8521
R8458 VDPWR.t767 VDPWR.t1139 73.8521
R8459 VDPWR.t326 VDPWR.t730 73.8521
R8460 VDPWR.t9 VDPWR 73.8521
R8461 VDPWR.t94 VDPWR.t65 72.1736
R8462 VDPWR.t44 VDPWR.t135 72.1736
R8463 VDPWR.t1108 VDPWR 72.1736
R8464 VDPWR VDPWR.t777 72.1736
R8465 VDPWR.n745 VDPWR.n744 70.6952
R8466 VDPWR.n748 VDPWR.n747 70.6952
R8467 VDPWR.t432 VDPWR.t400 68.8168
R8468 VDPWR.t1110 VDPWR.t161 68.8168
R8469 VDPWR.t333 VDPWR.t271 68.8168
R8470 VDPWR VDPWR.t356 68.8168
R8471 VDPWR VDPWR.t810 67.1383
R8472 VDPWR.t383 VDPWR.t767 67.1383
R8473 VDPWR.t1139 VDPWR.t142 67.1383
R8474 VDPWR.t730 VDPWR.t1027 67.1383
R8475 VDPWR.t966 VDPWR 67.1383
R8476 VDPWR.n545 VDPWR.t965 66.8398
R8477 VDPWR.n265 VDPWR.t189 66.8398
R8478 VDPWR.n2873 VDPWR.t15 66.8398
R8479 VDPWR.n2769 VDPWR.t268 66.8398
R8480 VDPWR.n7 VDPWR.t217 66.8398
R8481 VDPWR.t362 VDPWR.t379 65.4599
R8482 VDPWR VDPWR.t771 65.4599
R8483 VDPWR.t387 VDPWR 65.4599
R8484 VDPWR.n387 VDPWR.n379 64.4072
R8485 VDPWR.n399 VDPWR.n391 64.4072
R8486 VDPWR.t1006 VDPWR.t828 63.7814
R8487 VDPWR.t143 VDPWR.t83 63.7814
R8488 VDPWR.t766 VDPWR.t138 63.7814
R8489 VDPWR.n700 VDPWR.n699 63.3551
R8490 VDPWR.n684 VDPWR.n683 63.3551
R8491 VDPWR.n511 VDPWR.n510 63.3551
R8492 VDPWR.n495 VDPWR.n494 63.3551
R8493 VDPWR.n457 VDPWR.n456 63.3551
R8494 VDPWR.n441 VDPWR.n440 63.3551
R8495 VDPWR.n3162 VDPWR.n3161 63.3551
R8496 VDPWR.n3146 VDPWR.n3145 63.3551
R8497 VDPWR.n565 VDPWR.t856 63.3219
R8498 VDPWR.n540 VDPWR.t789 63.3219
R8499 VDPWR.n285 VDPWR.t236 63.3219
R8500 VDPWR.n260 VDPWR.t109 63.3219
R8501 VDPWR.n1967 VDPWR.t1018 63.3219
R8502 VDPWR.n1967 VDPWR.t935 63.3219
R8503 VDPWR.n2887 VDPWR.t1142 63.3219
R8504 VDPWR.n2776 VDPWR.t386 63.3219
R8505 VDPWR.n2625 VDPWR.t351 63.3219
R8506 VDPWR.n2625 VDPWR.t101 63.3219
R8507 VDPWR.n2647 VDPWR.t1030 63.3219
R8508 VDPWR.n2647 VDPWR.t222 63.3219
R8509 VDPWR.n27 VDPWR.t131 63.3219
R8510 VDPWR.n2 VDPWR.t113 63.3219
R8511 VDPWR.n716 VDPWR.n715 62.2257
R8512 VDPWR.n527 VDPWR.n526 62.2257
R8513 VDPWR.n463 VDPWR.n462 62.2257
R8514 VDPWR.n3168 VDPWR.n3167 62.2257
R8515 VDPWR VDPWR.t30 62.103
R8516 VDPWR VDPWR.t848 62.103
R8517 VDPWR.t816 VDPWR 62.103
R8518 VDPWR VDPWR.t960 62.103
R8519 VDPWR.n711 VDPWR.n710 61.6672
R8520 VDPWR.n714 VDPWR.n713 61.6672
R8521 VDPWR.n696 VDPWR.n695 61.6672
R8522 VDPWR.n699 VDPWR.n698 61.6672
R8523 VDPWR.n680 VDPWR.n679 61.6672
R8524 VDPWR.n683 VDPWR.n682 61.6672
R8525 VDPWR.n660 VDPWR.n659 61.6672
R8526 VDPWR.n662 VDPWR.n661 61.6672
R8527 VDPWR.n522 VDPWR.n521 61.6672
R8528 VDPWR.n525 VDPWR.n524 61.6672
R8529 VDPWR.n507 VDPWR.n506 61.6672
R8530 VDPWR.n510 VDPWR.n509 61.6672
R8531 VDPWR.n491 VDPWR.n490 61.6672
R8532 VDPWR.n494 VDPWR.n493 61.6672
R8533 VDPWR.n474 VDPWR.n473 61.6672
R8534 VDPWR.n477 VDPWR.n476 61.6672
R8535 VDPWR.n410 VDPWR.n409 61.6672
R8536 VDPWR.n413 VDPWR.n412 61.6672
R8537 VDPWR.n381 VDPWR.n380 61.6672
R8538 VDPWR.n393 VDPWR.n392 61.6672
R8539 VDPWR.n453 VDPWR.n452 61.6672
R8540 VDPWR.n456 VDPWR.n455 61.6672
R8541 VDPWR.n437 VDPWR.n436 61.6672
R8542 VDPWR.n440 VDPWR.n439 61.6672
R8543 VDPWR.n417 VDPWR.n416 61.6672
R8544 VDPWR.n419 VDPWR.n418 61.6672
R8545 VDPWR.n766 VDPWR.n765 61.6672
R8546 VDPWR.n769 VDPWR.n768 61.6672
R8547 VDPWR.n3158 VDPWR.n3157 61.6672
R8548 VDPWR.n3161 VDPWR.n3160 61.6672
R8549 VDPWR.n3142 VDPWR.n3141 61.6672
R8550 VDPWR.n3145 VDPWR.n3144 61.6672
R8551 VDPWR.n3125 VDPWR.n3124 61.6672
R8552 VDPWR.n3128 VDPWR.n3127 61.6672
R8553 VDPWR.n668 VDPWR.n657 61.4728
R8554 VDPWR.n479 VDPWR.n478 61.4728
R8555 VDPWR.n425 VDPWR.n414 61.4728
R8556 VDPWR.n3130 VDPWR.n3129 61.4728
R8557 VDPWR.n534 VDPWR.n533 61.346
R8558 VDPWR.n3174 VDPWR.n3173 61.346
R8559 VDPWR.n383 VDPWR.n379 60.9564
R8560 VDPWR.n384 VDPWR.n381 60.9564
R8561 VDPWR.n395 VDPWR.n391 60.9564
R8562 VDPWR.n396 VDPWR.n393 60.9564
R8563 VDPWR.t870 VDPWR.t51 60.4245
R8564 VDPWR.t293 VDPWR.t864 58.7461
R8565 VDPWR VDPWR.t1002 57.0676
R8566 VDPWR.t1017 VDPWR.t132 57.0676
R8567 VDPWR.t1063 VDPWR 57.0676
R8568 VDPWR.t495 VDPWR.t318 57.0676
R8569 VDPWR.t910 VDPWR 55.3892
R8570 VDPWR.t1089 VDPWR 55.3892
R8571 VDPWR VDPWR.t406 55.3892
R8572 VDPWR.t55 VDPWR 55.3892
R8573 VDPWR VDPWR.t1156 53.7107
R8574 VDPWR.t788 VDPWR 52.0323
R8575 VDPWR.t108 VDPWR 52.0323
R8576 VDPWR VDPWR.t1087 52.0323
R8577 VDPWR VDPWR.t825 52.0323
R8578 VDPWR VDPWR.t1013 52.0323
R8579 VDPWR VDPWR.t736 52.0323
R8580 VDPWR.t900 VDPWR 52.0323
R8581 VDPWR.t225 VDPWR.t1102 52.0323
R8582 VDPWR VDPWR.t16 52.0323
R8583 VDPWR VDPWR.t1158 52.0323
R8584 VDPWR VDPWR.t1006 52.0323
R8585 VDPWR VDPWR.t34 52.0323
R8586 VDPWR VDPWR.t1029 52.0323
R8587 VDPWR.t835 VDPWR 52.0323
R8588 VDPWR.t20 VDPWR 52.0323
R8589 VDPWR.t295 VDPWR 52.0323
R8590 VDPWR.t801 VDPWR 52.0323
R8591 VDPWR VDPWR.t324 52.0323
R8592 VDPWR VDPWR.t159 52.0323
R8593 VDPWR VDPWR.t124 52.0323
R8594 VDPWR VDPWR.t874 52.0323
R8595 VDPWR VDPWR.t757 52.0323
R8596 VDPWR VDPWR.t938 52.0323
R8597 VDPWR.t112 VDPWR 52.0323
R8598 VDPWR.n2050 VDPWR.t1249 50.5057
R8599 VDPWR.t857 VDPWR.t25 50.3539
R8600 VDPWR VDPWR.t687 50.3539
R8601 VDPWR.t354 VDPWR.t483 50.3539
R8602 VDPWR VDPWR.t967 50.3539
R8603 VDPWR VDPWR.t724 48.6754
R8604 VDPWR VDPWR.t605 48.6754
R8605 VDPWR VDPWR.t562 48.6754
R8606 VDPWR VDPWR.t553 48.6754
R8607 VDPWR.t637 VDPWR 48.6754
R8608 VDPWR VDPWR.t510 48.6754
R8609 VDPWR VDPWR.t733 48.6754
R8610 VDPWR.n2051 VDPWR.n1130 46.0805
R8611 VDPWR VDPWR.t28 45.3185
R8612 VDPWR VDPWR.t110 45.3185
R8613 VDPWR.t1067 VDPWR.t630 45.3185
R8614 VDPWR.t1134 VDPWR.t1047 45.3185
R8615 VDPWR VDPWR.t790 45.3185
R8616 VDPWR VDPWR.t229 45.3185
R8617 VDPWR VDPWR.t1038 45.3185
R8618 VDPWR VDPWR.t192 43.6401
R8619 VDPWR.t140 VDPWR 43.6401
R8620 VDPWR.n2783 VDPWR.t263 42.3555
R8621 VDPWR.n2348 VDPWR.t374 42.3555
R8622 VDPWR.n2438 VDPWR.t230 42.3555
R8623 VDPWR VDPWR.t979 41.9616
R8624 VDPWR VDPWR.t1010 41.9616
R8625 VDPWR.t874 VDPWR.t265 41.9616
R8626 VDPWR VDPWR.t208 41.9616
R8627 VDPWR.n1220 VDPWR.t826 41.5552
R8628 VDPWR.n1220 VDPWR.t164 41.5552
R8629 VDPWR.n1989 VDPWR.t1014 41.5552
R8630 VDPWR.n1989 VDPWR.t137 41.5552
R8631 VDPWR.n2829 VDPWR.t1159 41.5552
R8632 VDPWR.n2829 VDPWR.t985 41.5552
R8633 VDPWR.n936 VDPWR.t154 41.5552
R8634 VDPWR.n936 VDPWR.t391 41.5552
R8635 VDPWR.n2619 VDPWR.t82 41.5552
R8636 VDPWR.n2619 VDPWR.t786 41.5552
R8637 VDPWR.n2648 VDPWR.t144 41.5552
R8638 VDPWR.n2648 VDPWR.t323 41.5552
R8639 VDPWR.n2585 VDPWR.t770 41.5552
R8640 VDPWR.n2585 VDPWR.t787 41.5552
R8641 VDPWR.n2586 VDPWR.t148 41.5552
R8642 VDPWR.n2586 VDPWR.t784 41.5552
R8643 VDPWR.n915 VDPWR.t335 41.5552
R8644 VDPWR.n915 VDPWR.t1016 41.5552
R8645 VDPWR.n919 VDPWR.t975 41.5552
R8646 VDPWR.n919 VDPWR.t393 41.5552
R8647 VDPWR.t821 VDPWR.t339 40.7512
R8648 VDPWR.t218 VDPWR.t821 40.7512
R8649 VDPWR.t252 VDPWR.t218 40.7512
R8650 VDPWR.t823 VDPWR.t341 40.7512
R8651 VDPWR.t819 VDPWR.t823 40.7512
R8652 VDPWR.t343 VDPWR.t819 40.7512
R8653 VDPWR VDPWR.t1110 40.2832
R8654 VDPWR.t308 VDPWR.t53 38.6047
R8655 VDPWR.n385 VDPWR.n384 38.5759
R8656 VDPWR.n383 VDPWR.n382 38.5759
R8657 VDPWR.n397 VDPWR.n396 38.5759
R8658 VDPWR.n395 VDPWR.n394 38.5759
R8659 VDPWR VDPWR.t984 36.9263
R8660 VDPWR.t983 VDPWR.t92 36.9263
R8661 VDPWR.t220 VDPWR.t32 36.9263
R8662 VDPWR.n1981 VDPWR.t347 36.4455
R8663 VDPWR.n1291 VDPWR.t1088 36.1587
R8664 VDPWR.n1291 VDPWR.t41 36.1587
R8665 VDPWR.n1005 VDPWR.t901 36.1587
R8666 VDPWR.n1005 VDPWR.t955 36.1587
R8667 VDPWR.n2822 VDPWR.t17 36.1587
R8668 VDPWR.n2822 VDPWR.t332 36.1587
R8669 VDPWR.n825 VDPWR.t939 36.1587
R8670 VDPWR.n825 VDPWR.t79 36.1587
R8671 VDPWR.n799 VDPWR.t875 36.1587
R8672 VDPWR.n799 VDPWR.t39 36.1587
R8673 VDPWR.n2462 VDPWR.t125 36.1587
R8674 VDPWR.n2462 VDPWR.t52 36.1587
R8675 VDPWR.n2458 VDPWR.t160 36.1587
R8676 VDPWR.n2458 VDPWR.t64 36.1587
R8677 VDPWR.n2347 VDPWR.t802 36.1587
R8678 VDPWR.n2347 VDPWR.t8 36.1587
R8679 VDPWR.n2355 VDPWR.t296 36.1587
R8680 VDPWR.n2355 VDPWR.t301 36.1587
R8681 VDPWR.n2368 VDPWR.t97 36.1587
R8682 VDPWR.n2368 VDPWR.t808 36.1587
R8683 VDPWR.n2370 VDPWR.t836 36.1587
R8684 VDPWR.n2370 VDPWR.t141 36.1587
R8685 VDPWR.n2441 VDPWR.t224 36.1587
R8686 VDPWR.n2441 VDPWR.t923 36.1587
R8687 VDPWR.n821 VDPWR.t758 36.1587
R8688 VDPWR.n821 VDPWR.t963 36.1587
R8689 VDPWR.n1847 VDPWR.t27 35.4605
R8690 VDPWR.n1917 VDPWR.t66 35.4605
R8691 VDPWR.n2851 VDPWR.t191 35.4605
R8692 VDPWR.n2915 VDPWR.t921 35.4605
R8693 VDPWR.n2612 VDPWR.t139 35.4605
R8694 VDPWR.n2609 VDPWR.t284 35.4605
R8695 VDPWR.n2582 VDPWR.t199 35.4605
R8696 VDPWR.n2581 VDPWR.t818 35.4605
R8697 VDPWR.n913 VDPWR.t272 35.4605
R8698 VDPWR.n899 VDPWR.t863 35.4605
R8699 VDPWR.t1025 VDPWR.t755 35.2479
R8700 VDPWR.n1969 VDPWR.n1920 34.6358
R8701 VDPWR.n2531 VDPWR.n2530 34.6358
R8702 VDPWR.n2469 VDPWR.n2463 34.6358
R8703 VDPWR.n3079 VDPWR.n800 34.6358
R8704 VDPWR.n1866 VDPWR.n1211 34.6358
R8705 VDPWR.n1870 VDPWR.n1211 34.6358
R8706 VDPWR.n1881 VDPWR.n1209 34.6358
R8707 VDPWR.n1882 VDPWR.n1881 34.6358
R8708 VDPWR.n1969 VDPWR.n1968 34.6358
R8709 VDPWR.n1980 VDPWR.n1186 34.6358
R8710 VDPWR.n2854 VDPWR.n2850 34.6358
R8711 VDPWR.n2858 VDPWR.n967 34.6358
R8712 VDPWR.n2868 VDPWR.n2867 34.6358
R8713 VDPWR.n2641 VDPWR.n2621 34.6358
R8714 VDPWR.n2679 VDPWR.n2678 34.6358
R8715 VDPWR.n2675 VDPWR.n2610 34.6358
R8716 VDPWR.n2671 VDPWR.n2610 34.6358
R8717 VDPWR.n2671 VDPWR.n2670 34.6358
R8718 VDPWR.n2683 VDPWR.n2605 34.6358
R8719 VDPWR.n2567 VDPWR.n2566 34.6358
R8720 VDPWR.n2713 VDPWR.n2712 34.6358
R8721 VDPWR.n2712 VDPWR.n2579 34.6358
R8722 VDPWR.n2708 VDPWR.n2579 34.6358
R8723 VDPWR.n2706 VDPWR.n2705 34.6358
R8724 VDPWR.n2705 VDPWR.n2583 34.6358
R8725 VDPWR.n2701 VDPWR.n2583 34.6358
R8726 VDPWR.n3050 VDPWR.n892 34.6358
R8727 VDPWR.n912 VDPWR.n911 34.6358
R8728 VDPWR.n3027 VDPWR.n912 34.6358
R8729 VDPWR.n2385 VDPWR.n2369 34.6358
R8730 VDPWR.n2512 VDPWR.n2442 34.6358
R8731 VDPWR.n812 VDPWR.n808 34.6358
R8732 VDPWR.n2623 VDPWR.t359 34.4755
R8733 VDPWR.n2356 VDPWR.t1050 34.4755
R8734 VDPWR.n2789 VDPWR.n2788 33.6462
R8735 VDPWR.n2796 VDPWR.n2795 33.6462
R8736 VDPWR.n2813 VDPWR.n984 33.6462
R8737 VDPWR VDPWR.t258 33.5694
R8738 VDPWR.t128 VDPWR 33.5694
R8739 VDPWR.n2859 VDPWR.t1007 33.4905
R8740 VDPWR.n2623 VDPWR.t193 33.4905
R8741 VDPWR.n2356 VDPWR.t21 33.4905
R8742 VDPWR.n813 VDPWR.t249 33.4905
R8743 VDPWR.n979 VDPWR.t367 32.7439
R8744 VDPWR.n388 VDPWR.n387 32.5881
R8745 VDPWR.n400 VDPWR.n399 32.5881
R8746 VDPWR.n2634 VDPWR.t1026 32.5055
R8747 VDPWR.n2634 VDPWR.t99 32.5055
R8748 VDPWR.n2352 VDPWR.t353 32.5055
R8749 VDPWR.n2352 VDPWR.t913 32.5055
R8750 VDPWR.n1983 VDPWR.n1184 32.377
R8751 VDPWR.n2850 VDPWR.n969 32.2581
R8752 VDPWR.n1988 VDPWR.n1987 32.0005
R8753 VDPWR.t1126 VDPWR 31.891
R8754 VDPWR.n752 VDPWR.t373 31.6605
R8755 VDPWR.n2679 VDPWR.n2608 31.624
R8756 VDPWR.n2578 VDPWR.n2547 31.624
R8757 VDPWR.n3046 VDPWR.n894 31.624
R8758 VDPWR.n3041 VDPWR.n897 31.624
R8759 VDPWR.n143 VDPWR.n140 30.8711
R8760 VDPWR.n1876 VDPWR.n1875 30.8711
R8761 VDPWR.n2866 VDPWR.n2865 30.8711
R8762 VDPWR.n2817 VDPWR.n2816 30.7205
R8763 VDPWR.n1927 VDPWR.t48 30.5355
R8764 VDPWR.n1877 VDPWR.n1872 30.4946
R8765 VDPWR.n2714 VDPWR.n2578 30.4946
R8766 VDPWR.n3046 VDPWR.n3045 30.4946
R8767 VDPWR.n3041 VDPWR.n3040 30.4946
R8768 VDPWR.t26 VDPWR 30.2125
R8769 VDPWR VDPWR.t678 30.2125
R8770 VDPWR.t1118 VDPWR.t267 30.2125
R8771 VDPWR.t262 VDPWR.t1116 30.2125
R8772 VDPWR.t98 VDPWR.t350 30.2125
R8773 VDPWR.t214 VDPWR.t204 30.2125
R8774 VDPWR.n2431 VDPWR.n2430 29.3652
R8775 VDPWR.n2785 VDPWR.n2782 29.2576
R8776 VDPWR.n2875 VDPWR.n2871 29.1064
R8777 VDPWR.n723 VDPWR.t340 28.6596
R8778 VDPWR.n725 VDPWR.t344 28.6583
R8779 VDPWR.n642 VDPWR 28.5341
R8780 VDPWR.n362 VDPWR 28.5341
R8781 VDPWR.n886 VDPWR 28.5341
R8782 VDPWR.t212 VDPWR.t862 28.5341
R8783 VDPWR.t846 VDPWR 28.5341
R8784 VDPWR.n104 VDPWR 28.5341
R8785 VDPWR.n2626 VDPWR.t1133 28.4453
R8786 VDPWR.n570 VDPWR.t5 28.4453
R8787 VDPWR.n551 VDPWR.t288 28.4453
R8788 VDPWR.n290 VDPWR.t303 28.4453
R8789 VDPWR.n271 VDPWR.t286 28.4453
R8790 VDPWR.n795 VDPWR.t999 28.4453
R8791 VDPWR.n32 VDPWR.t207 28.4453
R8792 VDPWR.n13 VDPWR.t261 28.4453
R8793 VDPWR.n2461 VDPWR.t847 28.4433
R8794 VDPWR.n1981 VDPWR.t1005 27.5805
R8795 VDPWR.n1927 VDPWR.t933 27.5805
R8796 VDPWR.n1050 VDPWR.t1064 27.5805
R8797 VDPWR.n2178 VDPWR.t1020 27.5805
R8798 VDPWR.n2178 VDPWR.t259 27.5805
R8799 VDPWR.n2201 VDPWR.t403 27.5805
R8800 VDPWR.n2201 VDPWR.t413 27.5805
R8801 VDPWR.n2199 VDPWR.t395 27.5805
R8802 VDPWR.n2195 VDPWR.t401 27.5805
R8803 VDPWR.n2195 VDPWR.t423 27.5805
R8804 VDPWR.n1098 VDPWR.t425 27.5805
R8805 VDPWR.n1098 VDPWR.t397 27.5805
R8806 VDPWR.n1099 VDPWR.t411 27.5805
R8807 VDPWR.n1099 VDPWR.t421 27.5805
R8808 VDPWR.n1102 VDPWR.t257 27.5805
R8809 VDPWR.n1102 VDPWR.t417 27.5805
R8810 VDPWR.n2208 VDPWR.t405 27.5805
R8811 VDPWR.n2208 VDPWR.t415 27.5805
R8812 VDPWR.n2204 VDPWR.t407 27.5805
R8813 VDPWR.n2204 VDPWR.t409 27.5805
R8814 VDPWR.n1030 VDPWR.t1153 27.5805
R8815 VDPWR.n1030 VDPWR.t780 27.5805
R8816 VDPWR.n1040 VDPWR.t1070 27.5805
R8817 VDPWR.n1040 VDPWR.t1074 27.5805
R8818 VDPWR.n1038 VDPWR.t1076 27.5805
R8819 VDPWR.n1038 VDPWR.t1066 27.5805
R8820 VDPWR.n1035 VDPWR.t1068 27.5805
R8821 VDPWR.n1035 VDPWR.t1072 27.5805
R8822 VDPWR.n1033 VDPWR.t1155 27.5805
R8823 VDPWR.n1033 VDPWR.t1062 27.5805
R8824 VDPWR.n1064 VDPWR.t1056 27.5805
R8825 VDPWR.n1064 VDPWR.t1078 27.5805
R8826 VDPWR.n1061 VDPWR.t1060 27.5805
R8827 VDPWR.n1061 VDPWR.t1084 27.5805
R8828 VDPWR.n1058 VDPWR.t1086 27.5805
R8829 VDPWR.n1058 VDPWR.t1058 27.5805
R8830 VDPWR.n2823 VDPWR.t782 27.5805
R8831 VDPWR.n2823 VDPWR.t776 27.5805
R8832 VDPWR.n2815 VDPWR.t1109 27.5805
R8833 VDPWR.n2815 VDPWR.t778 27.5805
R8834 VDPWR.n2772 VDPWR.t1113 27.5805
R8835 VDPWR.n2772 VDPWR.t1115 27.5805
R8836 VDPWR.n1000 VDPWR.t1131 27.5805
R8837 VDPWR.n1000 VDPWR.t1123 27.5805
R8838 VDPWR.n2781 VDPWR.t1127 27.5805
R8839 VDPWR.n2781 VDPWR.t1117 27.5805
R8840 VDPWR.n997 VDPWR.t1125 27.5805
R8841 VDPWR.n996 VDPWR.t1129 27.5805
R8842 VDPWR.n996 VDPWR.t1103 27.5805
R8843 VDPWR.n2792 VDPWR.t1101 27.5805
R8844 VDPWR.n2792 VDPWR.t1111 27.5805
R8845 VDPWR.n983 VDPWR.t1105 27.5805
R8846 VDPWR.n983 VDPWR.t1107 27.5805
R8847 VDPWR.n2837 VDPWR.n2834 27.4829
R8848 VDPWR.n2860 VDPWR.n2858 27.4829
R8849 VDPWR.n2635 VDPWR.n2633 27.4829
R8850 VDPWR.n2701 VDPWR.n2700 27.4829
R8851 VDPWR.n3025 VDPWR.n3024 27.4829
R8852 VDPWR.n1499 VDPWR.n1498 27.0566
R8853 VDPWR.n2904 VDPWR.n2902 27.0566
R8854 VDPWR.n1916 VDPWR.t95 26.9729
R8855 VDPWR.n2636 VDPWR.t33 26.9729
R8856 VDPWR.n2642 VDPWR.t791 26.9729
R8857 VDPWR.t1013 VDPWR.t102 26.8556
R8858 VDPWR.n1866 VDPWR.n1865 26.7859
R8859 VDPWR.n645 VDPWR.n644 26.7299
R8860 VDPWR.n365 VDPWR.n364 26.7299
R8861 VDPWR.n107 VDPWR.n106 26.7299
R8862 VDPWR.n2684 VDPWR.n2683 26.7299
R8863 VDPWR.n139 VDPWR.t861 26.5955
R8864 VDPWR.n139 VDPWR.t243 26.5955
R8865 VDPWR.n1873 VDPWR.t937 26.5955
R8866 VDPWR.n1873 VDPWR.t941 26.5955
R8867 VDPWR.n1874 VDPWR.t907 26.5955
R8868 VDPWR.n1874 VDPWR.t1 26.5955
R8869 VDPWR.n1921 VDPWR.t993 26.5955
R8870 VDPWR.n1921 VDPWR.t995 26.5955
R8871 VDPWR.n1050 VDPWR.t1080 26.5955
R8872 VDPWR.n2199 VDPWR.t399 26.5955
R8873 VDPWR.n964 VDPWR.t54 26.5955
R8874 VDPWR.n964 VDPWR.t378 26.5955
R8875 VDPWR.n997 VDPWR.t1121 26.5955
R8876 VDPWR.n952 VDPWR.t811 26.5955
R8877 VDPWR.n952 VDPWR.t158 26.5955
R8878 VDPWR.n2607 VDPWR.t384 26.5955
R8879 VDPWR.n2607 VDPWR.t1140 26.5955
R8880 VDPWR.n2546 VDPWR.t1144 26.5955
R8881 VDPWR.n2546 VDPWR.t330 26.5955
R8882 VDPWR.n2545 VDPWR.t832 26.5955
R8883 VDPWR.n2545 VDPWR.t321 26.5955
R8884 VDPWR.n2603 VDPWR.t319 26.5955
R8885 VDPWR.n2603 VDPWR.t769 26.5955
R8886 VDPWR.n887 VDPWR.t327 26.5955
R8887 VDPWR.n887 VDPWR.t1028 26.5955
R8888 VDPWR.n893 VDPWR.t203 26.5955
R8889 VDPWR.n893 VDPWR.t270 26.5955
R8890 VDPWR.n896 VDPWR.t215 26.5955
R8891 VDPWR.n896 VDPWR.t37 26.5955
R8892 VDPWR.n2366 VDPWR.t809 26.5955
R8893 VDPWR.n2366 VDPWR.t806 26.5955
R8894 VDPWR.n856 VDPWR.n820 26.3341
R8895 VDPWR.n144 VDPWR.n143 25.977
R8896 VDPWR.n644 VDPWR.n643 25.6953
R8897 VDPWR.n364 VDPWR.n363 25.6953
R8898 VDPWR.n106 VDPWR.n105 25.6953
R8899 VDPWR.n610 VDPWR.n594 25.224
R8900 VDPWR.n606 VDPWR.n594 25.224
R8901 VDPWR.n615 VDPWR.n593 25.224
R8902 VDPWR.n611 VDPWR.n593 25.224
R8903 VDPWR.n617 VDPWR.n591 25.224
R8904 VDPWR.n617 VDPWR.n616 25.224
R8905 VDPWR.n635 VDPWR.n631 25.224
R8906 VDPWR.n330 VDPWR.n314 25.224
R8907 VDPWR.n326 VDPWR.n314 25.224
R8908 VDPWR.n335 VDPWR.n313 25.224
R8909 VDPWR.n331 VDPWR.n313 25.224
R8910 VDPWR.n337 VDPWR.n311 25.224
R8911 VDPWR.n337 VDPWR.n336 25.224
R8912 VDPWR.n355 VDPWR.n351 25.224
R8913 VDPWR.n247 VDPWR.n120 25.224
R8914 VDPWR.n247 VDPWR.n246 25.224
R8915 VDPWR.n245 VDPWR.n244 25.224
R8916 VDPWR.n244 VDPWR.n123 25.224
R8917 VDPWR.n240 VDPWR.n239 25.224
R8918 VDPWR.n239 VDPWR.n124 25.224
R8919 VDPWR.n235 VDPWR.n234 25.224
R8920 VDPWR.n234 VDPWR.n125 25.224
R8921 VDPWR.n230 VDPWR.n229 25.224
R8922 VDPWR.n229 VDPWR.n126 25.224
R8923 VDPWR.n225 VDPWR.n224 25.224
R8924 VDPWR.n224 VDPWR.n204 25.224
R8925 VDPWR.n220 VDPWR.n219 25.224
R8926 VDPWR.n219 VDPWR.n205 25.224
R8927 VDPWR.n215 VDPWR.n214 25.224
R8928 VDPWR.n214 VDPWR.n206 25.224
R8929 VDPWR.n210 VDPWR.n209 25.224
R8930 VDPWR.n209 VDPWR.n119 25.224
R8931 VDPWR.n183 VDPWR.n133 25.224
R8932 VDPWR.n179 VDPWR.n133 25.224
R8933 VDPWR.n188 VDPWR.n132 25.224
R8934 VDPWR.n184 VDPWR.n132 25.224
R8935 VDPWR.n193 VDPWR.n131 25.224
R8936 VDPWR.n189 VDPWR.n131 25.224
R8937 VDPWR.n198 VDPWR.n130 25.224
R8938 VDPWR.n194 VDPWR.n130 25.224
R8939 VDPWR.n200 VDPWR.n129 25.224
R8940 VDPWR.n200 VDPWR.n199 25.224
R8941 VDPWR.n159 VDPWR.n154 25.224
R8942 VDPWR.n155 VDPWR.n154 25.224
R8943 VDPWR.n164 VDPWR.n153 25.224
R8944 VDPWR.n160 VDPWR.n153 25.224
R8945 VDPWR.n169 VDPWR.n152 25.224
R8946 VDPWR.n165 VDPWR.n152 25.224
R8947 VDPWR.n171 VDPWR.n135 25.224
R8948 VDPWR.n171 VDPWR.n170 25.224
R8949 VDPWR.n72 VDPWR.n56 25.224
R8950 VDPWR.n68 VDPWR.n56 25.224
R8951 VDPWR.n77 VDPWR.n55 25.224
R8952 VDPWR.n73 VDPWR.n55 25.224
R8953 VDPWR.n79 VDPWR.n53 25.224
R8954 VDPWR.n79 VDPWR.n78 25.224
R8955 VDPWR.n97 VDPWR.n93 25.224
R8956 VDPWR.n2632 VDPWR.n2629 25.1912
R8957 VDPWR.n2430 VDPWR.n2349 25.1912
R8958 VDPWR.n2412 VDPWR.n2410 25.1912
R8959 VDPWR.n3080 VDPWR.n3079 25.1912
R8960 VDPWR.t986 VDPWR 25.1772
R8961 VDPWR VDPWR.t1150 25.1772
R8962 VDPWR.t388 VDPWR 25.1772
R8963 VDPWR.n725 VDPWR.n724 25.0224
R8964 VDPWR.n727 VDPWR.n726 25.0224
R8965 VDPWR.n723 VDPWR.n722 25.0224
R8966 VDPWR.n1107 VDPWR.n1106 24.0557
R8967 VDPWR.n2687 VDPWR.n2686 23.7181
R8968 VDPWR.n581 VDPWR.n564 23.7181
R8969 VDPWR.n640 VDPWR.n562 23.7181
R8970 VDPWR.n301 VDPWR.n284 23.7181
R8971 VDPWR.n360 VDPWR.n282 23.7181
R8972 VDPWR.n1498 VDPWR.n1297 23.7181
R8973 VDPWR.n1882 VDPWR.n1205 23.7181
R8974 VDPWR.n2738 VDPWR.n2735 23.7181
R8975 VDPWR.n2744 VDPWR.n2738 23.7181
R8976 VDPWR.n2902 VDPWR.n954 23.7181
R8977 VDPWR.n2633 VDPWR.n2632 23.7181
R8978 VDPWR.n2657 VDPWR.n2656 23.7181
R8979 VDPWR.n2567 VDPWR.n2565 23.7181
R8980 VDPWR.n2687 VDPWR.n2594 23.7181
R8981 VDPWR.n2530 VDPWR.n2433 23.7181
R8982 VDPWR.n2380 VDPWR.n2377 23.7181
R8983 VDPWR.n3097 VDPWR.n3096 23.7181
R8984 VDPWR.n43 VDPWR.n26 23.7181
R8985 VDPWR.n102 VDPWR.n24 23.7181
R8986 VDPWR.t1077 VDPWR.t589 23.4987
R8987 VDPWR.t991 VDPWR.t269 23.4987
R8988 VDPWR.t352 VDPWR.t300 23.4987
R8989 VDPWR.n808 VDPWR.n807 22.9652
R8990 VDPWR.n1990 VDPWR.n1988 22.9652
R8991 VDPWR.n2657 VDPWR.n2620 22.9652
R8992 VDPWR.n2649 VDPWR.n2613 22.9652
R8993 VDPWR.n2699 VDPWR.n2587 22.9652
R8994 VDPWR.n3023 VDPWR.n916 22.9652
R8995 VDPWR.n2817 VDPWR.n2814 22.6748
R8996 VDPWR.n2828 VDPWR.n981 22.5887
R8997 VDPWR.n2643 VDPWR.n2641 22.5887
R8998 VDPWR.n2637 VDPWR.n2621 22.5887
R8999 VDPWR.n2774 VDPWR.n1001 22.3091
R9000 VDPWR.n1982 VDPWR.n1980 22.2123
R9001 VDPWR.n1983 VDPWR.n1982 22.2123
R9002 VDPWR.n2824 VDPWR.n2821 22.2123
R9003 VDPWR.n2824 VDPWR.n981 22.2123
R9004 VDPWR.n2387 VDPWR.n2386 22.2123
R9005 VDPWR.n2381 VDPWR.n2369 22.2123
R9006 VDPWR.n2386 VDPWR.n2385 22.2123
R9007 VDPWR.n2381 VDPWR.n2380 22.2123
R9008 VDPWR.n2513 VDPWR.n2512 22.2123
R9009 VDPWR.n2668 VDPWR.n2613 21.8358
R9010 VDPWR.n2700 VDPWR.n2699 21.8358
R9011 VDPWR.n3024 VDPWR.n3023 21.8358
R9012 VDPWR.t360 VDPWR.t1124 21.8203
R9013 VDPWR.t1042 VDPWR.t1128 21.8203
R9014 VDPWR.n2812 VDPWR.t1104 21.8203
R9015 VDPWR.t231 VDPWR.t299 21.8203
R9016 VDPWR.n630 VDPWR.n564 21.4593
R9017 VDPWR.n350 VDPWR.n284 21.4593
R9018 VDPWR.n2656 VDPWR.n2649 21.4593
R9019 VDPWR.n2594 VDPWR.n2587 21.4593
R9020 VDPWR.n92 VDPWR.n26 21.4593
R9021 VDPWR.n2763 VDPWR.n1003 21.05
R9022 VDPWR.n2106 VDPWR.n2091 20.912
R9023 VDPWR.n2780 VDPWR.n1001 20.8462
R9024 VDPWR.n857 VDPWR.n856 20.4852
R9025 VDPWR.n2774 VDPWR.n2773 20.4805
R9026 VDPWR.n735 VDPWR.t252 20.3758
R9027 VDPWR.t341 VDPWR.n735 20.3758
R9028 VDPWR.n611 VDPWR.n610 20.3299
R9029 VDPWR.n616 VDPWR.n615 20.3299
R9030 VDPWR.n331 VDPWR.n330 20.3299
R9031 VDPWR.n336 VDPWR.n335 20.3299
R9032 VDPWR.n246 VDPWR.n245 20.3299
R9033 VDPWR.n240 VDPWR.n123 20.3299
R9034 VDPWR.n235 VDPWR.n124 20.3299
R9035 VDPWR.n230 VDPWR.n125 20.3299
R9036 VDPWR.n225 VDPWR.n126 20.3299
R9037 VDPWR.n220 VDPWR.n204 20.3299
R9038 VDPWR.n215 VDPWR.n205 20.3299
R9039 VDPWR.n210 VDPWR.n206 20.3299
R9040 VDPWR.n184 VDPWR.n183 20.3299
R9041 VDPWR.n189 VDPWR.n188 20.3299
R9042 VDPWR.n194 VDPWR.n193 20.3299
R9043 VDPWR.n199 VDPWR.n198 20.3299
R9044 VDPWR.n155 VDPWR.n129 20.3299
R9045 VDPWR.n160 VDPWR.n159 20.3299
R9046 VDPWR.n165 VDPWR.n164 20.3299
R9047 VDPWR.n170 VDPWR.n169 20.3299
R9048 VDPWR.n73 VDPWR.n72 20.3299
R9049 VDPWR.n78 VDPWR.n77 20.3299
R9050 VDPWR.t18 VDPWR.t184 20.1418
R9051 VDPWR.t989 VDPWR.t178 20.1418
R9052 VDPWR.t1114 VDPWR.t968 20.1418
R9053 VDPWR.t221 VDPWR.t81 20.1418
R9054 VDPWR.t196 VDPWR.t878 20.1418
R9055 VDPWR.n2782 VDPWR.n2780 20.1148
R9056 VDPWR.n2053 VDPWR.n1130 20.0749
R9057 VDPWR.n2463 VDPWR.n789 19.9534
R9058 VDPWR.n2742 VDPWR.n2741 19.9237
R9059 VDPWR.n650 VDPWR.n649 19.8181
R9060 VDPWR.n370 VDPWR.n369 19.8181
R9061 VDPWR.n112 VDPWR.n111 19.8181
R9062 VDPWR.n2784 VDPWR.n998 19.7491
R9063 VDPWR.n2790 VDPWR.n2789 19.7491
R9064 VDPWR.n646 VDPWR.n645 19.6946
R9065 VDPWR.n366 VDPWR.n365 19.6946
R9066 VDPWR.n108 VDPWR.n107 19.6946
R9067 VDPWR.n1966 VDPWR.n1922 19.577
R9068 VDPWR.n2315 VDPWR.n1026 19.2067
R9069 VDPWR.n2226 VDPWR.n2225 18.7808
R9070 VDPWR.n1829 VDPWR.n1827 18.7591
R9071 VDPWR.t1143 VDPWR.t377 18.4634
R9072 VDPWR.t322 VDPWR.t816 18.4634
R9073 VDPWR.n1918 VDPWR.n1186 18.4476
R9074 VDPWR.n2854 VDPWR.n2853 18.4476
R9075 VDPWR.n2676 VDPWR.n2675 18.4476
R9076 VDPWR.n2707 VDPWR.n2706 18.4476
R9077 VDPWR.n911 VDPWR.n900 18.4476
R9078 VDPWR.n3026 VDPWR.n3025 18.4476
R9079 VDPWR.n2821 VDPWR.n982 18.0711
R9080 VDPWR.n2405 VDPWR.n2404 18.0382
R9081 VDPWR.n1576 VDPWR.n1575 17.9678
R9082 VDPWR VDPWR.n2359 17.6841
R9083 VDPWR.n2184 VDPWR.n1103 17.612
R9084 VDPWR.n622 VDPWR.n591 17.3181
R9085 VDPWR.n634 VDPWR.n633 17.3181
R9086 VDPWR.n640 VDPWR.n539 17.3181
R9087 VDPWR.n342 VDPWR.n311 17.3181
R9088 VDPWR.n354 VDPWR.n353 17.3181
R9089 VDPWR.n360 VDPWR.n259 17.3181
R9090 VDPWR.n251 VDPWR.n119 17.3181
R9091 VDPWR.n175 VDPWR.n135 17.3181
R9092 VDPWR.n84 VDPWR.n53 17.3181
R9093 VDPWR.n96 VDPWR.n95 17.3181
R9094 VDPWR.n102 VDPWR.n1 17.3181
R9095 VDPWR.n606 VDPWR.n605 17.2853
R9096 VDPWR.n326 VDPWR.n325 17.2853
R9097 VDPWR.n68 VDPWR.n67 17.2853
R9098 VDPWR.n3052 VDPWR.n3051 16.9417
R9099 VDPWR.n2410 VDPWR.n2353 16.9417
R9100 VDPWR.t1130 VDPWR.t866 16.785
R9101 VDPWR.t438 VDPWR.t167 16.785
R9102 VDPWR.t480 VDPWR.t227 16.785
R9103 VDPWR.n1830 VDPWR.n1829 16.7729
R9104 VDPWR.n2173 VDPWR.n1108 16.7729
R9105 VDPWR.n1466 VDPWR.n1465 16.6847
R9106 VDPWR.n2939 VDPWR.n2938 16.5825
R9107 VDPWR.n631 VDPWR.n630 16.5652
R9108 VDPWR.n635 VDPWR.n634 16.5652
R9109 VDPWR.n351 VDPWR.n350 16.5652
R9110 VDPWR.n355 VDPWR.n354 16.5652
R9111 VDPWR.n93 VDPWR.n92 16.5652
R9112 VDPWR.n97 VDPWR.n96 16.5652
R9113 VDPWR.n2794 VDPWR.n2793 16.4576
R9114 VDPWR.n2670 VDPWR.n2669 16.1887
R9115 VDPWR.n2708 VDPWR.n2707 16.1887
R9116 VDPWR.n3039 VDPWR.n900 16.1887
R9117 VDPWR.n3027 VDPWR.n3026 16.1887
R9118 VDPWR.n250 VDPWR.n120 15.8123
R9119 VDPWR.n179 VDPWR.n178 15.8123
R9120 VDPWR.n732 VDPWR.n730 15.4172
R9121 VDPWR.n735 VDPWR.n732 15.4172
R9122 VDPWR.n731 VDPWR.n729 15.4172
R9123 VDPWR.n735 VDPWR.n731 15.4172
R9124 VDPWR.n2795 VDPWR.n2794 15.3605
R9125 VDPWR.n1107 VDPWR.n1105 15.2281
R9126 VDPWR.n1827 VDPWR.n1222 15.101
R9127 VDPWR.n2861 VDPWR.n965 15.0593
R9128 VDPWR.n2714 VDPWR.n2713 15.0593
R9129 VDPWR.n3045 VDPWR.n3044 15.0593
R9130 VDPWR.n3040 VDPWR.n3039 15.0593
R9131 VDPWR.n2406 VDPWR.n2353 15.0593
R9132 VDPWR.n2514 VDPWR.n2513 15.0593
R9133 VDPWR.n1435 VDPWR.n1434 14.9
R9134 VDPWR.n3097 VDPWR.n789 14.6829
R9135 VDPWR.n1994 VDPWR.n1182 14.6484
R9136 VDPWR.n644 VDPWR.n560 14.6078
R9137 VDPWR.n364 VDPWR.n280 14.6078
R9138 VDPWR.n106 VDPWR.n22 14.6078
R9139 VDPWR.n1481 VDPWR.n1297 14.5851
R9140 VDPWR.n1549 VDPWR.n1537 14.5851
R9141 VDPWR.n2853 VDPWR.n2852 14.3064
R9142 VDPWR.n2643 VDPWR.n2620 14.3064
R9143 VDPWR.n3019 VDPWR.n916 14.3064
R9144 VDPWR.n623 VDPWR.n622 14.2735
R9145 VDPWR.n582 VDPWR.n581 14.2735
R9146 VDPWR.n343 VDPWR.n342 14.2735
R9147 VDPWR.n302 VDPWR.n301 14.2735
R9148 VDPWR.n1948 VDPWR.n1936 14.2735
R9149 VDPWR.n2888 VDPWR.n954 14.2735
R9150 VDPWR.n3053 VDPWR.n885 14.2735
R9151 VDPWR.n3000 VDPWR.n2988 14.2735
R9152 VDPWR.n2526 VDPWR.n2433 14.2735
R9153 VDPWR.n3096 VDPWR.n3095 14.2735
R9154 VDPWR.n843 VDPWR.n831 14.2735
R9155 VDPWR.n85 VDPWR.n84 14.2735
R9156 VDPWR.n44 VDPWR.n43 14.2735
R9157 VDPWR.n1919 VDPWR.n1918 13.9299
R9158 VDPWR.n2264 VDPWR.n1075 13.8955
R9159 VDPWR.n2973 VDPWR.n929 13.8955
R9160 VDPWR.n651 VDPWR.n650 13.5534
R9161 VDPWR.n371 VDPWR.n370 13.5534
R9162 VDPWR.n113 VDPWR.n112 13.5534
R9163 VDPWR VDPWR.n571 13.4732
R9164 VDPWR VDPWR.n291 13.4732
R9165 VDPWR VDPWR.n33 13.4732
R9166 VDPWR.t984 VDPWR.t366 13.4281
R9167 VDPWR.t22 VDPWR.t501 13.4281
R9168 VDPWR.t358 VDPWR.t100 13.4281
R9169 VDPWR.t1049 VDPWR.t295 13.4281
R9170 VDPWR VDPWR.t1146 13.4281
R9171 VDPWR.n2767 VDPWR.n1003 12.9181
R9172 VDPWR.n175 VDPWR.n136 12.8005
R9173 VDPWR.n148 VDPWR.n136 12.8005
R9174 VDPWR.n148 VDPWR.n145 12.8005
R9175 VDPWR.n145 VDPWR.n144 12.8005
R9176 VDPWR.n1366 VDPWR.n1357 12.8005
R9177 VDPWR.n1699 VDPWR.n1690 12.8005
R9178 VDPWR.n1896 VDPWR.n1205 12.8005
R9179 VDPWR.n1621 VDPWR.n1620 12.8005
R9180 VDPWR.n2102 VDPWR.n2095 12.8005
R9181 VDPWR.n2565 VDPWR.n2556 12.8005
R9182 VDPWR.n3053 VDPWR.n3052 12.8005
R9183 VDPWR.n2837 VDPWR.n2836 12.3976
R9184 VDPWR.n3019 VDPWR.n3018 12.3912
R9185 VDPWR.n651 VDPWR.n539 12.0476
R9186 VDPWR.n371 VDPWR.n259 12.0476
R9187 VDPWR.n113 VDPWR.n1 12.0476
R9188 VDPWR.t16 VDPWR.t781 11.7496
R9189 VDPWR.t890 VDPWR.t250 11.7496
R9190 VDPWR.n814 VDPWR.n812 11.6993
R9191 VDPWR.n807 VDPWR.n800 11.6711
R9192 VDPWR.n587 VDPWR.n586 11.4366
R9193 VDPWR.n307 VDPWR.n306 11.4366
R9194 VDPWR.n49 VDPWR.n48 11.4366
R9195 VDPWR VDPWR.n535 11.4331
R9196 VDPWR VDPWR.n3175 11.4331
R9197 VDPWR.n389 VDPWR.n388 11.3235
R9198 VDPWR.n401 VDPWR.n400 11.3235
R9199 VDPWR.n2830 VDPWR.n2828 11.2946
R9200 VDPWR.n2669 VDPWR.n2668 11.2946
R9201 VDPWR.n643 VDPWR.n561 11.2937
R9202 VDPWR.n363 VDPWR.n281 11.2937
R9203 VDPWR.n105 VDPWR.n23 11.2937
R9204 VDPWR.n628 VDPWR.n627 11.2737
R9205 VDPWR.n348 VDPWR.n347 11.2737
R9206 VDPWR.n90 VDPWR.n89 11.2737
R9207 VDPWR.n2814 VDPWR.n2813 10.9719
R9208 VDPWR.n141 VDPWR.n140 10.9345
R9209 VDPWR.n2861 VDPWR.n2860 10.9181
R9210 VDPWR.n2052 VDPWR.n2051 10.912
R9211 VDPWR.n2744 VDPWR.n2743 10.5744
R9212 VDPWR.n2406 VDPWR.n2405 10.5417
R9213 VDPWR.n560 VDPWR.n559 10.1786
R9214 VDPWR.n280 VDPWR.n279 10.1786
R9215 VDPWR.n22 VDPWR.n21 10.1786
R9216 VDPWR.n2834 VDPWR.n980 10.1652
R9217 VDPWR.t979 VDPWR.t855 10.0712
R9218 VDPWR.t1010 VDPWR.t235 10.0712
R9219 VDPWR.t605 VDPWR.t759 10.0712
R9220 VDPWR.t208 VDPWR.t130 10.0712
R9221 VDPWR.n2107 VDPWR.n2106 9.8812
R9222 VDPWR.n2830 VDPWR.n980 9.78874
R9223 VDPWR.n2637 VDPWR.n2635 9.78874
R9224 VDPWR.n1519 VDPWR.n1518 9.73273
R9225 VDPWR.n1762 VDPWR.n1760 9.73273
R9226 VDPWR.n1840 VDPWR.n1839 9.73273
R9227 VDPWR.n1842 VDPWR.n1218 9.73273
R9228 VDPWR.n1846 VDPWR.n1218 9.73273
R9229 VDPWR.n1850 VDPWR.n1846 9.73273
R9230 VDPWR.n1850 VDPWR.n1849 9.73273
R9231 VDPWR.n2171 VDPWR.n1110 9.73273
R9232 VDPWR.n2216 VDPWR.n2215 9.73273
R9233 VDPWR.n2309 VDPWR.n2308 9.73273
R9234 VDPWR.n2908 VDPWR.n2907 9.73273
R9235 VDPWR.n2914 VDPWR.n2913 9.73273
R9236 VDPWR.n2917 VDPWR.n2914 9.73273
R9237 VDPWR.n2921 VDPWR.n948 9.73273
R9238 VDPWR.n2922 VDPWR.n2921 9.73273
R9239 VDPWR.n2923 VDPWR.n2922 9.73273
R9240 VDPWR.n2947 VDPWR.n2944 9.73273
R9241 VDPWR.n2951 VDPWR.n935 9.73273
R9242 VDPWR.n2480 VDPWR.n2479 9.73273
R9243 VDPWR.n2479 VDPWR.n2478 9.73273
R9244 VDPWR.n2220 VDPWR.n2219 9.71972
R9245 VDPWR.n2275 VDPWR.n2274 9.71972
R9246 VDPWR.n2173 VDPWR.n2172 9.71084
R9247 VDPWR.n2188 VDPWR.n2187 9.65296
R9248 VDPWR.n2243 VDPWR.n2242 9.65296
R9249 VDPWR.n2233 VDPWR.n2232 9.65296
R9250 VDPWR.n2230 VDPWR.n2200 9.65296
R9251 VDPWR.n2305 VDPWR.n2304 9.65296
R9252 VDPWR.n2302 VDPWR.n1036 9.65296
R9253 VDPWR.n2298 VDPWR.n2297 9.65296
R9254 VDPWR.n2281 VDPWR.n1059 9.65296
R9255 VDPWR.n600 VDPWR.n599 9.60526
R9256 VDPWR.n588 VDPWR.n587 9.60526
R9257 VDPWR.n553 VDPWR.n552 9.60526
R9258 VDPWR.n320 VDPWR.n319 9.60526
R9259 VDPWR.n308 VDPWR.n307 9.60526
R9260 VDPWR.n273 VDPWR.n272 9.60526
R9261 VDPWR.n62 VDPWR.n61 9.60526
R9262 VDPWR.n50 VDPWR.n49 9.60526
R9263 VDPWR.n15 VDPWR.n14 9.60526
R9264 VDPWR.n2742 VDPWR.n2739 9.6005
R9265 VDPWR.n2782 VDPWR.n999 9.56172
R9266 VDPWR.n2944 VDPWR.n937 9.52116
R9267 VDPWR.n1830 VDPWR.n1826 9.49016
R9268 VDPWR.n2285 VDPWR.n1057 9.35121
R9269 VDPWR.n250 VDPWR 9.30627
R9270 VDPWR.n590 VDPWR.n566 9.3005
R9271 VDPWR.n626 VDPWR.n625 9.3005
R9272 VDPWR.n623 VDPWR.n567 9.3005
R9273 VDPWR.n622 VDPWR.n620 9.3005
R9274 VDPWR.n619 VDPWR.n591 9.3005
R9275 VDPWR.n618 VDPWR.n617 9.3005
R9276 VDPWR.n616 VDPWR.n592 9.3005
R9277 VDPWR.n615 VDPWR.n614 9.3005
R9278 VDPWR.n613 VDPWR.n593 9.3005
R9279 VDPWR.n612 VDPWR.n611 9.3005
R9280 VDPWR.n610 VDPWR.n609 9.3005
R9281 VDPWR.n608 VDPWR.n594 9.3005
R9282 VDPWR.n607 VDPWR.n606 9.3005
R9283 VDPWR.n605 VDPWR.n604 9.3005
R9284 VDPWR.n603 VDPWR.n602 9.3005
R9285 VDPWR.n601 VDPWR.n597 9.3005
R9286 VDPWR.n573 VDPWR.n572 9.3005
R9287 VDPWR.n576 VDPWR.n568 9.3005
R9288 VDPWR.n585 VDPWR.n584 9.3005
R9289 VDPWR.n582 VDPWR.n569 9.3005
R9290 VDPWR.n581 VDPWR.n580 9.3005
R9291 VDPWR.n579 VDPWR.n564 9.3005
R9292 VDPWR.n630 VDPWR.n629 9.3005
R9293 VDPWR.n631 VDPWR.n563 9.3005
R9294 VDPWR.n636 VDPWR.n635 9.3005
R9295 VDPWR.n637 VDPWR.n562 9.3005
R9296 VDPWR.n640 VDPWR.n639 9.3005
R9297 VDPWR.n638 VDPWR.n539 9.3005
R9298 VDPWR.n652 VDPWR.n651 9.3005
R9299 VDPWR.n650 VDPWR.n538 9.3005
R9300 VDPWR.n649 VDPWR.n648 9.3005
R9301 VDPWR.n647 VDPWR.n646 9.3005
R9302 VDPWR.n645 VDPWR.n542 9.3005
R9303 VDPWR.n644 VDPWR.n547 9.3005
R9304 VDPWR.n559 VDPWR.n558 9.3005
R9305 VDPWR.n557 VDPWR.n556 9.3005
R9306 VDPWR.n554 VDPWR.n549 9.3005
R9307 VDPWR.n310 VDPWR.n286 9.3005
R9308 VDPWR.n346 VDPWR.n345 9.3005
R9309 VDPWR.n343 VDPWR.n287 9.3005
R9310 VDPWR.n342 VDPWR.n340 9.3005
R9311 VDPWR.n339 VDPWR.n311 9.3005
R9312 VDPWR.n338 VDPWR.n337 9.3005
R9313 VDPWR.n336 VDPWR.n312 9.3005
R9314 VDPWR.n335 VDPWR.n334 9.3005
R9315 VDPWR.n333 VDPWR.n313 9.3005
R9316 VDPWR.n332 VDPWR.n331 9.3005
R9317 VDPWR.n330 VDPWR.n329 9.3005
R9318 VDPWR.n328 VDPWR.n314 9.3005
R9319 VDPWR.n327 VDPWR.n326 9.3005
R9320 VDPWR.n325 VDPWR.n324 9.3005
R9321 VDPWR.n323 VDPWR.n322 9.3005
R9322 VDPWR.n321 VDPWR.n317 9.3005
R9323 VDPWR.n293 VDPWR.n292 9.3005
R9324 VDPWR.n296 VDPWR.n288 9.3005
R9325 VDPWR.n305 VDPWR.n304 9.3005
R9326 VDPWR.n302 VDPWR.n289 9.3005
R9327 VDPWR.n301 VDPWR.n300 9.3005
R9328 VDPWR.n299 VDPWR.n284 9.3005
R9329 VDPWR.n350 VDPWR.n349 9.3005
R9330 VDPWR.n351 VDPWR.n283 9.3005
R9331 VDPWR.n356 VDPWR.n355 9.3005
R9332 VDPWR.n357 VDPWR.n282 9.3005
R9333 VDPWR.n360 VDPWR.n359 9.3005
R9334 VDPWR.n358 VDPWR.n259 9.3005
R9335 VDPWR.n372 VDPWR.n371 9.3005
R9336 VDPWR.n370 VDPWR.n258 9.3005
R9337 VDPWR.n369 VDPWR.n368 9.3005
R9338 VDPWR.n367 VDPWR.n366 9.3005
R9339 VDPWR.n365 VDPWR.n262 9.3005
R9340 VDPWR.n364 VDPWR.n267 9.3005
R9341 VDPWR.n279 VDPWR.n278 9.3005
R9342 VDPWR.n277 VDPWR.n276 9.3005
R9343 VDPWR.n274 VDPWR.n269 9.3005
R9344 VDPWR.n143 VDPWR.n142 9.3005
R9345 VDPWR.n144 VDPWR.n138 9.3005
R9346 VDPWR.n145 VDPWR.n137 9.3005
R9347 VDPWR.n149 VDPWR.n148 9.3005
R9348 VDPWR.n150 VDPWR.n136 9.3005
R9349 VDPWR.n175 VDPWR.n174 9.3005
R9350 VDPWR.n173 VDPWR.n135 9.3005
R9351 VDPWR.n172 VDPWR.n171 9.3005
R9352 VDPWR.n170 VDPWR.n151 9.3005
R9353 VDPWR.n169 VDPWR.n168 9.3005
R9354 VDPWR.n167 VDPWR.n152 9.3005
R9355 VDPWR.n166 VDPWR.n165 9.3005
R9356 VDPWR.n164 VDPWR.n163 9.3005
R9357 VDPWR.n162 VDPWR.n153 9.3005
R9358 VDPWR.n161 VDPWR.n160 9.3005
R9359 VDPWR.n159 VDPWR.n158 9.3005
R9360 VDPWR.n157 VDPWR.n154 9.3005
R9361 VDPWR.n156 VDPWR.n155 9.3005
R9362 VDPWR.n129 VDPWR.n127 9.3005
R9363 VDPWR.n201 VDPWR.n200 9.3005
R9364 VDPWR.n199 VDPWR.n128 9.3005
R9365 VDPWR.n198 VDPWR.n197 9.3005
R9366 VDPWR.n196 VDPWR.n130 9.3005
R9367 VDPWR.n195 VDPWR.n194 9.3005
R9368 VDPWR.n193 VDPWR.n192 9.3005
R9369 VDPWR.n191 VDPWR.n131 9.3005
R9370 VDPWR.n190 VDPWR.n189 9.3005
R9371 VDPWR.n188 VDPWR.n187 9.3005
R9372 VDPWR.n186 VDPWR.n132 9.3005
R9373 VDPWR.n185 VDPWR.n184 9.3005
R9374 VDPWR.n183 VDPWR.n182 9.3005
R9375 VDPWR.n181 VDPWR.n133 9.3005
R9376 VDPWR.n180 VDPWR.n179 9.3005
R9377 VDPWR.n178 VDPWR.n177 9.3005
R9378 VDPWR.n252 VDPWR.n251 9.3005
R9379 VDPWR.n249 VDPWR.n120 9.3005
R9380 VDPWR.n248 VDPWR.n247 9.3005
R9381 VDPWR.n246 VDPWR.n121 9.3005
R9382 VDPWR.n245 VDPWR.n122 9.3005
R9383 VDPWR.n244 VDPWR.n243 9.3005
R9384 VDPWR.n242 VDPWR.n123 9.3005
R9385 VDPWR.n241 VDPWR.n240 9.3005
R9386 VDPWR.n239 VDPWR.n238 9.3005
R9387 VDPWR.n237 VDPWR.n124 9.3005
R9388 VDPWR.n236 VDPWR.n235 9.3005
R9389 VDPWR.n234 VDPWR.n233 9.3005
R9390 VDPWR.n232 VDPWR.n125 9.3005
R9391 VDPWR.n231 VDPWR.n230 9.3005
R9392 VDPWR.n229 VDPWR.n228 9.3005
R9393 VDPWR.n227 VDPWR.n126 9.3005
R9394 VDPWR.n226 VDPWR.n225 9.3005
R9395 VDPWR.n224 VDPWR.n223 9.3005
R9396 VDPWR.n222 VDPWR.n204 9.3005
R9397 VDPWR.n221 VDPWR.n220 9.3005
R9398 VDPWR.n219 VDPWR.n218 9.3005
R9399 VDPWR.n217 VDPWR.n205 9.3005
R9400 VDPWR.n216 VDPWR.n215 9.3005
R9401 VDPWR.n214 VDPWR.n213 9.3005
R9402 VDPWR.n212 VDPWR.n206 9.3005
R9403 VDPWR.n211 VDPWR.n210 9.3005
R9404 VDPWR.n209 VDPWR.n208 9.3005
R9405 VDPWR.n207 VDPWR.n119 9.3005
R9406 VDPWR.n1549 VDPWR.n1548 9.3005
R9407 VDPWR.n1550 VDPWR.n1549 9.3005
R9408 VDPWR.n1549 VDPWR.n1535 9.3005
R9409 VDPWR.n1369 VDPWR.n1368 9.3005
R9410 VDPWR.n1376 VDPWR.n1375 9.3005
R9411 VDPWR.n1378 VDPWR.n1348 9.3005
R9412 VDPWR.n1380 VDPWR.n1379 9.3005
R9413 VDPWR.n1389 VDPWR.n1388 9.3005
R9414 VDPWR.n1390 VDPWR.n1342 9.3005
R9415 VDPWR.n1393 VDPWR.n1392 9.3005
R9416 VDPWR.n1394 VDPWR.n1341 9.3005
R9417 VDPWR.n1396 VDPWR.n1395 9.3005
R9418 VDPWR.n1398 VDPWR.n1340 9.3005
R9419 VDPWR.n1400 VDPWR.n1399 9.3005
R9420 VDPWR.n1402 VDPWR.n1401 9.3005
R9421 VDPWR.n1404 VDPWR.n1338 9.3005
R9422 VDPWR.n1407 VDPWR.n1406 9.3005
R9423 VDPWR.n1408 VDPWR.n1337 9.3005
R9424 VDPWR.n1410 VDPWR.n1409 9.3005
R9425 VDPWR.n1412 VDPWR.n1335 9.3005
R9426 VDPWR.n1415 VDPWR.n1414 9.3005
R9427 VDPWR.n1413 VDPWR.n1329 9.3005
R9428 VDPWR.n1428 VDPWR.n1427 9.3005
R9429 VDPWR.n1432 VDPWR.n1431 9.3005
R9430 VDPWR.n1436 VDPWR.n1435 9.3005
R9431 VDPWR.n1438 VDPWR.n1437 9.3005
R9432 VDPWR.n1439 VDPWR.n1322 9.3005
R9433 VDPWR.n1442 VDPWR.n1441 9.3005
R9434 VDPWR.n1443 VDPWR.n1321 9.3005
R9435 VDPWR.n1445 VDPWR.n1444 9.3005
R9436 VDPWR.n1447 VDPWR.n1446 9.3005
R9437 VDPWR.n1451 VDPWR.n1314 9.3005
R9438 VDPWR.n1461 VDPWR.n1460 9.3005
R9439 VDPWR.n1462 VDPWR.n1313 9.3005
R9440 VDPWR.n1464 VDPWR.n1463 9.3005
R9441 VDPWR.n1465 VDPWR 9.3005
R9442 VDPWR.n1467 VDPWR.n1466 9.3005
R9443 VDPWR.n1469 VDPWR.n1468 9.3005
R9444 VDPWR.n1470 VDPWR.n1310 9.3005
R9445 VDPWR.n1472 VDPWR.n1471 9.3005
R9446 VDPWR.n1474 VDPWR.n1473 9.3005
R9447 VDPWR.n1475 VDPWR.n1308 9.3005
R9448 VDPWR.n1477 VDPWR.n1476 9.3005
R9449 VDPWR.n1478 VDPWR.n1307 9.3005
R9450 VDPWR.n1480 VDPWR.n1479 9.3005
R9451 VDPWR.n1487 VDPWR.n1486 9.3005
R9452 VDPWR.n1485 VDPWR.n1484 9.3005
R9453 VDPWR.n1481 VDPWR.n1298 9.3005
R9454 VDPWR.n1496 VDPWR.n1297 9.3005
R9455 VDPWR.n1498 VDPWR.n1497 9.3005
R9456 VDPWR.n1500 VDPWR.n1499 9.3005
R9457 VDPWR.n1502 VDPWR.n1501 9.3005
R9458 VDPWR.n1504 VDPWR.n1295 9.3005
R9459 VDPWR.n1508 VDPWR.n1507 9.3005
R9460 VDPWR.n1509 VDPWR.n1294 9.3005
R9461 VDPWR.n1511 VDPWR.n1510 9.3005
R9462 VDPWR.n1512 VDPWR.n1293 9.3005
R9463 VDPWR.n1514 VDPWR.n1513 9.3005
R9464 VDPWR.n1516 VDPWR.n1515 9.3005
R9465 VDPWR.n1518 VDPWR.n1517 9.3005
R9466 VDPWR.n1519 VDPWR.n1289 9.3005
R9467 VDPWR.n1577 VDPWR.n1576 9.3005
R9468 VDPWR.n1575 VDPWR.n1574 9.3005
R9469 VDPWR.n1573 VDPWR.n1572 9.3005
R9470 VDPWR.n1571 VDPWR.n1523 9.3005
R9471 VDPWR.n1570 VDPWR.n1569 9.3005
R9472 VDPWR.n1568 VDPWR.n1567 9.3005
R9473 VDPWR.n1566 VDPWR.n1525 9.3005
R9474 VDPWR.n1565 VDPWR.n1564 9.3005
R9475 VDPWR.n1563 VDPWR.n1526 9.3005
R9476 VDPWR.n1562 VDPWR.n1561 9.3005
R9477 VDPWR.n1560 VDPWR.n1527 9.3005
R9478 VDPWR.n1559 VDPWR.n1558 9.3005
R9479 VDPWR.n1537 VDPWR.n1529 9.3005
R9480 VDPWR.n1897 VDPWR.n1896 9.3005
R9481 VDPWR.n1896 VDPWR.n1198 9.3005
R9482 VDPWR.n1896 VDPWR.n1892 9.3005
R9483 VDPWR.n1702 VDPWR.n1701 9.3005
R9484 VDPWR.n1704 VDPWR.n1703 9.3005
R9485 VDPWR.n1709 VDPWR.n1708 9.3005
R9486 VDPWR.n1707 VDPWR.n1706 9.3005
R9487 VDPWR.n1719 VDPWR.n1718 9.3005
R9488 VDPWR.n1720 VDPWR.n1278 9.3005
R9489 VDPWR.n1723 VDPWR.n1722 9.3005
R9490 VDPWR.n1724 VDPWR.n1277 9.3005
R9491 VDPWR.n1726 VDPWR.n1725 9.3005
R9492 VDPWR.n1728 VDPWR.n1276 9.3005
R9493 VDPWR.n1730 VDPWR.n1729 9.3005
R9494 VDPWR.n1732 VDPWR.n1731 9.3005
R9495 VDPWR.n1734 VDPWR.n1274 9.3005
R9496 VDPWR.n1737 VDPWR.n1736 9.3005
R9497 VDPWR.n1738 VDPWR.n1273 9.3005
R9498 VDPWR.n1740 VDPWR.n1739 9.3005
R9499 VDPWR.n1742 VDPWR.n1271 9.3005
R9500 VDPWR.n1746 VDPWR.n1745 9.3005
R9501 VDPWR.n1744 VDPWR.n1264 9.3005
R9502 VDPWR.n1758 VDPWR.n1263 9.3005
R9503 VDPWR.n1760 VDPWR.n1759 9.3005
R9504 VDPWR.n1763 VDPWR.n1762 9.3005
R9505 VDPWR.n1768 VDPWR.n1256 9.3005
R9506 VDPWR.n1772 VDPWR.n1771 9.3005
R9507 VDPWR.n1773 VDPWR.n1255 9.3005
R9508 VDPWR.n1775 VDPWR.n1774 9.3005
R9509 VDPWR.n1777 VDPWR.n1250 9.3005
R9510 VDPWR.n1779 VDPWR.n1778 9.3005
R9511 VDPWR.n1242 VDPWR.n1241 9.3005
R9512 VDPWR.n1789 VDPWR.n1788 9.3005
R9513 VDPWR.n1790 VDPWR.n1240 9.3005
R9514 VDPWR.n1793 VDPWR.n1792 9.3005
R9515 VDPWR.n1797 VDPWR.n1238 9.3005
R9516 VDPWR.n1800 VDPWR.n1799 9.3005
R9517 VDPWR.n1802 VDPWR.n1801 9.3005
R9518 VDPWR.n1803 VDPWR.n1236 9.3005
R9519 VDPWR.n1806 VDPWR.n1805 9.3005
R9520 VDPWR.n1807 VDPWR.n1235 9.3005
R9521 VDPWR.n1809 VDPWR.n1808 9.3005
R9522 VDPWR.n1815 VDPWR.n1814 9.3005
R9523 VDPWR.n1813 VDPWR.n1812 9.3005
R9524 VDPWR.n1225 VDPWR.n1224 9.3005
R9525 VDPWR.n1825 VDPWR.n1824 9.3005
R9526 VDPWR.n1831 VDPWR.n1830 9.3005
R9527 VDPWR.n1837 VDPWR.n1836 9.3005
R9528 VDPWR.n1839 VDPWR.n1838 9.3005
R9529 VDPWR.n1840 VDPWR.n1219 9.3005
R9530 VDPWR.n1843 VDPWR.n1842 9.3005
R9531 VDPWR.n1844 VDPWR.n1218 9.3005
R9532 VDPWR.n1846 VDPWR.n1845 9.3005
R9533 VDPWR.n1851 VDPWR.n1850 9.3005
R9534 VDPWR.n1849 VDPWR.n1214 9.3005
R9535 VDPWR.n1865 VDPWR.n1864 9.3005
R9536 VDPWR.n1867 VDPWR.n1866 9.3005
R9537 VDPWR.n1868 VDPWR.n1211 9.3005
R9538 VDPWR.n1870 VDPWR.n1869 9.3005
R9539 VDPWR.n1872 VDPWR.n1210 9.3005
R9540 VDPWR.n1878 VDPWR.n1877 9.3005
R9541 VDPWR.n1879 VDPWR.n1209 9.3005
R9542 VDPWR.n1881 VDPWR.n1880 9.3005
R9543 VDPWR.n1883 VDPWR.n1882 9.3005
R9544 VDPWR.n1885 VDPWR.n1205 9.3005
R9545 VDPWR.n1948 VDPWR.n1947 9.3005
R9546 VDPWR.n1949 VDPWR.n1948 9.3005
R9547 VDPWR.n1948 VDPWR.n1934 9.3005
R9548 VDPWR.n1608 VDPWR.n1603 9.3005
R9549 VDPWR.n1607 VDPWR.n1601 9.3005
R9550 VDPWR.n1667 VDPWR.n1666 9.3005
R9551 VDPWR.n1665 VDPWR.n1664 9.3005
R9552 VDPWR.n1656 VDPWR.n1655 9.3005
R9553 VDPWR.n1654 VDPWR.n1626 9.3005
R9554 VDPWR.n1653 VDPWR.n1652 9.3005
R9555 VDPWR.n1651 VDPWR.n1650 9.3005
R9556 VDPWR.n1649 VDPWR.n1648 9.3005
R9557 VDPWR.n1647 VDPWR.n1646 9.3005
R9558 VDPWR.n1645 VDPWR.n1629 9.3005
R9559 VDPWR.n1643 VDPWR.n1642 9.3005
R9560 VDPWR.n1641 VDPWR.n1640 9.3005
R9561 VDPWR.n1638 VDPWR.n1631 9.3005
R9562 VDPWR.n1637 VDPWR.n1636 9.3005
R9563 VDPWR.n1635 VDPWR.n1634 9.3005
R9564 VDPWR.n1632 VDPWR.n1121 9.3005
R9565 VDPWR.n1125 VDPWR.n1122 9.3005
R9566 VDPWR.n2061 VDPWR.n2060 9.3005
R9567 VDPWR.n2058 VDPWR.n2057 9.3005
R9568 VDPWR.n2056 VDPWR.n1126 9.3005
R9569 VDPWR.n2054 VDPWR.n2053 9.3005
R9570 VDPWR.n2046 VDPWR.n1129 9.3005
R9571 VDPWR.n2045 VDPWR.n2044 9.3005
R9572 VDPWR.n2043 VDPWR.n1131 9.3005
R9573 VDPWR.n2042 VDPWR.n2041 9.3005
R9574 VDPWR.n2040 VDPWR.n2039 9.3005
R9575 VDPWR.n1142 VDPWR.n1135 9.3005
R9576 VDPWR.n1148 VDPWR.n1147 9.3005
R9577 VDPWR.n1149 VDPWR.n1140 9.3005
R9578 VDPWR.n2030 VDPWR.n2029 9.3005
R9579 VDPWR.n2028 VDPWR.n1141 9.3005
R9580 VDPWR.n2026 VDPWR.n2025 9.3005
R9581 VDPWR.n2024 VDPWR.n1151 9.3005
R9582 VDPWR.n2023 VDPWR.n2022 9.3005
R9583 VDPWR.n2021 VDPWR.n1152 9.3005
R9584 VDPWR.n2020 VDPWR.n2019 9.3005
R9585 VDPWR.n2018 VDPWR.n2017 9.3005
R9586 VDPWR.n2016 VDPWR.n2015 9.3005
R9587 VDPWR.n2014 VDPWR.n2013 9.3005
R9588 VDPWR.n2012 VDPWR.n1157 9.3005
R9589 VDPWR.n2011 VDPWR.n2010 9.3005
R9590 VDPWR.n1169 VDPWR.n1168 9.3005
R9591 VDPWR.n1176 VDPWR.n1175 9.3005
R9592 VDPWR.n1178 VDPWR.n1165 9.3005
R9593 VDPWR.n2002 VDPWR.n2001 9.3005
R9594 VDPWR.n2000 VDPWR.n1999 9.3005
R9595 VDPWR.n1998 VDPWR.n1997 9.3005
R9596 VDPWR.n1996 VDPWR.n1180 9.3005
R9597 VDPWR.n1994 VDPWR.n1993 9.3005
R9598 VDPWR.n1992 VDPWR.n1182 9.3005
R9599 VDPWR.n1991 VDPWR.n1990 9.3005
R9600 VDPWR.n1988 VDPWR.n1183 9.3005
R9601 VDPWR.n1986 VDPWR.n1985 9.3005
R9602 VDPWR.n1984 VDPWR.n1983 9.3005
R9603 VDPWR.n1982 VDPWR.n1185 9.3005
R9604 VDPWR.n1980 VDPWR 9.3005
R9605 VDPWR.n1912 VDPWR.n1186 9.3005
R9606 VDPWR.n1920 VDPWR.n1914 9.3005
R9607 VDPWR.n1970 VDPWR.n1969 9.3005
R9608 VDPWR.n1966 VDPWR.n1965 9.3005
R9609 VDPWR.n1963 VDPWR.n1922 9.3005
R9610 VDPWR.n1962 VDPWR.n1961 9.3005
R9611 VDPWR.n1959 VDPWR.n1923 9.3005
R9612 VDPWR.n1958 VDPWR.n1957 9.3005
R9613 VDPWR.n1936 VDPWR.n1929 9.3005
R9614 VDPWR.n1086 VDPWR.n1075 9.3005
R9615 VDPWR.n1084 VDPWR.n1075 9.3005
R9616 VDPWR.n1077 VDPWR.n1075 9.3005
R9617 VDPWR.n2106 VDPWR.n2105 9.3005
R9618 VDPWR.n2109 VDPWR.n2108 9.3005
R9619 VDPWR.n2115 VDPWR.n2114 9.3005
R9620 VDPWR.n2119 VDPWR.n2118 9.3005
R9621 VDPWR.n2120 VDPWR.n2084 9.3005
R9622 VDPWR.n2129 VDPWR.n2128 9.3005
R9623 VDPWR.n2130 VDPWR.n2083 9.3005
R9624 VDPWR.n2132 VDPWR.n2131 9.3005
R9625 VDPWR.n2134 VDPWR.n2133 9.3005
R9626 VDPWR.n2135 VDPWR.n2081 9.3005
R9627 VDPWR.n2138 VDPWR.n2137 9.3005
R9628 VDPWR.n2140 VDPWR.n2139 9.3005
R9629 VDPWR.n2143 VDPWR.n2142 9.3005
R9630 VDPWR.n2145 VDPWR.n2144 9.3005
R9631 VDPWR.n2146 VDPWR.n2078 9.3005
R9632 VDPWR.n2148 VDPWR.n2147 9.3005
R9633 VDPWR.n2150 VDPWR.n2149 9.3005
R9634 VDPWR.n2152 VDPWR.n2151 9.3005
R9635 VDPWR.n1113 VDPWR.n1112 9.3005
R9636 VDPWR.n2165 VDPWR.n2164 9.3005
R9637 VDPWR.n2168 VDPWR.n2167 9.3005
R9638 VDPWR.n2169 VDPWR.n1110 9.3005
R9639 VDPWR.n2171 VDPWR.n2170 9.3005
R9640 VDPWR.n2174 VDPWR.n2173 9.3005
R9641 VDPWR.n2176 VDPWR.n2175 9.3005
R9642 VDPWR.n2181 VDPWR.n2180 9.3005
R9643 VDPWR.n2182 VDPWR.n1103 9.3005
R9644 VDPWR.n2184 VDPWR.n2183 9.3005
R9645 VDPWR.n2187 VDPWR.n1101 9.3005
R9646 VDPWR.n2189 VDPWR.n2188 9.3005
R9647 VDPWR.n2191 VDPWR.n2190 9.3005
R9648 VDPWR.n2193 VDPWR.n1096 9.3005
R9649 VDPWR.n2244 VDPWR.n2243 9.3005
R9650 VDPWR.n2242 VDPWR.n2241 9.3005
R9651 VDPWR.n2234 VDPWR.n2233 9.3005
R9652 VDPWR.n2232 VDPWR.n2198 9.3005
R9653 VDPWR.n2230 VDPWR.n2229 9.3005
R9654 VDPWR.n2228 VDPWR.n2200 9.3005
R9655 VDPWR.n2227 VDPWR.n2226 9.3005
R9656 VDPWR.n2225 VDPWR.n2224 9.3005
R9657 VDPWR.n2223 VDPWR.n2222 9.3005
R9658 VDPWR.n2220 VDPWR.n2206 9.3005
R9659 VDPWR.n2219 VDPWR.n2218 9.3005
R9660 VDPWR.n2217 VDPWR.n2216 9.3005
R9661 VDPWR.n2215 VDPWR.n2214 9.3005
R9662 VDPWR.n2213 VDPWR.n2212 9.3005
R9663 VDPWR.n2326 VDPWR.n2325 9.3005
R9664 VDPWR.n2324 VDPWR.n2323 9.3005
R9665 VDPWR.n1025 VDPWR.n1020 9.3005
R9666 VDPWR.n2318 VDPWR.n2317 9.3005
R9667 VDPWR.n2315 VDPWR.n2314 9.3005
R9668 VDPWR.n2313 VDPWR.n1026 9.3005
R9669 VDPWR.n2312 VDPWR.n2311 9.3005
R9670 VDPWR.n2309 VDPWR.n1027 9.3005
R9671 VDPWR.n2308 VDPWR.n2307 9.3005
R9672 VDPWR.n2306 VDPWR.n2305 9.3005
R9673 VDPWR.n2304 VDPWR.n1032 9.3005
R9674 VDPWR.n2302 VDPWR.n2301 9.3005
R9675 VDPWR.n2300 VDPWR.n1036 9.3005
R9676 VDPWR.n2299 VDPWR.n2298 9.3005
R9677 VDPWR.n2297 VDPWR.n2296 9.3005
R9678 VDPWR.n1053 VDPWR.n1052 9.3005
R9679 VDPWR.n1056 VDPWR.n1055 9.3005
R9680 VDPWR.n2286 VDPWR.n2285 9.3005
R9681 VDPWR.n2283 VDPWR.n1049 9.3005
R9682 VDPWR.n2281 VDPWR.n2280 9.3005
R9683 VDPWR.n2279 VDPWR.n1059 9.3005
R9684 VDPWR.n2278 VDPWR.n2277 9.3005
R9685 VDPWR.n2275 VDPWR.n1060 9.3005
R9686 VDPWR.n2274 VDPWR.n2273 9.3005
R9687 VDPWR.n2272 VDPWR.n2271 9.3005
R9688 VDPWR.n2270 VDPWR.n2269 9.3005
R9689 VDPWR.n2268 VDPWR.n2267 9.3005
R9690 VDPWR.n2266 VDPWR.n1067 9.3005
R9691 VDPWR.n2264 VDPWR.n2263 9.3005
R9692 VDPWR.n2974 VDPWR.n2973 9.3005
R9693 VDPWR.n2973 VDPWR.n928 9.3005
R9694 VDPWR.n2973 VDPWR.n2969 9.3005
R9695 VDPWR.n2738 VDPWR.n2737 9.3005
R9696 VDPWR.n2745 VDPWR.n2744 9.3005
R9697 VDPWR.n2750 VDPWR.n2749 9.3005
R9698 VDPWR.n2749 VDPWR.n2748 9.3005
R9699 VDPWR.n2760 VDPWR.n2759 9.3005
R9700 VDPWR.n2761 VDPWR.n1004 9.3005
R9701 VDPWR.n2764 VDPWR.n2763 9.3005
R9702 VDPWR.n2765 VDPWR.n1003 9.3005
R9703 VDPWR.n2767 VDPWR.n2766 9.3005
R9704 VDPWR.n2771 VDPWR.n1002 9.3005
R9705 VDPWR.n2775 VDPWR.n2774 9.3005
R9706 VDPWR.n2778 VDPWR.n2777 9.3005
R9707 VDPWR.n2780 VDPWR.n2779 9.3005
R9708 VDPWR.n2786 VDPWR.n2785 9.3005
R9709 VDPWR.n2788 VDPWR.n2787 9.3005
R9710 VDPWR.n2789 VDPWR.n993 9.3005
R9711 VDPWR.n2797 VDPWR.n2796 9.3005
R9712 VDPWR.n2795 VDPWR.n985 9.3005
R9713 VDPWR.n2809 VDPWR.n984 9.3005
R9714 VDPWR.n2813 VDPWR.n2810 9.3005
R9715 VDPWR.n2818 VDPWR.n2817 9.3005
R9716 VDPWR.n2819 VDPWR.n982 9.3005
R9717 VDPWR.n2821 VDPWR.n2820 9.3005
R9718 VDPWR.n2825 VDPWR.n2824 9.3005
R9719 VDPWR.n2826 VDPWR.n981 9.3005
R9720 VDPWR.n2828 VDPWR.n2827 9.3005
R9721 VDPWR.n2831 VDPWR.n2830 9.3005
R9722 VDPWR.n2832 VDPWR.n980 9.3005
R9723 VDPWR.n2834 VDPWR.n2833 9.3005
R9724 VDPWR.n2838 VDPWR.n2837 9.3005
R9725 VDPWR.n2839 VDPWR.n969 9.3005
R9726 VDPWR.n2850 VDPWR.n2849 9.3005
R9727 VDPWR.n2855 VDPWR.n2854 9.3005
R9728 VDPWR.n2856 VDPWR.n967 9.3005
R9729 VDPWR.n2858 VDPWR.n2857 9.3005
R9730 VDPWR.n2860 VDPWR.n966 9.3005
R9731 VDPWR.n2862 VDPWR.n2861 9.3005
R9732 VDPWR.n2863 VDPWR.n965 9.3005
R9733 VDPWR.n2865 VDPWR.n2864 9.3005
R9734 VDPWR.n2867 VDPWR.n963 9.3005
R9735 VDPWR.n2869 VDPWR.n2868 9.3005
R9736 VDPWR.n2871 VDPWR.n2870 9.3005
R9737 VDPWR.n2876 VDPWR.n2875 9.3005
R9738 VDPWR.n2883 VDPWR.n2882 9.3005
R9739 VDPWR.n2886 VDPWR.n959 9.3005
R9740 VDPWR.n2892 VDPWR.n2891 9.3005
R9741 VDPWR.n2888 VDPWR.n955 9.3005
R9742 VDPWR.n2900 VDPWR.n954 9.3005
R9743 VDPWR.n2902 VDPWR.n2901 9.3005
R9744 VDPWR.n2905 VDPWR.n2904 9.3005
R9745 VDPWR.n2907 VDPWR.n2906 9.3005
R9746 VDPWR.n2908 VDPWR.n951 9.3005
R9747 VDPWR.n2911 VDPWR.n2910 9.3005
R9748 VDPWR.n2913 VDPWR.n2912 9.3005
R9749 VDPWR.n2914 VDPWR.n949 9.3005
R9750 VDPWR.n2918 VDPWR.n2917 9.3005
R9751 VDPWR.n2919 VDPWR.n948 9.3005
R9752 VDPWR.n2921 VDPWR.n2920 9.3005
R9753 VDPWR.n2922 VDPWR.n947 9.3005
R9754 VDPWR.n2924 VDPWR.n2923 9.3005
R9755 VDPWR.n2937 VDPWR.n2936 9.3005
R9756 VDPWR.n2939 VDPWR.n938 9.3005
R9757 VDPWR.n2942 VDPWR.n2941 9.3005
R9758 VDPWR.n2944 VDPWR.n2943 9.3005
R9759 VDPWR.n2948 VDPWR.n2947 9.3005
R9760 VDPWR.n2949 VDPWR.n935 9.3005
R9761 VDPWR.n2951 VDPWR.n2950 9.3005
R9762 VDPWR.n2954 VDPWR.n2953 9.3005
R9763 VDPWR.n2955 VDPWR.n934 9.3005
R9764 VDPWR.n2957 VDPWR.n2956 9.3005
R9765 VDPWR.n2958 VDPWR.n933 9.3005
R9766 VDPWR.n2961 VDPWR.n2960 9.3005
R9767 VDPWR.n2962 VDPWR.n929 9.3005
R9768 VDPWR.n3001 VDPWR.n3000 9.3005
R9769 VDPWR.n3000 VDPWR.n2996 9.3005
R9770 VDPWR.n3000 VDPWR.n2993 9.3005
R9771 VDPWR.n2568 VDPWR.n2567 9.3005
R9772 VDPWR.n2566 VDPWR.n2548 9.3005
R9773 VDPWR.n2578 VDPWR.n2577 9.3005
R9774 VDPWR.n2715 VDPWR.n2714 9.3005
R9775 VDPWR.n2713 VDPWR.n2544 9.3005
R9776 VDPWR.n2712 VDPWR.n2711 9.3005
R9777 VDPWR.n2710 VDPWR.n2579 9.3005
R9778 VDPWR.n2709 VDPWR.n2708 9.3005
R9779 VDPWR.n2706 VDPWR.n2580 9.3005
R9780 VDPWR.n2705 VDPWR.n2704 9.3005
R9781 VDPWR.n2703 VDPWR.n2583 9.3005
R9782 VDPWR.n2702 VDPWR.n2701 9.3005
R9783 VDPWR.n2700 VDPWR.n2584 9.3005
R9784 VDPWR.n2699 VDPWR.n2698 9.3005
R9785 VDPWR.n2697 VDPWR.n2587 9.3005
R9786 VDPWR.n2594 VDPWR.n2588 9.3005
R9787 VDPWR.n2687 VDPWR.n2602 9.3005
R9788 VDPWR.n2687 VDPWR.n2593 9.3005
R9789 VDPWR.n2688 VDPWR.n2687 9.3005
R9790 VDPWR.n2686 VDPWR.n2604 9.3005
R9791 VDPWR.n2683 VDPWR.n2682 9.3005
R9792 VDPWR.n2681 VDPWR.n2605 9.3005
R9793 VDPWR.n2680 VDPWR.n2679 9.3005
R9794 VDPWR.n2678 VDPWR.n2606 9.3005
R9795 VDPWR.n2675 VDPWR.n2674 9.3005
R9796 VDPWR.n2673 VDPWR.n2610 9.3005
R9797 VDPWR.n2672 VDPWR.n2671 9.3005
R9798 VDPWR.n2670 VDPWR.n2611 9.3005
R9799 VDPWR.n2668 VDPWR.n2667 9.3005
R9800 VDPWR.n2614 VDPWR.n2613 9.3005
R9801 VDPWR.n2651 VDPWR.n2649 9.3005
R9802 VDPWR.n2656 VDPWR.n2655 9.3005
R9803 VDPWR.n2658 VDPWR.n2657 9.3005
R9804 VDPWR.n2657 VDPWR.n2646 9.3005
R9805 VDPWR.n2645 VDPWR.n2620 9.3005
R9806 VDPWR.n2644 VDPWR.n2643 9.3005
R9807 VDPWR.n2641 VDPWR.n2640 9.3005
R9808 VDPWR.n2639 VDPWR.n2621 9.3005
R9809 VDPWR.n2638 VDPWR.n2637 9.3005
R9810 VDPWR.n2635 VDPWR.n2622 9.3005
R9811 VDPWR.n2632 VDPWR.n2631 9.3005
R9812 VDPWR.n2630 VDPWR.n2629 9.3005
R9813 VDPWR.n3062 VDPWR.n3061 9.3005
R9814 VDPWR.n3060 VDPWR.n3059 9.3005
R9815 VDPWR.n885 VDPWR.n880 9.3005
R9816 VDPWR.n3054 VDPWR.n3053 9.3005
R9817 VDPWR.n3050 VDPWR.n3049 9.3005
R9818 VDPWR.n3048 VDPWR.n892 9.3005
R9819 VDPWR.n3047 VDPWR.n3046 9.3005
R9820 VDPWR.n3045 VDPWR.n895 9.3005
R9821 VDPWR.n3044 VDPWR.n3043 9.3005
R9822 VDPWR.n3042 VDPWR.n3041 9.3005
R9823 VDPWR.n3040 VDPWR.n898 9.3005
R9824 VDPWR.n3039 VDPWR.n3038 9.3005
R9825 VDPWR.n911 VDPWR.n910 9.3005
R9826 VDPWR.n912 VDPWR.n907 9.3005
R9827 VDPWR.n3028 VDPWR.n3027 9.3005
R9828 VDPWR.n3025 VDPWR.n908 9.3005
R9829 VDPWR.n3024 VDPWR.n914 9.3005
R9830 VDPWR.n3023 VDPWR.n3022 9.3005
R9831 VDPWR.n3021 VDPWR.n916 9.3005
R9832 VDPWR.n3020 VDPWR.n3019 9.3005
R9833 VDPWR.n3018 VDPWR.n3017 9.3005
R9834 VDPWR.n3016 VDPWR.n3015 9.3005
R9835 VDPWR.n3013 VDPWR.n918 9.3005
R9836 VDPWR.n3012 VDPWR.n3011 9.3005
R9837 VDPWR.n3010 VDPWR.n920 9.3005
R9838 VDPWR.n2988 VDPWR.n921 9.3005
R9839 VDPWR.n843 VDPWR.n842 9.3005
R9840 VDPWR.n843 VDPWR.n835 9.3005
R9841 VDPWR.n844 VDPWR.n843 9.3005
R9842 VDPWR.n2380 VDPWR.n2379 9.3005
R9843 VDPWR.n2382 VDPWR.n2381 9.3005
R9844 VDPWR.n2383 VDPWR.n2369 9.3005
R9845 VDPWR.n2385 VDPWR.n2384 9.3005
R9846 VDPWR.n2386 VDPWR.n2367 9.3005
R9847 VDPWR.n2388 VDPWR.n2387 9.3005
R9848 VDPWR.n2397 VDPWR.n2396 9.3005
R9849 VDPWR.n2400 VDPWR.n2358 9.3005
R9850 VDPWR.n2402 VDPWR.n2401 9.3005
R9851 VDPWR.n2404 VDPWR.n2403 9.3005
R9852 VDPWR.n2405 VDPWR.n2354 9.3005
R9853 VDPWR.n2407 VDPWR.n2406 9.3005
R9854 VDPWR.n2408 VDPWR.n2353 9.3005
R9855 VDPWR.n2410 VDPWR.n2409 9.3005
R9856 VDPWR.n2413 VDPWR.n2412 9.3005
R9857 VDPWR.n2414 VDPWR.n2351 9.3005
R9858 VDPWR.n2416 VDPWR.n2415 9.3005
R9859 VDPWR.n2418 VDPWR.n2350 9.3005
R9860 VDPWR.n2423 VDPWR.n2422 9.3005
R9861 VDPWR.n2425 VDPWR.n2349 9.3005
R9862 VDPWR.n2430 VDPWR.n2429 9.3005
R9863 VDPWR.n2532 VDPWR.n2531 9.3005
R9864 VDPWR.n2530 VDPWR.n2529 9.3005
R9865 VDPWR.n2528 VDPWR.n2433 9.3005
R9866 VDPWR.n2527 VDPWR.n2526 9.3005
R9867 VDPWR.n2524 VDPWR.n2523 9.3005
R9868 VDPWR.n2522 VDPWR.n2521 9.3005
R9869 VDPWR.n2520 VDPWR.n2435 9.3005
R9870 VDPWR.n2518 VDPWR.n2517 9.3005
R9871 VDPWR.n2516 VDPWR.n2515 9.3005
R9872 VDPWR.n2514 VDPWR.n2439 9.3005
R9873 VDPWR.n2513 VDPWR.n2440 9.3005
R9874 VDPWR.n2512 VDPWR.n2511 9.3005
R9875 VDPWR.n2443 VDPWR.n2442 9.3005
R9876 VDPWR.n2451 VDPWR.n2448 9.3005
R9877 VDPWR.n2493 VDPWR.n2492 9.3005
R9878 VDPWR.n2490 VDPWR.n2489 9.3005
R9879 VDPWR.n2488 VDPWR.n2454 9.3005
R9880 VDPWR.n2487 VDPWR.n2486 9.3005
R9881 VDPWR.n2484 VDPWR.n2455 9.3005
R9882 VDPWR.n2483 VDPWR.n2482 9.3005
R9883 VDPWR.n2481 VDPWR.n2480 9.3005
R9884 VDPWR.n2479 VDPWR.n2457 9.3005
R9885 VDPWR.n2478 VDPWR.n2477 9.3005
R9886 VDPWR.n2469 VDPWR.n2468 9.3005
R9887 VDPWR.n2463 VDPWR.n787 9.3005
R9888 VDPWR.n3098 VDPWR.n3097 9.3005
R9889 VDPWR.n3096 VDPWR.n790 9.3005
R9890 VDPWR.n3095 VDPWR.n3094 9.3005
R9891 VDPWR.n3093 VDPWR.n3092 9.3005
R9892 VDPWR.n3089 VDPWR.n3088 9.3005
R9893 VDPWR.n3087 VDPWR.n793 9.3005
R9894 VDPWR.n3086 VDPWR.n3085 9.3005
R9895 VDPWR.n3084 VDPWR.n794 9.3005
R9896 VDPWR.n3083 VDPWR.n3082 9.3005
R9897 VDPWR.n3081 VDPWR.n3080 9.3005
R9898 VDPWR.n3079 VDPWR.n3078 9.3005
R9899 VDPWR.n3077 VDPWR.n800 9.3005
R9900 VDPWR.n808 VDPWR.n801 9.3005
R9901 VDPWR.n812 VDPWR.n811 9.3005
R9902 VDPWR.n866 VDPWR.n865 9.3005
R9903 VDPWR.n863 VDPWR.n862 9.3005
R9904 VDPWR.n861 VDPWR.n815 9.3005
R9905 VDPWR.n860 VDPWR.n859 9.3005
R9906 VDPWR.n858 VDPWR.n816 9.3005
R9907 VDPWR.n856 VDPWR.n855 9.3005
R9908 VDPWR.n853 VDPWR.n852 9.3005
R9909 VDPWR.n851 VDPWR.n850 9.3005
R9910 VDPWR.n849 VDPWR.n826 9.3005
R9911 VDPWR.n831 VDPWR.n827 9.3005
R9912 VDPWR.n52 VDPWR.n28 9.3005
R9913 VDPWR.n88 VDPWR.n87 9.3005
R9914 VDPWR.n85 VDPWR.n29 9.3005
R9915 VDPWR.n84 VDPWR.n82 9.3005
R9916 VDPWR.n81 VDPWR.n53 9.3005
R9917 VDPWR.n80 VDPWR.n79 9.3005
R9918 VDPWR.n78 VDPWR.n54 9.3005
R9919 VDPWR.n77 VDPWR.n76 9.3005
R9920 VDPWR.n75 VDPWR.n55 9.3005
R9921 VDPWR.n74 VDPWR.n73 9.3005
R9922 VDPWR.n72 VDPWR.n71 9.3005
R9923 VDPWR.n70 VDPWR.n56 9.3005
R9924 VDPWR.n69 VDPWR.n68 9.3005
R9925 VDPWR.n67 VDPWR.n66 9.3005
R9926 VDPWR.n65 VDPWR.n64 9.3005
R9927 VDPWR.n63 VDPWR.n59 9.3005
R9928 VDPWR.n35 VDPWR.n34 9.3005
R9929 VDPWR.n38 VDPWR.n30 9.3005
R9930 VDPWR.n47 VDPWR.n46 9.3005
R9931 VDPWR.n44 VDPWR.n31 9.3005
R9932 VDPWR.n43 VDPWR.n42 9.3005
R9933 VDPWR.n41 VDPWR.n26 9.3005
R9934 VDPWR.n92 VDPWR.n91 9.3005
R9935 VDPWR.n93 VDPWR.n25 9.3005
R9936 VDPWR.n98 VDPWR.n97 9.3005
R9937 VDPWR.n99 VDPWR.n24 9.3005
R9938 VDPWR.n102 VDPWR.n101 9.3005
R9939 VDPWR.n100 VDPWR.n1 9.3005
R9940 VDPWR.n114 VDPWR.n113 9.3005
R9941 VDPWR.n112 VDPWR.n0 9.3005
R9942 VDPWR.n111 VDPWR.n110 9.3005
R9943 VDPWR.n109 VDPWR.n108 9.3005
R9944 VDPWR.n107 VDPWR.n4 9.3005
R9945 VDPWR.n106 VDPWR.n9 9.3005
R9946 VDPWR.n21 VDPWR.n20 9.3005
R9947 VDPWR.n19 VDPWR.n18 9.3005
R9948 VDPWR.n16 VDPWR.n11 9.3005
R9949 VDPWR.n1520 VDPWR.n1519 9.09802
R9950 VDPWR.n2317 VDPWR.n2316 9.09802
R9951 VDPWR.n2311 VDPWR.n1029 9.09802
R9952 VDPWR.n2311 VDPWR.n2310 9.09802
R9953 VDPWR.n2923 VDPWR.n939 9.09802
R9954 VDPWR.n2941 VDPWR.n2940 9.09802
R9955 VDPWR.n2222 VDPWR.n2207 9.02345
R9956 VDPWR.n1052 VDPWR.n1051 9.02345
R9957 VDPWR.n2284 VDPWR.n2283 9.02345
R9958 VDPWR.n1841 VDPWR.n1840 8.99224
R9959 VDPWR.n823 VDPWR.n820 8.9761
R9960 VDPWR.n2907 VDPWR.n953 8.88645
R9961 VDPWR.n2788 VDPWR.n998 8.77764
R9962 VDPWR.n2222 VDPWR.n2221 8.60378
R9963 VDPWR.n2277 VDPWR.n2276 8.60378
R9964 VDPWR.n1431 VDPWR.n1428 8.44958
R9965 VDPWR.n1760 VDPWR.n1263 8.44958
R9966 VDPWR.n1825 VDPWR.n1224 8.44958
R9967 VDPWR.n2001 VDPWR.n1178 8.44958
R9968 VDPWR.n2058 VDPWR.n1126 8.44958
R9969 VDPWR.n2167 VDPWR.n1110 8.44958
R9970 VDPWR.t331 VDPWR.t775 8.39273
R9971 VDPWR.n2282 VDPWR.n2281 8.28902
R9972 VDPWR.n1872 VDPWR.n1871 8.28285
R9973 VDPWR.n2677 VDPWR.n2676 8.28285
R9974 VDPWR.n671 VDPWR.n657 8.23557
R9975 VDPWR.n428 VDPWR.n414 8.23557
R9976 VDPWR.n2791 VDPWR.n2790 8.04621
R9977 VDPWR.n2274 VDPWR.n1065 8.04017
R9978 VDPWR.n1766 VDPWR.n1257 7.98741
R9979 VDPWR.n2480 VDPWR 7.93438
R9980 VDPWR.n2678 VDPWR.n2677 7.90638
R9981 VDPWR.n2686 VDPWR.n2684 7.90638
R9982 VDPWR.n1518 VDPWR.n1516 7.75995
R9983 VDPWR.n2001 VDPWR.n2000 7.75995
R9984 VDPWR.n2215 VDPWR.n2212 7.75995
R9985 VDPWR.n2317 VDPWR.n1025 7.75995
R9986 VDPWR.n2271 VDPWR.n2270 7.75995
R9987 VDPWR.n2953 VDPWR.n2951 7.75995
R9988 VDPWR.n2484 VDPWR.n2483 7.75995
R9989 VDPWR.n2203 VDPWR.n2202 7.65952
R9990 VDPWR.n718 VDPWR.n717 7.54407
R9991 VDPWR.n702 VDPWR.n701 7.54407
R9992 VDPWR.n686 VDPWR.n685 7.54407
R9993 VDPWR.n670 VDPWR.n669 7.54407
R9994 VDPWR.n529 VDPWR.n528 7.54407
R9995 VDPWR.n513 VDPWR.n512 7.54407
R9996 VDPWR.n497 VDPWR.n496 7.54407
R9997 VDPWR.n481 VDPWR.n480 7.54407
R9998 VDPWR.n459 VDPWR.n458 7.54407
R9999 VDPWR.n443 VDPWR.n442 7.54407
R10000 VDPWR.n427 VDPWR.n426 7.54407
R10001 VDPWR.n3170 VDPWR.n3169 7.54407
R10002 VDPWR.n3132 VDPWR.n3131 7.54407
R10003 VDPWR.n465 VDPWR.n464 7.54307
R10004 VDPWR.n3164 VDPWR.n3163 7.54307
R10005 VDPWR.n3148 VDPWR.n3147 7.54307
R10006 VDPWR.n2910 VDPWR.n2909 7.51124
R10007 VDPWR.n2515 VDPWR.n2514 7.49704
R10008 VDPWR.n1108 VDPWR.n1105 7.28326
R10009 VDPWR.n1106 VDPWR.n1104 7.23528
R10010 VDPWR.n2017 VDPWR.n2016 7.21067
R10011 VDPWR.n2026 VDPWR.n1151 7.21067
R10012 VDPWR.n2142 VDPWR.n2140 7.21067
R10013 VDPWR.n2186 VDPWR.n2185 7.17134
R10014 VDPWR.n1502 VDPWR.n1296 7.12524
R10015 VDPWR.n537 VDPWR.n532 7.10511
R10016 VDPWR.n2231 VDPWR.n2230 7.03001
R10017 VDPWR.n546 VDPWR.n543 6.8005
R10018 VDPWR.n266 VDPWR.n263 6.8005
R10019 VDPWR.n8 VDPWR.n5 6.8005
R10020 VDPWR.n1871 VDPWR.n1870 6.77697
R10021 VDPWR.n1990 VDPWR.n1182 6.77697
R10022 VDPWR.n3051 VDPWR.n3050 6.77697
R10023 VDPWR.n858 VDPWR.n857 6.73838
R10024 VDPWR.t136 VDPWR.t6 6.71428
R10025 VDPWR.t918 VDPWR.t348 6.71428
R10026 VDPWR.t1015 VDPWR.t9 6.71428
R10027 VDPWR.t807 VDPWR.t805 6.71428
R10028 VDPWR.t229 VDPWR.t223 6.71428
R10029 VDPWR.n1431 VDPWR.n1327 6.66496
R10030 VDPWR.n1762 VDPWR.n1761 6.66496
R10031 VDPWR.n1826 VDPWR.n1825 6.66496
R10032 VDPWR.n1836 VDPWR.n1834 6.66496
R10033 VDPWR.n1127 VDPWR.n1126 6.66496
R10034 VDPWR.n2172 VDPWR.n2171 6.66496
R10035 VDPWR.n2478 VDPWR.n2459 6.66496
R10036 VDPWR.n1396 VDPWR.n1341 6.52104
R10037 VDPWR.n1726 VDPWR.n1277 6.52104
R10038 VDPWR.n2135 VDPWR.n2134 6.52104
R10039 VDPWR.n2041 VDPWR.n2040 6.52104
R10040 VDPWR.n1650 VDPWR.n1649 6.52104
R10041 VDPWR.n2188 VDPWR.n1100 6.50542
R10042 VDPWR.n2304 VDPWR.n2303 6.50542
R10043 VDPWR.n1261 VDPWR.n1260 6.48583
R10044 VDPWR.n2475 VDPWR.n2474 6.48583
R10045 VDPWR.n2471 VDPWR.n2470 6.46951
R10046 VDPWR.n2865 VDPWR.n965 6.4005
R10047 VDPWR.n2387 VDPWR 6.4005
R10048 VDPWR.n2470 VDPWR.n2469 6.4005
R10049 VDPWR.n749 VDPWR.n748 6.37981
R10050 VDPWR.n745 VDPWR.n743 6.37981
R10051 VDPWR.n737 VDPWR.n736 6.37981
R10052 VDPWR.n734 VDPWR.n733 6.37981
R10053 VDPWR.n2771 VDPWR.n2768 6.3005
R10054 VDPWR.n720 VDPWR.n656 6.18087
R10055 VDPWR.n3177 VDPWR.n3172 6.12434
R10056 VDPWR.n714 VDPWR.n705 6.02403
R10057 VDPWR.n661 VDPWR.n658 6.02403
R10058 VDPWR.n525 VDPWR.n516 6.02403
R10059 VDPWR.n477 VDPWR.n468 6.02403
R10060 VDPWR.n413 VDPWR.n404 6.02403
R10061 VDPWR.n418 VDPWR.n415 6.02403
R10062 VDPWR.n769 VDPWR.n760 6.02403
R10063 VDPWR.n3128 VDPWR.n3119 6.02403
R10064 VDPWR.n2741 VDPWR.n2740 5.97436
R10065 VDPWR.n1259 VDPWR.n1258 5.8885
R10066 VDPWR.n2473 VDPWR.n2472 5.8885
R10067 VDPWR.n2796 VDPWR.n2791 5.85193
R10068 VDPWR.n3177 VDPWR.n3176 5.75618
R10069 VDPWR.n2233 VDPWR.n2196 5.66607
R10070 VDPWR.n1052 VDPWR.n1041 5.66607
R10071 VDPWR.n1439 VDPWR.n1438 5.66204
R10072 VDPWR.n1441 VDPWR.n1439 5.66204
R10073 VDPWR.n1445 VDPWR.n1321 5.66204
R10074 VDPWR.n1446 VDPWR.n1445 5.66204
R10075 VDPWR.n1446 VDPWR.n1314 5.66204
R10076 VDPWR.n1461 VDPWR.n1314 5.66204
R10077 VDPWR.n1462 VDPWR.n1461 5.66204
R10078 VDPWR.n1463 VDPWR.n1462 5.66204
R10079 VDPWR.n1470 VDPWR.n1469 5.66204
R10080 VDPWR.n1471 VDPWR.n1470 5.66204
R10081 VDPWR.n1475 VDPWR.n1474 5.66204
R10082 VDPWR.n1476 VDPWR.n1475 5.66204
R10083 VDPWR.n1476 VDPWR.n1307 5.66204
R10084 VDPWR.n1480 VDPWR.n1307 5.66204
R10085 VDPWR.n1486 VDPWR.n1480 5.66204
R10086 VDPWR.n1486 VDPWR.n1485 5.66204
R10087 VDPWR.n1399 VDPWR.n1398 5.66204
R10088 VDPWR.n1406 VDPWR.n1337 5.66204
R10089 VDPWR.n1410 VDPWR.n1337 5.66204
R10090 VDPWR.n1414 VDPWR.n1412 5.66204
R10091 VDPWR.n1414 VDPWR.n1413 5.66204
R10092 VDPWR.n1572 VDPWR.n1571 5.66204
R10093 VDPWR.n1571 VDPWR.n1570 5.66204
R10094 VDPWR.n1567 VDPWR.n1566 5.66204
R10095 VDPWR.n1566 VDPWR.n1565 5.66204
R10096 VDPWR.n1565 VDPWR.n1526 5.66204
R10097 VDPWR.n1561 VDPWR.n1526 5.66204
R10098 VDPWR.n1561 VDPWR.n1560 5.66204
R10099 VDPWR.n1560 VDPWR.n1559 5.66204
R10100 VDPWR.n1729 VDPWR.n1728 5.66204
R10101 VDPWR.n1736 VDPWR.n1273 5.66204
R10102 VDPWR.n1740 VDPWR.n1273 5.66204
R10103 VDPWR.n1745 VDPWR.n1742 5.66204
R10104 VDPWR.n1745 VDPWR.n1744 5.66204
R10105 VDPWR.n1775 VDPWR.n1255 5.66204
R10106 VDPWR.n1778 VDPWR.n1777 5.66204
R10107 VDPWR.n1778 VDPWR.n1241 5.66204
R10108 VDPWR.n1789 VDPWR.n1241 5.66204
R10109 VDPWR.n1790 VDPWR.n1789 5.66204
R10110 VDPWR.n1803 VDPWR.n1802 5.66204
R10111 VDPWR.n1805 VDPWR.n1235 5.66204
R10112 VDPWR.n1809 VDPWR.n1235 5.66204
R10113 VDPWR.n1814 VDPWR.n1809 5.66204
R10114 VDPWR.n1814 VDPWR.n1813 5.66204
R10115 VDPWR.n2013 VDPWR.n2012 5.66204
R10116 VDPWR.n2012 VDPWR.n2011 5.66204
R10117 VDPWR.n1176 VDPWR.n1168 5.66204
R10118 VDPWR.n2022 VDPWR.n2021 5.66204
R10119 VDPWR.n2021 VDPWR.n2020 5.66204
R10120 VDPWR.n1148 VDPWR.n1142 5.66204
R10121 VDPWR.n1149 VDPWR.n1148 5.66204
R10122 VDPWR.n2029 VDPWR.n2028 5.66204
R10123 VDPWR.n1638 VDPWR.n1637 5.66204
R10124 VDPWR.n1637 VDPWR.n1634 5.66204
R10125 VDPWR.n1632 VDPWR.n1125 5.66204
R10126 VDPWR.n2060 VDPWR.n1125 5.66204
R10127 VDPWR.n1646 VDPWR.n1645 5.66204
R10128 VDPWR.n2146 VDPWR.n2145 5.66204
R10129 VDPWR.n2147 VDPWR.n2146 5.66204
R10130 VDPWR.n2151 VDPWR.n2150 5.66204
R10131 VDPWR.n2151 VDPWR.n1112 5.66204
R10132 VDPWR.n2165 VDPWR.n1112 5.66204
R10133 VDPWR.n535 VDPWR 5.6325
R10134 VDPWR.n3175 VDPWR 5.6325
R10135 VDPWR.n1792 VDPWR.n1239 5.48759
R10136 VDPWR.n1768 VDPWR.n1767 5.42606
R10137 VDPWR.n1797 VDPWR.n1796 5.42606
R10138 VDPWR.n1833 VDPWR.n1222 5.3712
R10139 VDPWR.n1438 VDPWR.n1323 5.29281
R10140 VDPWR.n1463 VDPWR.n1312 5.29281
R10141 VDPWR.n1469 VDPWR.n1311 5.29281
R10142 VDPWR.n1485 VDPWR.n1482 5.29281
R10143 VDPWR.n1398 VDPWR.n1397 5.29281
R10144 VDPWR.n1399 VDPWR.n1339 5.29281
R10145 VDPWR.n1406 VDPWR.n1405 5.29281
R10146 VDPWR.n1413 VDPWR.n1328 5.29281
R10147 VDPWR.n1572 VDPWR.n1521 5.29281
R10148 VDPWR.n1559 VDPWR.n1528 5.29281
R10149 VDPWR.n1728 VDPWR.n1727 5.29281
R10150 VDPWR.n1729 VDPWR.n1275 5.29281
R10151 VDPWR.n1736 VDPWR.n1735 5.29281
R10152 VDPWR.n1744 VDPWR.n1743 5.29281
R10153 VDPWR.n1771 VDPWR.n1769 5.29281
R10154 VDPWR.n1791 VDPWR.n1790 5.29281
R10155 VDPWR.n1799 VDPWR.n1798 5.29281
R10156 VDPWR.n1813 VDPWR.n1810 5.29281
R10157 VDPWR.n2013 VDPWR.n1156 5.29281
R10158 VDPWR.n1177 VDPWR.n1176 5.29281
R10159 VDPWR.n2022 VDPWR.n1153 5.29281
R10160 VDPWR.n1142 VDPWR.n1134 5.29281
R10161 VDPWR.n2028 VDPWR.n2027 5.29281
R10162 VDPWR.n1639 VDPWR.n1638 5.29281
R10163 VDPWR.n2060 VDPWR.n2059 5.29281
R10164 VDPWR.n1646 VDPWR.n1628 5.29281
R10165 VDPWR.n1645 VDPWR.n1644 5.29281
R10166 VDPWR.n2137 VDPWR.n2136 5.29281
R10167 VDPWR.n2137 VDPWR.n2080 5.29281
R10168 VDPWR.n2166 VDPWR.n2165 5.29281
R10169 VDPWR.n2871 VDPWR.n962 5.27109
R10170 VDPWR.n2531 VDPWR.n2431 5.27109
R10171 VDPWR.n2095 VDPWR.n2094 5.25888
R10172 VDPWR.n2194 VDPWR.n2193 5.2464
R10173 VDPWR.n1039 VDPWR.n1036 5.2464
R10174 VDPWR.n1836 VDPWR.n1835 5.18397
R10175 VDPWR.n1849 VDPWR.n1848 5.18397
R10176 VDPWR.n2219 VDPWR.n2209 5.18397
R10177 VDPWR.n2910 VDPWR.n950 5.18397
R10178 VDPWR.n2916 VDPWR.n948 5.18397
R10179 VDPWR.n717 VDPWR.n716 5.18145
R10180 VDPWR.n701 VDPWR.n700 5.18145
R10181 VDPWR.n685 VDPWR.n684 5.18145
R10182 VDPWR.n669 VDPWR.n668 5.18145
R10183 VDPWR.n528 VDPWR.n527 5.18145
R10184 VDPWR.n512 VDPWR.n511 5.18145
R10185 VDPWR.n496 VDPWR.n495 5.18145
R10186 VDPWR.n480 VDPWR.n479 5.18145
R10187 VDPWR.n464 VDPWR.n463 5.18145
R10188 VDPWR.n458 VDPWR.n457 5.18145
R10189 VDPWR.n442 VDPWR.n441 5.18145
R10190 VDPWR.n426 VDPWR.n425 5.18145
R10191 VDPWR.n3169 VDPWR.n3168 5.18145
R10192 VDPWR.n3163 VDPWR.n3162 5.18145
R10193 VDPWR.n3147 VDPWR.n3146 5.18145
R10194 VDPWR.n3131 VDPWR.n3130 5.18145
R10195 VDPWR.n2192 VDPWR.n2191 5.14148
R10196 VDPWR.n2785 VDPWR.n2784 5.1205
R10197 VDPWR.n2308 VDPWR.n1031 5.103
R10198 VDPWR.n1063 VDPWR.n1062 5.03657
R10199 VDPWR.t133 VDPWR.t346 5.03584
R10200 VDPWR.t134 VDPWR.t1004 5.03584
R10201 VDPWR.t562 VDPWR.t254 5.03584
R10202 VDPWR.t797 VDPWR.t785 5.03584
R10203 VDPWR.t334 VDPWR.t294 5.03584
R10204 VDPWR.n824 VDPWR.n822 4.98336
R10205 VDPWR.n2874 VDPWR.n961 4.9005
R10206 VDPWR.n699 VDPWR.n691 4.89462
R10207 VDPWR.n675 VDPWR.n673 4.89462
R10208 VDPWR.n510 VDPWR.n502 4.89462
R10209 VDPWR.n486 VDPWR.n484 4.89462
R10210 VDPWR.n456 VDPWR.n448 4.89462
R10211 VDPWR.n432 VDPWR.n430 4.89462
R10212 VDPWR.n3161 VDPWR.n3153 4.89462
R10213 VDPWR.n3137 VDPWR.n3135 4.89462
R10214 VDPWR.n3133 VDPWR.n3118 4.72727
R10215 VDPWR.n2108 VDPWR.n2107 4.69218
R10216 VDPWR.n602 VDPWR.n601 4.67352
R10217 VDPWR.n625 VDPWR.n590 4.67352
R10218 VDPWR.n322 VDPWR.n321 4.67352
R10219 VDPWR.n345 VDPWR.n310 4.67352
R10220 VDPWR.n1959 VDPWR.n1958 4.67352
R10221 VDPWR.n2891 VDPWR.n2886 4.67352
R10222 VDPWR.n2761 VDPWR.n2760 4.67352
R10223 VDPWR.n3061 VDPWR.n3060 4.67352
R10224 VDPWR.n3013 VDPWR.n3012 4.67352
R10225 VDPWR.n3012 VDPWR.n920 4.67352
R10226 VDPWR.n2416 VDPWR.n2351 4.67352
R10227 VDPWR.n2422 VDPWR.n2418 4.67352
R10228 VDPWR.n2401 VDPWR.n2400 4.67352
R10229 VDPWR.n2521 VDPWR.n2520 4.67352
R10230 VDPWR.n3089 VDPWR.n793 4.67352
R10231 VDPWR.n3085 VDPWR.n3084 4.67352
R10232 VDPWR.n3084 VDPWR.n3083 4.67352
R10233 VDPWR.n863 VDPWR.n815 4.67352
R10234 VDPWR.n859 VDPWR.n815 4.67352
R10235 VDPWR.n859 VDPWR.n858 4.67352
R10236 VDPWR.n852 VDPWR.n851 4.67352
R10237 VDPWR.n851 VDPWR.n826 4.67352
R10238 VDPWR.n64 VDPWR.n63 4.67352
R10239 VDPWR.n87 VDPWR.n52 4.67352
R10240 VDPWR.n751 VDPWR.n750 4.6505
R10241 VDPWR.n1968 VDPWR.n1915 4.62124
R10242 VDPWR.n2633 VDPWR.n2624 4.62124
R10243 VDPWR.n1764 VDPWR.n1261 4.62124
R10244 VDPWR.n1766 VDPWR.n1765 4.62124
R10245 VDPWR.n1795 VDPWR.n1794 4.62124
R10246 VDPWR.n2104 VDPWR.n2095 4.62124
R10247 VDPWR.n2476 VDPWR.n2475 4.62124
R10248 VDPWR.n2470 VDPWR.n2460 4.62124
R10249 VDPWR.n2743 VDPWR.n2739 4.5918
R10250 VDPWR.n1961 VDPWR.n1960 4.57193
R10251 VDPWR.n3014 VDPWR.n3013 4.57193
R10252 VDPWR.n2913 VDPWR.n950 4.54926
R10253 VDPWR.n2917 VDPWR.n2916 4.54926
R10254 VDPWR.n2946 VDPWR.n2945 4.54926
R10255 VDPWR.n2945 VDPWR.n935 4.54926
R10256 VDPWR.n2180 VDPWR.n2177 4.52113
R10257 VDPWR.n2868 VDPWR.n962 4.51815
R10258 VDPWR.n2696 VDPWR.n2695 4.51401
R10259 VDPWR.n2690 VDPWR.n2689 4.51401
R10260 VDPWR.n2666 VDPWR.n2665 4.51401
R10261 VDPWR.n2660 VDPWR.n2659 4.51401
R10262 VDPWR.n2510 VDPWR.n2509 4.51401
R10263 VDPWR.n2449 VDPWR.n2446 4.51401
R10264 VDPWR.n1490 VDPWR.n1302 4.51401
R10265 VDPWR.n1495 VDPWR.n1494 4.51401
R10266 VDPWR.n1454 VDPWR.n1319 4.51401
R10267 VDPWR.n1459 VDPWR.n1458 4.51401
R10268 VDPWR.n1421 VDPWR.n1333 4.51401
R10269 VDPWR.n1426 VDPWR.n1425 4.51401
R10270 VDPWR.n1374 VDPWR.n1373 4.51401
R10271 VDPWR.n1387 VDPWR.n1386 4.51401
R10272 VDPWR.n1557 VDPWR.n1556 4.51401
R10273 VDPWR.n1547 VDPWR.n1546 4.51401
R10274 VDPWR.n1586 VDPWR.n1287 4.51401
R10275 VDPWR.n1522 VDPWR.n1290 4.51401
R10276 VDPWR.n1818 VDPWR.n1230 4.51401
R10277 VDPWR.n1823 VDPWR.n1822 4.51401
R10278 VDPWR.n1782 VDPWR.n1248 4.51401
R10279 VDPWR.n1787 VDPWR.n1786 4.51401
R10280 VDPWR.n1752 VDPWR.n1269 4.51401
R10281 VDPWR.n1757 VDPWR.n1756 4.51401
R10282 VDPWR.n1712 VDPWR.n1677 4.51401
R10283 VDPWR.n1717 VDPWR.n1716 4.51401
R10284 VDPWR.n1887 VDPWR.n1886 4.51401
R10285 VDPWR.n1898 VDPWR.n1195 4.51401
R10286 VDPWR.n1856 VDPWR.n1217 4.51401
R10287 VDPWR.n1861 VDPWR.n1212 4.51401
R10288 VDPWR.n2009 VDPWR.n2008 4.51401
R10289 VDPWR.n2004 VDPWR.n2003 4.51401
R10290 VDPWR.n2038 VDPWR.n2037 4.51401
R10291 VDPWR.n2032 VDPWR.n2031 4.51401
R10292 VDPWR.n2070 VDPWR.n1119 4.51401
R10293 VDPWR.n1124 VDPWR.n1123 4.51401
R10294 VDPWR.n1670 VDPWR.n1598 4.51401
R10295 VDPWR.n1661 VDPWR.n1657 4.51401
R10296 VDPWR.n1956 VDPWR.n1955 4.51401
R10297 VDPWR.n1946 VDPWR.n1945 4.51401
R10298 VDPWR.n1188 VDPWR.n1187 4.51401
R10299 VDPWR.n1972 VDPWR.n1971 4.51401
R10300 VDPWR.n2329 VDPWR.n1015 4.51401
R10301 VDPWR.n2320 VDPWR.n2319 4.51401
R10302 VDPWR.n2247 VDPWR.n1094 4.51401
R10303 VDPWR.n2240 VDPWR.n2239 4.51401
R10304 VDPWR.n2157 VDPWR.n2075 4.51401
R10305 VDPWR.n2161 VDPWR.n1111 4.51401
R10306 VDPWR.n2113 VDPWR.n2112 4.51401
R10307 VDPWR.n2127 VDPWR.n2126 4.51401
R10308 VDPWR.n1078 VDPWR.n1076 4.51401
R10309 VDPWR.n1088 VDPWR.n1087 4.51401
R10310 VDPWR.n1043 VDPWR.n1037 4.51401
R10311 VDPWR.n2288 VDPWR.n2287 4.51401
R10312 VDPWR.n2881 VDPWR.n2880 4.51401
R10313 VDPWR.n2899 VDPWR.n2898 4.51401
R10314 VDPWR.n2842 VDPWR.n976 4.51401
R10315 VDPWR.n2846 VDPWR.n968 4.51401
R10316 VDPWR.n2803 VDPWR.n991 4.51401
R10317 VDPWR.n2808 VDPWR.n2807 4.51401
R10318 VDPWR.n2753 VDPWR.n2721 4.51401
R10319 VDPWR.n2758 VDPWR.n2757 4.51401
R10320 VDPWR.n2964 VDPWR.n2963 4.51401
R10321 VDPWR.n2975 VDPWR.n925 4.51401
R10322 VDPWR.n2930 VDPWR.n945 4.51401
R10323 VDPWR.n2935 VDPWR.n2934 4.51401
R10324 VDPWR.n903 VDPWR.n901 4.51401
R10325 VDPWR.n3030 VDPWR.n3029 4.51401
R10326 VDPWR.n3065 VDPWR.n875 4.51401
R10327 VDPWR.n3056 VDPWR.n3055 4.51401
R10328 VDPWR.n2464 VDPWR.n785 4.51401
R10329 VDPWR.n788 VDPWR.n784 4.51401
R10330 VDPWR.n2569 VDPWR.n2549 4.51401
R10331 VDPWR.n2717 VDPWR.n2716 4.51401
R10332 VDPWR.n3009 VDPWR.n3008 4.51401
R10333 VDPWR.n3003 VDPWR.n3002 4.51401
R10334 VDPWR.n2424 VDPWR.n2344 4.51401
R10335 VDPWR.n2346 VDPWR.n2342 4.51401
R10336 VDPWR.n2391 VDPWR.n2365 4.51401
R10337 VDPWR.n2393 VDPWR.n2361 4.51401
R10338 VDPWR.n848 VDPWR.n847 4.51401
R10339 VDPWR.n841 VDPWR.n772 4.51401
R10340 VDPWR.n3076 VDPWR.n3075 4.51401
R10341 VDPWR.n806 VDPWR.n804 4.51401
R10342 VDPWR.n2193 VDPWR.n2192 4.51198
R10343 VDPWR.n2277 VDPWR.n1063 4.51198
R10344 VDPWR.n537 VDPWR.n536 4.5005
R10345 VDPWR.n1534 VDPWR.n1530 4.5005
R10346 VDPWR.n1552 VDPWR.n1551 4.5005
R10347 VDPWR.n1544 VDPWR.n1536 4.5005
R10348 VDPWR.n1371 VDPWR.n1370 4.5005
R10349 VDPWR.n1382 VDPWR.n1381 4.5005
R10350 VDPWR.n1345 VDPWR.n1344 4.5005
R10351 VDPWR.n1420 VDPWR.n1419 4.5005
R10352 VDPWR.n1418 VDPWR.n1417 4.5005
R10353 VDPWR.n1336 VDPWR.n1330 4.5005
R10354 VDPWR.n1453 VDPWR.n1452 4.5005
R10355 VDPWR.n1450 VDPWR.n1449 4.5005
R10356 VDPWR.n1316 VDPWR.n1315 4.5005
R10357 VDPWR.n1489 VDPWR.n1488 4.5005
R10358 VDPWR.n1306 VDPWR.n1305 4.5005
R10359 VDPWR.n1483 VDPWR.n1299 4.5005
R10360 VDPWR.n1585 VDPWR.n1584 4.5005
R10361 VDPWR.n1583 VDPWR.n1582 4.5005
R10362 VDPWR.n1579 VDPWR.n1578 4.5005
R10363 VDPWR.n1890 VDPWR.n1889 4.5005
R10364 VDPWR.n1891 VDPWR.n1197 4.5005
R10365 VDPWR.n1900 VDPWR.n1899 4.5005
R10366 VDPWR.n1711 VDPWR.n1710 4.5005
R10367 VDPWR.n1681 VDPWR.n1680 4.5005
R10368 VDPWR.n1281 VDPWR.n1280 4.5005
R10369 VDPWR.n1751 VDPWR.n1750 4.5005
R10370 VDPWR.n1749 VDPWR.n1748 4.5005
R10371 VDPWR.n1272 VDPWR.n1265 4.5005
R10372 VDPWR.n1781 VDPWR.n1780 4.5005
R10373 VDPWR.n1254 VDPWR.n1253 4.5005
R10374 VDPWR.n1251 VDPWR.n1243 4.5005
R10375 VDPWR.n1817 VDPWR.n1816 4.5005
R10376 VDPWR.n1234 VDPWR.n1233 4.5005
R10377 VDPWR.n1811 VDPWR.n1226 4.5005
R10378 VDPWR.n1855 VDPWR.n1854 4.5005
R10379 VDPWR.n1853 VDPWR.n1852 4.5005
R10380 VDPWR.n1863 VDPWR.n1862 4.5005
R10381 VDPWR.n1933 VDPWR.n1930 4.5005
R10382 VDPWR.n1951 VDPWR.n1950 4.5005
R10383 VDPWR.n1943 VDPWR.n1935 4.5005
R10384 VDPWR.n1669 VDPWR.n1668 4.5005
R10385 VDPWR.n1658 VDPWR.n1600 4.5005
R10386 VDPWR.n1663 VDPWR.n1662 4.5005
R10387 VDPWR.n2069 VDPWR.n2068 4.5005
R10388 VDPWR.n2067 VDPWR.n2066 4.5005
R10389 VDPWR.n2063 VDPWR.n2062 4.5005
R10390 VDPWR.n1143 VDPWR.n1136 4.5005
R10391 VDPWR.n1146 VDPWR.n1145 4.5005
R10392 VDPWR.n1144 VDPWR.n1139 4.5005
R10393 VDPWR.n1160 VDPWR.n1159 4.5005
R10394 VDPWR.n1173 VDPWR.n1172 4.5005
R10395 VDPWR.n1174 VDPWR.n1164 4.5005
R10396 VDPWR.n1979 VDPWR.n1978 4.5005
R10397 VDPWR.n1911 VDPWR.n1189 4.5005
R10398 VDPWR.n1913 VDPWR.n1910 4.5005
R10399 VDPWR.n2262 VDPWR.n2261 4.5005
R10400 VDPWR.n1083 VDPWR.n1079 4.5005
R10401 VDPWR.n1085 VDPWR.n1082 4.5005
R10402 VDPWR.n2110 VDPWR.n2089 4.5005
R10403 VDPWR.n2122 VDPWR.n2121 4.5005
R10404 VDPWR.n2086 VDPWR.n2085 4.5005
R10405 VDPWR.n2156 VDPWR.n2155 4.5005
R10406 VDPWR.n2154 VDPWR.n2153 4.5005
R10407 VDPWR.n2163 VDPWR.n2162 4.5005
R10408 VDPWR.n2246 VDPWR.n2245 4.5005
R10409 VDPWR.n2235 VDPWR.n1097 4.5005
R10410 VDPWR.n2238 VDPWR.n2197 4.5005
R10411 VDPWR.n2328 VDPWR.n2327 4.5005
R10412 VDPWR.n1021 VDPWR.n1017 4.5005
R10413 VDPWR.n2322 VDPWR.n2321 4.5005
R10414 VDPWR.n2295 VDPWR.n2294 4.5005
R10415 VDPWR.n1044 VDPWR.n1042 4.5005
R10416 VDPWR.n1054 VDPWR.n1048 4.5005
R10417 VDPWR.n2967 VDPWR.n2966 4.5005
R10418 VDPWR.n2968 VDPWR.n927 4.5005
R10419 VDPWR.n2977 VDPWR.n2976 4.5005
R10420 VDPWR.n2752 VDPWR.n2751 4.5005
R10421 VDPWR.n2725 VDPWR.n2724 4.5005
R10422 VDPWR.n2747 VDPWR.n1007 4.5005
R10423 VDPWR.n2802 VDPWR.n2801 4.5005
R10424 VDPWR.n2800 VDPWR.n2799 4.5005
R10425 VDPWR.n994 VDPWR.n986 4.5005
R10426 VDPWR.n2841 VDPWR.n2840 4.5005
R10427 VDPWR.n977 VDPWR.n970 4.5005
R10428 VDPWR.n2848 VDPWR.n2847 4.5005
R10429 VDPWR.n2878 VDPWR.n2877 4.5005
R10430 VDPWR.n2894 VDPWR.n2893 4.5005
R10431 VDPWR.n960 VDPWR.n956 4.5005
R10432 VDPWR.n2929 VDPWR.n2928 4.5005
R10433 VDPWR.n2927 VDPWR.n2926 4.5005
R10434 VDPWR.n941 VDPWR.n940 4.5005
R10435 VDPWR.n2571 VDPWR.n2570 4.5005
R10436 VDPWR.n2576 VDPWR.n2575 4.5005
R10437 VDPWR.n2543 VDPWR.n2542 4.5005
R10438 VDPWR.n2598 VDPWR.n2589 4.5005
R10439 VDPWR.n2600 VDPWR.n2599 4.5005
R10440 VDPWR.n2601 VDPWR.n2592 4.5005
R10441 VDPWR.n2650 VDPWR.n2615 4.5005
R10442 VDPWR.n2653 VDPWR.n2652 4.5005
R10443 VDPWR.n2654 VDPWR.n2618 4.5005
R10444 VDPWR.n3064 VDPWR.n3063 4.5005
R10445 VDPWR.n881 VDPWR.n877 4.5005
R10446 VDPWR.n3058 VDPWR.n3057 4.5005
R10447 VDPWR.n3037 VDPWR.n3036 4.5005
R10448 VDPWR.n904 VDPWR.n902 4.5005
R10449 VDPWR.n909 VDPWR.n906 4.5005
R10450 VDPWR.n2992 VDPWR.n922 4.5005
R10451 VDPWR.n2995 VDPWR.n2994 4.5005
R10452 VDPWR.n2986 VDPWR.n2985 4.5005
R10453 VDPWR.n846 VDPWR.n845 4.5005
R10454 VDPWR.n829 VDPWR.n828 4.5005
R10455 VDPWR.n840 VDPWR.n839 4.5005
R10456 VDPWR.n2390 VDPWR.n2389 4.5005
R10457 VDPWR.n2363 VDPWR.n2360 4.5005
R10458 VDPWR.n2395 VDPWR.n2394 4.5005
R10459 VDPWR.n2427 VDPWR.n2426 4.5005
R10460 VDPWR.n2428 VDPWR.n2345 4.5005
R10461 VDPWR.n2534 VDPWR.n2533 4.5005
R10462 VDPWR.n2447 VDPWR.n2444 4.5005
R10463 VDPWR.n2497 VDPWR.n2496 4.5005
R10464 VDPWR.n2495 VDPWR.n2494 4.5005
R10465 VDPWR.n2466 VDPWR.n2465 4.5005
R10466 VDPWR.n2467 VDPWR.n786 4.5005
R10467 VDPWR.n3100 VDPWR.n3099 4.5005
R10468 VDPWR.n809 VDPWR.n802 4.5005
R10469 VDPWR.n810 VDPWR.n805 4.5005
R10470 VDPWR.n868 VDPWR.n867 4.5005
R10471 VDPWR.n2048 VDPWR.n1130 4.49637
R10472 VDPWR.n2243 VDPWR.n2194 4.40706
R10473 VDPWR.n2298 VDPWR.n1039 4.40706
R10474 VDPWR.n759 VDPWR.n758 4.38372
R10475 VDPWR.n601 VDPWR.n600 4.36875
R10476 VDPWR.n625 VDPWR.n624 4.36875
R10477 VDPWR.n584 VDPWR.n583 4.36875
R10478 VDPWR.n554 VDPWR.n553 4.36875
R10479 VDPWR.n321 VDPWR.n320 4.36875
R10480 VDPWR.n345 VDPWR.n344 4.36875
R10481 VDPWR.n304 VDPWR.n303 4.36875
R10482 VDPWR.n274 VDPWR.n273 4.36875
R10483 VDPWR.n1958 VDPWR.n1928 4.36875
R10484 VDPWR.n2180 VDPWR.n2179 4.36875
R10485 VDPWR.n2762 VDPWR.n2761 4.36875
R10486 VDPWR.n3015 VDPWR.n917 4.36875
R10487 VDPWR.n2987 VDPWR.n920 4.36875
R10488 VDPWR.n2411 VDPWR.n2351 4.36875
R10489 VDPWR.n2418 VDPWR.n2417 4.36875
R10490 VDPWR.n2401 VDPWR.n2357 4.36875
R10491 VDPWR.n2525 VDPWR.n2524 4.36875
R10492 VDPWR.n2521 VDPWR.n2434 4.36875
R10493 VDPWR.n2518 VDPWR.n2437 4.36875
R10494 VDPWR.n3092 VDPWR.n792 4.36875
R10495 VDPWR.n864 VDPWR.n863 4.36875
R10496 VDPWR.n830 VDPWR.n826 4.36875
R10497 VDPWR.n63 VDPWR.n62 4.36875
R10498 VDPWR.n87 VDPWR.n86 4.36875
R10499 VDPWR.n46 VDPWR.n45 4.36875
R10500 VDPWR.n16 VDPWR.n15 4.36875
R10501 VDPWR.n2405 VDPWR 4.3525
R10502 VDPWR.n1835 VDPWR.n1221 4.33769
R10503 VDPWR.n2093 VDPWR.n2092 4.29023
R10504 VDPWR.n2890 VDPWR.n2889 4.26717
R10505 VDPWR.n1968 VDPWR.n1966 4.14168
R10506 VDPWR.n3172 VDPWR.n3171 4.06613
R10507 VDPWR.n720 VDPWR.n719 4.05291
R10508 VDPWR.n1434 VDPWR.n1326 4.02033
R10509 VDPWR.n1357 VDPWR.n1353 4.02033
R10510 VDPWR.n1357 VDPWR.n1356 4.02033
R10511 VDPWR.n1366 VDPWR.n1360 4.02033
R10512 VDPWR.n1366 VDPWR.n1365 4.02033
R10513 VDPWR.n1549 VDPWR.n1540 4.02033
R10514 VDPWR.n1549 VDPWR.n1543 4.02033
R10515 VDPWR.n1690 VDPWR.n1686 4.02033
R10516 VDPWR.n1690 VDPWR.n1689 4.02033
R10517 VDPWR.n1699 VDPWR.n1693 4.02033
R10518 VDPWR.n1699 VDPWR.n1698 4.02033
R10519 VDPWR.n1896 VDPWR.n1208 4.02033
R10520 VDPWR.n1896 VDPWR.n1895 4.02033
R10521 VDPWR.n2048 VDPWR.n1128 4.02033
R10522 VDPWR.n1621 VDPWR.n1606 4.02033
R10523 VDPWR.n1621 VDPWR.n1612 4.02033
R10524 VDPWR.n1620 VDPWR.n1615 4.02033
R10525 VDPWR.n1620 VDPWR.n1619 4.02033
R10526 VDPWR.n1948 VDPWR.n1939 4.02033
R10527 VDPWR.n1948 VDPWR.n1942 4.02033
R10528 VDPWR.n2102 VDPWR.n2098 4.02033
R10529 VDPWR.n2102 VDPWR.n2101 4.02033
R10530 VDPWR.n1075 VDPWR.n1071 4.02033
R10531 VDPWR.n1075 VDPWR.n1074 4.02033
R10532 VDPWR.n2735 VDPWR.n2731 4.02033
R10533 VDPWR.n2735 VDPWR.n2734 4.02033
R10534 VDPWR.n2973 VDPWR.n932 4.02033
R10535 VDPWR.n2973 VDPWR.n2972 4.02033
R10536 VDPWR.n2556 VDPWR.n2552 4.02033
R10537 VDPWR.n2556 VDPWR.n2555 4.02033
R10538 VDPWR.n2687 VDPWR.n2597 4.02033
R10539 VDPWR.n3052 VDPWR.n891 4.02033
R10540 VDPWR.n3000 VDPWR.n2991 4.02033
R10541 VDPWR.n3000 VDPWR.n2999 4.02033
R10542 VDPWR.n2377 VDPWR.n2373 4.02033
R10543 VDPWR.n2377 VDPWR.n2376 4.02033
R10544 VDPWR.n843 VDPWR.n834 4.02033
R10545 VDPWR.n843 VDPWR.n838 4.02033
R10546 VDPWR.n2242 VDPWR.n2196 3.98739
R10547 VDPWR.n2297 VDPWR.n1041 3.98739
R10548 VDPWR.n1848 VDPWR.n1213 3.91455
R10549 VDPWR.n2519 VDPWR.n2518 3.86082
R10550 VDPWR.n1767 VDPWR.n1766 3.78037
R10551 VDPWR.n1796 VDPWR.n1795 3.78037
R10552 VDPWR.n1761 VDPWR.n1261 3.75517
R10553 VDPWR.n1828 VDPWR.n1827 3.75222
R10554 VDPWR.n1795 VDPWR.n1239 3.69446
R10555 VDPWR.n2475 VDPWR.n2459 3.66983
R10556 VDPWR.n724 VDPWR.t824 3.61217
R10557 VDPWR.n724 VDPWR.t820 3.61217
R10558 VDPWR.n726 VDPWR.t253 3.61217
R10559 VDPWR.n726 VDPWR.t342 3.61217
R10560 VDPWR.n722 VDPWR.t822 3.61217
R10561 VDPWR.n722 VDPWR.t219 3.61217
R10562 VDPWR.n2421 VDPWR.n2420 3.55606
R10563 VDPWR.n2092 VDPWR.n2091 3.53179
R10564 VDPWR.n2836 VDPWR.n969 3.4812
R10565 VDPWR.n1379 VDPWR.n1378 3.47425
R10566 VDPWR.n1390 VDPWR.n1389 3.47425
R10567 VDPWR.n1392 VDPWR.n1390 3.47425
R10568 VDPWR.n1511 VDPWR.n1294 3.47425
R10569 VDPWR.n1512 VDPWR.n1511 3.47425
R10570 VDPWR.n1513 VDPWR.n1512 3.47425
R10571 VDPWR.n1708 VDPWR.n1707 3.47425
R10572 VDPWR.n1720 VDPWR.n1719 3.47425
R10573 VDPWR.n1722 VDPWR.n1720 3.47425
R10574 VDPWR.n1997 VDPWR.n1996 3.47425
R10575 VDPWR.n2046 VDPWR.n2045 3.47425
R10576 VDPWR.n2045 VDPWR.n1131 3.47425
R10577 VDPWR.n1666 VDPWR.n1665 3.47425
R10578 VDPWR.n1655 VDPWR.n1654 3.47425
R10579 VDPWR.n1654 VDPWR.n1653 3.47425
R10580 VDPWR.n2129 VDPWR.n2084 3.47425
R10581 VDPWR.n2130 VDPWR.n2129 3.47425
R10582 VDPWR.n2131 VDPWR.n2130 3.47425
R10583 VDPWR.n2325 VDPWR.n2324 3.47425
R10584 VDPWR.n2267 VDPWR.n2266 3.47425
R10585 VDPWR.n2957 VDPWR.n934 3.47425
R10586 VDPWR.n2958 VDPWR.n2957 3.47425
R10587 VDPWR.n2960 VDPWR.n2958 3.47425
R10588 VDPWR.n2490 VDPWR.n2454 3.47425
R10589 VDPWR.n3178 VDPWR.n3177 3.44037
R10590 VDPWR.n2691 VDPWR.n2690 3.43925
R10591 VDPWR.n2695 VDPWR.n2694 3.43925
R10592 VDPWR.n2661 VDPWR.n2660 3.43925
R10593 VDPWR.n2665 VDPWR.n2664 3.43925
R10594 VDPWR.n1494 VDPWR.n1493 3.43925
R10595 VDPWR.n1491 VDPWR.n1490 3.43925
R10596 VDPWR.n1458 VDPWR.n1457 3.43925
R10597 VDPWR.n1455 VDPWR.n1454 3.43925
R10598 VDPWR.n1425 VDPWR.n1424 3.43925
R10599 VDPWR.n1422 VDPWR.n1421 3.43925
R10600 VDPWR.n1386 VDPWR.n1385 3.43925
R10601 VDPWR.n1373 VDPWR.n1372 3.43925
R10602 VDPWR.n1546 VDPWR.n1545 3.43925
R10603 VDPWR.n1556 VDPWR.n1555 3.43925
R10604 VDPWR.n1290 VDPWR.n1285 3.43925
R10605 VDPWR.n1587 VDPWR.n1586 3.43925
R10606 VDPWR.n1822 VDPWR.n1821 3.43925
R10607 VDPWR.n1819 VDPWR.n1818 3.43925
R10608 VDPWR.n1786 VDPWR.n1785 3.43925
R10609 VDPWR.n1783 VDPWR.n1782 3.43925
R10610 VDPWR.n1756 VDPWR.n1755 3.43925
R10611 VDPWR.n1753 VDPWR.n1752 3.43925
R10612 VDPWR.n1716 VDPWR.n1715 3.43925
R10613 VDPWR.n1713 VDPWR.n1712 3.43925
R10614 VDPWR.n1903 VDPWR.n1195 3.43925
R10615 VDPWR.n1887 VDPWR.n1194 3.43925
R10616 VDPWR.n1861 VDPWR.n1860 3.43925
R10617 VDPWR.n1857 VDPWR.n1856 3.43925
R10618 VDPWR.n2005 VDPWR.n2004 3.43925
R10619 VDPWR.n2008 VDPWR.n2007 3.43925
R10620 VDPWR.n2033 VDPWR.n2032 3.43925
R10621 VDPWR.n2037 VDPWR.n2036 3.43925
R10622 VDPWR.n1123 VDPWR.n1117 3.43925
R10623 VDPWR.n2071 VDPWR.n2070 3.43925
R10624 VDPWR.n1661 VDPWR.n1595 3.43925
R10625 VDPWR.n1671 VDPWR.n1670 3.43925
R10626 VDPWR.n1945 VDPWR.n1944 3.43925
R10627 VDPWR.n1955 VDPWR.n1954 3.43925
R10628 VDPWR.n1973 VDPWR.n1972 3.43925
R10629 VDPWR.n1975 VDPWR.n1188 3.43925
R10630 VDPWR.n2320 VDPWR.n1013 3.43925
R10631 VDPWR.n2330 VDPWR.n2329 3.43925
R10632 VDPWR.n2239 VDPWR.n1092 3.43925
R10633 VDPWR.n2248 VDPWR.n2247 3.43925
R10634 VDPWR.n2161 VDPWR.n2160 3.43925
R10635 VDPWR.n2158 VDPWR.n2157 3.43925
R10636 VDPWR.n2126 VDPWR.n2125 3.43925
R10637 VDPWR.n2112 VDPWR.n2111 3.43925
R10638 VDPWR.n2257 VDPWR.n1088 3.43925
R10639 VDPWR.n1080 VDPWR.n1078 3.43925
R10640 VDPWR.n2289 VDPWR.n2288 3.43925
R10641 VDPWR.n2291 VDPWR.n1043 3.43925
R10642 VDPWR.n2898 VDPWR.n2897 3.43925
R10643 VDPWR.n2880 VDPWR.n2879 3.43925
R10644 VDPWR.n2846 VDPWR.n2845 3.43925
R10645 VDPWR.n2843 VDPWR.n2842 3.43925
R10646 VDPWR.n2807 VDPWR.n2806 3.43925
R10647 VDPWR.n2804 VDPWR.n2803 3.43925
R10648 VDPWR.n2757 VDPWR.n2756 3.43925
R10649 VDPWR.n2754 VDPWR.n2753 3.43925
R10650 VDPWR.n2980 VDPWR.n925 3.43925
R10651 VDPWR.n2964 VDPWR.n924 3.43925
R10652 VDPWR.n2934 VDPWR.n2933 3.43925
R10653 VDPWR.n2931 VDPWR.n2930 3.43925
R10654 VDPWR.n3031 VDPWR.n3030 3.43925
R10655 VDPWR.n3033 VDPWR.n903 3.43925
R10656 VDPWR.n3056 VDPWR.n873 3.43925
R10657 VDPWR.n3066 VDPWR.n3065 3.43925
R10658 VDPWR.n3004 VDPWR.n3003 3.43925
R10659 VDPWR.n3008 VDPWR.n3007 3.43925
R10660 VDPWR.n2491 VDPWR.n2490 3.43649
R10661 VDPWR.n656 VDPWR.n655 3.4105
R10662 VDPWR.n2693 VDPWR.n2590 3.4105
R10663 VDPWR.n2692 VDPWR.n2591 3.4105
R10664 VDPWR.n2663 VDPWR.n2616 3.4105
R10665 VDPWR.n2662 VDPWR.n2617 3.4105
R10666 VDPWR.n1303 VDPWR.n1301 3.4105
R10667 VDPWR.n1304 VDPWR.n1300 3.4105
R10668 VDPWR.n1320 VDPWR.n1318 3.4105
R10669 VDPWR.n1448 VDPWR.n1317 3.4105
R10670 VDPWR.n1334 VDPWR.n1332 3.4105
R10671 VDPWR.n1416 VDPWR.n1331 3.4105
R10672 VDPWR.n1347 VDPWR.n1346 3.4105
R10673 VDPWR.n1384 VDPWR.n1383 3.4105
R10674 VDPWR.n1554 VDPWR.n1553 3.4105
R10675 VDPWR.n1533 VDPWR.n1532 3.4105
R10676 VDPWR.n1288 VDPWR.n1286 3.4105
R10677 VDPWR.n1581 VDPWR.n1580 3.4105
R10678 VDPWR.n1231 VDPWR.n1229 3.4105
R10679 VDPWR.n1232 VDPWR.n1227 3.4105
R10680 VDPWR.n1249 VDPWR.n1247 3.4105
R10681 VDPWR.n1252 VDPWR.n1244 3.4105
R10682 VDPWR.n1270 VDPWR.n1268 3.4105
R10683 VDPWR.n1747 VDPWR.n1266 3.4105
R10684 VDPWR.n1678 VDPWR.n1676 3.4105
R10685 VDPWR.n1679 VDPWR.n1282 3.4105
R10686 VDPWR.n1888 VDPWR.n1196 3.4105
R10687 VDPWR.n1902 VDPWR.n1901 3.4105
R10688 VDPWR.n1858 VDPWR.n1216 3.4105
R10689 VDPWR.n1859 VDPWR.n1215 3.4105
R10690 VDPWR.n1170 VDPWR.n1161 3.4105
R10691 VDPWR.n1171 VDPWR.n1163 3.4105
R10692 VDPWR.n2035 VDPWR.n1137 3.4105
R10693 VDPWR.n2034 VDPWR.n1138 3.4105
R10694 VDPWR.n1120 VDPWR.n1118 3.4105
R10695 VDPWR.n2065 VDPWR.n2064 3.4105
R10696 VDPWR.n1599 VDPWR.n1597 3.4105
R10697 VDPWR.n1660 VDPWR.n1659 3.4105
R10698 VDPWR.n1953 VDPWR.n1952 3.4105
R10699 VDPWR.n1932 VDPWR.n1931 3.4105
R10700 VDPWR.n1977 VDPWR.n1976 3.4105
R10701 VDPWR.n1909 VDPWR.n1190 3.4105
R10702 VDPWR.n1016 VDPWR.n1014 3.4105
R10703 VDPWR.n1023 VDPWR.n1022 3.4105
R10704 VDPWR.n1095 VDPWR.n1093 3.4105
R10705 VDPWR.n2237 VDPWR.n2236 3.4105
R10706 VDPWR.n2076 VDPWR.n2074 3.4105
R10707 VDPWR.n1115 VDPWR.n1114 3.4105
R10708 VDPWR.n2088 VDPWR.n2087 3.4105
R10709 VDPWR.n2124 VDPWR.n2123 3.4105
R10710 VDPWR.n2260 VDPWR.n2259 3.4105
R10711 VDPWR.n2258 VDPWR.n1081 3.4105
R10712 VDPWR.n2293 VDPWR.n2292 3.4105
R10713 VDPWR.n1047 VDPWR.n1045 3.4105
R10714 VDPWR.n958 VDPWR.n957 3.4105
R10715 VDPWR.n2896 VDPWR.n2895 3.4105
R10716 VDPWR.n978 VDPWR.n975 3.4105
R10717 VDPWR.n972 VDPWR.n971 3.4105
R10718 VDPWR.n992 VDPWR.n990 3.4105
R10719 VDPWR.n2798 VDPWR.n987 3.4105
R10720 VDPWR.n2722 VDPWR.n2720 3.4105
R10721 VDPWR.n2723 VDPWR.n1008 3.4105
R10722 VDPWR.n2965 VDPWR.n926 3.4105
R10723 VDPWR.n2979 VDPWR.n2978 3.4105
R10724 VDPWR.n946 VDPWR.n944 3.4105
R10725 VDPWR.n2925 VDPWR.n942 3.4105
R10726 VDPWR.n3035 VDPWR.n3034 3.4105
R10727 VDPWR.n3032 VDPWR.n905 3.4105
R10728 VDPWR.n876 VDPWR.n874 3.4105
R10729 VDPWR.n883 VDPWR.n882 3.4105
R10730 VDPWR.n3102 VDPWR.n784 3.4105
R10731 VDPWR.n3102 VDPWR.n785 3.4105
R10732 VDPWR.n3102 VDPWR.n783 3.4105
R10733 VDPWR.n3102 VDPWR.n3101 3.4105
R10734 VDPWR.n2508 VDPWR.n2446 3.4105
R10735 VDPWR.n2509 VDPWR.n2508 3.4105
R10736 VDPWR.n2508 VDPWR.n2498 3.4105
R10737 VDPWR.n2508 VDPWR.n2445 3.4105
R10738 VDPWR.n2719 VDPWR.n2718 3.4105
R10739 VDPWR.n2719 VDPWR.n2338 3.4105
R10740 VDPWR.n2718 VDPWR.n2717 3.4105
R10741 VDPWR.n2549 VDPWR.n2338 3.4105
R10742 VDPWR.n2573 VDPWR.n2572 3.4105
R10743 VDPWR.n2574 VDPWR.n2541 3.4105
R10744 VDPWR.n3006 VDPWR.n2983 3.4105
R10745 VDPWR.n3005 VDPWR.n2984 3.4105
R10746 VDPWR.n2536 VDPWR.n2342 3.4105
R10747 VDPWR.n2536 VDPWR.n2344 3.4105
R10748 VDPWR.n2536 VDPWR.n2341 3.4105
R10749 VDPWR.n2536 VDPWR.n2535 3.4105
R10750 VDPWR.n2393 VDPWR.n2392 3.4105
R10751 VDPWR.n2392 VDPWR.n2391 3.4105
R10752 VDPWR.n2392 VDPWR.n2364 3.4105
R10753 VDPWR.n2392 VDPWR.n2362 3.4105
R10754 VDPWR.n3074 VDPWR.n804 3.4105
R10755 VDPWR.n3075 VDPWR.n3074 3.4105
R10756 VDPWR.n3074 VDPWR.n803 3.4105
R10757 VDPWR.n3074 VDPWR.n869 3.4105
R10758 VDPWR.n3113 VDPWR.n771 3.4105
R10759 VDPWR.n847 VDPWR.n771 3.4105
R10760 VDPWR.n3114 VDPWR.n773 3.4105
R10761 VDPWR.n3114 VDPWR.n774 3.4105
R10762 VDPWR.n3114 VDPWR.n772 3.4105
R10763 VDPWR.t186 VDPWR.t788 3.35739
R10764 VDPWR.t964 VDPWR.t1162 3.35739
R10765 VDPWR.t176 VDPWR.t108 3.35739
R10766 VDPWR.t188 VDPWR.t72 3.35739
R10767 VDPWR.t906 VDPWR.t940 3.35739
R10768 VDPWR.t0 VDPWR.t46 3.35739
R10769 VDPWR.t385 VDPWR.t1122 3.35739
R10770 VDPWR.t833 VDPWR.t637 3.35739
R10771 VDPWR.t880 VDPWR.t112 3.35739
R10772 VDPWR.t216 VDPWR.t304 3.35739
R10773 VDPWR.n1376 VDPWR.n1350 3.2477
R10774 VDPWR.n1392 VDPWR.n1391 3.2477
R10775 VDPWR.n1504 VDPWR.n1503 3.2477
R10776 VDPWR.n1513 VDPWR.n1292 3.2477
R10777 VDPWR.n1704 VDPWR.n1683 3.2477
R10778 VDPWR.n1722 VDPWR.n1721 3.2477
R10779 VDPWR.n1996 VDPWR.n1995 3.2477
R10780 VDPWR.n2047 VDPWR.n2046 3.2477
R10781 VDPWR.n1602 VDPWR.n1601 3.2477
R10782 VDPWR.n1653 VDPWR.n1627 3.2477
R10783 VDPWR.n2115 VDPWR.n2090 3.2477
R10784 VDPWR.n2131 VDPWR.n2082 3.2477
R10785 VDPWR.n2324 VDPWR.n1019 3.2477
R10786 VDPWR.n2266 VDPWR.n2265 3.2477
R10787 VDPWR.n2952 VDPWR.n934 3.2477
R10788 VDPWR.n2960 VDPWR.n2959 3.2477
R10789 VDPWR.n2492 VDPWR.n2450 3.2477
R10790 VDPWR.n2486 VDPWR.n2485 3.2477
R10791 VDPWR.n478 VDPWR.n467 3.24308
R10792 VDPWR.n3129 VDPWR.n3118 3.24308
R10793 VDPWR.n691 VDPWR.n688 3.23917
R10794 VDPWR.n502 VDPWR.n499 3.23917
R10795 VDPWR.n448 VDPWR.n445 3.23917
R10796 VDPWR.n3153 VDPWR.n3150 3.23917
R10797 VDPWR.n675 VDPWR.n672 3.23136
R10798 VDPWR.n486 VDPWR.n483 3.23136
R10799 VDPWR.n432 VDPWR.n429 3.23136
R10800 VDPWR.n3137 VDPWR.n3134 3.23136
R10801 VDPWR.n462 VDPWR.n461 3.22655
R10802 VDPWR.n715 VDPWR.n704 3.22655
R10803 VDPWR.n526 VDPWR.n515 3.22655
R10804 VDPWR.n3167 VDPWR.n3166 3.22655
R10805 VDPWR.n2760 VDPWR.n1006 3.2005
R10806 VDPWR.n1258 VDPWR.n1257 3.151
R10807 VDPWR.n2191 VDPWR.n1100 3.14804
R10808 VDPWR.n2303 VDPWR.n2302 3.14804
R10809 VDPWR.n859 VDPWR.n819 3.12116
R10810 VDPWR.n1361 VDPWR.n1357 3.05586
R10811 VDPWR.n1694 VDPWR.n1690 3.05586
R10812 VDPWR.n1620 VDPWR.n1616 3.05586
R10813 VDPWR.n2103 VDPWR.n2102 3.05586
R10814 VDPWR.n2736 VDPWR.n2735 3.05586
R10815 VDPWR.n2560 VDPWR.n2556 3.05586
R10816 VDPWR.n2378 VDPWR.n2377 3.05586
R10817 VDPWR.n1366 VDPWR.n1362 3.04861
R10818 VDPWR.n1699 VDPWR.n1695 3.04861
R10819 VDPWR.n1884 VDPWR.n1205 3.04861
R10820 VDPWR.n1621 VDPWR.n1609 3.04861
R10821 VDPWR.n3052 VDPWR.n888 3.04861
R10822 VDPWR.n1434 VDPWR.n1433 3.04861
R10823 VDPWR.n1833 VDPWR.n1832 3.04861
R10824 VDPWR.n2055 VDPWR.n1128 3.04861
R10825 VDPWR.n1964 VDPWR.n1922 3.04861
R10826 VDPWR.n2749 VDPWR.n2746 3.04861
R10827 VDPWR.n854 VDPWR.n822 3.04861
R10828 VDPWR.n1441 VDPWR.n1440 3.01588
R10829 VDPWR.n1471 VDPWR.n1309 3.01588
R10830 VDPWR.n1411 VDPWR.n1410 3.01588
R10831 VDPWR.n1570 VDPWR.n1524 3.01588
R10832 VDPWR.n1741 VDPWR.n1740 3.01588
R10833 VDPWR.n1771 VDPWR.n1770 3.01588
R10834 VDPWR.n1776 VDPWR.n1775 3.01588
R10835 VDPWR.n1799 VDPWR.n1237 3.01588
R10836 VDPWR.n1804 VDPWR.n1803 3.01588
R10837 VDPWR.n2011 VDPWR.n1158 3.01588
R10838 VDPWR.n2020 VDPWR.n1154 3.01588
R10839 VDPWR.n1150 VDPWR.n1149 3.01588
R10840 VDPWR.n1634 VDPWR.n1633 3.01588
R10841 VDPWR.n2147 VDPWR.n2077 3.01588
R10842 VDPWR.n1875 VDPWR.n1209 3.01226
R10843 VDPWR.n2867 VDPWR.n2866 3.01226
R10844 VDPWR.n2608 VDPWR.n2605 3.01226
R10845 VDPWR.n2566 VDPWR.n2547 3.01226
R10846 VDPWR.n894 VDPWR.n892 3.01226
R10847 VDPWR.n3044 VDPWR.n897 3.01226
R10848 VDPWR.n1961 VDPWR.n1926 2.99733
R10849 VDPWR.n852 VDPWR.n824 2.99733
R10850 VDPWR.n1205 VDPWR.n1201 2.91308
R10851 VDPWR.n1205 VDPWR.n1204 2.91308
R10852 VDPWR.n2565 VDPWR.n2559 2.91308
R10853 VDPWR.n2565 VDPWR.n2564 2.91308
R10854 VDPWR.n1924 VDPWR.n1922 2.87861
R10855 VDPWR.n2210 VDPWR.n2209 2.8567
R10856 VDPWR.n709 VDPWR.n708 2.84665
R10857 VDPWR.n712 VDPWR.n708 2.84665
R10858 VDPWR.n707 VDPWR.n706 2.84665
R10859 VDPWR.n712 VDPWR.n707 2.84665
R10860 VDPWR.n694 VDPWR.n693 2.84665
R10861 VDPWR.n697 VDPWR.n693 2.84665
R10862 VDPWR.n692 VDPWR.n690 2.84665
R10863 VDPWR.n697 VDPWR.n692 2.84665
R10864 VDPWR.n678 VDPWR.n677 2.84665
R10865 VDPWR.n681 VDPWR.n677 2.84665
R10866 VDPWR.n676 VDPWR.n674 2.84665
R10867 VDPWR.n681 VDPWR.n676 2.84665
R10868 VDPWR.n664 VDPWR.n663 2.84665
R10869 VDPWR.n665 VDPWR.n664 2.84665
R10870 VDPWR.n667 VDPWR.n666 2.84665
R10871 VDPWR.n666 VDPWR.n665 2.84665
R10872 VDPWR.n520 VDPWR.n519 2.84665
R10873 VDPWR.n523 VDPWR.n519 2.84665
R10874 VDPWR.n518 VDPWR.n517 2.84665
R10875 VDPWR.n523 VDPWR.n518 2.84665
R10876 VDPWR.n505 VDPWR.n504 2.84665
R10877 VDPWR.n508 VDPWR.n504 2.84665
R10878 VDPWR.n503 VDPWR.n501 2.84665
R10879 VDPWR.n508 VDPWR.n503 2.84665
R10880 VDPWR.n489 VDPWR.n488 2.84665
R10881 VDPWR.n492 VDPWR.n488 2.84665
R10882 VDPWR.n487 VDPWR.n485 2.84665
R10883 VDPWR.n492 VDPWR.n487 2.84665
R10884 VDPWR.n472 VDPWR.n471 2.84665
R10885 VDPWR.n475 VDPWR.n471 2.84665
R10886 VDPWR.n470 VDPWR.n469 2.84665
R10887 VDPWR.n475 VDPWR.n470 2.84665
R10888 VDPWR.n406 VDPWR.n405 2.84665
R10889 VDPWR.n411 VDPWR.n406 2.84665
R10890 VDPWR.n408 VDPWR.n407 2.84665
R10891 VDPWR.n411 VDPWR.n407 2.84665
R10892 VDPWR.n386 VDPWR.n385 2.84665
R10893 VDPWR.n382 VDPWR.n378 2.84665
R10894 VDPWR.n398 VDPWR.n397 2.84665
R10895 VDPWR.n394 VDPWR.n390 2.84665
R10896 VDPWR.n451 VDPWR.n450 2.84665
R10897 VDPWR.n454 VDPWR.n450 2.84665
R10898 VDPWR.n449 VDPWR.n447 2.84665
R10899 VDPWR.n454 VDPWR.n449 2.84665
R10900 VDPWR.n435 VDPWR.n434 2.84665
R10901 VDPWR.n438 VDPWR.n434 2.84665
R10902 VDPWR.n433 VDPWR.n431 2.84665
R10903 VDPWR.n438 VDPWR.n433 2.84665
R10904 VDPWR.n421 VDPWR.n420 2.84665
R10905 VDPWR.n422 VDPWR.n421 2.84665
R10906 VDPWR.n424 VDPWR.n423 2.84665
R10907 VDPWR.n423 VDPWR.n422 2.84665
R10908 VDPWR.n764 VDPWR.n763 2.84665
R10909 VDPWR.n767 VDPWR.n763 2.84665
R10910 VDPWR.n762 VDPWR.n761 2.84665
R10911 VDPWR.n767 VDPWR.n762 2.84665
R10912 VDPWR.n3154 VDPWR.n3152 2.84665
R10913 VDPWR.n3159 VDPWR.n3154 2.84665
R10914 VDPWR.n3156 VDPWR.n3155 2.84665
R10915 VDPWR.n3159 VDPWR.n3155 2.84665
R10916 VDPWR.n3138 VDPWR.n3136 2.84665
R10917 VDPWR.n3143 VDPWR.n3138 2.84665
R10918 VDPWR.n3140 VDPWR.n3139 2.84665
R10919 VDPWR.n3143 VDPWR.n3139 2.84665
R10920 VDPWR.n3123 VDPWR.n3122 2.84665
R10921 VDPWR.n3126 VDPWR.n3122 2.84665
R10922 VDPWR.n3121 VDPWR.n3120 2.84665
R10923 VDPWR.n3126 VDPWR.n3121 2.84665
R10924 VDPWR.n1260 VDPWR.n1258 2.8165
R10925 VDPWR.n2474 VDPWR.n2472 2.8165
R10926 VDPWR.n1377 VDPWR.n1349 2.6965
R10927 VDPWR.n1705 VDPWR.n1682 2.6965
R10928 VDPWR.n1624 VDPWR.n1623 2.6965
R10929 VDPWR.n3060 VDPWR.n879 2.69256
R10930 VDPWR.n1440 VDPWR.n1321 2.64665
R10931 VDPWR.n1474 VDPWR.n1309 2.64665
R10932 VDPWR.n1412 VDPWR.n1411 2.64665
R10933 VDPWR.n1567 VDPWR.n1524 2.64665
R10934 VDPWR.n1742 VDPWR.n1741 2.64665
R10935 VDPWR.n1770 VDPWR.n1255 2.64665
R10936 VDPWR.n1777 VDPWR.n1776 2.64665
R10937 VDPWR.n1802 VDPWR.n1237 2.64665
R10938 VDPWR.n1805 VDPWR.n1804 2.64665
R10939 VDPWR.n1168 VDPWR.n1158 2.64665
R10940 VDPWR.n2029 VDPWR.n1150 2.64665
R10941 VDPWR.n1633 VDPWR.n1632 2.64665
R10942 VDPWR.n2141 VDPWR.n2079 2.64665
R10943 VDPWR.n2145 VDPWR.n2079 2.64665
R10944 VDPWR.n2150 VDPWR.n2077 2.64665
R10945 VDPWR.n1987 VDPWR.n1986 2.63579
R10946 VDPWR.n1326 VDPWR.n1324 2.63539
R10947 VDPWR.n1353 VDPWR.n1351 2.63539
R10948 VDPWR.n1356 VDPWR.n1354 2.63539
R10949 VDPWR.n1360 VDPWR.n1358 2.63539
R10950 VDPWR.n1365 VDPWR.n1363 2.63539
R10951 VDPWR.n1540 VDPWR.n1538 2.63539
R10952 VDPWR.n1543 VDPWR.n1541 2.63539
R10953 VDPWR.n1686 VDPWR.n1684 2.63539
R10954 VDPWR.n1689 VDPWR.n1687 2.63539
R10955 VDPWR.n1693 VDPWR.n1691 2.63539
R10956 VDPWR.n1698 VDPWR.n1696 2.63539
R10957 VDPWR.n1208 VDPWR.n1206 2.63539
R10958 VDPWR.n1895 VDPWR.n1893 2.63539
R10959 VDPWR.n1606 VDPWR.n1604 2.63539
R10960 VDPWR.n1612 VDPWR.n1610 2.63539
R10961 VDPWR.n1615 VDPWR.n1613 2.63539
R10962 VDPWR.n1619 VDPWR.n1617 2.63539
R10963 VDPWR.n1939 VDPWR.n1937 2.63539
R10964 VDPWR.n1942 VDPWR.n1940 2.63539
R10965 VDPWR.n2098 VDPWR.n2096 2.63539
R10966 VDPWR.n2101 VDPWR.n2099 2.63539
R10967 VDPWR.n1071 VDPWR.n1069 2.63539
R10968 VDPWR.n1074 VDPWR.n1072 2.63539
R10969 VDPWR.n2731 VDPWR.n2729 2.63539
R10970 VDPWR.n2734 VDPWR.n2732 2.63539
R10971 VDPWR.n932 VDPWR.n930 2.63539
R10972 VDPWR.n2972 VDPWR.n2970 2.63539
R10973 VDPWR.n2552 VDPWR.n2550 2.63539
R10974 VDPWR.n2555 VDPWR.n2553 2.63539
R10975 VDPWR.n2597 VDPWR.n2595 2.63539
R10976 VDPWR.n891 VDPWR.n889 2.63539
R10977 VDPWR.n2991 VDPWR.n2989 2.63539
R10978 VDPWR.n2999 VDPWR.n2997 2.63539
R10979 VDPWR.n819 VDPWR.n817 2.63539
R10980 VDPWR.n2373 VDPWR.n2371 2.63539
R10981 VDPWR.n2376 VDPWR.n2374 2.63539
R10982 VDPWR.n834 VDPWR.n832 2.63539
R10983 VDPWR.n838 VDPWR.n836 2.63539
R10984 VDPWR.n2232 VDPWR.n2231 2.62345
R10985 VDPWR.n1926 VDPWR.n1925 2.61352
R10986 VDPWR.n1034 VDPWR.n1031 2.56175
R10987 VDPWR.n577 VDPWR.n576 2.54018
R10988 VDPWR.n556 VDPWR.n555 2.54018
R10989 VDPWR.n297 VDPWR.n296 2.54018
R10990 VDPWR.n276 VDPWR.n275 2.54018
R10991 VDPWR.n796 VDPWR.n793 2.54018
R10992 VDPWR.n39 VDPWR.n38 2.54018
R10993 VDPWR.n18 VDPWR.n17 2.54018
R10994 VDPWR.n3083 VDPWR.n797 2.3878
R10995 VDPWR.n824 VDPWR.n823 2.37764
R10996 VDPWR.n1325 VDPWR.n1324 2.37495
R10997 VDPWR.n1355 VDPWR.n1354 2.37495
R10998 VDPWR.n1352 VDPWR.n1351 2.37495
R10999 VDPWR.n1364 VDPWR.n1363 2.37495
R11000 VDPWR.n1359 VDPWR.n1358 2.37495
R11001 VDPWR.n1542 VDPWR.n1541 2.37495
R11002 VDPWR.n1539 VDPWR.n1538 2.37495
R11003 VDPWR.n1688 VDPWR.n1687 2.37495
R11004 VDPWR.n1685 VDPWR.n1684 2.37495
R11005 VDPWR.n1697 VDPWR.n1696 2.37495
R11006 VDPWR.n1692 VDPWR.n1691 2.37495
R11007 VDPWR.n1894 VDPWR.n1893 2.37495
R11008 VDPWR.n1207 VDPWR.n1206 2.37495
R11009 VDPWR.n1611 VDPWR.n1610 2.37495
R11010 VDPWR.n1605 VDPWR.n1604 2.37495
R11011 VDPWR.n1618 VDPWR.n1617 2.37495
R11012 VDPWR.n1614 VDPWR.n1613 2.37495
R11013 VDPWR.n1941 VDPWR.n1940 2.37495
R11014 VDPWR.n1938 VDPWR.n1937 2.37495
R11015 VDPWR.n2100 VDPWR.n2099 2.37495
R11016 VDPWR.n2097 VDPWR.n2096 2.37495
R11017 VDPWR.n1073 VDPWR.n1072 2.37495
R11018 VDPWR.n1070 VDPWR.n1069 2.37495
R11019 VDPWR.n2733 VDPWR.n2732 2.37495
R11020 VDPWR.n2730 VDPWR.n2729 2.37495
R11021 VDPWR.n2971 VDPWR.n2970 2.37495
R11022 VDPWR.n931 VDPWR.n930 2.37495
R11023 VDPWR.n2554 VDPWR.n2553 2.37495
R11024 VDPWR.n2551 VDPWR.n2550 2.37495
R11025 VDPWR.n2596 VDPWR.n2595 2.37495
R11026 VDPWR.n890 VDPWR.n889 2.37495
R11027 VDPWR.n2998 VDPWR.n2997 2.37495
R11028 VDPWR.n2990 VDPWR.n2989 2.37495
R11029 VDPWR.n818 VDPWR.n817 2.37495
R11030 VDPWR.n2375 VDPWR.n2374 2.37495
R11031 VDPWR.n2372 VDPWR.n2371 2.37495
R11032 VDPWR.n837 VDPWR.n836 2.37495
R11033 VDPWR.n833 VDPWR.n832 2.37495
R11034 VDPWR.n602 VDPWR.n598 2.33701
R11035 VDPWR.n590 VDPWR.n589 2.33701
R11036 VDPWR.n576 VDPWR.n575 2.33701
R11037 VDPWR.n556 VDPWR.n550 2.33701
R11038 VDPWR.n322 VDPWR.n318 2.33701
R11039 VDPWR.n310 VDPWR.n309 2.33701
R11040 VDPWR.n296 VDPWR.n295 2.33701
R11041 VDPWR.n276 VDPWR.n270 2.33701
R11042 VDPWR.n1105 VDPWR.n1104 2.33701
R11043 VDPWR.n2886 VDPWR.n2885 2.33701
R11044 VDPWR.n3061 VDPWR.n878 2.33701
R11045 VDPWR.n2400 VDPWR.n2399 2.33701
R11046 VDPWR.n64 VDPWR.n60 2.33701
R11047 VDPWR.n52 VDPWR.n51 2.33701
R11048 VDPWR.n38 VDPWR.n37 2.33701
R11049 VDPWR.n18 VDPWR.n12 2.33701
R11050 VDPWR.n1434 VDPWR.n1327 2.32777
R11051 VDPWR.n1128 VDPWR.n1127 2.32777
R11052 VDPWR.n1834 VDPWR.n1833 2.28432
R11053 VDPWR.n2749 VDPWR.n2726 2.28407
R11054 VDPWR.n2749 VDPWR.n2728 2.28407
R11055 VDPWR.n2094 VDPWR.n2092 2.28374
R11056 VDPWR.n1155 VDPWR.n1154 2.27742
R11057 VDPWR.n1920 VDPWR.n1919 2.25932
R11058 VDPWR.n1986 VDPWR.n1184 2.25932
R11059 VDPWR.n2565 VDPWR.n2561 2.25293
R11060 VDPWR.n3090 VDPWR.n3089 2.23542
R11061 VDPWR.n2909 VDPWR.n2908 2.22199
R11062 VDPWR.n3118 VDPWR.n3117 2.16151
R11063 VDPWR.n402 VDPWR.n401 2.13883
R11064 VDPWR.n483 VDPWR.n482 2.13544
R11065 VDPWR.n584 VDPWR.n577 2.13383
R11066 VDPWR.n555 VDPWR.n554 2.13383
R11067 VDPWR.n304 VDPWR.n297 2.13383
R11068 VDPWR.n275 VDPWR.n274 2.13383
R11069 VDPWR.n3085 VDPWR.n796 2.13383
R11070 VDPWR.n46 VDPWR.n39 2.13383
R11071 VDPWR.n17 VDPWR.n16 2.13383
R11072 VDPWR.n1057 VDPWR.n1056 2.0932
R11073 VDPWR.n2740 VDPWR.n2739 2.07374
R11074 VDPWR.n2727 VDPWR.n1006 2.07374
R11075 VDPWR.n598 VDPWR.n596 2.03225
R11076 VDPWR.n589 VDPWR.n588 2.03225
R11077 VDPWR.n575 VDPWR.n574 2.03225
R11078 VDPWR.n550 VDPWR.n548 2.03225
R11079 VDPWR.n318 VDPWR.n316 2.03225
R11080 VDPWR.n309 VDPWR.n308 2.03225
R11081 VDPWR.n295 VDPWR.n294 2.03225
R11082 VDPWR.n270 VDPWR.n268 2.03225
R11083 VDPWR.n2885 VDPWR.n2884 2.03225
R11084 VDPWR.n2399 VDPWR.n2398 2.03225
R11085 VDPWR.n60 VDPWR.n58 2.03225
R11086 VDPWR.n51 VDPWR.n50 2.03225
R11087 VDPWR.n37 VDPWR.n36 2.03225
R11088 VDPWR.n12 VDPWR.n10 2.03225
R11089 VDPWR.n1201 VDPWR.n1199 2.01703
R11090 VDPWR.n1204 VDPWR.n1202 2.01703
R11091 VDPWR.n2559 VDPWR.n2557 2.01703
R11092 VDPWR.n2564 VDPWR.n2562 2.01703
R11093 VDPWR.n3092 VDPWR.n3091 1.98145
R11094 VDPWR.n798 VDPWR.n797 1.98145
R11095 VDPWR.n482 VDPWR.n467 1.95379
R11096 VDPWR.n2187 VDPWR.n2186 1.88902
R11097 VDPWR.n2305 VDPWR.n1034 1.88902
R11098 VDPWR.n1203 VDPWR.n1202 1.88416
R11099 VDPWR.n1200 VDPWR.n1199 1.88416
R11100 VDPWR.n2563 VDPWR.n2562 1.88416
R11101 VDPWR.n2558 VDPWR.n2557 1.88416
R11102 VDPWR.n1643 VDPWR.n1630 1.88325
R11103 VDPWR.n1403 VDPWR.n1402 1.88295
R11104 VDPWR.n1733 VDPWR.n1732 1.88295
R11105 VDPWR.n661 VDPWR.n657 1.88285
R11106 VDPWR.n478 VDPWR.n477 1.88285
R11107 VDPWR.n418 VDPWR.n414 1.88285
R11108 VDPWR.n3129 VDPWR.n3128 1.88285
R11109 VDPWR.n2852 VDPWR.n967 1.88285
R11110 VDPWR.n1377 VDPWR.n1376 1.85065
R11111 VDPWR.n1379 VDPWR.n1343 1.85065
R11112 VDPWR.n1507 VDPWR.n1506 1.85065
R11113 VDPWR.n1705 VDPWR.n1704 1.85065
R11114 VDPWR.n1707 VDPWR.n1279 1.85065
R11115 VDPWR.n1132 VDPWR.n1131 1.85065
R11116 VDPWR.n1624 VDPWR.n1601 1.85065
R11117 VDPWR.n1665 VDPWR.n1625 1.85065
R11118 VDPWR.n2118 VDPWR.n2117 1.85065
R11119 VDPWR.n2456 VDPWR.n2454 1.85065
R11120 VDPWR.n2793 VDPWR.n984 1.82907
R11121 VDPWR.n2628 VDPWR.n2627 1.82907
R11122 VDPWR.n1505 VDPWR.n1504 1.81289
R11123 VDPWR.n2116 VDPWR.n2115 1.81289
R11124 VDPWR.n2483 VDPWR 1.79885
R11125 VDPWR.n654 VDPWR.n653 1.753
R11126 VDPWR.n374 VDPWR.n373 1.753
R11127 VDPWR.n116 VDPWR.n115 1.753
R11128 VDPWR.n1997 VDPWR.n1181 1.73737
R11129 VDPWR.n2325 VDPWR.n1018 1.73737
R11130 VDPWR.n2267 VDPWR.n1068 1.73737
R11131 VDPWR.n2216 VDPWR.n2210 1.69306
R11132 VDPWR.n2271 VDPWR.n1065 1.69306
R11133 VDPWR.n3031 VDPWR.n870 1.69188
R11134 VDPWR.n3033 VDPWR.n870 1.69188
R11135 VDPWR.n2933 VDPWR.n2932 1.69188
R11136 VDPWR.n2932 VDPWR.n2931 1.69188
R11137 VDPWR.n2290 VDPWR.n2289 1.69188
R11138 VDPWR.n2291 VDPWR.n2290 1.69188
R11139 VDPWR.n1974 VDPWR.n1973 1.69188
R11140 VDPWR.n1975 VDPWR.n1974 1.69188
R11141 VDPWR.n1860 VDPWR.n1191 1.69188
R11142 VDPWR.n1857 VDPWR.n1191 1.69188
R11143 VDPWR.n1588 VDPWR.n1285 1.69188
R11144 VDPWR.n1588 VDPWR.n1587 1.69188
R11145 VDPWR.n3067 VDPWR.n873 1.69188
R11146 VDPWR.n3067 VDPWR.n3066 1.69188
R11147 VDPWR.n2897 VDPWR.n872 1.69188
R11148 VDPWR.n2879 VDPWR.n872 1.69188
R11149 VDPWR.n2331 VDPWR.n1013 1.69188
R11150 VDPWR.n2331 VDPWR.n2330 1.69188
R11151 VDPWR.n2006 VDPWR.n2005 1.69188
R11152 VDPWR.n2007 VDPWR.n2006 1.69188
R11153 VDPWR.n1821 VDPWR.n1820 1.69188
R11154 VDPWR.n1820 VDPWR.n1819 1.69188
R11155 VDPWR.n1493 VDPWR.n1492 1.69188
R11156 VDPWR.n1492 VDPWR.n1491 1.69188
R11157 VDPWR.n2661 VDPWR.n974 1.69188
R11158 VDPWR.n2664 VDPWR.n974 1.69188
R11159 VDPWR.n2845 VDPWR.n2844 1.69188
R11160 VDPWR.n2844 VDPWR.n2843 1.69188
R11161 VDPWR.n2249 VDPWR.n1092 1.69188
R11162 VDPWR.n2249 VDPWR.n2248 1.69188
R11163 VDPWR.n2033 VDPWR.n1091 1.69188
R11164 VDPWR.n2036 VDPWR.n1091 1.69188
R11165 VDPWR.n1785 VDPWR.n1784 1.69188
R11166 VDPWR.n1784 VDPWR.n1783 1.69188
R11167 VDPWR.n1457 VDPWR.n1456 1.69188
R11168 VDPWR.n1456 VDPWR.n1455 1.69188
R11169 VDPWR.n2756 VDPWR.n2755 1.69188
R11170 VDPWR.n2755 VDPWR.n2754 1.69188
R11171 VDPWR.n2125 VDPWR.n1009 1.69188
R11172 VDPWR.n2111 VDPWR.n1009 1.69188
R11173 VDPWR.n1672 VDPWR.n1595 1.69188
R11174 VDPWR.n1672 VDPWR.n1671 1.69188
R11175 VDPWR.n1715 VDPWR.n1714 1.69188
R11176 VDPWR.n1714 VDPWR.n1713 1.69188
R11177 VDPWR.n1385 VDPWR.n1283 1.69188
R11178 VDPWR.n1372 VDPWR.n1283 1.69188
R11179 VDPWR.n2719 VDPWR.n2337 1.69188
R11180 VDPWR.n3007 VDPWR.n2982 1.69188
R11181 VDPWR.n3004 VDPWR.n2982 1.69188
R11182 VDPWR.n2981 VDPWR.n924 1.69188
R11183 VDPWR.n2981 VDPWR.n2980 1.69188
R11184 VDPWR.n2256 VDPWR.n1080 1.69188
R11185 VDPWR.n2257 VDPWR.n2256 1.69188
R11186 VDPWR.n1954 VDPWR.n1089 1.69188
R11187 VDPWR.n1944 VDPWR.n1089 1.69188
R11188 VDPWR.n1904 VDPWR.n1194 1.69188
R11189 VDPWR.n1904 VDPWR.n1903 1.69188
R11190 VDPWR.n1555 VDPWR.n1531 1.69188
R11191 VDPWR.n1545 VDPWR.n1531 1.69188
R11192 VDPWR.n2691 VDPWR.n989 1.69188
R11193 VDPWR.n2694 VDPWR.n989 1.69188
R11194 VDPWR.n2806 VDPWR.n2805 1.69188
R11195 VDPWR.n2805 VDPWR.n2804 1.69188
R11196 VDPWR.n2160 VDPWR.n2159 1.69188
R11197 VDPWR.n2159 VDPWR.n2158 1.69188
R11198 VDPWR.n2072 VDPWR.n1117 1.69188
R11199 VDPWR.n2072 VDPWR.n2071 1.69188
R11200 VDPWR.n1755 VDPWR.n1754 1.69188
R11201 VDPWR.n1754 VDPWR.n1753 1.69188
R11202 VDPWR.n1424 VDPWR.n1423 1.69188
R11203 VDPWR.n1423 VDPWR.n1422 1.69188
R11204 VDPWR.t996 VDPWR 1.67895
R11205 VDPWR.t126 VDPWR 1.67895
R11206 VDPWR.n884 VDPWR.n879 1.67669
R11207 VDPWR.n1507 VDPWR.n1505 1.66186
R11208 VDPWR.n2118 VDPWR.n2116 1.66186
R11209 VDPWR.n2491 VDPWR.n2453 1.64857
R11210 VDPWR.n1378 VDPWR.n1377 1.6241
R11211 VDPWR.n1389 VDPWR.n1343 1.6241
R11212 VDPWR.n1506 VDPWR.n1294 1.6241
R11213 VDPWR.n1708 VDPWR.n1705 1.6241
R11214 VDPWR.n1719 VDPWR.n1279 1.6241
R11215 VDPWR.n1666 VDPWR.n1624 1.6241
R11216 VDPWR.n1655 VDPWR.n1625 1.6241
R11217 VDPWR.n2117 VDPWR.n2084 1.6241
R11218 VDPWR.n2486 VDPWR.n2456 1.6241
R11219 VDPWR.n1404 VDPWR.n1403 1.62167
R11220 VDPWR.n1734 VDPWR.n1733 1.62167
R11221 VDPWR.n1640 VDPWR.n1630 1.62136
R11222 VDPWR.n3172 VDPWR.n117 1.59405
R11223 VDPWR.n754 VDPWR.n753 1.57294
R11224 VDPWR.n747 VDPWR.t372 1.53603
R11225 VDPWR.n744 VDPWR.t372 1.53603
R11226 VDPWR.n531 VDPWR.n530 1.51493
R11227 VDPWR.n1181 VDPWR.n1179 1.51082
R11228 VDPWR.n2211 VDPWR.n1018 1.51082
R11229 VDPWR.n1068 VDPWR.n1066 1.51082
R11230 VDPWR.n758 VDPWR 1.48239
R11231 VDPWR.n573 VDPWR.n571 1.46504
R11232 VDPWR.n293 VDPWR.n291 1.46504
R11233 VDPWR.n35 VDPWR.n33 1.46504
R11234 VDPWR.n532 VDPWR.n253 1.42384
R11235 VDPWR.n646 VDPWR.n546 1.4005
R11236 VDPWR.n366 VDPWR.n266 1.4005
R11237 VDPWR.n2875 VDPWR.n2874 1.4005
R11238 VDPWR.n2768 VDPWR.n2767 1.4005
R11239 VDPWR.n108 VDPWR.n8 1.4005
R11240 VDPWR.n1133 VDPWR.n1132 1.39755
R11241 VDPWR.n2202 VDPWR.n2200 1.36443
R11242 VDPWR.n2283 VDPWR.n2282 1.36443
R11243 VDPWR.n758 VDPWR.n757 1.34339
R11244 VDPWR.n2883 VDPWR.n961 1.3232
R11245 VDPWR.n402 VDPWR.n389 1.28133
R11246 VDPWR.n1926 VDPWR.n1924 1.2502
R11247 VDPWR.n257 VDPWR.n256 1.16828
R11248 VDPWR.n3133 VDPWR.n3132 1.16528
R11249 VDPWR.n755 VDPWR.n118 1.15151
R11250 VDPWR.n703 VDPWR.n702 1.143
R11251 VDPWR.n687 VDPWR.n686 1.143
R11252 VDPWR.n514 VDPWR.n513 1.143
R11253 VDPWR.n498 VDPWR.n497 1.143
R11254 VDPWR.n460 VDPWR.n459 1.143
R11255 VDPWR.n444 VDPWR.n443 1.143
R11256 VDPWR.n3165 VDPWR.n3164 1.143
R11257 VDPWR.n3149 VDPWR.n3148 1.143
R11258 VDPWR.n719 VDPWR.n718 1.13925
R11259 VDPWR.n530 VDPWR.n529 1.13925
R11260 VDPWR.n466 VDPWR.n465 1.13925
R11261 VDPWR.n3171 VDPWR.n3170 1.13925
R11262 VDPWR.n3114 VDPWR.n3113 1.13717
R11263 VDPWR.n671 VDPWR.n670 1.13675
R11264 VDPWR.n482 VDPWR.n481 1.13675
R11265 VDPWR.n428 VDPWR.n427 1.13675
R11266 VDPWR.n715 VDPWR.n714 1.12991
R11267 VDPWR.n691 VDPWR.n689 1.12991
R11268 VDPWR.n683 VDPWR.n675 1.12991
R11269 VDPWR.n526 VDPWR.n525 1.12991
R11270 VDPWR.n502 VDPWR.n500 1.12991
R11271 VDPWR.n494 VDPWR.n486 1.12991
R11272 VDPWR.n462 VDPWR.n413 1.12991
R11273 VDPWR.n448 VDPWR.n446 1.12991
R11274 VDPWR.n440 VDPWR.n432 1.12991
R11275 VDPWR.n3167 VDPWR.n769 1.12991
R11276 VDPWR.n3153 VDPWR.n3151 1.12991
R11277 VDPWR.n3145 VDPWR.n3137 1.12991
R11278 VDPWR.n2472 VDPWR.n2471 1.11173
R11279 VDPWR.n2397 VDPWR.n2359 1.08324
R11280 VDPWR.n721 VDPWR.n720 1.06914
R11281 VDPWR.n595 VDPWR 1.06099
R11282 VDPWR.n315 VDPWR 1.06099
R11283 VDPWR.n57 VDPWR 1.06099
R11284 VDPWR.n1368 VDPWR.n1367 1.05773
R11285 VDPWR.n1701 VDPWR.n1700 1.05773
R11286 VDPWR.n1622 VDPWR.n1603 1.05773
R11287 VDPWR.n2452 VDPWR.n2451 1.05773
R11288 VDPWR.n2221 VDPWR.n2220 1.04968
R11289 VDPWR.n2276 VDPWR.n2275 1.04968
R11290 VDPWR.n2739 VDPWR.n2726 0.992049
R11291 VDPWR.n2728 VDPWR.n1006 0.992049
R11292 VDPWR.n3117 VDPWR.n117 0.973454
R11293 VDPWR.n2049 VDPWR.n1130 0.899674
R11294 VDPWR VDPWR.n118 0.891339
R11295 VDPWR.n756 VDPWR.n755 0.884173
R11296 VDPWR.n2176 VDPWR.n1104 0.863992
R11297 VDPWR.n376 VDPWR.n375 0.853
R11298 VDPWR.n3102 VDPWR.n782 0.853
R11299 VDPWR.n2508 VDPWR.n2507 0.853
R11300 VDPWR.n2537 VDPWR.n2536 0.853
R11301 VDPWR.n2392 VDPWR.n2339 0.853
R11302 VDPWR.n3074 VDPWR.n3073 0.853
R11303 VDPWR.n688 VDPWR.n687 0.849559
R11304 VDPWR.n445 VDPWR.n444 0.849559
R11305 VDPWR.n499 VDPWR.n498 0.849559
R11306 VDPWR.n531 VDPWR.n377 0.843267
R11307 VDPWR.n2422 VDPWR.n2421 0.813198
R11308 VDPWR.n2520 VDPWR.n2519 0.813198
R11309 VDPWR.n532 VDPWR.n531 0.810458
R11310 VDPWR VDPWR.n3116 0.778686
R11311 VDPWR.n822 VDPWR 0.777643
R11312 VDPWR.n739 VDPWR.n738 0.7755
R11313 VDPWR.n672 VDPWR.n671 0.770881
R11314 VDPWR.n429 VDPWR.n428 0.770881
R11315 VDPWR.n403 VDPWR.n402 0.767167
R11316 VDPWR.n375 VDPWR.n374 0.763912
R11317 VDPWR.n633 VDPWR.n562 0.753441
R11318 VDPWR.n353 VDPWR.n282 0.753441
R11319 VDPWR.n1877 VDPWR.n1876 0.753441
R11320 VDPWR.n95 VDPWR.n24 0.753441
R11321 VDPWR.n1842 VDPWR.n1841 0.740996
R11322 VDPWR.n461 VDPWR.n460 0.73614
R11323 VDPWR.n704 VDPWR.n703 0.717512
R11324 VDPWR.n515 VDPWR.n514 0.717512
R11325 VDPWR.n2938 VDPWR.n2937 0.706789
R11326 VDPWR.n758 VDPWR.n118 0.70421
R11327 VDPWR.n255 VDPWR 0.659186
R11328 VDPWR.n865 VDPWR.n814 0.65125
R11329 VDPWR.n1499 VDPWR.n1296 0.635211
R11330 VDPWR.n1576 VDPWR.n1520 0.635211
R11331 VDPWR.n1865 VDPWR.n1213 0.635211
R11332 VDPWR.n2185 VDPWR.n2184 0.635211
R11333 VDPWR.n2316 VDPWR.n2315 0.635211
R11334 VDPWR.n2310 VDPWR.n2309 0.635211
R11335 VDPWR.n2904 VDPWR.n2903 0.635211
R11336 VDPWR.n2937 VDPWR.n939 0.635211
R11337 VDPWR.n2940 VDPWR.n2939 0.635211
R11338 VDPWR.n2947 VDPWR.n2946 0.635211
R11339 VDPWR.n2226 VDPWR.n2203 0.630008
R11340 VDPWR.n1056 VDPWR.n1051 0.630008
R11341 VDPWR.n2285 VDPWR.n2284 0.630008
R11342 VDPWR.n656 VDPWR.n537 0.624567
R11343 VDPWR.n543 VDPWR.n541 0.6005
R11344 VDPWR.n263 VDPWR.n261 0.6005
R11345 VDPWR.n5 VDPWR.n3 0.6005
R11346 VDPWR.n2207 VDPWR.n2205 0.52509
R11347 VDPWR.n467 VDPWR.n466 0.518882
R11348 VDPWR.n655 VDPWR.n654 0.511794
R11349 VDPWR.n3178 VDPWR.n116 0.511794
R11350 VDPWR.n2336 VDPWR.n2335 0.500125
R11351 VDPWR.n1594 VDPWR.n1593 0.500125
R11352 VDPWR.n1675 VDPWR.n1674 0.500125
R11353 VDPWR.n1596 VDPWR.n1090 0.500125
R11354 VDPWR.n2540 VDPWR.n2539 0.500125
R11355 VDPWR.n2504 VDPWR.n2501 0.500125
R11356 VDPWR.n142 VDPWR.n141 0.465384
R11357 VDPWR.n654 VDPWR 0.460219
R11358 VDPWR.n374 VDPWR 0.460219
R11359 VDPWR.n116 VDPWR 0.460219
R11360 VDPWR.n3091 VDPWR.n3090 0.457643
R11361 VDPWR.n376 VDPWR.n257 0.45408
R11362 VDPWR.n719 VDPWR.n704 0.405788
R11363 VDPWR.n649 VDPWR.n541 0.4005
R11364 VDPWR.n369 VDPWR.n261 0.4005
R11365 VDPWR.n111 VDPWR.n3 0.4005
R11366 VDPWR.n2253 VDPWR.n1046 0.3805
R11367 VDPWR.n1908 VDPWR.n1907 0.3805
R11368 VDPWR.n1590 VDPWR.n1589 0.3805
R11369 VDPWR.n1011 VDPWR.n943 0.3805
R11370 VDPWR.n3072 VDPWR.n3071 0.3805
R11371 VDPWR.n3069 VDPWR.n3068 0.3805
R11372 VDPWR.n2252 VDPWR.n1012 0.3805
R11373 VDPWR.n1192 VDPWR.n1162 0.3805
R11374 VDPWR.n1591 VDPWR.n1228 0.3805
R11375 VDPWR.n2333 VDPWR.n2332 0.3805
R11376 VDPWR.n2499 VDPWR.n871 0.3805
R11377 VDPWR.n2251 VDPWR.n2250 0.3805
R11378 VDPWR.n1673 VDPWR.n1246 0.3805
R11379 VDPWR.n1592 VDPWR.n1245 0.3805
R11380 VDPWR.n2334 VDPWR.n973 0.3805
R11381 VDPWR.n2506 VDPWR.n2505 0.3805
R11382 VDPWR.n780 VDPWR.n776 0.3805
R11383 VDPWR.n3109 VDPWR.n3108 0.3805
R11384 VDPWR.n2255 VDPWR.n2254 0.3805
R11385 VDPWR.n1906 VDPWR.n1905 0.3805
R11386 VDPWR.n1284 VDPWR.n1193 0.3805
R11387 VDPWR.n1010 VDPWR.n923 0.3805
R11388 VDPWR.n3070 VDPWR.n775 0.3805
R11389 VDPWR.n3111 VDPWR.n3110 0.3805
R11390 VDPWR.n2504 VDPWR.n2503 0.3805
R11391 VDPWR.n2539 VDPWR.n2538 0.3805
R11392 VDPWR.n2073 VDPWR.n1090 0.3805
R11393 VDPWR.n1674 VDPWR.n1116 0.3805
R11394 VDPWR.n1593 VDPWR.n1267 0.3805
R11395 VDPWR.n2335 VDPWR.n988 0.3805
R11396 VDPWR.n687 VDPWR.n672 0.379066
R11397 VDPWR.n444 VDPWR.n429 0.379066
R11398 VDPWR.n498 VDPWR.n483 0.379066
R11399 VDPWR.n721 VDPWR.n253 0.375001
R11400 VDPWR.n377 VDPWR 0.36983
R11401 VDPWR.n1435 VDPWR.n1323 0.369731
R11402 VDPWR.n1465 VDPWR.n1312 0.369731
R11403 VDPWR.n1466 VDPWR.n1311 0.369731
R11404 VDPWR.n1482 VDPWR.n1481 0.369731
R11405 VDPWR.n1397 VDPWR.n1396 0.369731
R11406 VDPWR.n1402 VDPWR.n1339 0.369731
R11407 VDPWR.n1405 VDPWR.n1404 0.369731
R11408 VDPWR.n1428 VDPWR.n1328 0.369731
R11409 VDPWR.n1575 VDPWR.n1521 0.369731
R11410 VDPWR.n1537 VDPWR.n1528 0.369731
R11411 VDPWR.n1727 VDPWR.n1726 0.369731
R11412 VDPWR.n1732 VDPWR.n1275 0.369731
R11413 VDPWR.n1735 VDPWR.n1734 0.369731
R11414 VDPWR.n1743 VDPWR.n1263 0.369731
R11415 VDPWR.n1769 VDPWR.n1768 0.369731
R11416 VDPWR.n1792 VDPWR.n1791 0.369731
R11417 VDPWR.n1798 VDPWR.n1797 0.369731
R11418 VDPWR.n1810 VDPWR.n1224 0.369731
R11419 VDPWR.n2016 VDPWR.n1156 0.369731
R11420 VDPWR.n1178 VDPWR.n1177 0.369731
R11421 VDPWR.n1153 VDPWR.n1151 0.369731
R11422 VDPWR.n2017 VDPWR.n1155 0.369731
R11423 VDPWR.n2040 VDPWR.n1134 0.369731
R11424 VDPWR.n2027 VDPWR.n2026 0.369731
R11425 VDPWR.n1640 VDPWR.n1639 0.369731
R11426 VDPWR.n2059 VDPWR.n2058 0.369731
R11427 VDPWR.n1649 VDPWR.n1628 0.369731
R11428 VDPWR.n1644 VDPWR.n1643 0.369731
R11429 VDPWR.n2136 VDPWR.n2135 0.369731
R11430 VDPWR.n2140 VDPWR.n2080 0.369731
R11431 VDPWR.n2142 VDPWR.n2141 0.369731
R11432 VDPWR.n2167 VDPWR.n2166 0.369731
R11433 VDPWR.n530 VDPWR.n515 0.360095
R11434 VDPWR.n703 VDPWR.n688 0.348599
R11435 VDPWR.n460 VDPWR.n445 0.348599
R11436 VDPWR.n514 VDPWR.n499 0.348599
R11437 VDPWR.n1028 VDPWR.n1026 0.317855
R11438 VDPWR.n1029 VDPWR.n1028 0.317855
R11439 VDPWR.n751 VDPWR.n739 0.310024
R11440 VDPWR.n605 VDPWR.n596 0.305262
R11441 VDPWR.n624 VDPWR.n623 0.305262
R11442 VDPWR.n574 VDPWR.n573 0.305262
R11443 VDPWR.n583 VDPWR.n582 0.305262
R11444 VDPWR.n559 VDPWR.n548 0.305262
R11445 VDPWR.n325 VDPWR.n316 0.305262
R11446 VDPWR.n344 VDPWR.n343 0.305262
R11447 VDPWR.n294 VDPWR.n293 0.305262
R11448 VDPWR.n303 VDPWR.n302 0.305262
R11449 VDPWR.n279 VDPWR.n268 0.305262
R11450 VDPWR.n750 VDPWR.n740 0.305262
R11451 VDPWR.n1936 VDPWR.n1928 0.305262
R11452 VDPWR.n2179 VDPWR.n1103 0.305262
R11453 VDPWR.n2884 VDPWR.n2883 0.305262
R11454 VDPWR.n2889 VDPWR.n2888 0.305262
R11455 VDPWR.n2763 VDPWR.n2762 0.305262
R11456 VDPWR.n2629 VDPWR.n2628 0.305262
R11457 VDPWR.n885 VDPWR.n884 0.305262
R11458 VDPWR.n3018 VDPWR.n917 0.305262
R11459 VDPWR.n2988 VDPWR.n2987 0.305262
R11460 VDPWR.n2412 VDPWR.n2411 0.305262
R11461 VDPWR.n2417 VDPWR.n2416 0.305262
R11462 VDPWR.n2420 VDPWR.n2349 0.305262
R11463 VDPWR.n2398 VDPWR.n2397 0.305262
R11464 VDPWR.n2404 VDPWR.n2357 0.305262
R11465 VDPWR.n2526 VDPWR.n2525 0.305262
R11466 VDPWR.n2524 VDPWR.n2434 0.305262
R11467 VDPWR.n2515 VDPWR.n2437 0.305262
R11468 VDPWR.n3095 VDPWR.n792 0.305262
R11469 VDPWR.n3080 VDPWR.n798 0.305262
R11470 VDPWR.n865 VDPWR.n864 0.305262
R11471 VDPWR.n831 VDPWR.n830 0.305262
R11472 VDPWR.n67 VDPWR.n58 0.305262
R11473 VDPWR.n86 VDPWR.n85 0.305262
R11474 VDPWR.n36 VDPWR.n35 0.305262
R11475 VDPWR.n45 VDPWR.n44 0.305262
R11476 VDPWR.n21 VDPWR.n10 0.305262
R11477 VDPWR.n2392 VDPWR.n2343 0.297373
R11478 VDPWR.n384 VDPWR.t772 0.27666
R11479 VDPWR.t772 VDPWR.n383 0.27666
R11480 VDPWR.n396 VDPWR.t119 0.27666
R11481 VDPWR.t119 VDPWR.n395 0.27666
R11482 VDPWR.n756 VDPWR.n721 0.262659
R11483 VDPWR.n738 VDPWR.n729 0.2565
R11484 VDPWR.n2773 VDPWR.n2771 0.25148
R11485 VDPWR.n2816 VDPWR.n982 0.246654
R11486 VDPWR.n256 VDPWR 0.245332
R11487 VDPWR.n2561 VDPWR 0.237784
R11488 VDPWR.n1886 VDPWR.n1884 0.231913
R11489 VDPWR.n1368 VDPWR.n1350 0.227049
R11490 VDPWR.n1391 VDPWR.n1341 0.227049
R11491 VDPWR.n1503 VDPWR.n1502 0.227049
R11492 VDPWR.n1516 VDPWR.n1292 0.227049
R11493 VDPWR.n1701 VDPWR.n1683 0.227049
R11494 VDPWR.n1721 VDPWR.n1277 0.227049
R11495 VDPWR.n2000 VDPWR.n1179 0.227049
R11496 VDPWR.n1995 VDPWR.n1994 0.227049
R11497 VDPWR.n2041 VDPWR.n1133 0.227049
R11498 VDPWR.n1603 VDPWR.n1602 0.227049
R11499 VDPWR.n1650 VDPWR.n1627 0.227049
R11500 VDPWR.n2108 VDPWR.n2090 0.227049
R11501 VDPWR.n2134 VDPWR.n2082 0.227049
R11502 VDPWR.n2212 VDPWR.n2211 0.227049
R11503 VDPWR.n1025 VDPWR.n1019 0.227049
R11504 VDPWR.n2270 VDPWR.n1066 0.227049
R11505 VDPWR.n2265 VDPWR.n2264 0.227049
R11506 VDPWR.n2953 VDPWR.n2952 0.227049
R11507 VDPWR.n2959 VDPWR.n929 0.227049
R11508 VDPWR.n2451 VDPWR.n2450 0.227049
R11509 VDPWR.n2485 VDPWR.n2484 0.227049
R11510 VDPWR.n1832 VDPWR 0.217591
R11511 VDPWR.n1839 VDPWR.n1221 0.21207
R11512 VDPWR.n2903 VDPWR.n953 0.21207
R11513 VDPWR.n2941 VDPWR.n937 0.21207
R11514 VDPWR.n2502 VDPWR 0.209323
R11515 VDPWR.n3166 VDPWR.n3165 0.209134
R11516 VDPWR.n3150 VDPWR.n3149 0.206276
R11517 VDPWR.n3107 VDPWR 0.206051
R11518 VDPWR.n2627 VDPWR.n878 0.203675
R11519 VDPWR.n2561 VDPWR 0.200023
R11520 VDPWR.n3116 VDPWR.n770 0.197315
R11521 VDPWR.n3103 VDPWR.n770 0.196829
R11522 VDPWR.n3107 VDPWR.n3106 0.196829
R11523 VDPWR.n2343 VDPWR.n779 0.195044
R11524 VDPWR.n2502 VDPWR.n778 0.195044
R11525 VDPWR.n2777 VDPWR.n1001 0.194439
R11526 VDPWR.n3176 VDPWR 0.189894
R11527 VDPWR.n1970 VDPWR.n1915 0.180304
R11528 VDPWR.n2624 VDPWR.n2622 0.180304
R11529 VDPWR.n1433 VDPWR 0.17983
R11530 VDPWR VDPWR.n2055 0.17983
R11531 VDPWR VDPWR.n1964 0.17983
R11532 VDPWR.n2746 VDPWR 0.17983
R11533 VDPWR VDPWR.n854 0.17983
R11534 VDPWR.n1362 VDPWR 0.179485
R11535 VDPWR.n1695 VDPWR 0.179485
R11536 VDPWR.n1884 VDPWR 0.179485
R11537 VDPWR VDPWR.n1609 0.179485
R11538 VDPWR.n1964 VDPWR 0.179485
R11539 VDPWR.n888 VDPWR 0.179485
R11540 VDPWR.n854 VDPWR 0.179485
R11541 VDPWR.n739 VDPWR.n728 0.176553
R11542 VDPWR VDPWR.n1361 0.172576
R11543 VDPWR VDPWR.n1694 0.172576
R11544 VDPWR.n1616 VDPWR 0.172576
R11545 VDPWR VDPWR.n2103 0.172576
R11546 VDPWR VDPWR.n2736 0.172576
R11547 VDPWR VDPWR.n2560 0.172576
R11548 VDPWR VDPWR.n2378 0.172576
R11549 VDPWR.n536 VDPWR 0.163379
R11550 VDPWR.n2932 VDPWR.n870 0.1603
R11551 VDPWR.n3067 VDPWR.n872 0.1603
R11552 VDPWR.n2844 VDPWR.n974 0.1603
R11553 VDPWR.n2755 VDPWR.n2719 0.1603
R11554 VDPWR.n2982 VDPWR.n2981 0.1603
R11555 VDPWR.n2805 VDPWR.n989 0.1603
R11556 VDPWR.n1765 VDPWR 0.158169
R11557 VDPWR.n1794 VDPWR 0.158169
R11558 VDPWR.n2460 VDPWR 0.158169
R11559 VDPWR.n203 VDPWR.n202 0.155911
R11560 VDPWR.n2177 VDPWR.n2176 0.152881
R11561 VDPWR.n3134 VDPWR.n3133 0.152187
R11562 VDPWR.n757 VDPWR.n756 0.150053
R11563 VDPWR.n3073 VDPWR.n3072 0.14385
R11564 VDPWR.n3068 VDPWR.n782 0.14385
R11565 VDPWR.n2507 VDPWR.n2499 0.14385
R11566 VDPWR.n2540 VDPWR.n2339 0.14385
R11567 VDPWR.n3113 VDPWR.n775 0.14385
R11568 VDPWR.n2538 VDPWR.n2537 0.14385
R11569 VDPWR.n2746 VDPWR.n2721 0.143027
R11570 VDPWR.n2290 VDPWR.n943 0.142675
R11571 VDPWR.n2332 VDPWR.n2331 0.142675
R11572 VDPWR.n2249 VDPWR.n973 0.142675
R11573 VDPWR.n2336 VDPWR.n1009 0.142675
R11574 VDPWR.n2256 VDPWR.n923 0.142675
R11575 VDPWR.n2159 VDPWR.n988 0.142675
R11576 VDPWR.n1362 VDPWR 0.14207
R11577 VDPWR.n1695 VDPWR 0.14207
R11578 VDPWR.n1609 VDPWR 0.14207
R11579 VDPWR VDPWR.n888 0.14207
R11580 VDPWR.n1433 VDPWR 0.141725
R11581 VDPWR.n1832 VDPWR 0.141725
R11582 VDPWR.n2055 VDPWR 0.141725
R11583 VDPWR.n1764 VDPWR 0.120408
R11584 VDPWR.n2104 VDPWR 0.120408
R11585 VDPWR VDPWR.n2476 0.120408
R11586 VDPWR.n1589 VDPWR.n1191 0.12035
R11587 VDPWR.n1820 VDPWR.n1228 0.12035
R11588 VDPWR.n1784 VDPWR.n1245 0.12035
R11589 VDPWR.n1714 VDPWR.n1594 0.12035
R11590 VDPWR.n1904 VDPWR.n1193 0.12035
R11591 VDPWR.n1754 VDPWR.n1267 0.12035
R11592 VDPWR.n587 VDPWR.n566 0.120292
R11593 VDPWR.n626 VDPWR.n567 0.120292
R11594 VDPWR.n619 VDPWR.n618 0.120292
R11595 VDPWR.n618 VDPWR.n592 0.120292
R11596 VDPWR.n614 VDPWR.n613 0.120292
R11597 VDPWR.n613 VDPWR.n612 0.120292
R11598 VDPWR.n609 VDPWR.n608 0.120292
R11599 VDPWR.n608 VDPWR.n607 0.120292
R11600 VDPWR.n604 VDPWR.n603 0.120292
R11601 VDPWR.n603 VDPWR.n597 0.120292
R11602 VDPWR.n599 VDPWR.n597 0.120292
R11603 VDPWR.n572 VDPWR.n568 0.120292
R11604 VDPWR.n585 VDPWR.n569 0.120292
R11605 VDPWR.n636 VDPWR.n563 0.120292
R11606 VDPWR.n637 VDPWR.n636 0.120292
R11607 VDPWR.n652 VDPWR.n538 0.120292
R11608 VDPWR.n648 VDPWR.n647 0.120292
R11609 VDPWR.n647 VDPWR.n542 0.120292
R11610 VDPWR.n558 VDPWR.n557 0.120292
R11611 VDPWR.n557 VDPWR.n549 0.120292
R11612 VDPWR.n552 VDPWR.n549 0.120292
R11613 VDPWR.n307 VDPWR.n286 0.120292
R11614 VDPWR.n346 VDPWR.n287 0.120292
R11615 VDPWR.n339 VDPWR.n338 0.120292
R11616 VDPWR.n338 VDPWR.n312 0.120292
R11617 VDPWR.n334 VDPWR.n333 0.120292
R11618 VDPWR.n333 VDPWR.n332 0.120292
R11619 VDPWR.n329 VDPWR.n328 0.120292
R11620 VDPWR.n328 VDPWR.n327 0.120292
R11621 VDPWR.n324 VDPWR.n323 0.120292
R11622 VDPWR.n323 VDPWR.n317 0.120292
R11623 VDPWR.n319 VDPWR.n317 0.120292
R11624 VDPWR.n292 VDPWR.n288 0.120292
R11625 VDPWR.n305 VDPWR.n289 0.120292
R11626 VDPWR.n356 VDPWR.n283 0.120292
R11627 VDPWR.n357 VDPWR.n356 0.120292
R11628 VDPWR.n372 VDPWR.n258 0.120292
R11629 VDPWR.n368 VDPWR.n367 0.120292
R11630 VDPWR.n367 VDPWR.n262 0.120292
R11631 VDPWR.n278 VDPWR.n277 0.120292
R11632 VDPWR.n277 VDPWR.n269 0.120292
R11633 VDPWR.n272 VDPWR.n269 0.120292
R11634 VDPWR.n1375 VDPWR.n1369 0.120292
R11635 VDPWR.n1388 VDPWR.n1342 0.120292
R11636 VDPWR.n1393 VDPWR.n1342 0.120292
R11637 VDPWR.n1394 VDPWR.n1393 0.120292
R11638 VDPWR.n1395 VDPWR.n1340 0.120292
R11639 VDPWR.n1400 VDPWR.n1340 0.120292
R11640 VDPWR.n1401 VDPWR.n1400 0.120292
R11641 VDPWR.n1407 VDPWR.n1338 0.120292
R11642 VDPWR.n1408 VDPWR.n1407 0.120292
R11643 VDPWR.n1409 VDPWR.n1408 0.120292
R11644 VDPWR.n1437 VDPWR.n1436 0.120292
R11645 VDPWR.n1437 VDPWR.n1322 0.120292
R11646 VDPWR.n1442 VDPWR.n1322 0.120292
R11647 VDPWR.n1443 VDPWR.n1442 0.120292
R11648 VDPWR.n1444 VDPWR.n1443 0.120292
R11649 VDPWR.n1464 VDPWR.n1313 0.120292
R11650 VDPWR VDPWR.n1464 0.120292
R11651 VDPWR.n1468 VDPWR.n1467 0.120292
R11652 VDPWR.n1468 VDPWR.n1310 0.120292
R11653 VDPWR.n1472 VDPWR.n1310 0.120292
R11654 VDPWR.n1473 VDPWR.n1472 0.120292
R11655 VDPWR.n1473 VDPWR.n1308 0.120292
R11656 VDPWR.n1477 VDPWR.n1308 0.120292
R11657 VDPWR.n1478 VDPWR.n1477 0.120292
R11658 VDPWR.n1479 VDPWR.n1478 0.120292
R11659 VDPWR.n1501 VDPWR.n1295 0.120292
R11660 VDPWR.n1508 VDPWR.n1295 0.120292
R11661 VDPWR.n1509 VDPWR.n1508 0.120292
R11662 VDPWR.n1510 VDPWR.n1509 0.120292
R11663 VDPWR.n1510 VDPWR.n1293 0.120292
R11664 VDPWR.n1514 VDPWR.n1293 0.120292
R11665 VDPWR.n1515 VDPWR.n1514 0.120292
R11666 VDPWR.n1574 VDPWR.n1573 0.120292
R11667 VDPWR.n1573 VDPWR.n1523 0.120292
R11668 VDPWR.n1569 VDPWR.n1523 0.120292
R11669 VDPWR.n1569 VDPWR.n1568 0.120292
R11670 VDPWR.n1568 VDPWR.n1525 0.120292
R11671 VDPWR.n1564 VDPWR.n1525 0.120292
R11672 VDPWR.n1564 VDPWR.n1563 0.120292
R11673 VDPWR.n1563 VDPWR.n1562 0.120292
R11674 VDPWR.n1562 VDPWR.n1527 0.120292
R11675 VDPWR.n1558 VDPWR.n1527 0.120292
R11676 VDPWR.n1703 VDPWR.n1702 0.120292
R11677 VDPWR.n1718 VDPWR.n1278 0.120292
R11678 VDPWR.n1723 VDPWR.n1278 0.120292
R11679 VDPWR.n1724 VDPWR.n1723 0.120292
R11680 VDPWR.n1725 VDPWR.n1276 0.120292
R11681 VDPWR.n1730 VDPWR.n1276 0.120292
R11682 VDPWR.n1731 VDPWR.n1730 0.120292
R11683 VDPWR.n1737 VDPWR.n1274 0.120292
R11684 VDPWR.n1738 VDPWR.n1737 0.120292
R11685 VDPWR.n1739 VDPWR.n1738 0.120292
R11686 VDPWR.n1772 VDPWR.n1256 0.120292
R11687 VDPWR.n1773 VDPWR.n1772 0.120292
R11688 VDPWR.n1774 VDPWR.n1773 0.120292
R11689 VDPWR.n1788 VDPWR.n1240 0.120292
R11690 VDPWR.n1793 VDPWR.n1240 0.120292
R11691 VDPWR.n1800 VDPWR.n1238 0.120292
R11692 VDPWR.n1801 VDPWR.n1800 0.120292
R11693 VDPWR.n1801 VDPWR.n1236 0.120292
R11694 VDPWR.n1806 VDPWR.n1236 0.120292
R11695 VDPWR.n1807 VDPWR.n1806 0.120292
R11696 VDPWR.n1808 VDPWR.n1807 0.120292
R11697 VDPWR.n1838 VDPWR.n1219 0.120292
R11698 VDPWR.n1843 VDPWR.n1219 0.120292
R11699 VDPWR.n1844 VDPWR.n1843 0.120292
R11700 VDPWR.n1845 VDPWR.n1844 0.120292
R11701 VDPWR.n1868 VDPWR.n1867 0.120292
R11702 VDPWR.n1869 VDPWR.n1868 0.120292
R11703 VDPWR.n1869 VDPWR.n1210 0.120292
R11704 VDPWR.n1878 VDPWR.n1210 0.120292
R11705 VDPWR.n1879 VDPWR.n1878 0.120292
R11706 VDPWR.n1880 VDPWR.n1879 0.120292
R11707 VDPWR.n1608 VDPWR.n1607 0.120292
R11708 VDPWR.n1656 VDPWR.n1626 0.120292
R11709 VDPWR.n1652 VDPWR.n1626 0.120292
R11710 VDPWR.n1652 VDPWR.n1651 0.120292
R11711 VDPWR.n1648 VDPWR.n1647 0.120292
R11712 VDPWR.n1647 VDPWR.n1629 0.120292
R11713 VDPWR.n1642 VDPWR.n1629 0.120292
R11714 VDPWR.n1641 VDPWR.n1631 0.120292
R11715 VDPWR.n1636 VDPWR.n1631 0.120292
R11716 VDPWR.n1636 VDPWR.n1635 0.120292
R11717 VDPWR.n2054 VDPWR.n1129 0.120292
R11718 VDPWR.n2044 VDPWR.n1129 0.120292
R11719 VDPWR.n2044 VDPWR.n2043 0.120292
R11720 VDPWR.n2043 VDPWR.n2042 0.120292
R11721 VDPWR.n2030 VDPWR.n1141 0.120292
R11722 VDPWR.n2025 VDPWR.n1141 0.120292
R11723 VDPWR.n2024 VDPWR.n2023 0.120292
R11724 VDPWR.n2023 VDPWR.n1152 0.120292
R11725 VDPWR.n2019 VDPWR.n1152 0.120292
R11726 VDPWR.n2019 VDPWR.n2018 0.120292
R11727 VDPWR.n2015 VDPWR.n2014 0.120292
R11728 VDPWR.n2014 VDPWR.n1157 0.120292
R11729 VDPWR.n2010 VDPWR.n1157 0.120292
R11730 VDPWR.n1999 VDPWR.n1998 0.120292
R11731 VDPWR.n1998 VDPWR.n1180 0.120292
R11732 VDPWR.n1993 VDPWR.n1180 0.120292
R11733 VDPWR.n1991 VDPWR.n1183 0.120292
R11734 VDPWR.n1985 VDPWR.n1984 0.120292
R11735 VDPWR.n1984 VDPWR.n1185 0.120292
R11736 VDPWR.n1962 VDPWR.n1923 0.120292
R11737 VDPWR.n1957 VDPWR.n1923 0.120292
R11738 VDPWR.n2114 VDPWR.n2109 0.120292
R11739 VDPWR.n2128 VDPWR.n2083 0.120292
R11740 VDPWR.n2132 VDPWR.n2083 0.120292
R11741 VDPWR.n2133 VDPWR.n2132 0.120292
R11742 VDPWR.n2138 VDPWR.n2081 0.120292
R11743 VDPWR.n2139 VDPWR.n2138 0.120292
R11744 VDPWR.n2144 VDPWR.n2143 0.120292
R11745 VDPWR.n2144 VDPWR.n2078 0.120292
R11746 VDPWR.n2148 VDPWR.n2078 0.120292
R11747 VDPWR.n2149 VDPWR.n2148 0.120292
R11748 VDPWR.n2182 VDPWR.n2181 0.120292
R11749 VDPWR.n2183 VDPWR.n1101 0.120292
R11750 VDPWR.n2189 VDPWR.n1101 0.120292
R11751 VDPWR.n2190 VDPWR.n2189 0.120292
R11752 VDPWR.n2234 VDPWR.n2198 0.120292
R11753 VDPWR.n2229 VDPWR.n2198 0.120292
R11754 VDPWR.n2229 VDPWR.n2228 0.120292
R11755 VDPWR.n2228 VDPWR.n2227 0.120292
R11756 VDPWR.n2224 VDPWR.n2223 0.120292
R11757 VDPWR.n2223 VDPWR.n2206 0.120292
R11758 VDPWR.n2218 VDPWR.n2206 0.120292
R11759 VDPWR.n2218 VDPWR.n2217 0.120292
R11760 VDPWR.n2312 VDPWR.n1027 0.120292
R11761 VDPWR.n2307 VDPWR.n1027 0.120292
R11762 VDPWR.n2307 VDPWR.n2306 0.120292
R11763 VDPWR.n2306 VDPWR.n1032 0.120292
R11764 VDPWR.n2301 VDPWR.n1032 0.120292
R11765 VDPWR.n2301 VDPWR.n2300 0.120292
R11766 VDPWR.n2300 VDPWR.n2299 0.120292
R11767 VDPWR.n2286 VDPWR.n1049 0.120292
R11768 VDPWR.n2280 VDPWR.n1049 0.120292
R11769 VDPWR.n2280 VDPWR.n2279 0.120292
R11770 VDPWR.n2279 VDPWR.n2278 0.120292
R11771 VDPWR.n2278 VDPWR.n1060 0.120292
R11772 VDPWR.n2273 VDPWR.n1060 0.120292
R11773 VDPWR.n2273 VDPWR.n2272 0.120292
R11774 VDPWR.n2269 VDPWR.n2268 0.120292
R11775 VDPWR.n2268 VDPWR.n1067 0.120292
R11776 VDPWR.n2764 VDPWR.n1004 0.120292
R11777 VDPWR.n2766 VDPWR.n2765 0.120292
R11778 VDPWR.n2766 VDPWR.n1002 0.120292
R11779 VDPWR.n2775 VDPWR.n1002 0.120292
R11780 VDPWR.n2778 VDPWR.n2775 0.120292
R11781 VDPWR.n2779 VDPWR.n2778 0.120292
R11782 VDPWR.n2786 VDPWR.n999 0.120292
R11783 VDPWR.n2787 VDPWR.n2786 0.120292
R11784 VDPWR.n2819 VDPWR.n2818 0.120292
R11785 VDPWR.n2826 VDPWR.n2825 0.120292
R11786 VDPWR.n2833 VDPWR.n2832 0.120292
R11787 VDPWR.n2856 VDPWR.n2855 0.120292
R11788 VDPWR.n2862 VDPWR.n966 0.120292
R11789 VDPWR.n2863 VDPWR.n2862 0.120292
R11790 VDPWR.n2864 VDPWR.n2863 0.120292
R11791 VDPWR.n2864 VDPWR.n963 0.120292
R11792 VDPWR.n2869 VDPWR.n963 0.120292
R11793 VDPWR.n2906 VDPWR.n2905 0.120292
R11794 VDPWR.n2906 VDPWR.n951 0.120292
R11795 VDPWR.n2911 VDPWR.n951 0.120292
R11796 VDPWR.n2912 VDPWR.n2911 0.120292
R11797 VDPWR.n2912 VDPWR.n949 0.120292
R11798 VDPWR.n2918 VDPWR.n949 0.120292
R11799 VDPWR.n2919 VDPWR.n2918 0.120292
R11800 VDPWR.n2920 VDPWR.n2919 0.120292
R11801 VDPWR.n2942 VDPWR.n938 0.120292
R11802 VDPWR.n2943 VDPWR.n2942 0.120292
R11803 VDPWR.n2949 VDPWR.n2948 0.120292
R11804 VDPWR.n2950 VDPWR.n2949 0.120292
R11805 VDPWR.n2955 VDPWR.n2954 0.120292
R11806 VDPWR.n2956 VDPWR.n2955 0.120292
R11807 VDPWR.n2956 VDPWR.n933 0.120292
R11808 VDPWR.n2961 VDPWR.n933 0.120292
R11809 VDPWR.n2715 VDPWR.n2544 0.120292
R11810 VDPWR.n2711 VDPWR.n2544 0.120292
R11811 VDPWR.n2711 VDPWR.n2710 0.120292
R11812 VDPWR.n2710 VDPWR.n2709 0.120292
R11813 VDPWR.n2709 VDPWR.n2580 0.120292
R11814 VDPWR.n2704 VDPWR.n2580 0.120292
R11815 VDPWR.n2704 VDPWR.n2703 0.120292
R11816 VDPWR.n2703 VDPWR.n2702 0.120292
R11817 VDPWR.n2702 VDPWR.n2584 0.120292
R11818 VDPWR.n2698 VDPWR.n2584 0.120292
R11819 VDPWR.n2698 VDPWR.n2697 0.120292
R11820 VDPWR.n2682 VDPWR.n2681 0.120292
R11821 VDPWR.n2681 VDPWR.n2680 0.120292
R11822 VDPWR.n2680 VDPWR.n2606 0.120292
R11823 VDPWR.n2674 VDPWR.n2606 0.120292
R11824 VDPWR.n2674 VDPWR.n2673 0.120292
R11825 VDPWR.n2673 VDPWR.n2672 0.120292
R11826 VDPWR.n2672 VDPWR.n2611 0.120292
R11827 VDPWR.n2667 VDPWR.n2611 0.120292
R11828 VDPWR.n2646 VDPWR.n2645 0.120292
R11829 VDPWR.n2645 VDPWR.n2644 0.120292
R11830 VDPWR.n2639 VDPWR.n2638 0.120292
R11831 VDPWR.n2638 VDPWR.n2622 0.120292
R11832 VDPWR.n3049 VDPWR.n3048 0.120292
R11833 VDPWR.n3048 VDPWR.n3047 0.120292
R11834 VDPWR.n3043 VDPWR.n895 0.120292
R11835 VDPWR.n3043 VDPWR.n3042 0.120292
R11836 VDPWR.n3042 VDPWR.n898 0.120292
R11837 VDPWR.n3028 VDPWR.n908 0.120292
R11838 VDPWR.n914 VDPWR.n908 0.120292
R11839 VDPWR.n3022 VDPWR.n914 0.120292
R11840 VDPWR.n3022 VDPWR.n3021 0.120292
R11841 VDPWR.n3021 VDPWR.n3020 0.120292
R11842 VDPWR.n3017 VDPWR.n3016 0.120292
R11843 VDPWR.n3016 VDPWR.n918 0.120292
R11844 VDPWR.n2384 VDPWR.n2367 0.120292
R11845 VDPWR.n2402 VDPWR.n2358 0.120292
R11846 VDPWR.n2407 VDPWR.n2354 0.120292
R11847 VDPWR.n2408 VDPWR.n2407 0.120292
R11848 VDPWR.n2414 VDPWR.n2413 0.120292
R11849 VDPWR.n2423 VDPWR.n2350 0.120292
R11850 VDPWR.n2522 VDPWR.n2435 0.120292
R11851 VDPWR.n2517 VDPWR.n2435 0.120292
R11852 VDPWR.n2517 VDPWR.n2516 0.120292
R11853 VDPWR.n2489 VDPWR.n2488 0.120292
R11854 VDPWR.n2488 VDPWR.n2487 0.120292
R11855 VDPWR.n2487 VDPWR.n2455 0.120292
R11856 VDPWR.n2482 VDPWR.n2481 0.120292
R11857 VDPWR.n2481 VDPWR.n2457 0.120292
R11858 VDPWR.n3088 VDPWR.n3087 0.120292
R11859 VDPWR.n3087 VDPWR.n3086 0.120292
R11860 VDPWR.n3086 VDPWR.n794 0.120292
R11861 VDPWR.n3082 VDPWR.n3081 0.120292
R11862 VDPWR.n861 VDPWR.n860 0.120292
R11863 VDPWR.n860 VDPWR.n816 0.120292
R11864 VDPWR.n49 VDPWR.n28 0.120292
R11865 VDPWR.n88 VDPWR.n29 0.120292
R11866 VDPWR.n81 VDPWR.n80 0.120292
R11867 VDPWR.n80 VDPWR.n54 0.120292
R11868 VDPWR.n76 VDPWR.n75 0.120292
R11869 VDPWR.n75 VDPWR.n74 0.120292
R11870 VDPWR.n71 VDPWR.n70 0.120292
R11871 VDPWR.n70 VDPWR.n69 0.120292
R11872 VDPWR.n66 VDPWR.n65 0.120292
R11873 VDPWR.n65 VDPWR.n59 0.120292
R11874 VDPWR.n61 VDPWR.n59 0.120292
R11875 VDPWR.n34 VDPWR.n30 0.120292
R11876 VDPWR.n47 VDPWR.n31 0.120292
R11877 VDPWR.n98 VDPWR.n25 0.120292
R11878 VDPWR.n99 VDPWR.n98 0.120292
R11879 VDPWR.n114 VDPWR.n0 0.120292
R11880 VDPWR.n110 VDPWR.n109 0.120292
R11881 VDPWR.n109 VDPWR.n4 0.120292
R11882 VDPWR.n20 VDPWR.n19 0.120292
R11883 VDPWR.n19 VDPWR.n11 0.120292
R11884 VDPWR.n14 VDPWR.n11 0.120292
R11885 VDPWR.n2335 VDPWR.n2334 0.120125
R11886 VDPWR.n2334 VDPWR.n2333 0.120125
R11887 VDPWR.n2333 VDPWR.n1011 0.120125
R11888 VDPWR.n1011 VDPWR.n1010 0.120125
R11889 VDPWR.n1593 VDPWR.n1592 0.120125
R11890 VDPWR.n1592 VDPWR.n1591 0.120125
R11891 VDPWR.n1591 VDPWR.n1590 0.120125
R11892 VDPWR.n1590 VDPWR.n1284 0.120125
R11893 VDPWR.n1674 VDPWR.n1673 0.120125
R11894 VDPWR.n1673 VDPWR.n1192 0.120125
R11895 VDPWR.n1907 VDPWR.n1192 0.120125
R11896 VDPWR.n1907 VDPWR.n1906 0.120125
R11897 VDPWR.n2251 VDPWR.n1090 0.120125
R11898 VDPWR.n2252 VDPWR.n2251 0.120125
R11899 VDPWR.n2253 VDPWR.n2252 0.120125
R11900 VDPWR.n2254 VDPWR.n2253 0.120125
R11901 VDPWR.n2539 VDPWR.n871 0.120125
R11902 VDPWR.n3069 VDPWR.n871 0.120125
R11903 VDPWR.n3071 VDPWR.n3069 0.120125
R11904 VDPWR.n3071 VDPWR.n3070 0.120125
R11905 VDPWR.n2505 VDPWR.n2504 0.120125
R11906 VDPWR.n2505 VDPWR.n776 0.120125
R11907 VDPWR.n3109 VDPWR.n776 0.120125
R11908 VDPWR.n3110 VDPWR.n3109 0.120125
R11909 VDPWR.n627 VDPWR.n566 0.11899
R11910 VDPWR.n347 VDPWR.n286 0.11899
R11911 VDPWR.n89 VDPWR.n28 0.11899
R11912 VDPWR.n3115 VDPWR.n771 0.116902
R11913 VDPWR.n2053 VDPWR.n2052 0.113774
R11914 VDPWR.n2052 VDPWR.n2047 0.113774
R11915 VDPWR.n757 VDPWR.n117 0.113371
R11916 VDPWR.n461 VDPWR.n403 0.1125
R11917 VDPWR.n1558 VDPWR.n1557 0.112479
R11918 VDPWR.n1076 VDPWR.n1067 0.112479
R11919 VDPWR.n2963 VDPWR.n2961 0.112479
R11920 VDPWR.n3010 VDPWR.n3009 0.112479
R11921 VDPWR.n849 VDPWR.n848 0.112479
R11922 VDPWR.n1974 VDPWR.n1046 0.1086
R11923 VDPWR.n2006 VDPWR.n1012 0.1086
R11924 VDPWR.n2250 VDPWR.n1091 0.1086
R11925 VDPWR.n1672 VDPWR.n1596 0.1086
R11926 VDPWR.n2255 VDPWR.n1089 0.1086
R11927 VDPWR.n2073 VDPWR.n2072 0.1086
R11928 VDPWR.n1444 VDPWR.n1319 0.107271
R11929 VDPWR.n1774 VDPWR.n1248 0.107271
R11930 VDPWR.n2039 VDPWR.n2038 0.107271
R11931 VDPWR.n2190 VDPWR.n1094 0.107271
R11932 VDPWR.n2833 VDPWR.n976 0.107271
R11933 VDPWR.n2667 VDPWR.n2666 0.107271
R11934 VDPWR.n3104 VDPWR.n779 0.10625
R11935 VDPWR.n3105 VDPWR.n778 0.10625
R11936 VDPWR.n2225 VDPWR.n2205 0.105418
R11937 VDPWR.n1062 VDPWR.n1059 0.105418
R11938 VDPWR.n1361 VDPWR 0.105238
R11939 VDPWR.n1694 VDPWR 0.105238
R11940 VDPWR.n1616 VDPWR 0.105238
R11941 VDPWR.n2103 VDPWR 0.105238
R11942 VDPWR.n2736 VDPWR 0.105238
R11943 VDPWR.n2560 VDPWR 0.105238
R11944 VDPWR.n2378 VDPWR 0.105238
R11945 VDPWR.n377 VDPWR.n254 0.103147
R11946 VDPWR.n1960 VDPWR.n1959 0.102087
R11947 VDPWR.n2891 VDPWR.n2890 0.102087
R11948 VDPWR.n3015 VDPWR.n3014 0.102087
R11949 VDPWR.n572 VDPWR 0.0981562
R11950 VDPWR.n292 VDPWR 0.0981562
R11951 VDPWR VDPWR.n1338 0.0981562
R11952 VDPWR.n1432 VDPWR 0.0981562
R11953 VDPWR.n1467 VDPWR 0.0981562
R11954 VDPWR.n1496 VDPWR 0.0981562
R11955 VDPWR VDPWR.n1274 0.0981562
R11956 VDPWR.n1759 VDPWR 0.0981562
R11957 VDPWR VDPWR.n1238 0.0981562
R11958 VDPWR.n1824 VDPWR 0.0981562
R11959 VDPWR.n1838 VDPWR 0.0981562
R11960 VDPWR VDPWR.n1641 0.0981562
R11961 VDPWR VDPWR.n2056 0.0981562
R11962 VDPWR VDPWR.n2054 0.0981562
R11963 VDPWR VDPWR.n2024 0.0981562
R11964 VDPWR.n2015 VDPWR 0.0981562
R11965 VDPWR VDPWR.n2002 0.0981562
R11966 VDPWR VDPWR.n1991 0.0981562
R11967 VDPWR VDPWR.n1962 0.0981562
R11968 VDPWR.n2143 VDPWR 0.0981562
R11969 VDPWR.n2169 VDPWR 0.0981562
R11970 VDPWR.n2175 VDPWR 0.0981562
R11971 VDPWR.n2181 VDPWR 0.0981562
R11972 VDPWR.n2224 VDPWR 0.0981562
R11973 VDPWR VDPWR.n2312 0.0981562
R11974 VDPWR VDPWR.n1004 0.0981562
R11975 VDPWR.n2825 VDPWR 0.0981562
R11976 VDPWR VDPWR.n966 0.0981562
R11977 VDPWR.n2646 VDPWR 0.0981562
R11978 VDPWR.n2382 VDPWR 0.0981562
R11979 VDPWR VDPWR.n2350 0.0981562
R11980 VDPWR VDPWR.n2522 0.0981562
R11981 VDPWR.n2440 VDPWR 0.0981562
R11982 VDPWR.n3088 VDPWR 0.0981562
R11983 VDPWR VDPWR.n3077 0.0981562
R11984 VDPWR VDPWR.n849 0.0981562
R11985 VDPWR.n34 VDPWR 0.0981562
R11986 VDPWR.n3103 VDPWR.n3102 0.0977722
R11987 VDPWR.n2508 VDPWR.n779 0.0977722
R11988 VDPWR.n2536 VDPWR.n2343 0.0977722
R11989 VDPWR.n3074 VDPWR.n770 0.0977722
R11990 VDPWR.n2832 VDPWR 0.0968542
R11991 VDPWR VDPWR.n3010 0.0968542
R11992 VDPWR.n628 VDPWR 0.0955521
R11993 VDPWR.n348 VDPWR 0.0955521
R11994 VDPWR.n90 VDPWR 0.0955521
R11995 VDPWR.n2695 VDPWR.n2589 0.0950946
R11996 VDPWR.n2690 VDPWR.n2592 0.0950946
R11997 VDPWR.n2665 VDPWR.n2615 0.0950946
R11998 VDPWR.n2660 VDPWR.n2618 0.0950946
R11999 VDPWR.n2509 VDPWR.n2444 0.0950946
R12000 VDPWR.n2494 VDPWR.n2446 0.0950946
R12001 VDPWR.n1490 VDPWR.n1489 0.0950946
R12002 VDPWR.n1494 VDPWR.n1299 0.0950946
R12003 VDPWR.n1454 VDPWR.n1453 0.0950946
R12004 VDPWR.n1458 VDPWR.n1316 0.0950946
R12005 VDPWR.n1421 VDPWR.n1420 0.0950946
R12006 VDPWR.n1425 VDPWR.n1330 0.0950946
R12007 VDPWR.n1373 VDPWR.n1371 0.0950946
R12008 VDPWR.n1386 VDPWR.n1345 0.0950946
R12009 VDPWR.n1556 VDPWR.n1530 0.0950946
R12010 VDPWR.n1546 VDPWR.n1544 0.0950946
R12011 VDPWR.n1586 VDPWR.n1585 0.0950946
R12012 VDPWR.n1579 VDPWR.n1290 0.0950946
R12013 VDPWR.n1818 VDPWR.n1817 0.0950946
R12014 VDPWR.n1822 VDPWR.n1226 0.0950946
R12015 VDPWR.n1782 VDPWR.n1781 0.0950946
R12016 VDPWR.n1786 VDPWR.n1243 0.0950946
R12017 VDPWR.n1752 VDPWR.n1751 0.0950946
R12018 VDPWR.n1756 VDPWR.n1265 0.0950946
R12019 VDPWR.n1712 VDPWR.n1711 0.0950946
R12020 VDPWR.n1716 VDPWR.n1281 0.0950946
R12021 VDPWR.n1889 VDPWR.n1887 0.0950946
R12022 VDPWR.n1900 VDPWR.n1195 0.0950946
R12023 VDPWR.n1856 VDPWR.n1855 0.0950946
R12024 VDPWR.n1862 VDPWR.n1861 0.0950946
R12025 VDPWR.n2008 VDPWR.n1160 0.0950946
R12026 VDPWR.n2004 VDPWR.n1164 0.0950946
R12027 VDPWR.n2037 VDPWR.n1136 0.0950946
R12028 VDPWR.n2032 VDPWR.n1139 0.0950946
R12029 VDPWR.n2070 VDPWR.n2069 0.0950946
R12030 VDPWR.n2063 VDPWR.n1123 0.0950946
R12031 VDPWR.n1670 VDPWR.n1669 0.0950946
R12032 VDPWR.n1662 VDPWR.n1661 0.0950946
R12033 VDPWR.n1955 VDPWR.n1930 0.0950946
R12034 VDPWR.n1945 VDPWR.n1943 0.0950946
R12035 VDPWR.n1978 VDPWR.n1188 0.0950946
R12036 VDPWR.n1972 VDPWR.n1910 0.0950946
R12037 VDPWR.n2329 VDPWR.n2328 0.0950946
R12038 VDPWR.n2321 VDPWR.n2320 0.0950946
R12039 VDPWR.n2247 VDPWR.n2246 0.0950946
R12040 VDPWR.n2239 VDPWR.n2238 0.0950946
R12041 VDPWR.n2157 VDPWR.n2156 0.0950946
R12042 VDPWR.n2162 VDPWR.n2161 0.0950946
R12043 VDPWR.n2112 VDPWR.n2110 0.0950946
R12044 VDPWR.n2126 VDPWR.n2086 0.0950946
R12045 VDPWR.n2261 VDPWR.n1078 0.0950946
R12046 VDPWR.n1088 VDPWR.n1082 0.0950946
R12047 VDPWR.n2294 VDPWR.n1043 0.0950946
R12048 VDPWR.n2288 VDPWR.n1048 0.0950946
R12049 VDPWR.n2880 VDPWR.n2878 0.0950946
R12050 VDPWR.n2898 VDPWR.n956 0.0950946
R12051 VDPWR.n2842 VDPWR.n2841 0.0950946
R12052 VDPWR.n2847 VDPWR.n2846 0.0950946
R12053 VDPWR.n2803 VDPWR.n2802 0.0950946
R12054 VDPWR.n2807 VDPWR.n986 0.0950946
R12055 VDPWR.n2753 VDPWR.n2752 0.0950946
R12056 VDPWR.n2757 VDPWR.n1007 0.0950946
R12057 VDPWR.n2966 VDPWR.n2964 0.0950946
R12058 VDPWR.n2977 VDPWR.n925 0.0950946
R12059 VDPWR.n2930 VDPWR.n2929 0.0950946
R12060 VDPWR.n2934 VDPWR.n941 0.0950946
R12061 VDPWR.n3036 VDPWR.n903 0.0950946
R12062 VDPWR.n3030 VDPWR.n906 0.0950946
R12063 VDPWR.n3065 VDPWR.n3064 0.0950946
R12064 VDPWR.n3057 VDPWR.n3056 0.0950946
R12065 VDPWR.n2465 VDPWR.n785 0.0950946
R12066 VDPWR.n3100 VDPWR.n784 0.0950946
R12067 VDPWR.n2571 VDPWR.n2549 0.0950946
R12068 VDPWR.n2717 VDPWR.n2542 0.0950946
R12069 VDPWR.n3008 VDPWR.n922 0.0950946
R12070 VDPWR.n3003 VDPWR.n2985 0.0950946
R12071 VDPWR.n2426 VDPWR.n2344 0.0950946
R12072 VDPWR.n2534 VDPWR.n2342 0.0950946
R12073 VDPWR.n2391 VDPWR.n2390 0.0950946
R12074 VDPWR.n2394 VDPWR.n2393 0.0950946
R12075 VDPWR.n847 VDPWR.n846 0.0950946
R12076 VDPWR.n839 VDPWR.n772 0.0950946
R12077 VDPWR.n3075 VDPWR.n802 0.0950946
R12078 VDPWR.n868 VDPWR.n804 0.0950946
R12079 VDPWR VDPWR.n2104 0.0930646
R12080 VDPWR.n586 VDPWR.n568 0.0916458
R12081 VDPWR.n306 VDPWR.n288 0.0916458
R12082 VDPWR.n48 VDPWR.n30 0.0916458
R12083 VDPWR.n3104 VDPWR.n3103 0.0913766
R12084 VDPWR.n3106 VDPWR.n3105 0.0913766
R12085 VDPWR.n3171 VDPWR.n759 0.08675
R12086 VDPWR.n1974 VDPWR.n1908 0.086275
R12087 VDPWR.n2006 VDPWR.n1162 0.086275
R12088 VDPWR.n1246 VDPWR.n1091 0.086275
R12089 VDPWR.n1675 VDPWR.n1672 0.086275
R12090 VDPWR.n1905 VDPWR.n1089 0.086275
R12091 VDPWR.n2072 VDPWR.n1116 0.086275
R12092 VDPWR.n3149 VDPWR.n3134 0.0848934
R12093 VDPWR.n3165 VDPWR.n3150 0.0844041
R12094 VDPWR.n1374 VDPWR.n1370 0.0838333
R12095 VDPWR.n1387 VDPWR.n1344 0.0838333
R12096 VDPWR.n1419 VDPWR.n1418 0.0838333
R12097 VDPWR.n1450 VDPWR.n1315 0.0838333
R12098 VDPWR.n1488 VDPWR.n1302 0.0838333
R12099 VDPWR.n1584 VDPWR.n1583 0.0838333
R12100 VDPWR.n1547 VDPWR.n1536 0.0838333
R12101 VDPWR.n1710 VDPWR.n1677 0.0838333
R12102 VDPWR.n1717 VDPWR.n1280 0.0838333
R12103 VDPWR.n1750 VDPWR.n1749 0.0838333
R12104 VDPWR.n1254 VDPWR.n1251 0.0838333
R12105 VDPWR.n1816 VDPWR.n1230 0.0838333
R12106 VDPWR.n1854 VDPWR.n1853 0.0838333
R12107 VDPWR.n1899 VDPWR.n1898 0.0838333
R12108 VDPWR.n1668 VDPWR.n1598 0.0838333
R12109 VDPWR.n1663 VDPWR.n1657 0.0838333
R12110 VDPWR.n2068 VDPWR.n2067 0.0838333
R12111 VDPWR.n1146 VDPWR.n1144 0.0838333
R12112 VDPWR.n2009 VDPWR.n1159 0.0838333
R12113 VDPWR.n1946 VDPWR.n1935 0.0838333
R12114 VDPWR.n2113 VDPWR.n2089 0.0838333
R12115 VDPWR.n2127 VDPWR.n2085 0.0838333
R12116 VDPWR.n2155 VDPWR.n2154 0.0838333
R12117 VDPWR.n2197 VDPWR.n1097 0.0838333
R12118 VDPWR.n2327 VDPWR.n1015 0.0838333
R12119 VDPWR.n2295 VDPWR.n1042 0.0838333
R12120 VDPWR.n1087 VDPWR.n1085 0.0838333
R12121 VDPWR.n2751 VDPWR.n2721 0.0838333
R12122 VDPWR.n2801 VDPWR.n2800 0.0838333
R12123 VDPWR.n2848 VDPWR.n970 0.0838333
R12124 VDPWR.n2881 VDPWR.n2877 0.0838333
R12125 VDPWR.n2928 VDPWR.n2927 0.0838333
R12126 VDPWR.n2976 VDPWR.n2975 0.0838333
R12127 VDPWR.n2570 VDPWR.n2569 0.0838333
R12128 VDPWR.n2716 VDPWR.n2543 0.0838333
R12129 VDPWR.n2654 VDPWR.n2653 0.0838333
R12130 VDPWR.n3063 VDPWR.n875 0.0838333
R12131 VDPWR.n3037 VDPWR.n902 0.0838333
R12132 VDPWR.n3002 VDPWR.n2986 0.0838333
R12133 VDPWR.n2389 VDPWR.n2365 0.0838333
R12134 VDPWR.n2395 VDPWR.n2361 0.0838333
R12135 VDPWR.n2496 VDPWR.n2495 0.0838333
R12136 VDPWR.n841 VDPWR.n840 0.0838333
R12137 VDPWR.n777 VDPWR 0.08275
R12138 VDPWR.n781 VDPWR 0.08275
R12139 VDPWR.n2500 VDPWR 0.08275
R12140 VDPWR.n3112 VDPWR 0.08275
R12141 VDPWR.n2340 VDPWR 0.08275
R12142 VDPWR VDPWR.n1915 0.082648
R12143 VDPWR VDPWR.n2624 0.082648
R12144 VDPWR VDPWR.n1764 0.082648
R12145 VDPWR.n1765 VDPWR 0.082648
R12146 VDPWR.n1794 VDPWR 0.082648
R12147 VDPWR.n2476 VDPWR 0.082648
R12148 VDPWR VDPWR.n2460 0.082648
R12149 VDPWR.n1427 VDPWR.n1426 0.0812292
R12150 VDPWR.n1460 VDPWR.n1459 0.0812292
R12151 VDPWR.n1483 VDPWR.n1298 0.0812292
R12152 VDPWR.n1578 VDPWR.n1289 0.0812292
R12153 VDPWR.n1551 VDPWR.n1550 0.0812292
R12154 VDPWR.n1758 VDPWR.n1757 0.0812292
R12155 VDPWR.n1787 VDPWR.n1242 0.0812292
R12156 VDPWR.n1811 VDPWR.n1225 0.0812292
R12157 VDPWR.n1863 VDPWR.n1214 0.0812292
R12158 VDPWR.n1891 VDPWR.n1198 0.0812292
R12159 VDPWR.n2057 VDPWR.n1124 0.0812292
R12160 VDPWR.n2031 VDPWR.n1140 0.0812292
R12161 VDPWR.n1174 VDPWR.n1165 0.0812292
R12162 VDPWR.n1913 VDPWR.n1912 0.0812292
R12163 VDPWR.n1950 VDPWR.n1949 0.0812292
R12164 VDPWR.n2168 VDPWR.n1111 0.0812292
R12165 VDPWR.n2241 VDPWR.n2240 0.0812292
R12166 VDPWR.n2322 VDPWR.n1020 0.0812292
R12167 VDPWR.n1054 VDPWR.n1053 0.0812292
R12168 VDPWR.n1084 VDPWR.n1083 0.0812292
R12169 VDPWR.n2809 VDPWR.n2808 0.0812292
R12170 VDPWR.n2849 VDPWR.n968 0.0812292
R12171 VDPWR.n960 VDPWR.n955 0.0812292
R12172 VDPWR.n2924 VDPWR.n940 0.0812292
R12173 VDPWR.n2968 VDPWR.n928 0.0812292
R12174 VDPWR.n2689 VDPWR.n2688 0.0812292
R12175 VDPWR.n3058 VDPWR.n880 0.0812292
R12176 VDPWR.n910 VDPWR.n909 0.0812292
R12177 VDPWR.n2996 VDPWR.n2995 0.0812292
R12178 VDPWR.n2529 VDPWR.n2346 0.0812292
R12179 VDPWR.n2493 VDPWR.n2449 0.0812292
R12180 VDPWR.n3099 VDPWR.n3098 0.0812292
R12181 VDPWR.n835 VDPWR.n829 0.0812292
R12182 VDPWR.n536 VDPWR 0.0800455
R12183 VDPWR.n1415 VDPWR.n1336 0.0760208
R12184 VDPWR.n1487 VDPWR.n1306 0.0760208
R12185 VDPWR.n1746 VDPWR.n1272 0.0760208
R12186 VDPWR.n1815 VDPWR.n1234 0.0760208
R12187 VDPWR.n1867 VDPWR.n1212 0.0760208
R12188 VDPWR.n2062 VDPWR.n1122 0.0760208
R12189 VDPWR.n1173 VDPWR.n1169 0.0760208
R12190 VDPWR.n1971 VDPWR.n1970 0.0760208
R12191 VDPWR.n2163 VDPWR.n1113 0.0760208
R12192 VDPWR.n2326 VDPWR.n1017 0.0760208
R12193 VDPWR.n2287 VDPWR.n2286 0.0760208
R12194 VDPWR.n2797 VDPWR.n994 0.0760208
R12195 VDPWR.n2893 VDPWR.n959 0.0760208
R12196 VDPWR.n2935 VDPWR.n938 0.0760208
R12197 VDPWR.n2602 VDPWR.n2601 0.0760208
R12198 VDPWR.n3062 VDPWR.n877 0.0760208
R12199 VDPWR.n3029 VDPWR.n3028 0.0760208
R12200 VDPWR.n862 VDPWR.n806 0.0760208
R12201 VDPWR.n1908 VDPWR.n1191 0.074525
R12202 VDPWR.n1820 VDPWR.n1162 0.074525
R12203 VDPWR.n1784 VDPWR.n1246 0.074525
R12204 VDPWR.n1714 VDPWR.n1675 0.074525
R12205 VDPWR.n1905 VDPWR.n1904 0.074525
R12206 VDPWR.n1754 VDPWR.n1116 0.074525
R12207 VDPWR.n753 VDPWR 0.0710357
R12208 VDPWR.n1381 VDPWR.n1348 0.0708125
R12209 VDPWR.n1452 VDPWR.n1447 0.0708125
R12210 VDPWR.n1709 VDPWR.n1681 0.0708125
R12211 VDPWR.n1780 VDPWR.n1250 0.0708125
R12212 VDPWR.n1845 VDPWR.n1217 0.0708125
R12213 VDPWR.n1667 VDPWR.n1600 0.0708125
R12214 VDPWR.n1143 VDPWR.n1135 0.0708125
R12215 VDPWR.n1187 VDPWR.n1185 0.0708125
R12216 VDPWR.n2121 VDPWR.n2119 0.0708125
R12217 VDPWR.n2245 VDPWR.n1096 0.0708125
R12218 VDPWR.n2299 VDPWR.n1037 0.0708125
R12219 VDPWR.n2750 VDPWR.n2725 0.0708125
R12220 VDPWR.n2840 VDPWR.n2838 0.0708125
R12221 VDPWR.n2920 VDPWR.n945 0.0708125
R12222 VDPWR.n2576 VDPWR.n2548 0.0708125
R12223 VDPWR.n2650 VDPWR.n2614 0.0708125
R12224 VDPWR.n901 VDPWR.n898 0.0708125
R12225 VDPWR.n3077 VDPWR.n3076 0.0708125
R12226 VDPWR.n2599 VDPWR.n2590 0.0680676
R12227 VDPWR.n2599 VDPWR.n2591 0.0680676
R12228 VDPWR.n2652 VDPWR.n2616 0.0680676
R12229 VDPWR.n2652 VDPWR.n2617 0.0680676
R12230 VDPWR.n2498 VDPWR.n2497 0.0680676
R12231 VDPWR.n2497 VDPWR.n2445 0.0680676
R12232 VDPWR.n1305 VDPWR.n1303 0.0680676
R12233 VDPWR.n1305 VDPWR.n1304 0.0680676
R12234 VDPWR.n1449 VDPWR.n1320 0.0680676
R12235 VDPWR.n1449 VDPWR.n1448 0.0680676
R12236 VDPWR.n1417 VDPWR.n1334 0.0680676
R12237 VDPWR.n1417 VDPWR.n1416 0.0680676
R12238 VDPWR.n1382 VDPWR.n1347 0.0680676
R12239 VDPWR.n1383 VDPWR.n1382 0.0680676
R12240 VDPWR.n1553 VDPWR.n1552 0.0680676
R12241 VDPWR.n1552 VDPWR.n1533 0.0680676
R12242 VDPWR.n1582 VDPWR.n1288 0.0680676
R12243 VDPWR.n1582 VDPWR.n1581 0.0680676
R12244 VDPWR.n1233 VDPWR.n1231 0.0680676
R12245 VDPWR.n1233 VDPWR.n1232 0.0680676
R12246 VDPWR.n1253 VDPWR.n1249 0.0680676
R12247 VDPWR.n1253 VDPWR.n1252 0.0680676
R12248 VDPWR.n1748 VDPWR.n1270 0.0680676
R12249 VDPWR.n1748 VDPWR.n1747 0.0680676
R12250 VDPWR.n1680 VDPWR.n1678 0.0680676
R12251 VDPWR.n1680 VDPWR.n1679 0.0680676
R12252 VDPWR.n1888 VDPWR.n1197 0.0680676
R12253 VDPWR.n1901 VDPWR.n1197 0.0680676
R12254 VDPWR.n1852 VDPWR.n1216 0.0680676
R12255 VDPWR.n1852 VDPWR.n1215 0.0680676
R12256 VDPWR.n1172 VDPWR.n1170 0.0680676
R12257 VDPWR.n1172 VDPWR.n1171 0.0680676
R12258 VDPWR.n1145 VDPWR.n1137 0.0680676
R12259 VDPWR.n1145 VDPWR.n1138 0.0680676
R12260 VDPWR.n2066 VDPWR.n1120 0.0680676
R12261 VDPWR.n2066 VDPWR.n2065 0.0680676
R12262 VDPWR.n1658 VDPWR.n1599 0.0680676
R12263 VDPWR.n1660 VDPWR.n1658 0.0680676
R12264 VDPWR.n1952 VDPWR.n1951 0.0680676
R12265 VDPWR.n1951 VDPWR.n1932 0.0680676
R12266 VDPWR.n1977 VDPWR.n1189 0.0680676
R12267 VDPWR.n1909 VDPWR.n1189 0.0680676
R12268 VDPWR.n1021 VDPWR.n1016 0.0680676
R12269 VDPWR.n1023 VDPWR.n1021 0.0680676
R12270 VDPWR.n2235 VDPWR.n1095 0.0680676
R12271 VDPWR.n2237 VDPWR.n2235 0.0680676
R12272 VDPWR.n2153 VDPWR.n2076 0.0680676
R12273 VDPWR.n2153 VDPWR.n1114 0.0680676
R12274 VDPWR.n2122 VDPWR.n2088 0.0680676
R12275 VDPWR.n2123 VDPWR.n2122 0.0680676
R12276 VDPWR.n2260 VDPWR.n1079 0.0680676
R12277 VDPWR.n1081 VDPWR.n1079 0.0680676
R12278 VDPWR.n2293 VDPWR.n1044 0.0680676
R12279 VDPWR.n1047 VDPWR.n1044 0.0680676
R12280 VDPWR.n2894 VDPWR.n958 0.0680676
R12281 VDPWR.n2895 VDPWR.n2894 0.0680676
R12282 VDPWR.n978 VDPWR.n977 0.0680676
R12283 VDPWR.n977 VDPWR.n971 0.0680676
R12284 VDPWR.n2799 VDPWR.n992 0.0680676
R12285 VDPWR.n2799 VDPWR.n2798 0.0680676
R12286 VDPWR.n2724 VDPWR.n2722 0.0680676
R12287 VDPWR.n2724 VDPWR.n2723 0.0680676
R12288 VDPWR.n2965 VDPWR.n927 0.0680676
R12289 VDPWR.n2978 VDPWR.n927 0.0680676
R12290 VDPWR.n2926 VDPWR.n946 0.0680676
R12291 VDPWR.n2926 VDPWR.n2925 0.0680676
R12292 VDPWR.n3035 VDPWR.n904 0.0680676
R12293 VDPWR.n905 VDPWR.n904 0.0680676
R12294 VDPWR.n881 VDPWR.n876 0.0680676
R12295 VDPWR.n883 VDPWR.n881 0.0680676
R12296 VDPWR.n786 VDPWR.n783 0.0680676
R12297 VDPWR.n3101 VDPWR.n786 0.0680676
R12298 VDPWR.n2575 VDPWR.n2573 0.0680676
R12299 VDPWR.n2575 VDPWR.n2574 0.0680676
R12300 VDPWR.n2994 VDPWR.n2983 0.0680676
R12301 VDPWR.n2994 VDPWR.n2984 0.0680676
R12302 VDPWR.n2345 VDPWR.n2341 0.0680676
R12303 VDPWR.n2535 VDPWR.n2345 0.0680676
R12304 VDPWR.n2364 VDPWR.n2363 0.0680676
R12305 VDPWR.n2363 VDPWR.n2362 0.0680676
R12306 VDPWR.n828 VDPWR.n773 0.0680676
R12307 VDPWR.n828 VDPWR.n774 0.0680676
R12308 VDPWR.n805 VDPWR.n803 0.0680676
R12309 VDPWR.n869 VDPWR.n805 0.0680676
R12310 VDPWR.n1409 VDPWR.n1333 0.0656042
R12311 VDPWR.n1739 VDPWR.n1269 0.0656042
R12312 VDPWR.n1635 VDPWR.n1119 0.0656042
R12313 VDPWR.n2149 VDPWR.n2075 0.0656042
R12314 VDPWR.n2787 VDPWR.n991 0.0656042
R12315 VDPWR.n2697 VDPWR.n2696 0.0656042
R12316 VDPWR.n2424 VDPWR.n2423 0.0656042
R12317 VDPWR.n718 VDPWR 0.06425
R12318 VDPWR.n702 VDPWR 0.06425
R12319 VDPWR.n686 VDPWR 0.06425
R12320 VDPWR.n670 VDPWR 0.06425
R12321 VDPWR.n529 VDPWR 0.06425
R12322 VDPWR.n513 VDPWR 0.06425
R12323 VDPWR.n497 VDPWR 0.06425
R12324 VDPWR.n481 VDPWR 0.06425
R12325 VDPWR.n465 VDPWR 0.06425
R12326 VDPWR.n389 VDPWR 0.06425
R12327 VDPWR.n401 VDPWR 0.06425
R12328 VDPWR.n459 VDPWR 0.06425
R12329 VDPWR.n443 VDPWR 0.06425
R12330 VDPWR.n427 VDPWR 0.06425
R12331 VDPWR.n3170 VDPWR 0.06425
R12332 VDPWR.n3164 VDPWR 0.06425
R12333 VDPWR.n3148 VDPWR 0.06425
R12334 VDPWR.n3132 VDPWR 0.06425
R12335 VDPWR.n256 VDPWR.n253 0.061697
R12336 VDPWR.n754 VDPWR 0.0615066
R12337 VDPWR.n620 VDPWR 0.0603958
R12338 VDPWR VDPWR.n619 0.0603958
R12339 VDPWR.n614 VDPWR 0.0603958
R12340 VDPWR.n609 VDPWR 0.0603958
R12341 VDPWR.n604 VDPWR 0.0603958
R12342 VDPWR.n580 VDPWR 0.0603958
R12343 VDPWR VDPWR.n579 0.0603958
R12344 VDPWR VDPWR.n563 0.0603958
R12345 VDPWR.n639 VDPWR 0.0603958
R12346 VDPWR VDPWR.n638 0.0603958
R12347 VDPWR.n648 VDPWR 0.0603958
R12348 VDPWR.n558 VDPWR 0.0603958
R12349 VDPWR.n340 VDPWR 0.0603958
R12350 VDPWR VDPWR.n339 0.0603958
R12351 VDPWR.n334 VDPWR 0.0603958
R12352 VDPWR.n329 VDPWR 0.0603958
R12353 VDPWR.n324 VDPWR 0.0603958
R12354 VDPWR.n300 VDPWR 0.0603958
R12355 VDPWR VDPWR.n299 0.0603958
R12356 VDPWR VDPWR.n283 0.0603958
R12357 VDPWR.n359 VDPWR 0.0603958
R12358 VDPWR VDPWR.n358 0.0603958
R12359 VDPWR.n368 VDPWR 0.0603958
R12360 VDPWR.n278 VDPWR 0.0603958
R12361 VDPWR.n1369 VDPWR 0.0603958
R12362 VDPWR.n1395 VDPWR 0.0603958
R12363 VDPWR.n1436 VDPWR 0.0603958
R12364 VDPWR.n1497 VDPWR 0.0603958
R12365 VDPWR.n1500 VDPWR 0.0603958
R12366 VDPWR.n1501 VDPWR 0.0603958
R12367 VDPWR.n1574 VDPWR 0.0603958
R12368 VDPWR.n1702 VDPWR 0.0603958
R12369 VDPWR.n1725 VDPWR 0.0603958
R12370 VDPWR.n1763 VDPWR 0.0603958
R12371 VDPWR VDPWR.n1256 0.0603958
R12372 VDPWR.n1831 VDPWR 0.0603958
R12373 VDPWR.n1837 VDPWR 0.0603958
R12374 VDPWR.n1883 VDPWR 0.0603958
R12375 VDPWR VDPWR.n1608 0.0603958
R12376 VDPWR.n1648 VDPWR 0.0603958
R12377 VDPWR.n2039 VDPWR 0.0603958
R12378 VDPWR.n1999 VDPWR 0.0603958
R12379 VDPWR VDPWR.n1992 0.0603958
R12380 VDPWR.n1985 VDPWR 0.0603958
R12381 VDPWR.n1965 VDPWR 0.0603958
R12382 VDPWR VDPWR.n1963 0.0603958
R12383 VDPWR.n1957 VDPWR 0.0603958
R12384 VDPWR.n2105 VDPWR 0.0603958
R12385 VDPWR.n2109 VDPWR 0.0603958
R12386 VDPWR VDPWR.n2081 0.0603958
R12387 VDPWR.n2170 VDPWR 0.0603958
R12388 VDPWR.n2174 VDPWR 0.0603958
R12389 VDPWR.n2183 VDPWR 0.0603958
R12390 VDPWR.n2217 VDPWR 0.0603958
R12391 VDPWR.n2214 VDPWR 0.0603958
R12392 VDPWR VDPWR.n2213 0.0603958
R12393 VDPWR VDPWR.n2318 0.0603958
R12394 VDPWR.n2314 VDPWR 0.0603958
R12395 VDPWR VDPWR.n2313 0.0603958
R12396 VDPWR.n2272 VDPWR 0.0603958
R12397 VDPWR.n2269 VDPWR 0.0603958
R12398 VDPWR.n2737 VDPWR 0.0603958
R12399 VDPWR.n2745 VDPWR 0.0603958
R12400 VDPWR.n2765 VDPWR 0.0603958
R12401 VDPWR VDPWR.n999 0.0603958
R12402 VDPWR.n2810 VDPWR 0.0603958
R12403 VDPWR.n2818 VDPWR 0.0603958
R12404 VDPWR.n2820 VDPWR 0.0603958
R12405 VDPWR VDPWR.n2826 0.0603958
R12406 VDPWR.n2827 VDPWR 0.0603958
R12407 VDPWR.n2831 VDPWR 0.0603958
R12408 VDPWR VDPWR.n2856 0.0603958
R12409 VDPWR.n2857 VDPWR 0.0603958
R12410 VDPWR VDPWR.n2869 0.0603958
R12411 VDPWR.n2870 VDPWR 0.0603958
R12412 VDPWR.n2870 VDPWR 0.0603958
R12413 VDPWR.n2876 VDPWR 0.0603958
R12414 VDPWR.n2882 VDPWR 0.0603958
R12415 VDPWR.n2900 VDPWR 0.0603958
R12416 VDPWR.n2901 VDPWR 0.0603958
R12417 VDPWR.n2905 VDPWR 0.0603958
R12418 VDPWR.n2948 VDPWR 0.0603958
R12419 VDPWR.n2954 VDPWR 0.0603958
R12420 VDPWR.n2568 VDPWR 0.0603958
R12421 VDPWR.n2604 VDPWR 0.0603958
R12422 VDPWR.n2682 VDPWR 0.0603958
R12423 VDPWR.n2640 VDPWR 0.0603958
R12424 VDPWR.n2640 VDPWR 0.0603958
R12425 VDPWR VDPWR.n2639 0.0603958
R12426 VDPWR.n2631 VDPWR 0.0603958
R12427 VDPWR VDPWR.n2630 0.0603958
R12428 VDPWR VDPWR.n3054 0.0603958
R12429 VDPWR.n3049 VDPWR 0.0603958
R12430 VDPWR.n3047 VDPWR 0.0603958
R12431 VDPWR.n895 VDPWR 0.0603958
R12432 VDPWR.n3017 VDPWR 0.0603958
R12433 VDPWR.n3011 VDPWR 0.0603958
R12434 VDPWR.n2379 VDPWR 0.0603958
R12435 VDPWR.n2383 VDPWR 0.0603958
R12436 VDPWR.n2384 VDPWR 0.0603958
R12437 VDPWR.n2388 VDPWR 0.0603958
R12438 VDPWR VDPWR.n2402 0.0603958
R12439 VDPWR.n2403 VDPWR 0.0603958
R12440 VDPWR VDPWR.n2354 0.0603958
R12441 VDPWR VDPWR.n2408 0.0603958
R12442 VDPWR.n2409 VDPWR 0.0603958
R12443 VDPWR.n2413 VDPWR 0.0603958
R12444 VDPWR VDPWR.n2414 0.0603958
R12445 VDPWR.n2415 VDPWR 0.0603958
R12446 VDPWR.n2529 VDPWR 0.0603958
R12447 VDPWR VDPWR.n2528 0.0603958
R12448 VDPWR VDPWR.n2527 0.0603958
R12449 VDPWR.n2523 VDPWR 0.0603958
R12450 VDPWR.n2439 VDPWR 0.0603958
R12451 VDPWR VDPWR.n2440 0.0603958
R12452 VDPWR.n2511 VDPWR 0.0603958
R12453 VDPWR.n2511 VDPWR 0.0603958
R12454 VDPWR.n2482 VDPWR 0.0603958
R12455 VDPWR VDPWR.n2457 0.0603958
R12456 VDPWR.n2477 VDPWR 0.0603958
R12457 VDPWR.n790 VDPWR 0.0603958
R12458 VDPWR.n3094 VDPWR 0.0603958
R12459 VDPWR VDPWR.n3093 0.0603958
R12460 VDPWR VDPWR.n794 0.0603958
R12461 VDPWR.n3082 VDPWR 0.0603958
R12462 VDPWR.n3078 VDPWR 0.0603958
R12463 VDPWR VDPWR.n861 0.0603958
R12464 VDPWR.n855 VDPWR 0.0603958
R12465 VDPWR VDPWR.n853 0.0603958
R12466 VDPWR.n850 VDPWR 0.0603958
R12467 VDPWR.n82 VDPWR 0.0603958
R12468 VDPWR VDPWR.n81 0.0603958
R12469 VDPWR.n76 VDPWR 0.0603958
R12470 VDPWR.n71 VDPWR 0.0603958
R12471 VDPWR.n66 VDPWR 0.0603958
R12472 VDPWR.n42 VDPWR 0.0603958
R12473 VDPWR VDPWR.n41 0.0603958
R12474 VDPWR VDPWR.n25 0.0603958
R12475 VDPWR.n101 VDPWR 0.0603958
R12476 VDPWR VDPWR.n100 0.0603958
R12477 VDPWR.n110 VDPWR 0.0603958
R12478 VDPWR.n20 VDPWR 0.0603958
R12479 VDPWR.n3115 VDPWR.n3114 0.0600933
R12480 VDPWR.n561 VDPWR 0.0590938
R12481 VDPWR.n281 VDPWR 0.0590938
R12482 VDPWR.n23 VDPWR 0.0590938
R12483 VDPWR.n3166 VDPWR.n759 0.0589638
R12484 VDPWR.n1911 VDPWR 0.0577917
R12485 VDPWR.n2758 VDPWR 0.0577917
R12486 VDPWR.n810 VDPWR 0.0577917
R12487 VDPWR.n2693 VDPWR.n2692 0.0574697
R12488 VDPWR.n2663 VDPWR.n2662 0.0574697
R12489 VDPWR.n1301 VDPWR.n1300 0.0574697
R12490 VDPWR.n1318 VDPWR.n1317 0.0574697
R12491 VDPWR.n1332 VDPWR.n1331 0.0574697
R12492 VDPWR.n1384 VDPWR.n1346 0.0574697
R12493 VDPWR.n1554 VDPWR.n1532 0.0574697
R12494 VDPWR.n1580 VDPWR.n1286 0.0574697
R12495 VDPWR.n1229 VDPWR.n1227 0.0574697
R12496 VDPWR.n1247 VDPWR.n1244 0.0574697
R12497 VDPWR.n1268 VDPWR.n1266 0.0574697
R12498 VDPWR.n1676 VDPWR.n1282 0.0574697
R12499 VDPWR.n1902 VDPWR.n1196 0.0574697
R12500 VDPWR.n1859 VDPWR.n1858 0.0574697
R12501 VDPWR.n1163 VDPWR.n1161 0.0574697
R12502 VDPWR.n2035 VDPWR.n2034 0.0574697
R12503 VDPWR.n2064 VDPWR.n1118 0.0574697
R12504 VDPWR.n1659 VDPWR.n1597 0.0574697
R12505 VDPWR.n1953 VDPWR.n1931 0.0574697
R12506 VDPWR.n1976 VDPWR.n1190 0.0574697
R12507 VDPWR.n1022 VDPWR.n1014 0.0574697
R12508 VDPWR.n2236 VDPWR.n1093 0.0574697
R12509 VDPWR.n2074 VDPWR.n1115 0.0574697
R12510 VDPWR.n2124 VDPWR.n2087 0.0574697
R12511 VDPWR.n2259 VDPWR.n2258 0.0574697
R12512 VDPWR.n2292 VDPWR.n1045 0.0574697
R12513 VDPWR.n2896 VDPWR.n957 0.0574697
R12514 VDPWR.n975 VDPWR.n972 0.0574697
R12515 VDPWR.n990 VDPWR.n987 0.0574697
R12516 VDPWR.n2720 VDPWR.n1008 0.0574697
R12517 VDPWR.n2979 VDPWR.n926 0.0574697
R12518 VDPWR.n944 VDPWR.n942 0.0574697
R12519 VDPWR.n3034 VDPWR.n3032 0.0574697
R12520 VDPWR.n882 VDPWR.n874 0.0574697
R12521 VDPWR.n2572 VDPWR.n2338 0.0574697
R12522 VDPWR.n2718 VDPWR.n2541 0.0574697
R12523 VDPWR.n3006 VDPWR.n3005 0.0574697
R12524 VDPWR.n1335 VDPWR.n1333 0.0551875
R12525 VDPWR.n1271 VDPWR.n1269 0.0551875
R12526 VDPWR.n1121 VDPWR.n1119 0.0551875
R12527 VDPWR.n2152 VDPWR.n2075 0.0551875
R12528 VDPWR.n993 VDPWR.n991 0.0551875
R12529 VDPWR.n2696 VDPWR.n2588 0.0551875
R12530 VDPWR.n2425 VDPWR.n2424 0.0551875
R12531 VDPWR.n752 VDPWR.n751 0.0540714
R12532 VDPWR.n466 VDPWR.n403 0.054
R12533 VDPWR.n1534 VDPWR 0.0538854
R12534 VDPWR.n2533 VDPWR 0.0538854
R12535 VDPWR VDPWR.n2467 0.0538854
R12536 VDPWR.n3176 VDPWR 0.0535303
R12537 VDPWR.n3116 VDPWR.n3115 0.0529556
R12538 VDPWR.n653 VDPWR 0.0525833
R12539 VDPWR.n373 VDPWR 0.0525833
R12540 VDPWR VDPWR.n1956 0.0525833
R12541 VDPWR.n2600 VDPWR 0.0525833
R12542 VDPWR.n2428 VDPWR 0.0525833
R12543 VDPWR.n2466 VDPWR 0.0525833
R12544 VDPWR.n115 VDPWR 0.0525833
R12545 VDPWR.n2290 VDPWR.n1046 0.0522
R12546 VDPWR.n2331 VDPWR.n1012 0.0522
R12547 VDPWR.n2250 VDPWR.n2249 0.0522
R12548 VDPWR.n1596 VDPWR.n1009 0.0522
R12549 VDPWR.n2256 VDPWR.n2255 0.0522
R12550 VDPWR.n2159 VDPWR.n2073 0.0522
R12551 VDPWR.n2507 VDPWR.n2506 0.051025
R12552 VDPWR VDPWR.n754 0.0500269
R12553 VDPWR.n1381 VDPWR.n1380 0.0499792
R12554 VDPWR.n1452 VDPWR.n1451 0.0499792
R12555 VDPWR.n1517 VDPWR.n1287 0.0499792
R12556 VDPWR.n1706 VDPWR.n1681 0.0499792
R12557 VDPWR.n1780 VDPWR.n1779 0.0499792
R12558 VDPWR.n1851 VDPWR.n1217 0.0499792
R12559 VDPWR.n1664 VDPWR.n1600 0.0499792
R12560 VDPWR.n1147 VDPWR.n1143 0.0499792
R12561 VDPWR VDPWR.n1187 0.0499792
R12562 VDPWR.n2121 VDPWR.n2120 0.0499792
R12563 VDPWR.n2245 VDPWR.n2244 0.0499792
R12564 VDPWR.n2296 VDPWR.n1037 0.0499792
R12565 VDPWR.n2748 VDPWR.n2725 0.0499792
R12566 VDPWR.n2840 VDPWR.n2839 0.0499792
R12567 VDPWR.n947 VDPWR.n945 0.0499792
R12568 VDPWR.n2577 VDPWR.n2576 0.0499792
R12569 VDPWR.n2651 VDPWR.n2650 0.0499792
R12570 VDPWR.n3038 VDPWR.n901 0.0499792
R12571 VDPWR.n2396 VDPWR.n2360 0.0499792
R12572 VDPWR.n2448 VDPWR.n2447 0.0499792
R12573 VDPWR.n3076 VDPWR.n801 0.0499792
R12574 VDPWR VDPWR.n2510 0.047375
R12575 VDPWR.n653 VDPWR.n652 0.0460729
R12576 VDPWR.n373 VDPWR.n372 0.0460729
R12577 VDPWR.n115 VDPWR.n114 0.0460729
R12578 VDPWR.n3108 VDPWR.n777 0.0460404
R12579 VDPWR.n781 VDPWR.n780 0.0460404
R12580 VDPWR.n3112 VDPWR.n3111 0.0460404
R12581 VDPWR.n2501 VDPWR.n2500 0.0454816
R12582 VDPWR.n1336 VDPWR.n1329 0.0447708
R12583 VDPWR.n1484 VDPWR.n1306 0.0447708
R12584 VDPWR.n1535 VDPWR.n1534 0.0447708
R12585 VDPWR.n1272 VDPWR.n1264 0.0447708
R12586 VDPWR.n1812 VDPWR.n1234 0.0447708
R12587 VDPWR.n1892 VDPWR.n1890 0.0447708
R12588 VDPWR.n2062 VDPWR.n2061 0.0447708
R12589 VDPWR.n1175 VDPWR.n1173 0.0447708
R12590 VDPWR.n1971 VDPWR.n1914 0.0447708
R12591 VDPWR.n1934 VDPWR.n1933 0.0447708
R12592 VDPWR.n2164 VDPWR.n2163 0.0447708
R12593 VDPWR.n2323 VDPWR.n1017 0.0447708
R12594 VDPWR.n2262 VDPWR.n1077 0.0447708
R12595 VDPWR.n994 VDPWR.n985 0.0447708
R12596 VDPWR.n2893 VDPWR.n2892 0.0447708
R12597 VDPWR.n2969 VDPWR.n2967 0.0447708
R12598 VDPWR.n2601 VDPWR.n2593 0.0447708
R12599 VDPWR.n3059 VDPWR.n877 0.0447708
R12600 VDPWR.n3029 VDPWR.n907 0.0447708
R12601 VDPWR.n2993 VDPWR.n2992 0.0447708
R12602 VDPWR.n2533 VDPWR.n2532 0.0447708
R12603 VDPWR.n2467 VDPWR.n787 0.0447708
R12604 VDPWR.n866 VDPWR.n806 0.0447708
R12605 VDPWR.n845 VDPWR.n844 0.0447708
R12606 VDPWR.n2503 VDPWR.n2340 0.0446687
R12607 VDPWR.n2590 VDPWR.n2589 0.0410405
R12608 VDPWR.n2592 VDPWR.n2591 0.0410405
R12609 VDPWR.n2616 VDPWR.n2615 0.0410405
R12610 VDPWR.n2618 VDPWR.n2617 0.0410405
R12611 VDPWR.n2498 VDPWR.n2444 0.0410405
R12612 VDPWR.n2494 VDPWR.n2445 0.0410405
R12613 VDPWR.n1489 VDPWR.n1303 0.0410405
R12614 VDPWR.n1304 VDPWR.n1299 0.0410405
R12615 VDPWR.n1453 VDPWR.n1320 0.0410405
R12616 VDPWR.n1448 VDPWR.n1316 0.0410405
R12617 VDPWR.n1420 VDPWR.n1334 0.0410405
R12618 VDPWR.n1416 VDPWR.n1330 0.0410405
R12619 VDPWR.n1371 VDPWR.n1347 0.0410405
R12620 VDPWR.n1383 VDPWR.n1345 0.0410405
R12621 VDPWR.n1553 VDPWR.n1530 0.0410405
R12622 VDPWR.n1544 VDPWR.n1533 0.0410405
R12623 VDPWR.n1585 VDPWR.n1288 0.0410405
R12624 VDPWR.n1581 VDPWR.n1579 0.0410405
R12625 VDPWR.n1817 VDPWR.n1231 0.0410405
R12626 VDPWR.n1232 VDPWR.n1226 0.0410405
R12627 VDPWR.n1781 VDPWR.n1249 0.0410405
R12628 VDPWR.n1252 VDPWR.n1243 0.0410405
R12629 VDPWR.n1751 VDPWR.n1270 0.0410405
R12630 VDPWR.n1747 VDPWR.n1265 0.0410405
R12631 VDPWR.n1711 VDPWR.n1678 0.0410405
R12632 VDPWR.n1679 VDPWR.n1281 0.0410405
R12633 VDPWR.n1889 VDPWR.n1888 0.0410405
R12634 VDPWR.n1901 VDPWR.n1900 0.0410405
R12635 VDPWR.n1855 VDPWR.n1216 0.0410405
R12636 VDPWR.n1862 VDPWR.n1215 0.0410405
R12637 VDPWR.n1170 VDPWR.n1160 0.0410405
R12638 VDPWR.n1171 VDPWR.n1164 0.0410405
R12639 VDPWR.n1137 VDPWR.n1136 0.0410405
R12640 VDPWR.n1139 VDPWR.n1138 0.0410405
R12641 VDPWR.n2069 VDPWR.n1120 0.0410405
R12642 VDPWR.n2065 VDPWR.n2063 0.0410405
R12643 VDPWR.n1669 VDPWR.n1599 0.0410405
R12644 VDPWR.n1662 VDPWR.n1660 0.0410405
R12645 VDPWR.n1952 VDPWR.n1930 0.0410405
R12646 VDPWR.n1943 VDPWR.n1932 0.0410405
R12647 VDPWR.n1978 VDPWR.n1977 0.0410405
R12648 VDPWR.n1910 VDPWR.n1909 0.0410405
R12649 VDPWR.n2328 VDPWR.n1016 0.0410405
R12650 VDPWR.n2321 VDPWR.n1023 0.0410405
R12651 VDPWR.n2246 VDPWR.n1095 0.0410405
R12652 VDPWR.n2238 VDPWR.n2237 0.0410405
R12653 VDPWR.n2156 VDPWR.n2076 0.0410405
R12654 VDPWR.n2162 VDPWR.n1114 0.0410405
R12655 VDPWR.n2110 VDPWR.n2088 0.0410405
R12656 VDPWR.n2123 VDPWR.n2086 0.0410405
R12657 VDPWR.n2261 VDPWR.n2260 0.0410405
R12658 VDPWR.n1082 VDPWR.n1081 0.0410405
R12659 VDPWR.n2294 VDPWR.n2293 0.0410405
R12660 VDPWR.n1048 VDPWR.n1047 0.0410405
R12661 VDPWR.n2878 VDPWR.n958 0.0410405
R12662 VDPWR.n2895 VDPWR.n956 0.0410405
R12663 VDPWR.n2841 VDPWR.n978 0.0410405
R12664 VDPWR.n2847 VDPWR.n971 0.0410405
R12665 VDPWR.n2802 VDPWR.n992 0.0410405
R12666 VDPWR.n2798 VDPWR.n986 0.0410405
R12667 VDPWR.n2752 VDPWR.n2722 0.0410405
R12668 VDPWR.n2723 VDPWR.n1007 0.0410405
R12669 VDPWR.n2966 VDPWR.n2965 0.0410405
R12670 VDPWR.n2978 VDPWR.n2977 0.0410405
R12671 VDPWR.n2929 VDPWR.n946 0.0410405
R12672 VDPWR.n2925 VDPWR.n941 0.0410405
R12673 VDPWR.n3036 VDPWR.n3035 0.0410405
R12674 VDPWR.n906 VDPWR.n905 0.0410405
R12675 VDPWR.n3064 VDPWR.n876 0.0410405
R12676 VDPWR.n3057 VDPWR.n883 0.0410405
R12677 VDPWR.n2465 VDPWR.n783 0.0410405
R12678 VDPWR.n3101 VDPWR.n3100 0.0410405
R12679 VDPWR.n2573 VDPWR.n2571 0.0410405
R12680 VDPWR.n2574 VDPWR.n2542 0.0410405
R12681 VDPWR.n2983 VDPWR.n922 0.0410405
R12682 VDPWR.n2985 VDPWR.n2984 0.0410405
R12683 VDPWR.n2426 VDPWR.n2341 0.0410405
R12684 VDPWR.n2535 VDPWR.n2534 0.0410405
R12685 VDPWR.n2390 VDPWR.n2364 0.0410405
R12686 VDPWR.n2394 VDPWR.n2362 0.0410405
R12687 VDPWR.n846 VDPWR.n773 0.0410405
R12688 VDPWR.n839 VDPWR.n774 0.0410405
R12689 VDPWR.n803 VDPWR.n802 0.0410405
R12690 VDPWR.n869 VDPWR.n868 0.0410405
R12691 VDPWR.n1589 VDPWR.n1588 0.04045
R12692 VDPWR.n1492 VDPWR.n1228 0.04045
R12693 VDPWR.n1456 VDPWR.n1245 0.04045
R12694 VDPWR.n1594 VDPWR.n1283 0.04045
R12695 VDPWR.n1531 VDPWR.n1193 0.04045
R12696 VDPWR.n1423 VDPWR.n1267 0.04045
R12697 VDPWR.n255 VDPWR.n254 0.0403788
R12698 VDPWR VDPWR.n376 0.0403708
R12699 VDPWR.n1426 VDPWR.n1329 0.0395625
R12700 VDPWR.n1459 VDPWR.n1313 0.0395625
R12701 VDPWR.n1484 VDPWR.n1483 0.0395625
R12702 VDPWR.n1578 VDPWR.n1577 0.0395625
R12703 VDPWR.n1551 VDPWR.n1535 0.0395625
R12704 VDPWR.n1757 VDPWR.n1264 0.0395625
R12705 VDPWR.n1788 VDPWR.n1787 0.0395625
R12706 VDPWR.n1812 VDPWR.n1811 0.0395625
R12707 VDPWR.n1864 VDPWR.n1863 0.0395625
R12708 VDPWR.n1892 VDPWR.n1891 0.0395625
R12709 VDPWR.n2061 VDPWR.n1124 0.0395625
R12710 VDPWR.n2031 VDPWR.n2030 0.0395625
R12711 VDPWR.n1175 VDPWR.n1174 0.0395625
R12712 VDPWR.n1914 VDPWR.n1913 0.0395625
R12713 VDPWR.n1950 VDPWR.n1934 0.0395625
R12714 VDPWR.n2164 VDPWR.n1111 0.0395625
R12715 VDPWR.n2240 VDPWR.n2234 0.0395625
R12716 VDPWR.n2323 VDPWR.n2322 0.0395625
R12717 VDPWR.n1055 VDPWR.n1054 0.0395625
R12718 VDPWR.n1083 VDPWR.n1077 0.0395625
R12719 VDPWR.n2808 VDPWR.n985 0.0395625
R12720 VDPWR.n2855 VDPWR.n968 0.0395625
R12721 VDPWR.n2892 VDPWR.n960 0.0395625
R12722 VDPWR.n2936 VDPWR.n940 0.0395625
R12723 VDPWR.n2969 VDPWR.n2968 0.0395625
R12724 VDPWR.n2689 VDPWR.n2593 0.0395625
R12725 VDPWR.n2659 VDPWR.n2658 0.0395625
R12726 VDPWR.n3059 VDPWR.n3058 0.0395625
R12727 VDPWR.n909 VDPWR.n907 0.0395625
R12728 VDPWR.n2995 VDPWR.n2993 0.0395625
R12729 VDPWR.n2532 VDPWR.n2346 0.0395625
R12730 VDPWR.n2489 VDPWR.n2449 0.0395625
R12731 VDPWR.n3099 VDPWR.n787 0.0395625
R12732 VDPWR.n867 VDPWR.n866 0.0395625
R12733 VDPWR.n844 VDPWR.n829 0.0395625
R12734 VDPWR.n580 VDPWR 0.0382604
R12735 VDPWR.n300 VDPWR 0.0382604
R12736 VDPWR.n42 VDPWR 0.0382604
R12737 VDPWR.n2492 VDPWR.n2491 0.0382581
R12738 VDPWR.n755 VDPWR 0.0376452
R12739 VDPWR VDPWR.n595 0.0369583
R12740 VDPWR VDPWR.n315 0.0369583
R12741 VDPWR VDPWR.n57 0.0369583
R12742 VDPWR.n2506 VDPWR 0.036925
R12743 VDPWR.n3108 VDPWR 0.0366988
R12744 VDPWR.n780 VDPWR 0.0366988
R12745 VDPWR.n3111 VDPWR 0.0366988
R12746 VDPWR VDPWR.n2501 0.0362546
R12747 VDPWR.n2503 VDPWR 0.0356084
R12748 VDPWR.n1380 VDPWR.n1344 0.0343542
R12749 VDPWR.n1451 VDPWR.n1450 0.0343542
R12750 VDPWR.n1548 VDPWR.n1547 0.0343542
R12751 VDPWR.n1706 VDPWR.n1280 0.0343542
R12752 VDPWR.n1779 VDPWR.n1254 0.0343542
R12753 VDPWR.n1854 VDPWR.n1851 0.0343542
R12754 VDPWR.n1898 VDPWR.n1897 0.0343542
R12755 VDPWR.n1664 VDPWR.n1663 0.0343542
R12756 VDPWR.n1147 VDPWR.n1146 0.0343542
R12757 VDPWR.n1947 VDPWR.n1946 0.0343542
R12758 VDPWR.n2120 VDPWR.n2085 0.0343542
R12759 VDPWR.n2244 VDPWR.n1097 0.0343542
R12760 VDPWR.n2296 VDPWR.n2295 0.0343542
R12761 VDPWR.n1087 VDPWR.n1086 0.0343542
R12762 VDPWR.n2839 VDPWR.n970 0.0343542
R12763 VDPWR.n2928 VDPWR.n947 0.0343542
R12764 VDPWR.n2975 VDPWR.n2974 0.0343542
R12765 VDPWR.n2577 VDPWR.n2543 0.0343542
R12766 VDPWR.n2653 VDPWR.n2651 0.0343542
R12767 VDPWR.n3038 VDPWR.n3037 0.0343542
R12768 VDPWR.n3002 VDPWR.n3001 0.0343542
R12769 VDPWR.n2396 VDPWR.n2395 0.0343542
R12770 VDPWR.n2496 VDPWR.n2448 0.0343542
R12771 VDPWR.n809 VDPWR.n801 0.0343542
R12772 VDPWR.n842 VDPWR.n841 0.0343542
R12773 VDPWR VDPWR.n1500 0.0330521
R12774 VDPWR VDPWR.n2745 0.0330521
R12775 VDPWR VDPWR.n2819 0.0330521
R12776 VDPWR.n2901 VDPWR 0.0330521
R12777 VDPWR VDPWR.n2382 0.0330521
R12778 VDPWR.n3094 VDPWR 0.0330521
R12779 VDPWR.n620 VDPWR 0.03175
R12780 VDPWR.n639 VDPWR 0.03175
R12781 VDPWR.n340 VDPWR 0.03175
R12782 VDPWR.n359 VDPWR 0.03175
R12783 VDPWR.n142 VDPWR.n138 0.03175
R12784 VDPWR.n173 VDPWR.n172 0.03175
R12785 VDPWR.n172 VDPWR.n151 0.03175
R12786 VDPWR.n168 VDPWR.n167 0.03175
R12787 VDPWR.n167 VDPWR.n166 0.03175
R12788 VDPWR.n163 VDPWR.n162 0.03175
R12789 VDPWR.n162 VDPWR.n161 0.03175
R12790 VDPWR.n158 VDPWR.n157 0.03175
R12791 VDPWR.n157 VDPWR.n156 0.03175
R12792 VDPWR.n201 VDPWR.n128 0.03175
R12793 VDPWR.n197 VDPWR.n196 0.03175
R12794 VDPWR.n196 VDPWR.n195 0.03175
R12795 VDPWR.n192 VDPWR.n191 0.03175
R12796 VDPWR.n191 VDPWR.n190 0.03175
R12797 VDPWR.n187 VDPWR.n186 0.03175
R12798 VDPWR.n186 VDPWR.n185 0.03175
R12799 VDPWR.n182 VDPWR.n181 0.03175
R12800 VDPWR.n181 VDPWR.n180 0.03175
R12801 VDPWR VDPWR.n1432 0.03175
R12802 VDPWR VDPWR.n1496 0.03175
R12803 VDPWR.n1497 VDPWR 0.03175
R12804 VDPWR.n1759 VDPWR 0.03175
R12805 VDPWR VDPWR.n1763 0.03175
R12806 VDPWR.n1824 VDPWR 0.03175
R12807 VDPWR VDPWR.n1883 0.03175
R12808 VDPWR.n2056 VDPWR 0.03175
R12809 VDPWR.n2002 VDPWR 0.03175
R12810 VDPWR.n1965 VDPWR 0.03175
R12811 VDPWR VDPWR.n2169 0.03175
R12812 VDPWR.n2170 VDPWR 0.03175
R12813 VDPWR.n2214 VDPWR 0.03175
R12814 VDPWR.n2318 VDPWR 0.03175
R12815 VDPWR.n2737 VDPWR 0.03175
R12816 VDPWR.n2810 VDPWR 0.03175
R12817 VDPWR VDPWR.n2876 0.03175
R12818 VDPWR VDPWR.n2900 0.03175
R12819 VDPWR VDPWR.n2598 0.03175
R12820 VDPWR VDPWR.n2604 0.03175
R12821 VDPWR.n2409 VDPWR 0.03175
R12822 VDPWR VDPWR.n2427 0.03175
R12823 VDPWR.n2528 VDPWR 0.03175
R12824 VDPWR.n2527 VDPWR 0.03175
R12825 VDPWR VDPWR.n2443 0.03175
R12826 VDPWR.n2477 VDPWR 0.03175
R12827 VDPWR VDPWR.n2464 0.03175
R12828 VDPWR VDPWR.n790 0.03175
R12829 VDPWR.n811 VDPWR 0.03175
R12830 VDPWR.n853 VDPWR 0.03175
R12831 VDPWR.n82 VDPWR 0.03175
R12832 VDPWR.n101 VDPWR 0.03175
R12833 VDPWR.n1555 VDPWR.n1554 0.0292489
R12834 VDPWR.n1545 VDPWR.n1532 0.0292489
R12835 VDPWR.n1196 VDPWR.n1194 0.0292489
R12836 VDPWR.n1903 VDPWR.n1902 0.0292489
R12837 VDPWR.n1954 VDPWR.n1953 0.0292489
R12838 VDPWR.n1944 VDPWR.n1931 0.0292489
R12839 VDPWR.n2259 VDPWR.n1080 0.0292489
R12840 VDPWR.n2258 VDPWR.n2257 0.0292489
R12841 VDPWR.n926 VDPWR.n924 0.0292489
R12842 VDPWR.n2980 VDPWR.n2979 0.0292489
R12843 VDPWR.n3034 VDPWR.n3033 0.0292489
R12844 VDPWR.n3032 VDPWR.n3031 0.0292489
R12845 VDPWR.n2931 VDPWR.n944 0.0292489
R12846 VDPWR.n2933 VDPWR.n942 0.0292489
R12847 VDPWR.n2292 VDPWR.n2291 0.0292489
R12848 VDPWR.n2289 VDPWR.n1045 0.0292489
R12849 VDPWR.n1976 VDPWR.n1975 0.0292489
R12850 VDPWR.n1973 VDPWR.n1190 0.0292489
R12851 VDPWR.n1858 VDPWR.n1857 0.0292489
R12852 VDPWR.n1860 VDPWR.n1859 0.0292489
R12853 VDPWR.n1587 VDPWR.n1286 0.0292489
R12854 VDPWR.n1580 VDPWR.n1285 0.0292489
R12855 VDPWR.n3066 VDPWR.n874 0.0292489
R12856 VDPWR.n882 VDPWR.n873 0.0292489
R12857 VDPWR.n2879 VDPWR.n957 0.0292489
R12858 VDPWR.n2897 VDPWR.n2896 0.0292489
R12859 VDPWR.n2330 VDPWR.n1014 0.0292489
R12860 VDPWR.n1022 VDPWR.n1013 0.0292489
R12861 VDPWR.n2007 VDPWR.n1161 0.0292489
R12862 VDPWR.n2005 VDPWR.n1163 0.0292489
R12863 VDPWR.n1819 VDPWR.n1229 0.0292489
R12864 VDPWR.n1821 VDPWR.n1227 0.0292489
R12865 VDPWR.n1491 VDPWR.n1301 0.0292489
R12866 VDPWR.n1493 VDPWR.n1300 0.0292489
R12867 VDPWR.n2664 VDPWR.n2663 0.0292489
R12868 VDPWR.n2662 VDPWR.n2661 0.0292489
R12869 VDPWR.n2843 VDPWR.n975 0.0292489
R12870 VDPWR.n2845 VDPWR.n972 0.0292489
R12871 VDPWR.n2248 VDPWR.n1093 0.0292489
R12872 VDPWR.n2236 VDPWR.n1092 0.0292489
R12873 VDPWR.n2036 VDPWR.n2035 0.0292489
R12874 VDPWR.n2034 VDPWR.n2033 0.0292489
R12875 VDPWR.n1783 VDPWR.n1247 0.0292489
R12876 VDPWR.n1785 VDPWR.n1244 0.0292489
R12877 VDPWR.n1455 VDPWR.n1318 0.0292489
R12878 VDPWR.n1457 VDPWR.n1317 0.0292489
R12879 VDPWR.n2754 VDPWR.n2720 0.0292489
R12880 VDPWR.n2756 VDPWR.n1008 0.0292489
R12881 VDPWR.n2111 VDPWR.n2087 0.0292489
R12882 VDPWR.n2125 VDPWR.n2124 0.0292489
R12883 VDPWR.n1671 VDPWR.n1597 0.0292489
R12884 VDPWR.n1659 VDPWR.n1595 0.0292489
R12885 VDPWR.n1713 VDPWR.n1676 0.0292489
R12886 VDPWR.n1715 VDPWR.n1282 0.0292489
R12887 VDPWR.n1372 VDPWR.n1346 0.0292489
R12888 VDPWR.n1385 VDPWR.n1384 0.0292489
R12889 VDPWR.n2541 VDPWR.n2337 0.0292489
R12890 VDPWR.n2572 VDPWR.n2337 0.0292489
R12891 VDPWR.n3007 VDPWR.n3006 0.0292489
R12892 VDPWR.n3005 VDPWR.n3004 0.0292489
R12893 VDPWR.n2694 VDPWR.n2693 0.0292489
R12894 VDPWR.n2692 VDPWR.n2691 0.0292489
R12895 VDPWR.n2804 VDPWR.n990 0.0292489
R12896 VDPWR.n2806 VDPWR.n987 0.0292489
R12897 VDPWR.n2158 VDPWR.n2074 0.0292489
R12898 VDPWR.n2160 VDPWR.n1115 0.0292489
R12899 VDPWR.n2071 VDPWR.n1118 0.0292489
R12900 VDPWR.n2064 VDPWR.n1117 0.0292489
R12901 VDPWR.n1753 VDPWR.n1268 0.0292489
R12902 VDPWR.n1755 VDPWR.n1266 0.0292489
R12903 VDPWR.n1422 VDPWR.n1332 0.0292489
R12904 VDPWR.n1424 VDPWR.n1331 0.0292489
R12905 VDPWR.n586 VDPWR.n585 0.0291458
R12906 VDPWR.n306 VDPWR.n305 0.0291458
R12907 VDPWR.n1419 VDPWR.n1335 0.0291458
R12908 VDPWR.n1479 VDPWR.n1302 0.0291458
R12909 VDPWR.n1750 VDPWR.n1271 0.0291458
R12910 VDPWR.n1808 VDPWR.n1230 0.0291458
R12911 VDPWR.n2068 VDPWR.n1121 0.0291458
R12912 VDPWR.n2010 VDPWR.n2009 0.0291458
R12913 VDPWR.n2155 VDPWR.n2152 0.0291458
R12914 VDPWR.n2213 VDPWR.n1015 0.0291458
R12915 VDPWR.n2801 VDPWR.n993 0.0291458
R12916 VDPWR.n2882 VDPWR.n2881 0.0291458
R12917 VDPWR.n2630 VDPWR.n875 0.0291458
R12918 VDPWR.n48 VDPWR.n47 0.0291458
R12919 VDPWR.n753 VDPWR.n752 0.0281786
R12920 VDPWR.n1979 VDPWR 0.0265417
R12921 VDPWR.n2747 VDPWR 0.0265417
R12922 VDPWR VDPWR.n809 0.0265417
R12923 VDPWR.n202 VDPWR.n127 0.0249565
R12924 VDPWR.n727 VDPWR.n725 0.0247347
R12925 VDPWR.n1375 VDPWR.n1374 0.0239375
R12926 VDPWR.n1703 VDPWR.n1677 0.0239375
R12927 VDPWR.n1607 VDPWR.n1598 0.0239375
R12928 VDPWR.n2114 VDPWR.n2113 0.0239375
R12929 VDPWR VDPWR.n2831 0.0239375
R12930 VDPWR.n2569 VDPWR.n2568 0.0239375
R12931 VDPWR.n3011 VDPWR 0.0239375
R12932 VDPWR.n2367 VDPWR.n2365 0.0239375
R12933 VDPWR.n655 VDPWR 0.0236148
R12934 VDPWR VDPWR.n3178 0.0236148
R12935 VDPWR.n728 VDPWR.n723 0.0234592
R12936 VDPWR.n1010 VDPWR 0.022975
R12937 VDPWR.n1284 VDPWR 0.022975
R12938 VDPWR.n1906 VDPWR 0.022975
R12939 VDPWR.n2254 VDPWR 0.022975
R12940 VDPWR.n3070 VDPWR 0.022975
R12941 VDPWR.n3110 VDPWR 0.022975
R12942 VDPWR VDPWR.n567 0.0226354
R12943 VDPWR VDPWR.n592 0.0226354
R12944 VDPWR.n612 VDPWR 0.0226354
R12945 VDPWR.n607 VDPWR 0.0226354
R12946 VDPWR.n599 VDPWR 0.0226354
R12947 VDPWR VDPWR.n569 0.0226354
R12948 VDPWR.n579 VDPWR 0.0226354
R12949 VDPWR.n629 VDPWR 0.0226354
R12950 VDPWR VDPWR.n637 0.0226354
R12951 VDPWR.n638 VDPWR 0.0226354
R12952 VDPWR VDPWR.n538 0.0226354
R12953 VDPWR VDPWR.n542 0.0226354
R12954 VDPWR VDPWR.n547 0.0226354
R12955 VDPWR.n552 VDPWR 0.0226354
R12956 VDPWR VDPWR.n287 0.0226354
R12957 VDPWR VDPWR.n312 0.0226354
R12958 VDPWR.n332 VDPWR 0.0226354
R12959 VDPWR.n327 VDPWR 0.0226354
R12960 VDPWR.n319 VDPWR 0.0226354
R12961 VDPWR VDPWR.n289 0.0226354
R12962 VDPWR.n299 VDPWR 0.0226354
R12963 VDPWR.n349 VDPWR 0.0226354
R12964 VDPWR VDPWR.n357 0.0226354
R12965 VDPWR.n358 VDPWR 0.0226354
R12966 VDPWR VDPWR.n258 0.0226354
R12967 VDPWR VDPWR.n262 0.0226354
R12968 VDPWR VDPWR.n267 0.0226354
R12969 VDPWR.n272 VDPWR 0.0226354
R12970 VDPWR VDPWR.n1394 0.0226354
R12971 VDPWR.n1401 VDPWR 0.0226354
R12972 VDPWR.n1427 VDPWR 0.0226354
R12973 VDPWR.n1515 VDPWR 0.0226354
R12974 VDPWR.n1517 VDPWR 0.0226354
R12975 VDPWR.n1577 VDPWR 0.0226354
R12976 VDPWR.n1522 VDPWR 0.0226354
R12977 VDPWR VDPWR.n1529 0.0226354
R12978 VDPWR.n1548 VDPWR 0.0226354
R12979 VDPWR VDPWR.n1724 0.0226354
R12980 VDPWR.n1731 VDPWR 0.0226354
R12981 VDPWR VDPWR.n1758 0.0226354
R12982 VDPWR VDPWR.n1793 0.0226354
R12983 VDPWR VDPWR.n1831 0.0226354
R12984 VDPWR VDPWR.n1837 0.0226354
R12985 VDPWR.n1864 VDPWR 0.0226354
R12986 VDPWR VDPWR.n1212 0.0226354
R12987 VDPWR.n1880 VDPWR 0.0226354
R12988 VDPWR.n1885 VDPWR 0.0226354
R12989 VDPWR.n1897 VDPWR 0.0226354
R12990 VDPWR.n1651 VDPWR 0.0226354
R12991 VDPWR.n1642 VDPWR 0.0226354
R12992 VDPWR.n2057 VDPWR 0.0226354
R12993 VDPWR.n2042 VDPWR 0.0226354
R12994 VDPWR.n2025 VDPWR 0.0226354
R12995 VDPWR.n2018 VDPWR 0.0226354
R12996 VDPWR.n1993 VDPWR 0.0226354
R12997 VDPWR.n1992 VDPWR 0.0226354
R12998 VDPWR.n1963 VDPWR 0.0226354
R12999 VDPWR VDPWR.n1929 0.0226354
R13000 VDPWR.n1947 VDPWR 0.0226354
R13001 VDPWR.n2105 VDPWR 0.0226354
R13002 VDPWR.n2133 VDPWR 0.0226354
R13003 VDPWR.n2139 VDPWR 0.0226354
R13004 VDPWR VDPWR.n2168 0.0226354
R13005 VDPWR VDPWR.n2174 0.0226354
R13006 VDPWR.n2175 VDPWR 0.0226354
R13007 VDPWR VDPWR.n2182 0.0226354
R13008 VDPWR.n2227 VDPWR 0.0226354
R13009 VDPWR.n2314 VDPWR 0.0226354
R13010 VDPWR.n2313 VDPWR 0.0226354
R13011 VDPWR.n1055 VDPWR 0.0226354
R13012 VDPWR.n2287 VDPWR 0.0226354
R13013 VDPWR.n2263 VDPWR 0.0226354
R13014 VDPWR.n1086 VDPWR 0.0226354
R13015 VDPWR.n2748 VDPWR 0.0226354
R13016 VDPWR.n2759 VDPWR 0.0226354
R13017 VDPWR VDPWR.n2764 0.0226354
R13018 VDPWR.n2779 VDPWR 0.0226354
R13019 VDPWR VDPWR.n2809 0.0226354
R13020 VDPWR.n2820 VDPWR 0.0226354
R13021 VDPWR.n2827 VDPWR 0.0226354
R13022 VDPWR.n2857 VDPWR 0.0226354
R13023 VDPWR.n2936 VDPWR 0.0226354
R13024 VDPWR VDPWR.n2935 0.0226354
R13025 VDPWR.n2943 VDPWR 0.0226354
R13026 VDPWR.n2962 VDPWR 0.0226354
R13027 VDPWR.n2974 VDPWR 0.0226354
R13028 VDPWR VDPWR.n2588 0.0226354
R13029 VDPWR.n2688 VDPWR 0.0226354
R13030 VDPWR.n2655 VDPWR 0.0226354
R13031 VDPWR.n2658 VDPWR 0.0226354
R13032 VDPWR.n2644 VDPWR 0.0226354
R13033 VDPWR.n3054 VDPWR 0.0226354
R13034 VDPWR.n3020 VDPWR 0.0226354
R13035 VDPWR VDPWR.n918 0.0226354
R13036 VDPWR VDPWR.n921 0.0226354
R13037 VDPWR.n3001 VDPWR 0.0226354
R13038 VDPWR.n2379 VDPWR 0.0226354
R13039 VDPWR VDPWR.n2383 0.0226354
R13040 VDPWR.n2403 VDPWR 0.0226354
R13041 VDPWR.n2415 VDPWR 0.0226354
R13042 VDPWR VDPWR.n2425 0.0226354
R13043 VDPWR.n2429 VDPWR 0.0226354
R13044 VDPWR.n2523 VDPWR 0.0226354
R13045 VDPWR.n2516 VDPWR 0.0226354
R13046 VDPWR VDPWR.n2439 0.0226354
R13047 VDPWR VDPWR.n2455 0.0226354
R13048 VDPWR.n2468 VDPWR 0.0226354
R13049 VDPWR.n3093 VDPWR 0.0226354
R13050 VDPWR.n3081 VDPWR 0.0226354
R13051 VDPWR.n3078 VDPWR 0.0226354
R13052 VDPWR.n862 VDPWR 0.0226354
R13053 VDPWR VDPWR.n816 0.0226354
R13054 VDPWR.n855 VDPWR 0.0226354
R13055 VDPWR.n850 VDPWR 0.0226354
R13056 VDPWR VDPWR.n827 0.0226354
R13057 VDPWR.n842 VDPWR 0.0226354
R13058 VDPWR VDPWR.n29 0.0226354
R13059 VDPWR VDPWR.n54 0.0226354
R13060 VDPWR.n74 VDPWR 0.0226354
R13061 VDPWR.n69 VDPWR 0.0226354
R13062 VDPWR.n61 VDPWR 0.0226354
R13063 VDPWR VDPWR.n31 0.0226354
R13064 VDPWR.n41 VDPWR 0.0226354
R13065 VDPWR.n91 VDPWR 0.0226354
R13066 VDPWR VDPWR.n99 0.0226354
R13067 VDPWR.n100 VDPWR 0.0226354
R13068 VDPWR VDPWR.n0 0.0226354
R13069 VDPWR VDPWR.n4 0.0226354
R13070 VDPWR VDPWR.n9 0.0226354
R13071 VDPWR.n14 VDPWR 0.0226354
R13072 VDPWR.n248 VDPWR.n121 0.0226154
R13073 VDPWR.n243 VDPWR.n242 0.0226154
R13074 VDPWR.n238 VDPWR.n237 0.0226154
R13075 VDPWR.n233 VDPWR.n232 0.0226154
R13076 VDPWR.n228 VDPWR.n227 0.0226154
R13077 VDPWR.n223 VDPWR.n222 0.0226154
R13078 VDPWR.n218 VDPWR.n217 0.0226154
R13079 VDPWR.n213 VDPWR.n212 0.0226154
R13080 VDPWR.n208 VDPWR.n207 0.0226154
R13081 VDPWR.n3105 VDPWR.n3104 0.0218125
R13082 VDPWR VDPWR.n1183 0.0213333
R13083 VDPWR.n2950 VDPWR 0.0213333
R13084 VDPWR.n2659 VDPWR 0.0213333
R13085 VDPWR.n2631 VDPWR 0.0213333
R13086 VDPWR.n867 VDPWR 0.0213333
R13087 VDPWR VDPWR.n1495 0.0200312
R13088 VDPWR VDPWR.n1823 0.0200312
R13089 VDPWR.n2003 VDPWR 0.0200312
R13090 VDPWR.n2319 VDPWR 0.0200312
R13091 VDPWR VDPWR.n2899 0.0200312
R13092 VDPWR.n3055 VDPWR 0.0200312
R13093 VDPWR VDPWR.n788 0.0200312
R13094 VDPWR VDPWR.n248 0.0185288
R13095 VDPWR.n243 VDPWR 0.0185288
R13096 VDPWR.n238 VDPWR 0.0185288
R13097 VDPWR.n233 VDPWR 0.0185288
R13098 VDPWR.n223 VDPWR 0.0185288
R13099 VDPWR.n218 VDPWR 0.0185288
R13100 VDPWR.n213 VDPWR 0.0185288
R13101 VDPWR.n208 VDPWR 0.0185288
R13102 VDPWR.n2932 VDPWR.n943 0.018125
R13103 VDPWR.n2332 VDPWR.n872 0.018125
R13104 VDPWR.n2844 VDPWR.n973 0.018125
R13105 VDPWR.n2755 VDPWR.n2336 0.018125
R13106 VDPWR.n2981 VDPWR.n923 0.018125
R13107 VDPWR.n2805 VDPWR.n988 0.018125
R13108 VDPWR.n3072 VDPWR.n870 0.01695
R13109 VDPWR.n3068 VDPWR.n3067 0.01695
R13110 VDPWR.n2499 VDPWR.n974 0.01695
R13111 VDPWR.n2719 VDPWR.n2540 0.01695
R13112 VDPWR.n2982 VDPWR.n775 0.01695
R13113 VDPWR.n2538 VDPWR.n989 0.01695
R13114 VDPWR VDPWR.n137 0.016125
R13115 VDPWR.n149 VDPWR 0.016125
R13116 VDPWR.n150 VDPWR 0.016125
R13117 VDPWR.n174 VDPWR 0.016125
R13118 VDPWR VDPWR.n173 0.016125
R13119 VDPWR.n168 VDPWR 0.016125
R13120 VDPWR.n163 VDPWR 0.016125
R13121 VDPWR.n158 VDPWR 0.016125
R13122 VDPWR VDPWR.n127 0.016125
R13123 VDPWR.n197 VDPWR 0.016125
R13124 VDPWR.n192 VDPWR 0.016125
R13125 VDPWR.n187 VDPWR 0.016125
R13126 VDPWR.n182 VDPWR 0.016125
R13127 VDPWR.n177 VDPWR 0.016125
R13128 VDPWR VDPWR.n1522 0.016125
R13129 VDPWR.n1890 VDPWR 0.016125
R13130 VDPWR.n1933 VDPWR 0.016125
R13131 VDPWR VDPWR.n2262 0.016125
R13132 VDPWR.n2967 VDPWR 0.016125
R13133 VDPWR.n2992 VDPWR 0.016125
R13134 VDPWR.n845 VDPWR 0.016125
R13135 VDPWR.n203 VDPWR 0.0137212
R13136 VDPWR.n1370 VDPWR.n1348 0.0135208
R13137 VDPWR.n1447 VDPWR.n1319 0.0135208
R13138 VDPWR.n1710 VDPWR.n1709 0.0135208
R13139 VDPWR.n1250 VDPWR.n1248 0.0135208
R13140 VDPWR.n1668 VDPWR.n1667 0.0135208
R13141 VDPWR.n2038 VDPWR.n1135 0.0135208
R13142 VDPWR.n2119 VDPWR.n2089 0.0135208
R13143 VDPWR.n1096 VDPWR.n1094 0.0135208
R13144 VDPWR.n2751 VDPWR.n2750 0.0135208
R13145 VDPWR.n2838 VDPWR.n976 0.0135208
R13146 VDPWR.n2570 VDPWR.n2548 0.0135208
R13147 VDPWR.n2666 VDPWR.n2614 0.0135208
R13148 VDPWR.n2389 VDPWR.n2388 0.0135208
R13149 VDPWR.n2510 VDPWR.n2443 0.0135208
R13150 VDPWR.n3117 VDPWR 0.0122968
R13151 VDPWR.n1584 VDPWR 0.0122188
R13152 VDPWR VDPWR.n1979 0.0122188
R13153 VDPWR VDPWR.n2747 0.0122188
R13154 VDPWR VDPWR.n249 0.0115577
R13155 VDPWR VDPWR.n121 0.0115577
R13156 VDPWR.n122 VDPWR 0.0115577
R13157 VDPWR.n242 VDPWR 0.0115577
R13158 VDPWR VDPWR.n241 0.0115577
R13159 VDPWR.n237 VDPWR 0.0115577
R13160 VDPWR VDPWR.n236 0.0115577
R13161 VDPWR.n232 VDPWR 0.0115577
R13162 VDPWR VDPWR.n231 0.0115577
R13163 VDPWR.n227 VDPWR 0.0115577
R13164 VDPWR VDPWR.n226 0.0115577
R13165 VDPWR.n222 VDPWR 0.0115577
R13166 VDPWR VDPWR.n221 0.0115577
R13167 VDPWR.n217 VDPWR 0.0115577
R13168 VDPWR VDPWR.n216 0.0115577
R13169 VDPWR.n212 VDPWR 0.0115577
R13170 VDPWR VDPWR.n211 0.0115577
R13171 VDPWR.n207 VDPWR 0.0115577
R13172 VDPWR.n252 VDPWR 0.0115577
R13173 VDPWR VDPWR.n1287 0.0109167
R13174 VDPWR VDPWR.n2360 0.0109167
R13175 VDPWR.n2447 VDPWR 0.0109167
R13176 VDPWR VDPWR.n3107 0.00972152
R13177 VDPWR.n3106 VDPWR 0.00972152
R13178 VDPWR VDPWR.n778 0.00972152
R13179 VDPWR VDPWR.n2502 0.00972152
R13180 VDPWR.n375 VDPWR.n254 0.00887356
R13181 VDPWR.n137 VDPWR 0.00865217
R13182 VDPWR VDPWR.n149 0.00865217
R13183 VDPWR VDPWR.n150 0.00865217
R13184 VDPWR.n174 VDPWR 0.00865217
R13185 VDPWR.n177 VDPWR 0.00865217
R13186 VDPWR.n1418 VDPWR.n1415 0.0083125
R13187 VDPWR.n1488 VDPWR.n1487 0.0083125
R13188 VDPWR.n1557 VDPWR.n1529 0.0083125
R13189 VDPWR.n1749 VDPWR.n1746 0.0083125
R13190 VDPWR.n1816 VDPWR.n1815 0.0083125
R13191 VDPWR.n1886 VDPWR.n1885 0.0083125
R13192 VDPWR.n2067 VDPWR.n1122 0.0083125
R13193 VDPWR.n1169 VDPWR.n1159 0.0083125
R13194 VDPWR.n1956 VDPWR.n1929 0.0083125
R13195 VDPWR.n2154 VDPWR.n1113 0.0083125
R13196 VDPWR.n2327 VDPWR.n2326 0.0083125
R13197 VDPWR.n2263 VDPWR.n1076 0.0083125
R13198 VDPWR.n2800 VDPWR.n2797 0.0083125
R13199 VDPWR.n2877 VDPWR.n959 0.0083125
R13200 VDPWR.n2963 VDPWR.n2962 0.0083125
R13201 VDPWR.n2602 VDPWR.n2600 0.0083125
R13202 VDPWR.n3063 VDPWR.n3062 0.0083125
R13203 VDPWR.n3009 VDPWR.n921 0.0083125
R13204 VDPWR.n2429 VDPWR.n2428 0.0083125
R13205 VDPWR.n2468 VDPWR.n2466 0.0083125
R13206 VDPWR.n848 VDPWR.n827 0.0083125
R13207 VDPWR.n202 VDPWR.n201 0.00729348
R13208 VDPWR.n2598 VDPWR 0.00701042
R13209 VDPWR.n2427 VDPWR 0.00701042
R13210 VDPWR.n2464 VDPWR 0.00701042
R13211 VDPWR VDPWR.n151 0.00627446
R13212 VDPWR.n166 VDPWR 0.00627446
R13213 VDPWR.n161 VDPWR 0.00627446
R13214 VDPWR.n156 VDPWR 0.00627446
R13215 VDPWR VDPWR.n128 0.00627446
R13216 VDPWR.n195 VDPWR 0.00627446
R13217 VDPWR.n190 VDPWR 0.00627446
R13218 VDPWR.n185 VDPWR 0.00627446
R13219 VDPWR.n180 VDPWR 0.00627446
R13220 VDPWR VDPWR.n252 0.00626923
R13221 VDPWR.n138 VDPWR 0.00593478
R13222 VDPWR.n228 VDPWR.n203 0.00530769
R13223 VDPWR.n3073 VDPWR.n777 0.0052
R13224 VDPWR.n782 VDPWR.n781 0.0052
R13225 VDPWR.n2500 VDPWR.n2339 0.0052
R13226 VDPWR.n3113 VDPWR.n3112 0.0052
R13227 VDPWR.n2537 VDPWR.n2340 0.0052
R13228 VDPWR.n249 VDPWR 0.00458654
R13229 VDPWR VDPWR.n122 0.00458654
R13230 VDPWR.n241 VDPWR 0.00458654
R13231 VDPWR.n236 VDPWR 0.00458654
R13232 VDPWR.n231 VDPWR 0.00458654
R13233 VDPWR.n226 VDPWR 0.00458654
R13234 VDPWR.n221 VDPWR 0.00458654
R13235 VDPWR.n216 VDPWR 0.00458654
R13236 VDPWR.n211 VDPWR 0.00458654
R13237 VDPWR.n629 VDPWR.n628 0.00310417
R13238 VDPWR.n349 VDPWR.n348 0.00310417
R13239 VDPWR.n1388 VDPWR.n1387 0.00310417
R13240 VDPWR.n1460 VDPWR.n1315 0.00310417
R13241 VDPWR.n1495 VDPWR.n1298 0.00310417
R13242 VDPWR.n1583 VDPWR.n1289 0.00310417
R13243 VDPWR.n1550 VDPWR.n1536 0.00310417
R13244 VDPWR.n1718 VDPWR.n1717 0.00310417
R13245 VDPWR.n1251 VDPWR.n1242 0.00310417
R13246 VDPWR.n1823 VDPWR.n1225 0.00310417
R13247 VDPWR.n1853 VDPWR.n1214 0.00310417
R13248 VDPWR.n1899 VDPWR.n1198 0.00310417
R13249 VDPWR.n1657 VDPWR.n1656 0.00310417
R13250 VDPWR.n1144 VDPWR.n1140 0.00310417
R13251 VDPWR.n2003 VDPWR.n1165 0.00310417
R13252 VDPWR.n1912 VDPWR.n1911 0.00310417
R13253 VDPWR.n1949 VDPWR.n1935 0.00310417
R13254 VDPWR.n2128 VDPWR.n2127 0.00310417
R13255 VDPWR.n2241 VDPWR.n2197 0.00310417
R13256 VDPWR.n2319 VDPWR.n1020 0.00310417
R13257 VDPWR.n1053 VDPWR.n1042 0.00310417
R13258 VDPWR.n1085 VDPWR.n1084 0.00310417
R13259 VDPWR.n2759 VDPWR.n2758 0.00310417
R13260 VDPWR.n2849 VDPWR.n2848 0.00310417
R13261 VDPWR.n2899 VDPWR.n955 0.00310417
R13262 VDPWR.n2927 VDPWR.n2924 0.00310417
R13263 VDPWR.n2976 VDPWR.n928 0.00310417
R13264 VDPWR.n2716 VDPWR.n2715 0.00310417
R13265 VDPWR.n2655 VDPWR.n2654 0.00310417
R13266 VDPWR.n3055 VDPWR.n880 0.00310417
R13267 VDPWR.n910 VDPWR.n902 0.00310417
R13268 VDPWR.n2996 VDPWR.n2986 0.00310417
R13269 VDPWR.n2361 VDPWR.n2358 0.00310417
R13270 VDPWR.n2495 VDPWR.n2493 0.00310417
R13271 VDPWR.n3098 VDPWR.n788 0.00310417
R13272 VDPWR.n811 VDPWR.n810 0.00310417
R13273 VDPWR.n840 VDPWR.n835 0.00310417
R13274 VDPWR.n91 VDPWR.n90 0.00310417
R13275 VDPWR.n627 VDPWR.n626 0.00180208
R13276 VDPWR.n595 VDPWR 0.00180208
R13277 VDPWR.n561 VDPWR.n547 0.00180208
R13278 VDPWR.n347 VDPWR.n346 0.00180208
R13279 VDPWR.n315 VDPWR 0.00180208
R13280 VDPWR.n281 VDPWR.n267 0.00180208
R13281 VDPWR.n89 VDPWR.n88 0.00180208
R13282 VDPWR.n57 VDPWR 0.00180208
R13283 VDPWR.n23 VDPWR.n9 0.00180208
R13284 VDPWR.n728 VDPWR.n727 0.00177551
R13285 VDPWR.n257 VDPWR.n255 0.00105731
R13286 muxtest_0.x2.x2.GP1.n2 muxtest_0.x2.x2.GP1.t4 450.938
R13287 muxtest_0.x2.x2.GP1.n2 muxtest_0.x2.x2.GP1.t5 445.666
R13288 muxtest_0.x2.x2.GP1.n4 muxtest_0.x2.x2.GP1.n3 195.832
R13289 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n0 96.8352
R13290 muxtest_0.x2.x2.GP1.n3 muxtest_0.x2.x2.GP1.t3 26.5955
R13291 muxtest_0.x2.x2.GP1.n3 muxtest_0.x2.x2.GP1.t2 26.5955
R13292 muxtest_0.x2.x2.GP1.n0 muxtest_0.x2.x2.GP1.t1 24.9236
R13293 muxtest_0.x2.x2.GP1.n0 muxtest_0.x2.x2.GP1.t0 24.9236
R13294 muxtest_0.x2.x2.GP1.n5 muxtest_0.x2.x2.GP1.n4 13.1346
R13295 muxtest_0.x2.x2.GP1.n4 muxtest_0.x2.x2.GP1 12.2007
R13296 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n1 11.2645
R13297 muxtest_0.x2.x2.GP1.n1 muxtest_0.x2.x2.GP1 6.1445
R13298 muxtest_0.x2.x2.GP1.n1 muxtest_0.x2.x2.GP1 4.65505
R13299 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n2 3.07707
R13300 muxtest_0.x2.x2.GP1.n5 muxtest_0.x2.x2.GP1 2.0485
R13301 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n5 1.55202
R13302 ua[3].n10 ua[3].t4 26.3998
R13303 ua[3].n6 ua[3].t6 23.6581
R13304 ua[3].n1 ua[3].t3 23.6581
R13305 ua[3].n10 ua[3].t5 23.5483
R13306 ua[3].n8 ua[3].t8 23.3739
R13307 ua[3].n3 ua[3].t2 23.3739
R13308 ua[3].n11 ua[3].t10 12.9758
R13309 ua[3].n11 ua[3].t11 10.8618
R13310 ua[3].n6 ua[3].t1 10.7528
R13311 ua[3].n1 ua[3].t9 10.7528
R13312 ua[3].n5 ua[3].t0 10.6417
R13313 ua[3].n0 ua[3].t7 10.6417
R13314 ua[3].n15 ua[3] 4.48702
R13315 ua[3].n12 ua[3].n10 3.06895
R13316 ua[3].n12 ua[3].n11 2.14822
R13317 ua[3].n14 ua[3] 1.938
R13318 ua[3].n7 ua[3].n6 1.30064
R13319 ua[3].n2 ua[3].n1 1.30064
R13320 ua[3].n13 ua[3].n12 1.12636
R13321 ua[3] ua[3].n9 0.983856
R13322 ua[3] ua[3].n4 0.966624
R13323 ua[3].n8 ua[3].n7 0.726502
R13324 ua[3].n3 ua[3].n2 0.726502
R13325 ua[3].n17 ua[3].n16 0.683625
R13326 ua[3].n7 ua[3].n5 0.512491
R13327 ua[3].n2 ua[3].n0 0.512491
R13328 ua[3].n15 ua[3] 0.398
R13329 ua[3] ua[3].n15 0.398
R13330 ua[3].n16 ua[3] 0.37425
R13331 ua[3].n9 ua[3].n5 0.359663
R13332 ua[3].n4 ua[3].n0 0.359663
R13333 ua[3].n16 ua[3] 0.2705
R13334 ua[3].n9 ua[3].n8 0.216071
R13335 ua[3].n4 ua[3].n3 0.216071
R13336 ua[3].n14 ua[3].n13 0.148615
R13337 ua[3] ua[3].n14 0.146333
R13338 ua[3].n17 ua[3] 0.124875
R13339 ua[3].n13 ua[3] 0.0655
R13340 ua[3] ua[3].n17 0.063
R13341 ua[2].n6 ua[2].t2 23.6581
R13342 ua[2].n15 ua[2].t6 23.6581
R13343 ua[2].n22 ua[2].t4 23.6581
R13344 ua[2].n1 ua[2].t9 23.6581
R13345 ua[2].n5 ua[2].t3 23.3739
R13346 ua[2].n14 ua[2].t7 23.3739
R13347 ua[2].n21 ua[2].t5 23.3739
R13348 ua[2].n0 ua[2].t8 23.3739
R13349 ua[2].n28 ua[2] 21.5313
R13350 ua[2].n6 ua[2].t15 10.7528
R13351 ua[2].n15 ua[2].t1 10.7528
R13352 ua[2].n22 ua[2].t10 10.7528
R13353 ua[2].n1 ua[2].t12 10.7528
R13354 ua[2].n8 ua[2].t14 10.6417
R13355 ua[2].n17 ua[2].t0 10.6417
R13356 ua[2].n24 ua[2].t11 10.6417
R13357 ua[2].n3 ua[2].t13 10.6417
R13358 ua[2].n7 ua[2].n6 1.30064
R13359 ua[2].n16 ua[2].n15 1.30064
R13360 ua[2].n23 ua[2].n22 1.30064
R13361 ua[2].n2 ua[2].n1 1.30064
R13362 ua[2] ua[2].n4 0.983856
R13363 ua[2].n10 ua[2].n9 0.956356
R13364 ua[2].n26 ua[2].n25 0.946356
R13365 ua[2].n19 ua[2].n18 0.927606
R13366 ua[2].n7 ua[2].n5 0.726502
R13367 ua[2].n16 ua[2].n14 0.726502
R13368 ua[2].n23 ua[2].n21 0.726502
R13369 ua[2].n2 ua[2].n0 0.726502
R13370 ua[2].n11 ua[2] 0.681056
R13371 ua[2].n20 ua[2].n13 0.54925
R13372 ua[2].n27 ua[2].n20 0.54425
R13373 ua[2].n28 ua[2].n27 0.53675
R13374 ua[2].n8 ua[2].n7 0.512491
R13375 ua[2].n17 ua[2].n16 0.512491
R13376 ua[2].n24 ua[2].n23 0.512491
R13377 ua[2].n3 ua[2].n2 0.512491
R13378 ua[2].n9 ua[2].n8 0.359663
R13379 ua[2].n18 ua[2].n17 0.359663
R13380 ua[2].n25 ua[2].n24 0.359663
R13381 ua[2].n4 ua[2].n3 0.359663
R13382 ua[2].n9 ua[2].n5 0.216071
R13383 ua[2].n18 ua[2].n14 0.216071
R13384 ua[2].n25 ua[2].n21 0.216071
R13385 ua[2].n4 ua[2].n0 0.216071
R13386 ua[2].n20 ua[2] 0.18675
R13387 ua[2].n13 ua[2] 0.18425
R13388 ua[2].n27 ua[2] 0.16425
R13389 ua[2] ua[2].n28 0.163
R13390 ua[2].n12 ua[2] 0.135115
R13391 ua[2].n19 ua[2] 0.05675
R13392 ua[2] ua[2].n19 0.0561931
R13393 ua[2].n12 ua[2].n11 0.0530774
R13394 ua[2].n26 ua[2] 0.038
R13395 ua[2] ua[2].n26 0.0376287
R13396 ua[2].n10 ua[2] 0.028
R13397 ua[2] ua[2].n10 0.0266905
R13398 ua[2].n11 ua[2] 0.01175
R13399 ua[2].n13 ua[2].n12 0.006125
R13400 ringtest_0.x4.clknet_0_clk.n33 ringtest_0.x4.clknet_0_clk.n31 333.392
R13401 ringtest_0.x4.clknet_0_clk.n38 ringtest_0.x4.clknet_0_clk.n26 301.392
R13402 ringtest_0.x4.clknet_0_clk.n37 ringtest_0.x4.clknet_0_clk.n27 301.392
R13403 ringtest_0.x4.clknet_0_clk.n36 ringtest_0.x4.clknet_0_clk.n28 301.392
R13404 ringtest_0.x4.clknet_0_clk.n35 ringtest_0.x4.clknet_0_clk.n29 301.392
R13405 ringtest_0.x4.clknet_0_clk.n34 ringtest_0.x4.clknet_0_clk.n30 301.392
R13406 ringtest_0.x4.clknet_0_clk.n33 ringtest_0.x4.clknet_0_clk.n32 301.392
R13407 ringtest_0.x4.clknet_0_clk.n39 ringtest_0.x4.clknet_0_clk.n25 297.863
R13408 ringtest_0.x4.clknet_0_clk.n2 ringtest_0.x4.clknet_0_clk.n0 248.638
R13409 ringtest_0.x4.clknet_0_clk.n2 ringtest_0.x4.clknet_0_clk.n1 203.463
R13410 ringtest_0.x4.clknet_0_clk.n4 ringtest_0.x4.clknet_0_clk.n3 203.463
R13411 ringtest_0.x4.clknet_0_clk.n8 ringtest_0.x4.clknet_0_clk.n7 203.463
R13412 ringtest_0.x4.clknet_0_clk.n24 ringtest_0.x4.clknet_0_clk.n23 203.463
R13413 ringtest_0.x4.clknet_0_clk.n6 ringtest_0.x4.clknet_0_clk.n5 202.456
R13414 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n41 199.607
R13415 ringtest_0.x4.clknet_0_clk.n21 ringtest_0.x4.clknet_0_clk.n9 188.201
R13416 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.t46 184.768
R13417 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.t43 184.768
R13418 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.t42 184.768
R13419 ringtest_0.x4.clknet_0_clk.n15 ringtest_0.x4.clknet_0_clk.t45 184.768
R13420 ringtest_0.x4.clknet_0_clk.n10 ringtest_0.x4.clknet_0_clk.t41 184.768
R13421 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.t37 184.768
R13422 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.t40 184.768
R13423 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.t39 184.768
R13424 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n18 173.609
R13425 ringtest_0.x4.clknet_0_clk.n14 ringtest_0.x4.clknet_0_clk.n13 171.375
R13426 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.t38 146.208
R13427 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.t35 146.208
R13428 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.t34 146.208
R13429 ringtest_0.x4.clknet_0_clk.n15 ringtest_0.x4.clknet_0_clk.t36 146.208
R13430 ringtest_0.x4.clknet_0_clk.n10 ringtest_0.x4.clknet_0_clk.t33 146.208
R13431 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.t44 146.208
R13432 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.t32 146.208
R13433 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.t47 146.208
R13434 ringtest_0.x4.clknet_0_clk.n4 ringtest_0.x4.clknet_0_clk.n2 45.177
R13435 ringtest_0.x4.clknet_0_clk.n22 ringtest_0.x4.clknet_0_clk.n8 45.177
R13436 ringtest_0.x4.clknet_0_clk.n24 ringtest_0.x4.clknet_0_clk.n22 45.177
R13437 ringtest_0.x4.clknet_0_clk.n6 ringtest_0.x4.clknet_0_clk.n4 44.0476
R13438 ringtest_0.x4.clknet_0_clk.n8 ringtest_0.x4.clknet_0_clk.n6 44.0476
R13439 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.n17 40.6397
R13440 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.n16 40.6397
R13441 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.n15 40.6397
R13442 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.n10 40.6397
R13443 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.n11 40.6397
R13444 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.n12 40.6397
R13445 ringtest_0.x4.clknet_0_clk.n0 ringtest_0.x4.clknet_0_clk.t2 40.0005
R13446 ringtest_0.x4.clknet_0_clk.n0 ringtest_0.x4.clknet_0_clk.t15 40.0005
R13447 ringtest_0.x4.clknet_0_clk.n1 ringtest_0.x4.clknet_0_clk.t4 40.0005
R13448 ringtest_0.x4.clknet_0_clk.n1 ringtest_0.x4.clknet_0_clk.t6 40.0005
R13449 ringtest_0.x4.clknet_0_clk.n3 ringtest_0.x4.clknet_0_clk.t8 40.0005
R13450 ringtest_0.x4.clknet_0_clk.n3 ringtest_0.x4.clknet_0_clk.t10 40.0005
R13451 ringtest_0.x4.clknet_0_clk.n5 ringtest_0.x4.clknet_0_clk.t5 40.0005
R13452 ringtest_0.x4.clknet_0_clk.n5 ringtest_0.x4.clknet_0_clk.t7 40.0005
R13453 ringtest_0.x4.clknet_0_clk.n7 ringtest_0.x4.clknet_0_clk.t9 40.0005
R13454 ringtest_0.x4.clknet_0_clk.n7 ringtest_0.x4.clknet_0_clk.t11 40.0005
R13455 ringtest_0.x4.clknet_0_clk.n9 ringtest_0.x4.clknet_0_clk.t0 40.0005
R13456 ringtest_0.x4.clknet_0_clk.n9 ringtest_0.x4.clknet_0_clk.t13 40.0005
R13457 ringtest_0.x4.clknet_0_clk.n23 ringtest_0.x4.clknet_0_clk.t14 40.0005
R13458 ringtest_0.x4.clknet_0_clk.n23 ringtest_0.x4.clknet_0_clk.t12 40.0005
R13459 ringtest_0.x4.clknet_0_clk.n41 ringtest_0.x4.clknet_0_clk.t1 40.0005
R13460 ringtest_0.x4.clknet_0_clk.n41 ringtest_0.x4.clknet_0_clk.t3 40.0005
R13461 ringtest_0.x4.clknet_0_clk.n38 ringtest_0.x4.clknet_0_clk.n37 32.0005
R13462 ringtest_0.x4.clknet_0_clk.n37 ringtest_0.x4.clknet_0_clk.n36 32.0005
R13463 ringtest_0.x4.clknet_0_clk.n35 ringtest_0.x4.clknet_0_clk.n34 32.0005
R13464 ringtest_0.x4.clknet_0_clk.n34 ringtest_0.x4.clknet_0_clk.n33 32.0005
R13465 ringtest_0.x4.clknet_0_clk.n36 ringtest_0.x4.clknet_0_clk.n35 31.2005
R13466 ringtest_0.x4.clknet_0_clk.n31 ringtest_0.x4.clknet_0_clk.t27 27.5805
R13467 ringtest_0.x4.clknet_0_clk.n31 ringtest_0.x4.clknet_0_clk.t24 27.5805
R13468 ringtest_0.x4.clknet_0_clk.n26 ringtest_0.x4.clknet_0_clk.t23 27.5805
R13469 ringtest_0.x4.clknet_0_clk.n26 ringtest_0.x4.clknet_0_clk.t21 27.5805
R13470 ringtest_0.x4.clknet_0_clk.n25 ringtest_0.x4.clknet_0_clk.t26 27.5805
R13471 ringtest_0.x4.clknet_0_clk.n25 ringtest_0.x4.clknet_0_clk.t28 27.5805
R13472 ringtest_0.x4.clknet_0_clk.n27 ringtest_0.x4.clknet_0_clk.t25 27.5805
R13473 ringtest_0.x4.clknet_0_clk.n27 ringtest_0.x4.clknet_0_clk.t22 27.5805
R13474 ringtest_0.x4.clknet_0_clk.n28 ringtest_0.x4.clknet_0_clk.t18 27.5805
R13475 ringtest_0.x4.clknet_0_clk.n28 ringtest_0.x4.clknet_0_clk.t20 27.5805
R13476 ringtest_0.x4.clknet_0_clk.n29 ringtest_0.x4.clknet_0_clk.t30 27.5805
R13477 ringtest_0.x4.clknet_0_clk.n29 ringtest_0.x4.clknet_0_clk.t16 27.5805
R13478 ringtest_0.x4.clknet_0_clk.n30 ringtest_0.x4.clknet_0_clk.t17 27.5805
R13479 ringtest_0.x4.clknet_0_clk.n30 ringtest_0.x4.clknet_0_clk.t19 27.5805
R13480 ringtest_0.x4.clknet_0_clk.n32 ringtest_0.x4.clknet_0_clk.t29 27.5805
R13481 ringtest_0.x4.clknet_0_clk.n32 ringtest_0.x4.clknet_0_clk.t31 27.5805
R13482 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n14 25.9814
R13483 ringtest_0.x4.clknet_0_clk.n22 ringtest_0.x4.clknet_0_clk.n21 15.262
R13484 ringtest_0.x4.clknet_0_clk.n20 ringtest_0.x4.clknet_0_clk.n19 14.7771
R13485 ringtest_0.x4.clknet_0_clk.n40 ringtest_0.x4.clknet_0_clk.n24 13.177
R13486 ringtest_0.x4.clknet_0_clk.n39 ringtest_0.x4.clknet_0_clk.n38 10.4484
R13487 ringtest_0.x4.clknet_0_clk.n19 ringtest_0.x4.clknet_0_clk 10.3624
R13488 ringtest_0.x4.clknet_0_clk.n21 ringtest_0.x4.clknet_0_clk.n20 9.3005
R13489 ringtest_0.x4.clknet_0_clk.n19 ringtest_0.x4.clknet_0_clk 3.45447
R13490 ringtest_0.x4.clknet_0_clk.n40 ringtest_0.x4.clknet_0_clk 3.13183
R13491 ringtest_0.x4.clknet_0_clk.n14 ringtest_0.x4.clknet_0_clk 2.23542
R13492 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n39 1.75844
R13493 ringtest_0.x4.clknet_0_clk.n20 ringtest_0.x4.clknet_0_clk 1.5927
R13494 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n40 0.604792
R13495 ringtest_0.x4.net6.n3 ringtest_0.x4.net6.t13 323.342
R13496 ringtest_0.x4.net6.n0 ringtest_0.x4.net6.t4 323.342
R13497 ringtest_0.x4.net6.n1 ringtest_0.x4.net6.t2 260.322
R13498 ringtest_0.x4.net6.n8 ringtest_0.x4.net6.t5 241.536
R13499 ringtest_0.x4.net6.n17 ringtest_0.x4.net6.t1 222.679
R13500 ringtest_0.x4.net6.n12 ringtest_0.x4.net6.t14 212.081
R13501 ringtest_0.x4.net6.n13 ringtest_0.x4.net6.t7 212.081
R13502 ringtest_0.x4.net6.n3 ringtest_0.x4.net6.t6 194.809
R13503 ringtest_0.x4.net6.n0 ringtest_0.x4.net6.t8 194.809
R13504 ringtest_0.x4.net6.n5 ringtest_0.x4.net6.t10 183.505
R13505 ringtest_0.x4.net6.n1 ringtest_0.x4.net6.t12 175.169
R13506 ringtest_0.x4.net6.n8 ringtest_0.x4.net6.t11 169.237
R13507 ringtest_0.x4.net6 ringtest_0.x4.net6.n3 158.133
R13508 ringtest_0.x4.net6 ringtest_0.x4.net6.n0 158.133
R13509 ringtest_0.x4.net6 ringtest_0.x4.net6.n8 157.555
R13510 ringtest_0.x4.net6.n15 ringtest_0.x4.net6.n14 155.52
R13511 ringtest_0.x4.net6.n6 ringtest_0.x4.net6.n5 153.863
R13512 ringtest_0.x4.net6.n2 ringtest_0.x4.net6.n1 152
R13513 ringtest_0.x4.net6.n12 ringtest_0.x4.net6.t9 139.78
R13514 ringtest_0.x4.net6.n13 ringtest_0.x4.net6.t15 139.78
R13515 ringtest_0.x4.net6.n18 ringtest_0.x4.net6.t0 129.078
R13516 ringtest_0.x4.net6.n5 ringtest_0.x4.net6.t3 114.532
R13517 ringtest_0.x4.net6.n18 ringtest_0.x4.net6.n17 96.7191
R13518 ringtest_0.x4.net6.n11 ringtest_0.x4.net6 55.2785
R13519 ringtest_0.x4.net6.n14 ringtest_0.x4.net6.n13 37.246
R13520 ringtest_0.x4.net6.n14 ringtest_0.x4.net6.n12 24.1005
R13521 ringtest_0.x4.net6.n10 ringtest_0.x4.net6.n9 21.4124
R13522 ringtest_0.x4.net6.n16 ringtest_0.x4.net6.n15 21.1949
R13523 ringtest_0.x4.net6.n4 ringtest_0.x4.net6.n2 20.043
R13524 ringtest_0.x4.net6.n7 ringtest_0.x4.net6.n6 15.2615
R13525 ringtest_0.x4.net6.n17 ringtest_0.x4.net6.n16 12.4213
R13526 ringtest_0.x4.net6.n9 ringtest_0.x4.net6 12.3175
R13527 ringtest_0.x4.net6.n16 ringtest_0.x4.net6.n11 8.09819
R13528 ringtest_0.x4.net6.n11 ringtest_0.x4.net6.n10 7.53948
R13529 ringtest_0.x4.net6.n4 ringtest_0.x4.net6 7.39885
R13530 ringtest_0.x4.net6 ringtest_0.x4.net6.n18 5.84085
R13531 ringtest_0.x4.net6.n15 ringtest_0.x4.net6 5.4405
R13532 ringtest_0.x4.net6.n9 ringtest_0.x4.net6 4.10616
R13533 ringtest_0.x4.net6.n7 ringtest_0.x4.net6.n4 2.60421
R13534 ringtest_0.x4.net6.n10 ringtest_0.x4.net6.n7 2.43577
R13535 ringtest_0.x4.net6.n6 ringtest_0.x4.net6 1.97868
R13536 ringtest_0.x4.net6.n2 ringtest_0.x4.net6 1.55726
R13537 ringtest_0.x4.clknet_1_1__leaf_clk.n29 ringtest_0.x4.clknet_1_1__leaf_clk.n27 333.392
R13538 ringtest_0.x4.clknet_1_1__leaf_clk.n29 ringtest_0.x4.clknet_1_1__leaf_clk.n28 301.392
R13539 ringtest_0.x4.clknet_1_1__leaf_clk.n31 ringtest_0.x4.clknet_1_1__leaf_clk.n30 301.392
R13540 ringtest_0.x4.clknet_1_1__leaf_clk.n33 ringtest_0.x4.clknet_1_1__leaf_clk.n32 301.392
R13541 ringtest_0.x4.clknet_1_1__leaf_clk.n35 ringtest_0.x4.clknet_1_1__leaf_clk.n34 301.392
R13542 ringtest_0.x4.clknet_1_1__leaf_clk.n37 ringtest_0.x4.clknet_1_1__leaf_clk.n36 301.392
R13543 ringtest_0.x4.clknet_1_1__leaf_clk.n39 ringtest_0.x4.clknet_1_1__leaf_clk.n38 301.392
R13544 ringtest_0.x4.clknet_1_1__leaf_clk.n40 ringtest_0.x4.clknet_1_1__leaf_clk.n26 297.863
R13545 ringtest_0.x4.clknet_1_1__leaf_clk.n18 ringtest_0.x4.clknet_1_1__leaf_clk.t36 294.557
R13546 ringtest_0.x4.clknet_1_1__leaf_clk.n15 ringtest_0.x4.clknet_1_1__leaf_clk.t33 294.557
R13547 ringtest_0.x4.clknet_1_1__leaf_clk.n13 ringtest_0.x4.clknet_1_1__leaf_clk.t34 294.557
R13548 ringtest_0.x4.clknet_1_1__leaf_clk.n11 ringtest_0.x4.clknet_1_1__leaf_clk.t41 294.557
R13549 ringtest_0.x4.clknet_1_1__leaf_clk.n10 ringtest_0.x4.clknet_1_1__leaf_clk.t32 294.557
R13550 ringtest_0.x4.clknet_1_1__leaf_clk.n2 ringtest_0.x4.clknet_1_1__leaf_clk.n0 248.638
R13551 ringtest_0.x4.clknet_1_1__leaf_clk.n18 ringtest_0.x4.clknet_1_1__leaf_clk.t39 211.01
R13552 ringtest_0.x4.clknet_1_1__leaf_clk.n15 ringtest_0.x4.clknet_1_1__leaf_clk.t40 211.01
R13553 ringtest_0.x4.clknet_1_1__leaf_clk.n13 ringtest_0.x4.clknet_1_1__leaf_clk.t38 211.01
R13554 ringtest_0.x4.clknet_1_1__leaf_clk.n11 ringtest_0.x4.clknet_1_1__leaf_clk.t35 211.01
R13555 ringtest_0.x4.clknet_1_1__leaf_clk.n10 ringtest_0.x4.clknet_1_1__leaf_clk.t37 211.01
R13556 ringtest_0.x4.clknet_1_1__leaf_clk.n2 ringtest_0.x4.clknet_1_1__leaf_clk.n1 203.463
R13557 ringtest_0.x4.clknet_1_1__leaf_clk.n4 ringtest_0.x4.clknet_1_1__leaf_clk.n3 203.463
R13558 ringtest_0.x4.clknet_1_1__leaf_clk.n8 ringtest_0.x4.clknet_1_1__leaf_clk.n7 203.463
R13559 ringtest_0.x4.clknet_1_1__leaf_clk.n25 ringtest_0.x4.clknet_1_1__leaf_clk.n24 203.463
R13560 ringtest_0.x4.clknet_1_1__leaf_clk.n6 ringtest_0.x4.clknet_1_1__leaf_clk.n5 202.456
R13561 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n42 199.607
R13562 ringtest_0.x4.clknet_1_1__leaf_clk.n22 ringtest_0.x4.clknet_1_1__leaf_clk.n9 188.201
R13563 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n13 156.207
R13564 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n10 156.207
R13565 ringtest_0.x4.clknet_1_1__leaf_clk.n19 ringtest_0.x4.clknet_1_1__leaf_clk.n18 153.097
R13566 ringtest_0.x4.clknet_1_1__leaf_clk.n16 ringtest_0.x4.clknet_1_1__leaf_clk.n15 152.296
R13567 ringtest_0.x4.clknet_1_1__leaf_clk.n12 ringtest_0.x4.clknet_1_1__leaf_clk.n11 152.296
R13568 ringtest_0.x4.clknet_1_1__leaf_clk.n4 ringtest_0.x4.clknet_1_1__leaf_clk.n2 45.177
R13569 ringtest_0.x4.clknet_1_1__leaf_clk.n23 ringtest_0.x4.clknet_1_1__leaf_clk.n8 45.177
R13570 ringtest_0.x4.clknet_1_1__leaf_clk.n25 ringtest_0.x4.clknet_1_1__leaf_clk.n23 45.177
R13571 ringtest_0.x4.clknet_1_1__leaf_clk.n6 ringtest_0.x4.clknet_1_1__leaf_clk.n4 44.0476
R13572 ringtest_0.x4.clknet_1_1__leaf_clk.n8 ringtest_0.x4.clknet_1_1__leaf_clk.n6 44.0476
R13573 ringtest_0.x4.clknet_1_1__leaf_clk.n0 ringtest_0.x4.clknet_1_1__leaf_clk.t13 40.0005
R13574 ringtest_0.x4.clknet_1_1__leaf_clk.n0 ringtest_0.x4.clknet_1_1__leaf_clk.t14 40.0005
R13575 ringtest_0.x4.clknet_1_1__leaf_clk.n1 ringtest_0.x4.clknet_1_1__leaf_clk.t15 40.0005
R13576 ringtest_0.x4.clknet_1_1__leaf_clk.n1 ringtest_0.x4.clknet_1_1__leaf_clk.t12 40.0005
R13577 ringtest_0.x4.clknet_1_1__leaf_clk.n3 ringtest_0.x4.clknet_1_1__leaf_clk.t11 40.0005
R13578 ringtest_0.x4.clknet_1_1__leaf_clk.n3 ringtest_0.x4.clknet_1_1__leaf_clk.t10 40.0005
R13579 ringtest_0.x4.clknet_1_1__leaf_clk.n5 ringtest_0.x4.clknet_1_1__leaf_clk.t6 40.0005
R13580 ringtest_0.x4.clknet_1_1__leaf_clk.n5 ringtest_0.x4.clknet_1_1__leaf_clk.t8 40.0005
R13581 ringtest_0.x4.clknet_1_1__leaf_clk.n7 ringtest_0.x4.clknet_1_1__leaf_clk.t2 40.0005
R13582 ringtest_0.x4.clknet_1_1__leaf_clk.n7 ringtest_0.x4.clknet_1_1__leaf_clk.t4 40.0005
R13583 ringtest_0.x4.clknet_1_1__leaf_clk.n9 ringtest_0.x4.clknet_1_1__leaf_clk.t5 40.0005
R13584 ringtest_0.x4.clknet_1_1__leaf_clk.n9 ringtest_0.x4.clknet_1_1__leaf_clk.t7 40.0005
R13585 ringtest_0.x4.clknet_1_1__leaf_clk.n24 ringtest_0.x4.clknet_1_1__leaf_clk.t1 40.0005
R13586 ringtest_0.x4.clknet_1_1__leaf_clk.n24 ringtest_0.x4.clknet_1_1__leaf_clk.t9 40.0005
R13587 ringtest_0.x4.clknet_1_1__leaf_clk.n42 ringtest_0.x4.clknet_1_1__leaf_clk.t3 40.0005
R13588 ringtest_0.x4.clknet_1_1__leaf_clk.n42 ringtest_0.x4.clknet_1_1__leaf_clk.t0 40.0005
R13589 ringtest_0.x4.clknet_1_1__leaf_clk.n21 ringtest_0.x4.clknet_1_1__leaf_clk 34.5053
R13590 ringtest_0.x4.clknet_1_1__leaf_clk.n14 ringtest_0.x4.clknet_1_1__leaf_clk 33.8485
R13591 ringtest_0.x4.clknet_1_1__leaf_clk.n31 ringtest_0.x4.clknet_1_1__leaf_clk.n29 32.0005
R13592 ringtest_0.x4.clknet_1_1__leaf_clk.n33 ringtest_0.x4.clknet_1_1__leaf_clk.n31 32.0005
R13593 ringtest_0.x4.clknet_1_1__leaf_clk.n37 ringtest_0.x4.clknet_1_1__leaf_clk.n35 32.0005
R13594 ringtest_0.x4.clknet_1_1__leaf_clk.n39 ringtest_0.x4.clknet_1_1__leaf_clk.n37 32.0005
R13595 ringtest_0.x4.clknet_1_1__leaf_clk.n35 ringtest_0.x4.clknet_1_1__leaf_clk.n33 31.2005
R13596 ringtest_0.x4.clknet_1_1__leaf_clk.n27 ringtest_0.x4.clknet_1_1__leaf_clk.t19 27.5805
R13597 ringtest_0.x4.clknet_1_1__leaf_clk.n27 ringtest_0.x4.clknet_1_1__leaf_clk.t20 27.5805
R13598 ringtest_0.x4.clknet_1_1__leaf_clk.n28 ringtest_0.x4.clknet_1_1__leaf_clk.t21 27.5805
R13599 ringtest_0.x4.clknet_1_1__leaf_clk.n28 ringtest_0.x4.clknet_1_1__leaf_clk.t18 27.5805
R13600 ringtest_0.x4.clknet_1_1__leaf_clk.n30 ringtest_0.x4.clknet_1_1__leaf_clk.t17 27.5805
R13601 ringtest_0.x4.clknet_1_1__leaf_clk.n30 ringtest_0.x4.clknet_1_1__leaf_clk.t16 27.5805
R13602 ringtest_0.x4.clknet_1_1__leaf_clk.n32 ringtest_0.x4.clknet_1_1__leaf_clk.t28 27.5805
R13603 ringtest_0.x4.clknet_1_1__leaf_clk.n32 ringtest_0.x4.clknet_1_1__leaf_clk.t30 27.5805
R13604 ringtest_0.x4.clknet_1_1__leaf_clk.n34 ringtest_0.x4.clknet_1_1__leaf_clk.t24 27.5805
R13605 ringtest_0.x4.clknet_1_1__leaf_clk.n34 ringtest_0.x4.clknet_1_1__leaf_clk.t26 27.5805
R13606 ringtest_0.x4.clknet_1_1__leaf_clk.n36 ringtest_0.x4.clknet_1_1__leaf_clk.t27 27.5805
R13607 ringtest_0.x4.clknet_1_1__leaf_clk.n36 ringtest_0.x4.clknet_1_1__leaf_clk.t29 27.5805
R13608 ringtest_0.x4.clknet_1_1__leaf_clk.n26 ringtest_0.x4.clknet_1_1__leaf_clk.t25 27.5805
R13609 ringtest_0.x4.clknet_1_1__leaf_clk.n26 ringtest_0.x4.clknet_1_1__leaf_clk.t22 27.5805
R13610 ringtest_0.x4.clknet_1_1__leaf_clk.n38 ringtest_0.x4.clknet_1_1__leaf_clk.t23 27.5805
R13611 ringtest_0.x4.clknet_1_1__leaf_clk.n38 ringtest_0.x4.clknet_1_1__leaf_clk.t31 27.5805
R13612 ringtest_0.x4.clknet_1_1__leaf_clk.n23 ringtest_0.x4.clknet_1_1__leaf_clk.n22 15.262
R13613 ringtest_0.x4.clknet_1_1__leaf_clk.n20 ringtest_0.x4.clknet_1_1__leaf_clk.n19 13.8005
R13614 ringtest_0.x4.clknet_1_1__leaf_clk.n41 ringtest_0.x4.clknet_1_1__leaf_clk.n25 13.177
R13615 ringtest_0.x4.clknet_1_1__leaf_clk.n14 ringtest_0.x4.clknet_1_1__leaf_clk.n12 11.6482
R13616 ringtest_0.x4.clknet_1_1__leaf_clk.n22 ringtest_0.x4.clknet_1_1__leaf_clk.n21 10.8268
R13617 ringtest_0.x4.clknet_1_1__leaf_clk.n40 ringtest_0.x4.clknet_1_1__leaf_clk.n39 10.4484
R13618 ringtest_0.x4.clknet_1_1__leaf_clk.n17 ringtest_0.x4.clknet_1_1__leaf_clk.n16 9.3005
R13619 ringtest_0.x4.clknet_1_1__leaf_clk.n20 ringtest_0.x4.clknet_1_1__leaf_clk.n17 8.37704
R13620 ringtest_0.x4.clknet_1_1__leaf_clk.n21 ringtest_0.x4.clknet_1_1__leaf_clk 5.19349
R13621 ringtest_0.x4.clknet_1_1__leaf_clk.n17 ringtest_0.x4.clknet_1_1__leaf_clk.n14 3.99105
R13622 ringtest_0.x4.clknet_1_1__leaf_clk.n41 ringtest_0.x4.clknet_1_1__leaf_clk 3.13183
R13623 ringtest_0.x4.clknet_1_1__leaf_clk.n19 ringtest_0.x4.clknet_1_1__leaf_clk 3.10907
R13624 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n40 1.75844
R13625 ringtest_0.x4.clknet_1_1__leaf_clk.n16 ringtest_0.x4.clknet_1_1__leaf_clk 1.67435
R13626 ringtest_0.x4.clknet_1_1__leaf_clk.n12 ringtest_0.x4.clknet_1_1__leaf_clk 1.67435
R13627 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n20 0.693495
R13628 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n41 0.604792
R13629 ui_in[1].n10 ui_in[1].t8 327.99
R13630 ui_in[1].n3 ui_in[1].t1 293.969
R13631 ui_in[1].n6 ui_in[1].t7 256.07
R13632 ui_in[1].n0 ui_in[1].t0 212.081
R13633 ui_in[1].n1 ui_in[1].t2 212.081
R13634 ui_in[1].n10 ui_in[1].t9 199.457
R13635 ui_in[1].n2 ui_in[1].n1 182.929
R13636 ui_in[1] ui_in[1].n3 154.065
R13637 ui_in[1].n11 ui_in[1].n10 152
R13638 ui_in[1].n7 ui_in[1].n6 152
R13639 ui_in[1].n6 ui_in[1].t3 150.03
R13640 ui_in[1].n0 ui_in[1].t5 139.78
R13641 ui_in[1].n1 ui_in[1].t6 139.78
R13642 ui_in[1].n3 ui_in[1].t4 138.338
R13643 ui_in[1].n1 ui_in[1].n0 61.346
R13644 ui_in[1].n16 ui_in[1] 30.7401
R13645 ui_in[1].n5 ui_in[1] 17.455
R13646 ui_in[1].n14 ui_in[1].n13 14.6836
R13647 ui_in[1].n13 ui_in[1].n12 14.6704
R13648 ui_in[1].n4 ui_in[1] 13.8328
R13649 ui_in[1].n14 ui_in[1].n2 10.6811
R13650 ui_in[1].n7 ui_in[1].n5 10.4374
R13651 ui_in[1].n9 ui_in[1].n8 8.15776
R13652 ui_in[1].n12 ui_in[1] 6.61383
R13653 ui_in[1].n2 ui_in[1] 6.1445
R13654 ui_in[1].n4 ui_in[1] 5.16179
R13655 ui_in[1].n11 ui_in[1] 4.90717
R13656 ui_in[1].n9 ui_in[1].n4 4.65206
R13657 ui_in[1].n15 ui_in[1] 4.54217
R13658 ui_in[1].n8 ui_in[1] 3.93896
R13659 ui_in[1].n12 ui_in[1].n11 2.98717
R13660 ui_in[1].n5 ui_in[1] 2.16665
R13661 ui_in[1].n8 ui_in[1].n7 1.57588
R13662 ui_in[1].n13 ui_in[1].n9 0.79438
R13663 ui_in[1].n15 ui_in[1] 0.606561
R13664 ui_in[1] ui_in[1].n14 0.248606
R13665 ui_in[1] ui_in[1].n15 0.222091
R13666 ui_in[1] ui_in[1].n16 0.122375
R13667 ui_in[1].n16 ui_in[1] 0.121168
R13668 muxtest_0.x1.x3.GP1.n3 muxtest_0.x1.x3.GP1.t4 450.938
R13669 muxtest_0.x1.x3.GP1.n2 muxtest_0.x1.x3.GP1.t6 450.938
R13670 muxtest_0.x1.x3.GP1.n3 muxtest_0.x1.x3.GP1.t5 445.666
R13671 muxtest_0.x1.x3.GP1.n2 muxtest_0.x1.x3.GP1.t7 445.666
R13672 muxtest_0.x1.x3.GP1.n6 muxtest_0.x1.x3.GP1.n5 195.832
R13673 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n0 96.8352
R13674 muxtest_0.x1.x3.GP1.n5 muxtest_0.x1.x3.GP1.t2 26.5955
R13675 muxtest_0.x1.x3.GP1.n5 muxtest_0.x1.x3.GP1.t3 26.5955
R13676 muxtest_0.x1.x3.GP1.n0 muxtest_0.x1.x3.GP1.t1 24.9236
R13677 muxtest_0.x1.x3.GP1.n0 muxtest_0.x1.x3.GP1.t0 24.9236
R13678 muxtest_0.x1.x3.GP1.n4 muxtest_0.x1.x3.GP1 13.257
R13679 muxtest_0.x1.x3.GP1.n7 muxtest_0.x1.x3.GP1.n6 13.1346
R13680 muxtest_0.x1.x3.GP1.n6 muxtest_0.x1.x3.GP1 11.8965
R13681 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n1 11.2645
R13682 muxtest_0.x1.x3.GP1.n1 muxtest_0.x1.x3.GP1 6.1445
R13683 muxtest_0.x1.x3.GP1.n4 muxtest_0.x1.x3.GP1 5.31412
R13684 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n4 5.26828
R13685 muxtest_0.x1.x3.GP1.n1 muxtest_0.x1.x3.GP1 4.65505
R13686 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n2 3.07895
R13687 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n3 2.90754
R13688 muxtest_0.x1.x3.GP1.n7 muxtest_0.x1.x3.GP1 2.0485
R13689 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n7 1.55202
R13690 muxtest_0.x1.x3.GP4.n3 muxtest_0.x1.x3.GP4.t5 450.938
R13691 muxtest_0.x1.x3.GP4.n2 muxtest_0.x1.x3.GP4.t7 450.938
R13692 muxtest_0.x1.x3.GP4.n3 muxtest_0.x1.x3.GP4.t4 445.666
R13693 muxtest_0.x1.x3.GP4.n2 muxtest_0.x1.x3.GP4.t6 445.666
R13694 muxtest_0.x1.x3.GP4.n7 muxtest_0.x1.x3.GP4.n6 208.965
R13695 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n0 96.8352
R13696 muxtest_0.x1.x3.GP4.n6 muxtest_0.x1.x3.GP4.t2 26.5955
R13697 muxtest_0.x1.x3.GP4.n6 muxtest_0.x1.x3.GP4.t3 26.5955
R13698 muxtest_0.x1.x3.GP4.n0 muxtest_0.x1.x3.GP4.t1 24.9236
R13699 muxtest_0.x1.x3.GP4.n0 muxtest_0.x1.x3.GP4.t0 24.9236
R13700 muxtest_0.x1.x3.GP4.n4 muxtest_0.x1.x3.x4.GP 10.9863
R13701 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n5 10.2405
R13702 muxtest_0.x1.x1.gpo3 muxtest_0.x1.x3.GP4.n4 9.34192
R13703 muxtest_0.x1.x3.GP4.n5 muxtest_0.x1.x1.gpo3 7.73829
R13704 muxtest_0.x1.x3.GP4.n1 muxtest_0.x1.x1.x14.Y 6.1445
R13705 muxtest_0.x1.x3.GP4.n4 muxtest_0.x1.x2.x4.GP 5.84951
R13706 muxtest_0.x1.x3.GP4.n1 muxtest_0.x1.x1.x14.Y 4.65505
R13707 muxtest_0.x1.x2.x4.GP muxtest_0.x1.x3.GP4.n3 2.95993
R13708 muxtest_0.x1.x3.x4.GP muxtest_0.x1.x3.GP4.n2 2.95993
R13709 muxtest_0.x1.x3.GP4.n7 muxtest_0.x1.x1.x14.Y 2.0485
R13710 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n7 1.55202
R13711 muxtest_0.x1.x3.GP4.n5 muxtest_0.x1.x3.GP4.n1 1.0245
R13712 ringtest_0.x4._11_ ringtest_0.x4._11_.n0 623.909
R13713 ringtest_0.x4._11_.n24 ringtest_0.x4._11_.t6 334.723
R13714 ringtest_0.x4._11_.n5 ringtest_0.x4._11_.t5 334.723
R13715 ringtest_0.x4._11_.n18 ringtest_0.x4._11_.t19 261.887
R13716 ringtest_0.x4._11_.n14 ringtest_0.x4._11_.t14 256.07
R13717 ringtest_0.x4._11_.n8 ringtest_0.x4._11_.t10 241.536
R13718 ringtest_0.x4._11_.n3 ringtest_0.x4._11_.t13 241.536
R13719 ringtest_0.x4._11_.n1 ringtest_0.x4._11_.t12 231.835
R13720 ringtest_0.x4._11_.n21 ringtest_0.x4._11_.t8 230.363
R13721 ringtest_0.x4._11_ ringtest_0.x4._11_.n30 216.464
R13722 ringtest_0.x4._11_.n24 ringtest_0.x4._11_.t20 206.19
R13723 ringtest_0.x4._11_.n5 ringtest_0.x4._11_.t17 206.19
R13724 ringtest_0.x4._11_.n11 ringtest_0.x4._11_.t11 183.505
R13725 ringtest_0.x4._11_.n8 ringtest_0.x4._11_.t21 169.237
R13726 ringtest_0.x4._11_.n3 ringtest_0.x4._11_.t7 169.237
R13727 ringtest_0.x4._11_.n21 ringtest_0.x4._11_.t16 158.064
R13728 ringtest_0.x4._11_ ringtest_0.x4._11_.n3 157.555
R13729 ringtest_0.x4._11_ ringtest_0.x4._11_.n8 157.166
R13730 ringtest_0.x4._11_.n1 ringtest_0.x4._11_.t9 157.07
R13731 ringtest_0.x4._11_.n18 ringtest_0.x4._11_.t15 155.847
R13732 ringtest_0.x4._11_.n22 ringtest_0.x4._11_.n21 154.048
R13733 ringtest_0.x4._11_.n12 ringtest_0.x4._11_.n11 153.863
R13734 ringtest_0.x4._11_.n19 ringtest_0.x4._11_.n18 153.13
R13735 ringtest_0.x4._11_.n25 ringtest_0.x4._11_.n24 152
R13736 ringtest_0.x4._11_.n15 ringtest_0.x4._11_.n14 152
R13737 ringtest_0.x4._11_.n6 ringtest_0.x4._11_.n5 152
R13738 ringtest_0.x4._11_.n2 ringtest_0.x4._11_.n1 152
R13739 ringtest_0.x4._11_.n14 ringtest_0.x4._11_.t4 150.03
R13740 ringtest_0.x4._11_.n11 ringtest_0.x4._11_.t18 114.532
R13741 ringtest_0.x4._11_.n27 ringtest_0.x4._11_.n26 41.0809
R13742 ringtest_0.x4._11_.n30 ringtest_0.x4._11_.t0 38.5719
R13743 ringtest_0.x4._11_.n30 ringtest_0.x4._11_.t1 38.5719
R13744 ringtest_0.x4._11_.n0 ringtest_0.x4._11_.t3 26.5955
R13745 ringtest_0.x4._11_.n0 ringtest_0.x4._11_.t2 26.5955
R13746 ringtest_0.x4._11_.n17 ringtest_0.x4._11_.n16 25.2401
R13747 ringtest_0.x4._11_.n20 ringtest_0.x4._11_.n19 22.3199
R13748 ringtest_0.x4._11_.n10 ringtest_0.x4._11_.n9 21.8442
R13749 ringtest_0.x4._11_.n10 ringtest_0.x4._11_.n7 20.8523
R13750 ringtest_0.x4._11_.n28 ringtest_0.x4._11_.n27 13.7699
R13751 ringtest_0.x4._11_.n28 ringtest_0.x4._11_.n2 12.7179
R13752 ringtest_0.x4._11_.n4 ringtest_0.x4._11_ 12.3175
R13753 ringtest_0.x4._11_.n9 ringtest_0.x4._11_ 11.4531
R13754 ringtest_0.x4._11_.n7 ringtest_0.x4._11_.n4 11.4418
R13755 ringtest_0.x4._11_.n23 ringtest_0.x4._11_.n20 10.8618
R13756 ringtest_0.x4._11_.n7 ringtest_0.x4._11_.n6 10.3976
R13757 ringtest_0.x4._11_.n25 ringtest_0.x4._11_ 9.6005
R13758 ringtest_0.x4._11_.n29 ringtest_0.x4._11_ 9.6005
R13759 ringtest_0.x4._11_ ringtest_0.x4._11_.n22 9.39918
R13760 ringtest_0.x4._11_.n13 ringtest_0.x4._11_.n12 9.3005
R13761 ringtest_0.x4._11_.n29 ringtest_0.x4._11_.n28 9.3005
R13762 ringtest_0.x4._11_.n23 ringtest_0.x4._11_ 8.80957
R13763 ringtest_0.x4._11_.n6 ringtest_0.x4._11_ 8.22907
R13764 ringtest_0.x4._11_.n15 ringtest_0.x4._11_ 7.6805
R13765 ringtest_0.x4._11_.n16 ringtest_0.x4._11_.n15 4.6085
R13766 ringtest_0.x4._11_.n16 ringtest_0.x4._11_ 4.58918
R13767 ringtest_0.x4._11_.n22 ringtest_0.x4._11_ 4.3525
R13768 ringtest_0.x4._11_.n4 ringtest_0.x4._11_ 4.10616
R13769 ringtest_0.x4._11_.n9 ringtest_0.x4._11_ 3.81804
R13770 ringtest_0.x4._11_.n26 ringtest_0.x4._11_ 3.62717
R13771 ringtest_0.x4._11_.n19 ringtest_0.x4._11_ 3.2005
R13772 ringtest_0.x4._11_ ringtest_0.x4._11_.n29 3.2005
R13773 ringtest_0.x4._11_.n17 ringtest_0.x4._11_.n13 2.49494
R13774 ringtest_0.x4._11_.n2 ringtest_0.x4._11_ 2.3045
R13775 ringtest_0.x4._11_.n12 ringtest_0.x4._11_ 1.97868
R13776 ringtest_0.x4._11_.n13 ringtest_0.x4._11_.n10 1.71582
R13777 ringtest_0.x4._11_.n27 ringtest_0.x4._11_.n23 1.38649
R13778 ringtest_0.x4._11_.n26 ringtest_0.x4._11_.n25 1.2805
R13779 ringtest_0.x4._11_.n20 ringtest_0.x4._11_.n17 1.24753
R13780 ui_in[0].n5 ui_in[0].t7 327.99
R13781 ui_in[0].n9 ui_in[0].t4 293.969
R13782 ui_in[0].n3 ui_in[0].t5 261.887
R13783 ui_in[0].n0 ui_in[0].t8 212.081
R13784 ui_in[0].n1 ui_in[0].t6 212.081
R13785 ui_in[0].n5 ui_in[0].t1 199.457
R13786 ui_in[0].n2 ui_in[0].n1 183.185
R13787 ui_in[0].n3 ui_in[0].t9 155.847
R13788 ui_in[0] ui_in[0].n9 154.065
R13789 ui_in[0].n4 ui_in[0].n3 153.506
R13790 ui_in[0].n6 ui_in[0].n5 152
R13791 ui_in[0].n0 ui_in[0].t3 139.78
R13792 ui_in[0].n1 ui_in[0].t0 139.78
R13793 ui_in[0].n9 ui_in[0].t2 138.338
R13794 ui_in[0].n1 ui_in[0].n0 61.346
R13795 ui_in[0].n13 ui_in[0] 38.2119
R13796 ui_in[0].n10 ui_in[0] 13.4199
R13797 ui_in[0].n11 ui_in[0].n8 11.7395
R13798 ui_in[0].n12 ui_in[0].n11 11.5949
R13799 ui_in[0].n8 ui_in[0].n4 10.4004
R13800 ui_in[0].n12 ui_in[0].n2 9.68118
R13801 ui_in[0].n6 ui_in[0] 9.6005
R13802 ui_in[0].n2 ui_in[0] 5.8885
R13803 ui_in[0].n10 ui_in[0] 5.57469
R13804 ui_in[0].n13 ui_in[0] 4.74482
R13805 ui_in[0].n8 ui_in[0].n7 4.6505
R13806 ui_in[0].n11 ui_in[0].n10 4.6505
R13807 ui_in[0].n7 ui_in[0].n6 2.98717
R13808 ui_in[0].n4 ui_in[0] 2.82403
R13809 ui_in[0].n7 ui_in[0] 1.9205
R13810 ui_in[0] ui_in[0].n12 0.559212
R13811 ui_in[0] ui_in[0].n13 0.02675
R13812 muxtest_0.R3R4.n5 muxtest_0.R3R4.t3 26.3998
R13813 muxtest_0.R3R4.n0 muxtest_0.R3R4.t6 26.3998
R13814 muxtest_0.R3R4.n5 muxtest_0.R3R4.t2 23.5483
R13815 muxtest_0.R3R4.n0 muxtest_0.R3R4.t5 23.5483
R13816 muxtest_0.R3R4.n6 muxtest_0.R3R4.t9 12.9758
R13817 muxtest_0.R3R4.n1 muxtest_0.R3R4.t0 12.9758
R13818 muxtest_0.R3R4.n6 muxtest_0.R3R4.t8 10.8618
R13819 muxtest_0.R3R4.n1 muxtest_0.R3R4.t1 10.8618
R13820 muxtest_0.R3R4.n4 muxtest_0.R3R4.t7 10.5285
R13821 muxtest_0.R3R4.n11 muxtest_0.R3R4.n10 7.08509
R13822 muxtest_0.R3R4.n7 muxtest_0.R3R4.n5 3.06895
R13823 muxtest_0.R3R4.n2 muxtest_0.R3R4.n0 3.06895
R13824 muxtest_0.R3R4.n7 muxtest_0.R3R4.n6 2.14822
R13825 muxtest_0.R3R4.n2 muxtest_0.R3R4.n1 2.14822
R13826 muxtest_0.R3R4.n8 muxtest_0.R3R4.n7 1.12636
R13827 muxtest_0.R3R4.n3 muxtest_0.R3R4.n2 1.12636
R13828 muxtest_0.R3R4.n4 muxtest_0.R3R4.t4 1.06523
R13829 muxtest_0.R3R4.n12 muxtest_0.R3R4 0.893
R13830 muxtest_0.R3R4.n9 muxtest_0.R3R4 0.670143
R13831 muxtest_0.R3R4.n12 muxtest_0.R3R4.n11 0.40675
R13832 muxtest_0.R3R4.n10 muxtest_0.R3R4.n9 0.223714
R13833 muxtest_0.R3R4.n11 muxtest_0.R3R4.n4 0.183423
R13834 muxtest_0.R3R4 muxtest_0.R3R4.n3 0.148615
R13835 muxtest_0.R3R4.n9 muxtest_0.R3R4.n8 0.132418
R13836 muxtest_0.R3R4.n12 muxtest_0.R3R4 0.08425
R13837 muxtest_0.R3R4.n8 muxtest_0.R3R4 0.0655
R13838 muxtest_0.R3R4.n3 muxtest_0.R3R4 0.0655
R13839 muxtest_0.R3R4 muxtest_0.R3R4.n12 0.04425
R13840 muxtest_0.R3R4.n10 muxtest_0.R3R4 0.00907843
R13841 ui_in[4].n26 ui_in[4].t3 327.99
R13842 ui_in[4].n10 ui_in[4].t0 327.99
R13843 ui_in[4].n19 ui_in[4].t1 293.969
R13844 ui_in[4].n3 ui_in[4].t19 293.969
R13845 ui_in[4].n22 ui_in[4].t14 256.07
R13846 ui_in[4].n6 ui_in[4].t12 256.07
R13847 ui_in[4].n16 ui_in[4].t9 212.081
R13848 ui_in[4].n17 ui_in[4].t15 212.081
R13849 ui_in[4].n0 ui_in[4].t6 212.081
R13850 ui_in[4].n1 ui_in[4].t4 212.081
R13851 ui_in[4].n26 ui_in[4].t8 199.457
R13852 ui_in[4].n10 ui_in[4].t5 199.457
R13853 ui_in[4].n18 ui_in[4].n17 182.929
R13854 ui_in[4].n2 ui_in[4].n1 182.929
R13855 ui_in[4] ui_in[4].n19 154.065
R13856 ui_in[4] ui_in[4].n3 154.065
R13857 ui_in[4].n27 ui_in[4].n26 152
R13858 ui_in[4].n23 ui_in[4].n22 152
R13859 ui_in[4].n11 ui_in[4].n10 152
R13860 ui_in[4].n7 ui_in[4].n6 152
R13861 ui_in[4].n22 ui_in[4].t11 150.03
R13862 ui_in[4].n6 ui_in[4].t7 150.03
R13863 ui_in[4].n16 ui_in[4].t18 139.78
R13864 ui_in[4].n17 ui_in[4].t2 139.78
R13865 ui_in[4].n0 ui_in[4].t16 139.78
R13866 ui_in[4].n1 ui_in[4].t10 139.78
R13867 ui_in[4].n19 ui_in[4].t17 138.338
R13868 ui_in[4].n3 ui_in[4].t13 138.338
R13869 ui_in[4].n17 ui_in[4].n16 61.346
R13870 ui_in[4].n1 ui_in[4].n0 61.346
R13871 ui_in[4].n31 ui_in[4] 29.9743
R13872 ui_in[4].n21 ui_in[4] 17.455
R13873 ui_in[4].n5 ui_in[4] 17.455
R13874 ui_in[4].n30 ui_in[4].n29 14.6836
R13875 ui_in[4].n14 ui_in[4].n13 14.6836
R13876 ui_in[4].n29 ui_in[4].n28 14.6704
R13877 ui_in[4].n13 ui_in[4].n12 14.6704
R13878 ui_in[4].n20 ui_in[4] 13.8328
R13879 ui_in[4].n4 ui_in[4] 13.8328
R13880 ui_in[4].n31 ui_in[4] 12.499
R13881 ui_in[4].n30 ui_in[4].n18 10.6811
R13882 ui_in[4].n14 ui_in[4].n2 10.6811
R13883 ui_in[4].n23 ui_in[4].n21 10.4374
R13884 ui_in[4].n7 ui_in[4].n5 10.4374
R13885 ui_in[4].n25 ui_in[4].n24 8.15776
R13886 ui_in[4].n9 ui_in[4].n8 8.15776
R13887 ui_in[4].n28 ui_in[4] 6.61383
R13888 ui_in[4].n12 ui_in[4] 6.61383
R13889 ui_in[4].n18 ui_in[4] 6.1445
R13890 ui_in[4].n2 ui_in[4] 6.1445
R13891 ui_in[4].n20 ui_in[4] 5.16179
R13892 ui_in[4].n4 ui_in[4] 5.16179
R13893 ui_in[4].n27 ui_in[4] 4.90717
R13894 ui_in[4].n11 ui_in[4] 4.90717
R13895 ui_in[4].n25 ui_in[4].n20 4.65206
R13896 ui_in[4].n9 ui_in[4].n4 4.65206
R13897 ui_in[4].n24 ui_in[4] 3.93896
R13898 ui_in[4].n8 ui_in[4] 3.93896
R13899 ui_in[4].n28 ui_in[4].n27 2.98717
R13900 ui_in[4].n12 ui_in[4].n11 2.98717
R13901 ui_in[4].n21 ui_in[4] 2.16665
R13902 ui_in[4].n5 ui_in[4] 2.16665
R13903 ui_in[4].n24 ui_in[4].n23 1.57588
R13904 ui_in[4].n8 ui_in[4].n7 1.57588
R13905 ui_in[4].n29 ui_in[4].n25 0.79438
R13906 ui_in[4].n13 ui_in[4].n9 0.79438
R13907 ui_in[4] ui_in[4].n15 0.287559
R13908 ui_in[4] ui_in[4].n31 0.28675
R13909 ui_in[4] ui_in[4].n30 0.248606
R13910 ui_in[4] ui_in[4].n14 0.248606
R13911 ui_in[4].n15 ui_in[4] 0.11603
R13912 ui_in[4].n15 ui_in[4] 0.0460882
R13913 muxtest_0.R1R2.n0 muxtest_0.R1R2.t1 26.3998
R13914 muxtest_0.R1R2.n0 muxtest_0.R1R2.t0 23.5483
R13915 muxtest_0.R1R2.n1 muxtest_0.R1R2.t5 12.9758
R13916 muxtest_0.R1R2.n4 muxtest_0.R1R2.t3 10.8648
R13917 muxtest_0.R1R2.n1 muxtest_0.R1R2.t4 10.8618
R13918 muxtest_0.R1R2.n4 muxtest_0.R1R2.t2 10.5295
R13919 muxtest_0.R1R2.n2 muxtest_0.R1R2.n0 3.06895
R13920 muxtest_0.R1R2.n2 muxtest_0.R1R2.n1 2.14822
R13921 muxtest_0.R1R2.n3 muxtest_0.R1R2.n2 1.12636
R13922 muxtest_0.R1R2.n5 muxtest_0.R1R2 0.96675
R13923 muxtest_0.R1R2.n5 muxtest_0.R1R2.n4 0.494965
R13924 muxtest_0.R1R2 muxtest_0.R1R2.n3 0.132418
R13925 muxtest_0.R1R2.n5 muxtest_0.R1R2 0.06925
R13926 muxtest_0.R1R2.n3 muxtest_0.R1R2 0.0655
R13927 muxtest_0.R1R2 muxtest_0.R1R2.n5 0.04425
R13928 a_19289_13081.n0 a_19289_13081.t12 1681.78
R13929 a_19289_13081.n2 a_19289_13081.t7 1681.21
R13930 a_19289_13081.n1 a_19289_13081.t13 1681.21
R13931 a_19289_13081.n0 a_19289_13081.t2 1681.21
R13932 a_19289_13081.n13 a_19289_13081.t14 1681.21
R13933 a_19289_13081.n11 a_19289_13081.t10 1681.21
R13934 a_19289_13081.n9 a_19289_13081.t17 1681.21
R13935 a_19289_13081.n7 a_19289_13081.t9 1681.21
R13936 a_19289_13081.n3 a_19289_13081.t4 703.317
R13937 a_19289_13081.n7 a_19289_13081.t6 702.768
R13938 a_19289_13081.n5 a_19289_13081.t11 702.747
R13939 a_19289_13081.n4 a_19289_13081.t5 702.747
R13940 a_19289_13081.n3 a_19289_13081.t15 702.747
R13941 a_19289_13081.n12 a_19289_13081.t3 702.747
R13942 a_19289_13081.n10 a_19289_13081.t8 702.747
R13943 a_19289_13081.n8 a_19289_13081.t16 702.747
R13944 a_19289_13081.n6 a_19289_13081.t0 30.088
R13945 a_19289_13081.t1 a_19289_13081.n15 26.0464
R13946 a_19289_13081.n15 a_19289_13081.n2 20.0759
R13947 a_19289_13081.n6 a_19289_13081.n5 0.875353
R13948 a_19289_13081.n1 a_19289_13081.n0 0.576859
R13949 a_19289_13081.n2 a_19289_13081.n1 0.576859
R13950 a_19289_13081.n4 a_19289_13081.n3 0.570292
R13951 a_19289_13081.n5 a_19289_13081.n4 0.570292
R13952 a_19289_13081.n15 a_19289_13081.n14 0.267403
R13953 a_19289_13081.n14 a_19289_13081.n6 0.10833
R13954 a_19289_13081.n14 a_19289_13081.n13 0.0744583
R13955 a_19289_13081.n8 a_19289_13081.n7 0.0205
R13956 a_19289_13081.n9 a_19289_13081.n8 0.0205
R13957 a_19289_13081.n10 a_19289_13081.n9 0.0205
R13958 a_19289_13081.n11 a_19289_13081.n10 0.0205
R13959 a_19289_13081.n12 a_19289_13081.n11 0.0205
R13960 a_19289_13081.n13 a_19289_13081.n12 0.0205
R13961 ringtest_0.drv_out.n7 ringtest_0.drv_out.t21 184.768
R13962 ringtest_0.drv_out.n6 ringtest_0.drv_out.t20 184.768
R13963 ringtest_0.drv_out.n5 ringtest_0.drv_out.t23 184.768
R13964 ringtest_0.drv_out.n4 ringtest_0.drv_out.t22 184.768
R13965 ringtest_0.drv_out.n8 ringtest_0.drv_out.n7 171.375
R13966 ringtest_0.drv_out.n7 ringtest_0.drv_out.t25 146.208
R13967 ringtest_0.drv_out.n6 ringtest_0.drv_out.t24 146.208
R13968 ringtest_0.drv_out.n5 ringtest_0.drv_out.t27 146.208
R13969 ringtest_0.drv_out.n4 ringtest_0.drv_out.t26 146.208
R13970 ringtest_0.drv_out.n7 ringtest_0.drv_out.n6 40.6397
R13971 ringtest_0.drv_out.n6 ringtest_0.drv_out.n5 40.6397
R13972 ringtest_0.drv_out.n5 ringtest_0.drv_out.n4 40.6397
R13973 ringtest_0.drv_out.n0 ringtest_0.drv_out.t19 26.3998
R13974 ringtest_0.drv_out.n21 ringtest_0.drv_out.n20 26.0838
R13975 ringtest_0.drv_out.n21 ringtest_0.drv_out.n17 26.0838
R13976 ringtest_0.drv_out.n21 ringtest_0.drv_out.n19 26.0838
R13977 ringtest_0.drv_out.n21 ringtest_0.drv_out.n18 26.0838
R13978 ringtest_0.drv_out.n16 ringtest_0.drv_out.n12 24.902
R13979 ringtest_0.drv_out.n16 ringtest_0.drv_out.n14 24.902
R13980 ringtest_0.drv_out.n16 ringtest_0.drv_out.n13 24.902
R13981 ringtest_0.drv_out.n16 ringtest_0.drv_out.n15 24.902
R13982 ringtest_0.drv_out.n0 ringtest_0.drv_out.t0 23.5483
R13983 ringtest_0.drv_out.n1 ringtest_0.drv_out.t1 12.9758
R13984 ringtest_0.drv_out ringtest_0.drv_out.n8 12.3171
R13985 ringtest_0.drv_out.n1 ringtest_0.drv_out.t2 10.8618
R13986 ringtest_0.drv_out.n20 ringtest_0.drv_out.t10 6.6005
R13987 ringtest_0.drv_out.n20 ringtest_0.drv_out.t5 6.6005
R13988 ringtest_0.drv_out.n17 ringtest_0.drv_out.t6 6.6005
R13989 ringtest_0.drv_out.n17 ringtest_0.drv_out.t8 6.6005
R13990 ringtest_0.drv_out.n19 ringtest_0.drv_out.t3 6.6005
R13991 ringtest_0.drv_out.n19 ringtest_0.drv_out.t4 6.6005
R13992 ringtest_0.drv_out.n18 ringtest_0.drv_out.t7 6.6005
R13993 ringtest_0.drv_out.n18 ringtest_0.drv_out.t9 6.6005
R13994 ringtest_0.drv_out.n11 ringtest_0.drv_out 5.69273
R13995 ringtest_0.drv_out.n12 ringtest_0.drv_out.t17 3.61217
R13996 ringtest_0.drv_out.n12 ringtest_0.drv_out.t12 3.61217
R13997 ringtest_0.drv_out.n14 ringtest_0.drv_out.t13 3.61217
R13998 ringtest_0.drv_out.n14 ringtest_0.drv_out.t15 3.61217
R13999 ringtest_0.drv_out.n13 ringtest_0.drv_out.t14 3.61217
R14000 ringtest_0.drv_out.n13 ringtest_0.drv_out.t16 3.61217
R14001 ringtest_0.drv_out.n15 ringtest_0.drv_out.t18 3.61217
R14002 ringtest_0.drv_out.n15 ringtest_0.drv_out.t11 3.61217
R14003 ringtest_0.drv_out.n2 ringtest_0.drv_out.n0 3.06895
R14004 ringtest_0.drv_out.n11 ringtest_0.drv_out 2.87193
R14005 ringtest_0.drv_out.n8 ringtest_0.drv_out 2.23542
R14006 ringtest_0.drv_out.n2 ringtest_0.drv_out.n1 2.14822
R14007 ringtest_0.drv_out.n10 ringtest_0.drv_out 1.7806
R14008 ringtest_0.drv_out ringtest_0.drv_out.n10 1.54574
R14009 ringtest_0.drv_out.n9 ringtest_0.drv_out 1.25273
R14010 ringtest_0.drv_out.n3 ringtest_0.drv_out.n2 1.12636
R14011 ringtest_0.drv_out ringtest_0.drv_out.n22 0.461707
R14012 ringtest_0.drv_out.n9 ringtest_0.drv_out 0.316378
R14013 ringtest_0.drv_out ringtest_0.drv_out.n11 0.188041
R14014 ringtest_0.drv_out ringtest_0.drv_out.n3 0.138152
R14015 ringtest_0.drv_out.n22 ringtest_0.drv_out.n16 0.0921193
R14016 ringtest_0.drv_out.n22 ringtest_0.drv_out.n21 0.069392
R14017 ringtest_0.drv_out.n3 ringtest_0.drv_out 0.0655
R14018 ringtest_0.drv_out.n10 ringtest_0.drv_out.n9 0.0596216
R14019 ringtest_0.x4.net3.t3 ringtest_0.x4.net3.t4 395.01
R14020 ringtest_0.x4.net3 ringtest_0.x4.net3.t3 320.745
R14021 ringtest_0.x4.net3.n3 ringtest_0.x4.net3.t6 260.322
R14022 ringtest_0.x4.net3.n0 ringtest_0.x4.net3.t7 229.369
R14023 ringtest_0.x4.net3.n7 ringtest_0.x4.net3.t1 222.68
R14024 ringtest_0.x4.net3.n3 ringtest_0.x4.net3.t5 175.169
R14025 ringtest_0.x4.net3.n0 ringtest_0.x4.net3.t2 157.07
R14026 ringtest_0.x4.net3.n4 ringtest_0.x4.net3.n3 152
R14027 ringtest_0.x4.net3.n1 ringtest_0.x4.net3.n0 152
R14028 ringtest_0.x4.net3.n8 ringtest_0.x4.net3.t0 132.322
R14029 ringtest_0.x4.net3.n8 ringtest_0.x4.net3.n7 95.0273
R14030 ringtest_0.x4.net3.n5 ringtest_0.x4.net3 25.2581
R14031 ringtest_0.x4.net3.n5 ringtest_0.x4.net3 20.1696
R14032 ringtest_0.x4.net3.n7 ringtest_0.x4.net3.n6 12.7813
R14033 ringtest_0.x4.net3.n1 ringtest_0.x4.net3 12.0005
R14034 ringtest_0.x4.net3 ringtest_0.x4.net3.n4 11.2497
R14035 ringtest_0.x4.net3.n6 ringtest_0.x4.net3.n2 9.79203
R14036 ringtest_0.x4.net3.n6 ringtest_0.x4.net3.n5 5.9277
R14037 ringtest_0.x4.net3.n2 ringtest_0.x4.net3 4.53383
R14038 ringtest_0.x4.net3 ringtest_0.x4.net3.n8 2.70465
R14039 ringtest_0.x4.net3.n2 ringtest_0.x4.net3.n1 1.6005
R14040 ringtest_0.x4.net3.n4 ringtest_0.x4.net3 1.55726
R14041 ui_in[2].n2 ui_in[2].t0 450.938
R14042 ui_in[2].n2 ui_in[2].t6 445.666
R14043 ui_in[2].n0 ui_in[2].t7 377.486
R14044 ui_in[2].n0 ui_in[2].t1 374.202
R14045 ui_in[2].n5 ui_in[2].t2 212.081
R14046 ui_in[2].n6 ui_in[2].t3 212.081
R14047 ui_in[2].n7 ui_in[2].n6 183.441
R14048 ui_in[2].n5 ui_in[2].t4 139.78
R14049 ui_in[2].n6 ui_in[2].t5 139.78
R14050 ui_in[2].n6 ui_in[2].n5 61.346
R14051 ui_in[2].n4 ui_in[2].n1 12.4088
R14052 ui_in[2] ui_in[2].n7 11.4331
R14053 ui_in[2].n4 ui_in[2].n3 9.10647
R14054 ui_in[2].n8 ui_in[2].n4 8.98648
R14055 ui_in[2].n7 ui_in[2] 5.6325
R14056 ui_in[2].n8 ui_in[2] 5.02323
R14057 ui_in[2].n3 ui_in[2].n2 3.1748
R14058 ui_in[2] ui_in[2].n0 2.04102
R14059 ui_in[2] ui_in[2].n8 0.888758
R14060 ui_in[2].n1 ui_in[2] 0.412375
R14061 ui_in[2].n3 ui_in[2] 0.063625
R14062 ui_in[2].n1 ui_in[2] 0.061125
R14063 ringtest_0.x3.x2.GP4.n2 ringtest_0.x3.x2.GP4.t5 450.938
R14064 ringtest_0.x3.x2.GP4.n2 ringtest_0.x3.x2.GP4.t4 445.666
R14065 ringtest_0.x3.x2.GP4.n5 ringtest_0.x3.x2.GP4.n4 208.965
R14066 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n0 96.8352
R14067 ringtest_0.x3.x2.GP4.n4 ringtest_0.x3.x2.GP4.t3 26.5955
R14068 ringtest_0.x3.x2.GP4.n4 ringtest_0.x3.x2.GP4.t2 26.5955
R14069 ringtest_0.x3.x2.GP4.n0 ringtest_0.x3.x2.GP4.t1 24.9236
R14070 ringtest_0.x3.x2.GP4.n0 ringtest_0.x3.x2.GP4.t0 24.9236
R14071 ringtest_0.x3.x1.gpo3 ringtest_0.x3.x2.x4.GP 16.5032
R14072 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n3 10.2405
R14073 ringtest_0.x3.x2.GP4.n3 ringtest_0.x3.x1.gpo3 7.76481
R14074 ringtest_0.x3.x2.GP4.n1 ringtest_0.x3.x1.x14.Y 6.1445
R14075 ringtest_0.x3.x2.GP4.n1 ringtest_0.x3.x1.x14.Y 4.65505
R14076 ringtest_0.x3.x2.x4.GP ringtest_0.x3.x2.GP4.n2 2.95993
R14077 ringtest_0.x3.x2.GP4.n5 ringtest_0.x3.x1.x14.Y 2.0485
R14078 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n5 1.55202
R14079 ringtest_0.x3.x2.GP4.n3 ringtest_0.x3.x2.GP4.n1 1.0245
R14080 ringtest_0.counter7.n0 ringtest_0.counter7.t5 368.521
R14081 ringtest_0.counter7.n1 ringtest_0.counter7.t4 216.155
R14082 ringtest_0.counter7.n1 ringtest_0.counter7 78.8791
R14083 ringtest_0.counter7.n4 ringtest_0.counter7.t0 26.3998
R14084 ringtest_0.counter7.n4 ringtest_0.counter7.t1 23.5483
R14085 ringtest_0.counter7.n3 ringtest_0.counter7.n2 18.2765
R14086 ringtest_0.counter7.n5 ringtest_0.counter7.t3 12.9758
R14087 ringtest_0.counter7.n5 ringtest_0.counter7.t2 10.8618
R14088 ringtest_0.counter7 ringtest_0.counter7.n0 10.5563
R14089 ringtest_0.counter7.n0 ringtest_0.counter7 5.48477
R14090 ringtest_0.counter7.n2 ringtest_0.counter7 4.18512
R14091 ringtest_0.counter7.n6 ringtest_0.counter7.n4 3.06895
R14092 ringtest_0.counter7.n6 ringtest_0.counter7.n5 2.14822
R14093 ringtest_0.counter7 ringtest_0.counter7.n6 1.27287
R14094 ringtest_0.counter7.n3 ringtest_0.counter7 1.27059
R14095 ringtest_0.counter7.n2 ringtest_0.counter7.n1 0.985115
R14096 ringtest_0.counter7 ringtest_0.counter7.n3 0.647091
R14097 ua[1].n6 ua[1].t12 23.6581
R14098 ua[1].n12 ua[1].t7 23.6581
R14099 ua[1].n19 ua[1].t2 23.6581
R14100 ua[1].n1 ua[1].t1 23.6581
R14101 ua[1].n5 ua[1].t4 23.3739
R14102 ua[1].n11 ua[1].t13 23.3739
R14103 ua[1].n18 ua[1].t3 23.3739
R14104 ua[1].n0 ua[1].t0 23.3739
R14105 ua[1].n25 ua[1] 15.3856
R14106 ua[1].n6 ua[1].t8 10.7528
R14107 ua[1].n12 ua[1].t11 10.7528
R14108 ua[1].n19 ua[1].t15 10.7528
R14109 ua[1].n1 ua[1].t5 10.7528
R14110 ua[1].n8 ua[1].t9 10.6417
R14111 ua[1].n14 ua[1].t10 10.6417
R14112 ua[1].n21 ua[1].t14 10.6417
R14113 ua[1].n3 ua[1].t6 10.6417
R14114 ua[1].n7 ua[1].n6 1.30064
R14115 ua[1].n13 ua[1].n12 1.30064
R14116 ua[1].n20 ua[1].n19 1.30064
R14117 ua[1].n2 ua[1].n1 1.30064
R14118 ua[1] ua[1].n4 0.983856
R14119 ua[1].n23 ua[1].n22 0.946356
R14120 ua[1].n16 ua[1].n15 0.927606
R14121 ua[1].n10 ua[1].n9 0.925106
R14122 ua[1].n17 ua[1] 0.748625
R14123 ua[1].n7 ua[1].n5 0.726502
R14124 ua[1].n13 ua[1].n11 0.726502
R14125 ua[1].n20 ua[1].n18 0.726502
R14126 ua[1].n2 ua[1].n0 0.726502
R14127 ua[1].n24 ua[1].n17 0.54425
R14128 ua[1].n25 ua[1] 0.532375
R14129 ua[1].n8 ua[1].n7 0.512491
R14130 ua[1].n14 ua[1].n13 0.512491
R14131 ua[1].n21 ua[1].n20 0.512491
R14132 ua[1].n3 ua[1].n2 0.512491
R14133 ua[1].n9 ua[1].n8 0.359663
R14134 ua[1].n15 ua[1].n14 0.359663
R14135 ua[1].n22 ua[1].n21 0.359663
R14136 ua[1].n4 ua[1].n3 0.359663
R14137 ua[1].n9 ua[1].n5 0.216071
R14138 ua[1].n15 ua[1].n11 0.216071
R14139 ua[1].n22 ua[1].n18 0.216071
R14140 ua[1].n4 ua[1].n0 0.216071
R14141 ua[1].n17 ua[1] 0.20175
R14142 ua[1].n24 ua[1] 0.17925
R14143 ua[1] ua[1].n25 0.178
R14144 ua[1].n24 ua[1] 0.063
R14145 ua[1].n10 ua[1] 0.05925
R14146 ua[1].n16 ua[1] 0.05675
R14147 ua[1] ua[1].n16 0.0561931
R14148 ua[1] ua[1].n10 0.0561872
R14149 ua[1].n23 ua[1] 0.038
R14150 ua[1] ua[1].n23 0.0376287
R14151 ua[1] ua[1].n24 0.004875
R14152 ringtest_0.x4.clknet_1_0__leaf_clk.n25 ringtest_0.x4.clknet_1_0__leaf_clk.n23 333.392
R14153 ringtest_0.x4.clknet_1_0__leaf_clk.n25 ringtest_0.x4.clknet_1_0__leaf_clk.n24 301.392
R14154 ringtest_0.x4.clknet_1_0__leaf_clk.n27 ringtest_0.x4.clknet_1_0__leaf_clk.n26 301.392
R14155 ringtest_0.x4.clknet_1_0__leaf_clk.n29 ringtest_0.x4.clknet_1_0__leaf_clk.n28 301.392
R14156 ringtest_0.x4.clknet_1_0__leaf_clk.n22 ringtest_0.x4.clknet_1_0__leaf_clk.n4 301.392
R14157 ringtest_0.x4.clknet_1_0__leaf_clk.n31 ringtest_0.x4.clknet_1_0__leaf_clk.n30 301.392
R14158 ringtest_0.x4.clknet_1_0__leaf_clk.n21 ringtest_0.x4.clknet_1_0__leaf_clk.n5 297.863
R14159 ringtest_0.x4.clknet_1_0__leaf_clk.n2 ringtest_0.x4.clknet_1_0__leaf_clk.t32 294.557
R14160 ringtest_0.x4.clknet_1_0__leaf_clk.n0 ringtest_0.x4.clknet_1_0__leaf_clk.t38 294.557
R14161 ringtest_0.x4.clknet_1_0__leaf_clk.n41 ringtest_0.x4.clknet_1_0__leaf_clk.t35 294.557
R14162 ringtest_0.x4.clknet_1_0__leaf_clk.n38 ringtest_0.x4.clknet_1_0__leaf_clk.t33 294.557
R14163 ringtest_0.x4.clknet_1_0__leaf_clk.n36 ringtest_0.x4.clknet_1_0__leaf_clk.t36 294.557
R14164 ringtest_0.x4.clknet_1_0__leaf_clk.n34 ringtest_0.x4.clknet_1_0__leaf_clk.n33 287.303
R14165 ringtest_0.x4.clknet_1_0__leaf_clk.n8 ringtest_0.x4.clknet_1_0__leaf_clk.n6 248.638
R14166 ringtest_0.x4.clknet_1_0__leaf_clk.n2 ringtest_0.x4.clknet_1_0__leaf_clk.t37 211.01
R14167 ringtest_0.x4.clknet_1_0__leaf_clk.n0 ringtest_0.x4.clknet_1_0__leaf_clk.t41 211.01
R14168 ringtest_0.x4.clknet_1_0__leaf_clk.n41 ringtest_0.x4.clknet_1_0__leaf_clk.t34 211.01
R14169 ringtest_0.x4.clknet_1_0__leaf_clk.n38 ringtest_0.x4.clknet_1_0__leaf_clk.t40 211.01
R14170 ringtest_0.x4.clknet_1_0__leaf_clk.n36 ringtest_0.x4.clknet_1_0__leaf_clk.t39 211.01
R14171 ringtest_0.x4.clknet_1_0__leaf_clk.n8 ringtest_0.x4.clknet_1_0__leaf_clk.n7 203.463
R14172 ringtest_0.x4.clknet_1_0__leaf_clk.n10 ringtest_0.x4.clknet_1_0__leaf_clk.n9 203.463
R14173 ringtest_0.x4.clknet_1_0__leaf_clk.n14 ringtest_0.x4.clknet_1_0__leaf_clk.n13 203.463
R14174 ringtest_0.x4.clknet_1_0__leaf_clk.n16 ringtest_0.x4.clknet_1_0__leaf_clk.n15 203.463
R14175 ringtest_0.x4.clknet_1_0__leaf_clk.n18 ringtest_0.x4.clknet_1_0__leaf_clk.n17 203.463
R14176 ringtest_0.x4.clknet_1_0__leaf_clk.n12 ringtest_0.x4.clknet_1_0__leaf_clk.n11 202.456
R14177 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n19 199.607
R14178 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n2 156.207
R14179 ringtest_0.x4.clknet_1_0__leaf_clk.n37 ringtest_0.x4.clknet_1_0__leaf_clk.n36 153.097
R14180 ringtest_0.x4.clknet_1_0__leaf_clk.n39 ringtest_0.x4.clknet_1_0__leaf_clk.n38 152.296
R14181 ringtest_0.x4.clknet_1_0__leaf_clk.n1 ringtest_0.x4.clknet_1_0__leaf_clk.n0 152
R14182 ringtest_0.x4.clknet_1_0__leaf_clk.n42 ringtest_0.x4.clknet_1_0__leaf_clk.n41 152
R14183 ringtest_0.x4.clknet_1_0__leaf_clk.n10 ringtest_0.x4.clknet_1_0__leaf_clk.n8 45.177
R14184 ringtest_0.x4.clknet_1_0__leaf_clk.n16 ringtest_0.x4.clknet_1_0__leaf_clk.n14 45.177
R14185 ringtest_0.x4.clknet_1_0__leaf_clk.n18 ringtest_0.x4.clknet_1_0__leaf_clk.n16 45.177
R14186 ringtest_0.x4.clknet_1_0__leaf_clk.n12 ringtest_0.x4.clknet_1_0__leaf_clk.n10 44.0476
R14187 ringtest_0.x4.clknet_1_0__leaf_clk.n14 ringtest_0.x4.clknet_1_0__leaf_clk.n12 44.0476
R14188 ringtest_0.x4.clknet_1_0__leaf_clk.n6 ringtest_0.x4.clknet_1_0__leaf_clk.t8 40.0005
R14189 ringtest_0.x4.clknet_1_0__leaf_clk.n6 ringtest_0.x4.clknet_1_0__leaf_clk.t11 40.0005
R14190 ringtest_0.x4.clknet_1_0__leaf_clk.n7 ringtest_0.x4.clknet_1_0__leaf_clk.t13 40.0005
R14191 ringtest_0.x4.clknet_1_0__leaf_clk.n7 ringtest_0.x4.clknet_1_0__leaf_clk.t15 40.0005
R14192 ringtest_0.x4.clknet_1_0__leaf_clk.n9 ringtest_0.x4.clknet_1_0__leaf_clk.t10 40.0005
R14193 ringtest_0.x4.clknet_1_0__leaf_clk.n9 ringtest_0.x4.clknet_1_0__leaf_clk.t12 40.0005
R14194 ringtest_0.x4.clknet_1_0__leaf_clk.n11 ringtest_0.x4.clknet_1_0__leaf_clk.t14 40.0005
R14195 ringtest_0.x4.clknet_1_0__leaf_clk.n11 ringtest_0.x4.clknet_1_0__leaf_clk.t9 40.0005
R14196 ringtest_0.x4.clknet_1_0__leaf_clk.n13 ringtest_0.x4.clknet_1_0__leaf_clk.t1 40.0005
R14197 ringtest_0.x4.clknet_1_0__leaf_clk.n13 ringtest_0.x4.clknet_1_0__leaf_clk.t4 40.0005
R14198 ringtest_0.x4.clknet_1_0__leaf_clk.n15 ringtest_0.x4.clknet_1_0__leaf_clk.t6 40.0005
R14199 ringtest_0.x4.clknet_1_0__leaf_clk.n15 ringtest_0.x4.clknet_1_0__leaf_clk.t7 40.0005
R14200 ringtest_0.x4.clknet_1_0__leaf_clk.n17 ringtest_0.x4.clknet_1_0__leaf_clk.t3 40.0005
R14201 ringtest_0.x4.clknet_1_0__leaf_clk.n17 ringtest_0.x4.clknet_1_0__leaf_clk.t5 40.0005
R14202 ringtest_0.x4.clknet_1_0__leaf_clk.n19 ringtest_0.x4.clknet_1_0__leaf_clk.t0 40.0005
R14203 ringtest_0.x4.clknet_1_0__leaf_clk.n19 ringtest_0.x4.clknet_1_0__leaf_clk.t2 40.0005
R14204 ringtest_0.x4.clknet_1_0__leaf_clk.n27 ringtest_0.x4.clknet_1_0__leaf_clk.n25 32.0005
R14205 ringtest_0.x4.clknet_1_0__leaf_clk.n29 ringtest_0.x4.clknet_1_0__leaf_clk.n27 32.0005
R14206 ringtest_0.x4.clknet_1_0__leaf_clk.n32 ringtest_0.x4.clknet_1_0__leaf_clk.n22 32.0005
R14207 ringtest_0.x4.clknet_1_0__leaf_clk.n32 ringtest_0.x4.clknet_1_0__leaf_clk.n31 32.0005
R14208 ringtest_0.x4.clknet_1_0__leaf_clk.n31 ringtest_0.x4.clknet_1_0__leaf_clk.n29 31.2005
R14209 ringtest_0.x4.clknet_1_0__leaf_clk.n35 ringtest_0.x4.clknet_1_0__leaf_clk.n34 28.6283
R14210 ringtest_0.x4.clknet_1_0__leaf_clk.n3 ringtest_0.x4.clknet_1_0__leaf_clk 28.0697
R14211 ringtest_0.x4.clknet_1_0__leaf_clk.n23 ringtest_0.x4.clknet_1_0__leaf_clk.t19 27.5805
R14212 ringtest_0.x4.clknet_1_0__leaf_clk.n23 ringtest_0.x4.clknet_1_0__leaf_clk.t22 27.5805
R14213 ringtest_0.x4.clknet_1_0__leaf_clk.n24 ringtest_0.x4.clknet_1_0__leaf_clk.t24 27.5805
R14214 ringtest_0.x4.clknet_1_0__leaf_clk.n24 ringtest_0.x4.clknet_1_0__leaf_clk.t26 27.5805
R14215 ringtest_0.x4.clknet_1_0__leaf_clk.n26 ringtest_0.x4.clknet_1_0__leaf_clk.t21 27.5805
R14216 ringtest_0.x4.clknet_1_0__leaf_clk.n26 ringtest_0.x4.clknet_1_0__leaf_clk.t23 27.5805
R14217 ringtest_0.x4.clknet_1_0__leaf_clk.n28 ringtest_0.x4.clknet_1_0__leaf_clk.t25 27.5805
R14218 ringtest_0.x4.clknet_1_0__leaf_clk.n28 ringtest_0.x4.clknet_1_0__leaf_clk.t20 27.5805
R14219 ringtest_0.x4.clknet_1_0__leaf_clk.n4 ringtest_0.x4.clknet_1_0__leaf_clk.t30 27.5805
R14220 ringtest_0.x4.clknet_1_0__leaf_clk.n4 ringtest_0.x4.clknet_1_0__leaf_clk.t16 27.5805
R14221 ringtest_0.x4.clknet_1_0__leaf_clk.n5 ringtest_0.x4.clknet_1_0__leaf_clk.t27 27.5805
R14222 ringtest_0.x4.clknet_1_0__leaf_clk.n5 ringtest_0.x4.clknet_1_0__leaf_clk.t29 27.5805
R14223 ringtest_0.x4.clknet_1_0__leaf_clk.n33 ringtest_0.x4.clknet_1_0__leaf_clk.t17 27.5805
R14224 ringtest_0.x4.clknet_1_0__leaf_clk.n33 ringtest_0.x4.clknet_1_0__leaf_clk.t18 27.5805
R14225 ringtest_0.x4.clknet_1_0__leaf_clk.n30 ringtest_0.x4.clknet_1_0__leaf_clk.t28 27.5805
R14226 ringtest_0.x4.clknet_1_0__leaf_clk.n30 ringtest_0.x4.clknet_1_0__leaf_clk.t31 27.5805
R14227 ringtest_0.x4.clknet_1_0__leaf_clk.n43 ringtest_0.x4.clknet_1_0__leaf_clk.n42 27.3319
R14228 ringtest_0.x4.clknet_1_0__leaf_clk.n40 ringtest_0.x4.clknet_1_0__leaf_clk.n39 21.4985
R14229 ringtest_0.x4.clknet_1_0__leaf_clk.n3 ringtest_0.x4.clknet_1_0__leaf_clk.n1 21.401
R14230 ringtest_0.x4.clknet_1_0__leaf_clk.n34 ringtest_0.x4.clknet_1_0__leaf_clk.n32 14.0898
R14231 ringtest_0.x4.clknet_1_0__leaf_clk.n20 ringtest_0.x4.clknet_1_0__leaf_clk.n18 13.177
R14232 ringtest_0.x4.clknet_1_0__leaf_clk.n40 ringtest_0.x4.clknet_1_0__leaf_clk.n37 11.0654
R14233 ringtest_0.x4.clknet_1_0__leaf_clk.n22 ringtest_0.x4.clknet_1_0__leaf_clk.n21 10.4484
R14234 ringtest_0.x4.clknet_1_0__leaf_clk.n43 ringtest_0.x4.clknet_1_0__leaf_clk.n40 7.18319
R14235 ringtest_0.x4.clknet_1_0__leaf_clk.n35 ringtest_0.x4.clknet_1_0__leaf_clk.n3 5.63649
R14236 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n20 3.13183
R14237 ringtest_0.x4.clknet_1_0__leaf_clk.n37 ringtest_0.x4.clknet_1_0__leaf_clk 3.10907
R14238 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n43 2.66671
R14239 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n35 2.66671
R14240 ringtest_0.x4.clknet_1_0__leaf_clk.n42 ringtest_0.x4.clknet_1_0__leaf_clk 2.01193
R14241 ringtest_0.x4.clknet_1_0__leaf_clk.n21 ringtest_0.x4.clknet_1_0__leaf_clk 1.75844
R14242 ringtest_0.x4.clknet_1_0__leaf_clk.n39 ringtest_0.x4.clknet_1_0__leaf_clk 1.67435
R14243 ringtest_0.x4.clknet_1_0__leaf_clk.n1 ringtest_0.x4.clknet_1_0__leaf_clk 1.37896
R14244 ringtest_0.x4.clknet_1_0__leaf_clk.n20 ringtest_0.x4.clknet_1_0__leaf_clk 0.604792
R14245 ringtest_0.counter3.n0 ringtest_0.counter3.t3 368.521
R14246 ringtest_0.counter3.n1 ringtest_0.counter3.t2 216.155
R14247 ringtest_0.counter3.n1 ringtest_0.counter3 78.8791
R14248 ringtest_0.counter3.n4 ringtest_0.counter3.t1 26.3998
R14249 ringtest_0.counter3.n4 ringtest_0.counter3.t0 23.5483
R14250 ringtest_0.counter3.n3 ringtest_0.counter3.n2 17.5689
R14251 ringtest_0.counter3.n5 ringtest_0.counter3.t5 12.9693
R14252 ringtest_0.counter3.n5 ringtest_0.counter3.t4 10.8444
R14253 ringtest_0.counter3 ringtest_0.counter3.n0 10.5563
R14254 ringtest_0.counter3.n0 ringtest_0.counter3 5.48477
R14255 ringtest_0.counter3.n2 ringtest_0.counter3 4.18512
R14256 ringtest_0.counter3.n6 ringtest_0.counter3.n4 3.06895
R14257 ringtest_0.counter3.n6 ringtest_0.counter3.n5 2.14822
R14258 ringtest_0.counter3.n3 ringtest_0.counter3 1.28175
R14259 ringtest_0.counter3 ringtest_0.counter3.n6 1.25828
R14260 ringtest_0.counter3.n2 ringtest_0.counter3.n1 0.985115
R14261 ringtest_0.counter3 ringtest_0.counter3.n3 0.688
R14262 muxtest_0.x1.x3.GP2.n3 muxtest_0.x1.x3.GP2.t4 450.938
R14263 muxtest_0.x1.x3.GP2.n2 muxtest_0.x1.x3.GP2.t7 450.938
R14264 muxtest_0.x1.x3.GP2.n3 muxtest_0.x1.x3.GP2.t5 445.666
R14265 muxtest_0.x1.x3.GP2.n2 muxtest_0.x1.x3.GP2.t6 445.666
R14266 muxtest_0.x1.x3.GP2.n6 muxtest_0.x1.x3.GP2.n5 195.958
R14267 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n0 96.8352
R14268 muxtest_0.x1.x3.GP2.n5 muxtest_0.x1.x3.GP2.t2 26.5955
R14269 muxtest_0.x1.x3.GP2.n5 muxtest_0.x1.x3.GP2.t3 26.5955
R14270 muxtest_0.x1.x3.GP2.n0 muxtest_0.x1.x3.GP2.t0 24.9236
R14271 muxtest_0.x1.x3.GP2.n0 muxtest_0.x1.x3.GP2.t1 24.9236
R14272 muxtest_0.x1.x3.GP2.n4 muxtest_0.x1.x3.GP2 14.8953
R14273 muxtest_0.x1.x3.GP2.n7 muxtest_0.x1.x3.GP2.n6 13.0077
R14274 muxtest_0.x1.x3.GP2.n6 muxtest_0.x1.x3.GP2 11.8741
R14275 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n1 11.2645
R14276 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n4 8.64182
R14277 muxtest_0.x1.x3.GP2.n1 muxtest_0.x1.x3.GP2 6.1445
R14278 muxtest_0.x1.x3.GP2.n4 muxtest_0.x1.x3.GP2 5.75481
R14279 muxtest_0.x1.x3.GP2.n1 muxtest_0.x1.x3.GP2 4.65505
R14280 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n2 3.12276
R14281 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n3 2.94361
R14282 muxtest_0.x1.x3.GP2.n7 muxtest_0.x1.x3.GP2 2.0485
R14283 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n7 1.55202
R14284 muxtest_0.R5R6.n0 muxtest_0.R5R6.t0 26.3998
R14285 muxtest_0.R5R6.n0 muxtest_0.R5R6.t1 23.5483
R14286 muxtest_0.R5R6.n1 muxtest_0.R5R6.t4 12.9758
R14287 muxtest_0.R5R6.n1 muxtest_0.R5R6.t5 10.8618
R14288 muxtest_0.R5R6.n4 muxtest_0.R5R6.t3 10.55
R14289 muxtest_0.R5R6.n2 muxtest_0.R5R6.n0 3.06895
R14290 muxtest_0.R5R6.n2 muxtest_0.R5R6.n1 2.14822
R14291 muxtest_0.R5R6.n3 muxtest_0.R5R6.n2 1.12636
R14292 muxtest_0.R5R6.n4 muxtest_0.R5R6.t2 1.11543
R14293 muxtest_0.R5R6 muxtest_0.R5R6.n4 0.694875
R14294 muxtest_0.R5R6 muxtest_0.R5R6.n3 0.132418
R14295 muxtest_0.R5R6.n3 muxtest_0.R5R6 0.0655
R14296 ringtest_0.x4._16_.n12 ringtest_0.x4._16_.t1 339.418
R14297 ringtest_0.x4._16_ ringtest_0.x4._16_.t0 269.426
R14298 ringtest_0.x4._16_.n1 ringtest_0.x4._16_.t7 264.029
R14299 ringtest_0.x4._16_ ringtest_0.x4._16_.n5 241.976
R14300 ringtest_0.x4._16_.n3 ringtest_0.x4._16_.t3 241.536
R14301 ringtest_0.x4._16_.n5 ringtest_0.x4._16_.t8 241.536
R14302 ringtest_0.x4._16_.n1 ringtest_0.x4._16_.t2 206.19
R14303 ringtest_0.x4._16_.n4 ringtest_0.x4._16_.n3 171.332
R14304 ringtest_0.x4._16_.n3 ringtest_0.x4._16_.t9 169.237
R14305 ringtest_0.x4._16_.n5 ringtest_0.x4._16_.t4 169.237
R14306 ringtest_0.x4._16_.n2 ringtest_0.x4._16_.n1 160.96
R14307 ringtest_0.x4._16_.n9 ringtest_0.x4._16_.n8 153.165
R14308 ringtest_0.x4._16_.n8 ringtest_0.x4._16_.t6 144.548
R14309 ringtest_0.x4._16_.n8 ringtest_0.x4._16_.t5 128.482
R14310 ringtest_0.x4._16_.n7 ringtest_0.x4._16_.n2 21.45
R14311 ringtest_0.x4._16_.n7 ringtest_0.x4._16_.n6 16.7975
R14312 ringtest_0.x4._16_.n10 ringtest_0.x4._16_ 15.8161
R14313 ringtest_0.x4._16_.n11 ringtest_0.x4._16_.n10 14.0946
R14314 ringtest_0.x4._16_ ringtest_0.x4._16_.n0 11.2645
R14315 ringtest_0.x4._16_ ringtest_0.x4._16_.n9 9.55788
R14316 ringtest_0.x4._16_.n6 ringtest_0.x4._16_ 6.4005
R14317 ringtest_0.x4._16_.n0 ringtest_0.x4._16_ 6.1445
R14318 ringtest_0.x4._16_.n2 ringtest_0.x4._16_ 5.4405
R14319 ringtest_0.x4._16_.n0 ringtest_0.x4._16_ 4.63498
R14320 ringtest_0.x4._16_.n4 ringtest_0.x4._16_ 4.44132
R14321 ringtest_0.x4._16_.n11 ringtest_0.x4._16_ 4.3525
R14322 ringtest_0.x4._16_.n13 ringtest_0.x4._16_.n12 4.0914
R14323 ringtest_0.x4._16_ ringtest_0.x4._16_.n13 3.61789
R14324 ringtest_0.x4._16_.n9 ringtest_0.x4._16_ 3.29747
R14325 ringtest_0.x4._16_.n13 ringtest_0.x4._16_.n11 2.3045
R14326 ringtest_0.x4._16_.n12 ringtest_0.x4._16_ 1.74382
R14327 ringtest_0.x4._16_.n6 ringtest_0.x4._16_.n4 1.50638
R14328 ringtest_0.x4._16_.n10 ringtest_0.x4._16_.n7 1.38649
R14329 muxtest_0.x2.x2.GP2.n2 muxtest_0.x2.x2.GP2.t4 450.938
R14330 muxtest_0.x2.x2.GP2.n2 muxtest_0.x2.x2.GP2.t5 445.666
R14331 muxtest_0.x2.x2.GP2.n4 muxtest_0.x2.x2.GP2.n3 195.958
R14332 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n0 96.8352
R14333 muxtest_0.x2.x2.GP2.n3 muxtest_0.x2.x2.GP2.t3 26.5955
R14334 muxtest_0.x2.x2.GP2.n3 muxtest_0.x2.x2.GP2.t2 26.5955
R14335 muxtest_0.x2.x2.GP2.n0 muxtest_0.x2.x2.GP2.t0 24.9236
R14336 muxtest_0.x2.x2.GP2.n0 muxtest_0.x2.x2.GP2.t1 24.9236
R14337 muxtest_0.x2.x2.GP2.n5 muxtest_0.x2.x2.GP2.n4 13.0077
R14338 muxtest_0.x2.x2.GP2.n4 muxtest_0.x2.x2.GP2 11.995
R14339 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n1 11.2645
R14340 muxtest_0.x2.x2.GP2.n1 muxtest_0.x2.x2.GP2 6.1445
R14341 muxtest_0.x2.x2.GP2.n1 muxtest_0.x2.x2.GP2 4.65505
R14342 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n2 3.12839
R14343 muxtest_0.x2.x2.GP2.n5 muxtest_0.x2.x2.GP2 2.0485
R14344 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n5 1.55202
R14345 muxtest_0.R6R7.n0 muxtest_0.R6R7.t1 26.3998
R14346 muxtest_0.R6R7.n0 muxtest_0.R6R7.t0 23.5483
R14347 muxtest_0.R6R7.n4 muxtest_0.R6R7.t4 17.4454
R14348 muxtest_0.R6R7.n1 muxtest_0.R6R7.t3 12.9758
R14349 muxtest_0.R6R7.n1 muxtest_0.R6R7.t2 10.8618
R14350 muxtest_0.R6R7.n4 muxtest_0.R6R7.t5 10.5739
R14351 muxtest_0.R6R7.n2 muxtest_0.R6R7.n0 3.06895
R14352 muxtest_0.R6R7.n2 muxtest_0.R6R7.n1 2.14822
R14353 muxtest_0.R6R7.n3 muxtest_0.R6R7.n2 1.12636
R14354 muxtest_0.R6R7.n5 muxtest_0.R6R7 1.11925
R14355 muxtest_0.R6R7.n5 muxtest_0.R6R7.n4 0.370193
R14356 muxtest_0.R6R7 muxtest_0.R6R7.n3 0.138152
R14357 muxtest_0.R6R7.n5 muxtest_0.R6R7 0.073
R14358 muxtest_0.R6R7.n3 muxtest_0.R6R7 0.0655
R14359 muxtest_0.R6R7 muxtest_0.R6R7.n5 0.04925
R14360 ua[0].n6 ua[0].t3 26.3998
R14361 ua[0].n0 ua[0].t5 26.3998
R14362 ua[0].n6 ua[0].t2 23.5483
R14363 ua[0].n0 ua[0].t6 23.5483
R14364 ua[0].n7 ua[0].t0 12.9758
R14365 ua[0].n1 ua[0].t7 12.9758
R14366 ua[0].n5 ua[0] 12.8371
R14367 ua[0].n7 ua[0].t1 10.8618
R14368 ua[0].n1 ua[0].t8 10.8618
R14369 ua[0].n4 ua[0].t4 10.5739
R14370 ua[0].n8 ua[0].n6 3.06895
R14371 ua[0].n2 ua[0].n0 3.06895
R14372 ua[0].n8 ua[0].n7 2.14822
R14373 ua[0].n2 ua[0].n1 2.14822
R14374 ua[0].n4 ua[0] 1.39577
R14375 ua[0].n9 ua[0].n8 1.12636
R14376 ua[0].n3 ua[0].n2 1.12636
R14377 ua[0].n5 ua[0].n4 0.545106
R14378 ua[0] ua[0].n9 0.138152
R14379 ua[0] ua[0].n3 0.134513
R14380 ua[0].n9 ua[0] 0.0655
R14381 ua[0].n3 ua[0] 0.0655
R14382 ua[0] ua[0].n5 0.0579534
R14383 ua[0].n5 ua[0] 0.0532872
R14384 muxtest_0.R7R8.n5 muxtest_0.R7R8.t5 26.3998
R14385 muxtest_0.R7R8.n0 muxtest_0.R7R8.t4 26.3998
R14386 muxtest_0.R7R8.n5 muxtest_0.R7R8.t6 23.5483
R14387 muxtest_0.R7R8.n0 muxtest_0.R7R8.t3 23.5483
R14388 muxtest_0.R7R8.n6 muxtest_0.R7R8.t8 12.9758
R14389 muxtest_0.R7R8.n1 muxtest_0.R7R8.t1 12.9758
R14390 muxtest_0.R7R8.n6 muxtest_0.R7R8.t7 10.8618
R14391 muxtest_0.R7R8.n1 muxtest_0.R7R8.t0 10.8618
R14392 muxtest_0.R7R8.n4 muxtest_0.R7R8.t9 10.5709
R14393 muxtest_0.R7R8.n9 muxtest_0.R7R8 8.65896
R14394 muxtest_0.R7R8.n7 muxtest_0.R7R8.n5 3.06895
R14395 muxtest_0.R7R8.n2 muxtest_0.R7R8.n0 3.06895
R14396 muxtest_0.R7R8.n7 muxtest_0.R7R8.n6 2.14822
R14397 muxtest_0.R7R8.n2 muxtest_0.R7R8.n1 2.14822
R14398 muxtest_0.R7R8.n8 muxtest_0.R7R8.n7 1.12636
R14399 muxtest_0.R7R8.n3 muxtest_0.R7R8.n2 1.12636
R14400 muxtest_0.R7R8.n4 muxtest_0.R7R8.t2 1.01856
R14401 muxtest_0.R7R8 muxtest_0.R7R8.n9 0.32175
R14402 muxtest_0.R7R8.n9 muxtest_0.R7R8.n4 0.230945
R14403 muxtest_0.R7R8 muxtest_0.R7R8.n3 0.148615
R14404 muxtest_0.R7R8 muxtest_0.R7R8.n8 0.134513
R14405 muxtest_0.R7R8.n8 muxtest_0.R7R8 0.0655
R14406 muxtest_0.R7R8.n3 muxtest_0.R7R8 0.0655
R14407 ui_in[3].n18 ui_in[3].t0 327.99
R14408 ui_in[3].n5 ui_in[3].t19 327.99
R14409 ui_in[3].n22 ui_in[3].t4 293.969
R14410 ui_in[3].n9 ui_in[3].t17 293.969
R14411 ui_in[3].n16 ui_in[3].t11 261.887
R14412 ui_in[3].n3 ui_in[3].t10 261.887
R14413 ui_in[3].n13 ui_in[3].t5 212.081
R14414 ui_in[3].n14 ui_in[3].t8 212.081
R14415 ui_in[3].n0 ui_in[3].t18 212.081
R14416 ui_in[3].n1 ui_in[3].t3 212.081
R14417 ui_in[3].n18 ui_in[3].t14 199.457
R14418 ui_in[3].n5 ui_in[3].t9 199.457
R14419 ui_in[3].n15 ui_in[3].n14 183.185
R14420 ui_in[3].n2 ui_in[3].n1 183.185
R14421 ui_in[3].n16 ui_in[3].t7 155.847
R14422 ui_in[3].n3 ui_in[3].t6 155.847
R14423 ui_in[3] ui_in[3].n22 154.065
R14424 ui_in[3] ui_in[3].n9 154.065
R14425 ui_in[3].n17 ui_in[3].n16 153.506
R14426 ui_in[3].n4 ui_in[3].n3 153.506
R14427 ui_in[3].n19 ui_in[3].n18 152
R14428 ui_in[3].n6 ui_in[3].n5 152
R14429 ui_in[3].n13 ui_in[3].t13 139.78
R14430 ui_in[3].n14 ui_in[3].t16 139.78
R14431 ui_in[3].n0 ui_in[3].t2 139.78
R14432 ui_in[3].n1 ui_in[3].t12 139.78
R14433 ui_in[3].n22 ui_in[3].t1 138.338
R14434 ui_in[3].n9 ui_in[3].t15 138.338
R14435 ui_in[3].n14 ui_in[3].n13 61.346
R14436 ui_in[3].n1 ui_in[3].n0 61.346
R14437 ui_in[3].n26 ui_in[3] 35.166
R14438 ui_in[3].n23 ui_in[3] 13.4199
R14439 ui_in[3].n10 ui_in[3] 13.4199
R14440 ui_in[3].n26 ui_in[3] 12.2088
R14441 ui_in[3].n24 ui_in[3].n21 11.7395
R14442 ui_in[3].n11 ui_in[3].n8 11.7395
R14443 ui_in[3].n25 ui_in[3].n24 11.5949
R14444 ui_in[3].n12 ui_in[3].n11 11.5949
R14445 ui_in[3].n21 ui_in[3].n17 10.4004
R14446 ui_in[3].n8 ui_in[3].n4 10.4004
R14447 ui_in[3].n25 ui_in[3].n15 9.68118
R14448 ui_in[3].n12 ui_in[3].n2 9.68118
R14449 ui_in[3].n19 ui_in[3] 9.6005
R14450 ui_in[3].n6 ui_in[3] 9.6005
R14451 ui_in[3].n15 ui_in[3] 5.8885
R14452 ui_in[3].n2 ui_in[3] 5.8885
R14453 ui_in[3].n23 ui_in[3] 5.57469
R14454 ui_in[3].n10 ui_in[3] 5.57469
R14455 ui_in[3].n21 ui_in[3].n20 4.6505
R14456 ui_in[3].n24 ui_in[3].n23 4.6505
R14457 ui_in[3].n8 ui_in[3].n7 4.6505
R14458 ui_in[3].n11 ui_in[3].n10 4.6505
R14459 ui_in[3].n20 ui_in[3].n19 2.98717
R14460 ui_in[3].n7 ui_in[3].n6 2.98717
R14461 ui_in[3].n17 ui_in[3] 2.82403
R14462 ui_in[3].n4 ui_in[3] 2.82403
R14463 ui_in[3].n20 ui_in[3] 1.9205
R14464 ui_in[3].n7 ui_in[3] 1.9205
R14465 ui_in[3] ui_in[3].n25 0.559212
R14466 ui_in[3] ui_in[3].n12 0.559212
R14467 ui_in[3] ui_in[3].n26 0.47425
R14468 ringtest_0.x3.x2.GP1.n2 ringtest_0.x3.x2.GP1.t5 450.938
R14469 ringtest_0.x3.x2.GP1.n2 ringtest_0.x3.x2.GP1.t4 445.666
R14470 ringtest_0.x3.x2.GP1.n4 ringtest_0.x3.x2.GP1.n3 195.832
R14471 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n0 96.8352
R14472 ringtest_0.x3.x2.GP1.n3 ringtest_0.x3.x2.GP1.t3 26.5955
R14473 ringtest_0.x3.x2.GP1.n3 ringtest_0.x3.x2.GP1.t2 26.5955
R14474 ringtest_0.x3.x2.GP1.n0 ringtest_0.x3.x2.GP1.t1 24.9236
R14475 ringtest_0.x3.x2.GP1.n0 ringtest_0.x3.x2.GP1.t0 24.9236
R14476 ringtest_0.x3.x2.GP1.n5 ringtest_0.x3.x2.GP1.n4 13.1346
R14477 ringtest_0.x3.x2.GP1.n4 ringtest_0.x3.x2.GP1 12.2007
R14478 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n1 11.2645
R14479 ringtest_0.x3.x2.GP1.n1 ringtest_0.x3.x2.GP1 6.1445
R14480 ringtest_0.x3.x2.GP1.n1 ringtest_0.x3.x2.GP1 4.65505
R14481 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n2 3.07707
R14482 ringtest_0.x3.x2.GP1.n5 ringtest_0.x3.x2.GP1 2.0485
R14483 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n5 1.55202
R14484 ringtest_0.ring_out.n0 ringtest_0.ring_out.t13 844.321
R14485 ringtest_0.ring_out.n0 ringtest_0.ring_out.t12 354.322
R14486 ringtest_0.ring_out.n3 ringtest_0.ring_out.n1 243.68
R14487 ringtest_0.ring_out.n8 ringtest_0.ring_out.t10 212.081
R14488 ringtest_0.ring_out.n7 ringtest_0.ring_out.t11 212.081
R14489 ringtest_0.ring_out.n5 ringtest_0.ring_out.n4 206.249
R14490 ringtest_0.ring_out.n3 ringtest_0.ring_out.n2 205.28
R14491 ringtest_0.ring_out.n9 ringtest_0.ring_out.n8 184.806
R14492 ringtest_0.ring_out.n8 ringtest_0.ring_out.t14 139.78
R14493 ringtest_0.ring_out.n7 ringtest_0.ring_out.t15 139.78
R14494 ringtest_0.ring_out.n8 ringtest_0.ring_out.n7 61.346
R14495 ringtest_0.ring_out.n1 ringtest_0.ring_out.t2 26.5955
R14496 ringtest_0.ring_out.n1 ringtest_0.ring_out.t1 26.5955
R14497 ringtest_0.ring_out.n2 ringtest_0.ring_out.t7 26.5955
R14498 ringtest_0.ring_out.n2 ringtest_0.ring_out.t8 26.5955
R14499 ringtest_0.ring_out.n11 ringtest_0.ring_out.t5 26.3998
R14500 ringtest_0.ring_out ringtest_0.ring_out.n3 24.9955
R14501 ringtest_0.ring_out.n4 ringtest_0.ring_out.t9 24.9236
R14502 ringtest_0.ring_out.n4 ringtest_0.ring_out.t0 24.9236
R14503 ringtest_0.ring_out.n11 ringtest_0.ring_out.t6 23.5483
R14504 ringtest_0.ring_out.n10 ringtest_0.ring_out.n9 21.363
R14505 ringtest_0.ring_out ringtest_0.ring_out.n5 14.8576
R14506 ringtest_0.ring_out.n12 ringtest_0.ring_out.t4 12.9758
R14507 ringtest_0.ring_out.n6 ringtest_0.ring_out 10.9719
R14508 ringtest_0.ring_out.n12 ringtest_0.ring_out.t3 10.8618
R14509 ringtest_0.ring_out.n10 ringtest_0.ring_out.n6 9.53262
R14510 ringtest_0.ring_out.n6 ringtest_0.ring_out 4.57193
R14511 ringtest_0.ring_out.n13 ringtest_0.ring_out.n11 3.06895
R14512 ringtest_0.ring_out.n9 ringtest_0.ring_out 2.32777
R14513 ringtest_0.ring_out.n13 ringtest_0.ring_out.n12 2.14822
R14514 ringtest_0.ring_out ringtest_0.ring_out.n13 1.12636
R14515 ringtest_0.ring_out.n5 ringtest_0.ring_out 0.686214
R14516 ringtest_0.ring_out ringtest_0.ring_out.n10 0.631142
R14517 ringtest_0.ring_out ringtest_0.ring_out.n0 0.354518
R14518 ringtest_0.x3.x2.GP2.n2 ringtest_0.x3.x2.GP2.t4 450.938
R14519 ringtest_0.x3.x2.GP2.n2 ringtest_0.x3.x2.GP2.t5 445.666
R14520 ringtest_0.x3.x2.GP2.n4 ringtest_0.x3.x2.GP2.n3 195.958
R14521 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n0 96.8352
R14522 ringtest_0.x3.x2.GP2.n3 ringtest_0.x3.x2.GP2.t3 26.5955
R14523 ringtest_0.x3.x2.GP2.n3 ringtest_0.x3.x2.GP2.t2 26.5955
R14524 ringtest_0.x3.x2.GP2.n0 ringtest_0.x3.x2.GP2.t1 24.9236
R14525 ringtest_0.x3.x2.GP2.n0 ringtest_0.x3.x2.GP2.t0 24.9236
R14526 ringtest_0.x3.x2.GP2.n5 ringtest_0.x3.x2.GP2.n4 13.0077
R14527 ringtest_0.x3.x2.GP2.n4 ringtest_0.x3.x2.GP2 11.995
R14528 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n1 11.2645
R14529 ringtest_0.x3.x2.GP2.n1 ringtest_0.x3.x2.GP2 6.1445
R14530 ringtest_0.x3.x2.GP2.n1 ringtest_0.x3.x2.GP2 4.65505
R14531 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n2 3.12839
R14532 ringtest_0.x3.x2.GP2.n5 ringtest_0.x3.x2.GP2 2.0485
R14533 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n5 1.55202
R14534 muxtest_0.x2.x2.GP4.n2 muxtest_0.x2.x2.GP4.t4 450.938
R14535 muxtest_0.x2.x2.GP4.n2 muxtest_0.x2.x2.GP4.t5 445.666
R14536 muxtest_0.x2.x2.GP4.n5 muxtest_0.x2.x2.GP4.n4 208.965
R14537 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n0 96.8352
R14538 muxtest_0.x2.x2.GP4.n4 muxtest_0.x2.x2.GP4.t3 26.5955
R14539 muxtest_0.x2.x2.GP4.n4 muxtest_0.x2.x2.GP4.t2 26.5955
R14540 muxtest_0.x2.x2.GP4.n0 muxtest_0.x2.x2.GP4.t1 24.9236
R14541 muxtest_0.x2.x2.GP4.n0 muxtest_0.x2.x2.GP4.t0 24.9236
R14542 muxtest_0.x2.x1.gpo3 muxtest_0.x2.x2.x4.GP 16.5032
R14543 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n3 10.2405
R14544 muxtest_0.x2.x2.GP4.n3 muxtest_0.x2.x1.gpo3 7.76481
R14545 muxtest_0.x2.x2.GP4.n1 muxtest_0.x2.x1.x14.Y 6.1445
R14546 muxtest_0.x2.x2.GP4.n1 muxtest_0.x2.x1.x14.Y 4.65505
R14547 muxtest_0.x2.x2.x4.GP muxtest_0.x2.x2.GP4.n2 2.95993
R14548 muxtest_0.x2.x2.GP4.n5 muxtest_0.x2.x1.x14.Y 2.0485
R14549 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n5 1.55202
R14550 muxtest_0.x2.x2.GP4.n3 muxtest_0.x2.x2.GP4.n1 1.0245
R14551 muxtest_0.R4R5.n0 muxtest_0.R4R5.t1 26.3998
R14552 muxtest_0.R4R5.n0 muxtest_0.R4R5.t2 23.5483
R14553 muxtest_0.R4R5.n1 muxtest_0.R4R5.t5 12.9758
R14554 muxtest_0.R4R5.n1 muxtest_0.R4R5.t4 10.8618
R14555 muxtest_0.R4R5.n4 muxtest_0.R4R5.t0 10.8231
R14556 muxtest_0.R4R5.n4 muxtest_0.R4R5.t3 10.5739
R14557 muxtest_0.R4R5.n2 muxtest_0.R4R5.n0 3.06895
R14558 muxtest_0.R4R5.n2 muxtest_0.R4R5.n1 2.14822
R14559 muxtest_0.R4R5.n3 muxtest_0.R4R5.n2 1.12636
R14560 muxtest_0.R4R5 muxtest_0.R4R5.n4 0.790021
R14561 muxtest_0.R4R5 muxtest_0.R4R5.n3 0.134513
R14562 muxtest_0.R4R5.n3 muxtest_0.R4R5 0.0655
R14563 muxtest_0.R2R3.n0 muxtest_0.R2R3.t0 26.3998
R14564 muxtest_0.R2R3.n0 muxtest_0.R2R3.t1 23.5483
R14565 muxtest_0.R2R3.n1 muxtest_0.R2R3.t3 12.9758
R14566 muxtest_0.R2R3.n1 muxtest_0.R2R3.t2 10.8618
R14567 muxtest_0.R2R3.n4 muxtest_0.R2R3.t4 10.8167
R14568 muxtest_0.R2R3.n4 muxtest_0.R2R3.t5 10.5739
R14569 muxtest_0.R2R3.n2 muxtest_0.R2R3.n0 3.06895
R14570 muxtest_0.R2R3.n2 muxtest_0.R2R3.n1 2.14822
R14571 muxtest_0.R2R3.n3 muxtest_0.R2R3.n2 1.12636
R14572 muxtest_0.R2R3 muxtest_0.R2R3.n4 0.71627
R14573 muxtest_0.R2R3 muxtest_0.R2R3.n3 0.138152
R14574 muxtest_0.R2R3.n3 muxtest_0.R2R3 0.0655
R14575 ui_in[6].n0 ui_in[6].t0 212.081
R14576 ui_in[6].n1 ui_in[6].t1 212.081
R14577 ui_in[6] ui_in[6].n2 152.512
R14578 ui_in[6].n0 ui_in[6].t2 139.78
R14579 ui_in[6].n1 ui_in[6].t3 139.78
R14580 ui_in[6].n2 ui_in[6].n0 30.6732
R14581 ui_in[6].n2 ui_in[6].n1 30.6732
R14582 ui_in[6].n3 ui_in[6] 16.4378
R14583 ui_in[6] ui_in[6].n3 0.7505
R14584 ui_in[6].n3 ui_in[6] 0.0808571
R14585 ui_in[5].n0 ui_in[5].t0 260.322
R14586 ui_in[5].n0 ui_in[5].t1 175.169
R14587 ui_in[5].n1 ui_in[5].n0 153.13
R14588 ui_in[5].n3 ui_in[5] 19.5879
R14589 ui_in[5] ui_in[5].n1 9.86591
R14590 ui_in[5].n3 ui_in[5].n2 4.07076
R14591 ui_in[5].n1 ui_in[5] 3.2005
R14592 ui_in[5].n2 ui_in[5] 0.960321
R14593 ui_in[5].n2 ui_in[5] 0.392836
R14594 ui_in[5] ui_in[5].n3 0.0499792
C0 a_20318_32213# muxtest_0.x1.x3.GN4 0.134079f
C1 muxtest_0.x1.x3.GN2 a_19242_32347# 0.002395f
C2 ringtest_0.x4._24_ a_27065_5156# 0.012283f
C3 ringtest_0.x4._00_ a_22052_9116# 0.00938f
C4 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ui_in[3] 9.57e-20
C5 ringtest_0.x4.net7 a_27233_5058# 8.32e-20
C6 ringtest_0.x4.net1 a_21425_9686# 0.224922f
C7 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2 2.14737f
C8 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net6 0.323735f
C9 ringtest_0.ring_out ringtest_0.x3.x1.nSEL0 1.86e-21
C10 muxtest_0.x1.x3.GP3 ui_in[2] 1.6e-19
C11 a_23529_6422# ringtest_0.x4.net7 0.002934f
C12 ringtest_0.x4.clknet_1_1__leaf_clk a_24895_4790# 0.486375f
C13 ringtest_0.x4.net8 a_25393_5308# 0.084103f
C14 ringtest_0.x4._11_ a_24361_5340# 1.58e-19
C15 ringtest_0.x4._17_ a_23529_6422# 0.043588f
C16 a_21375_3867# VDPWR 0.272145f
C17 ringtest_0.x4.net10 ringtest_0.x4.net11 0.310558f
C18 a_16027_11759# ringtest_0.x3.x2.GP1 9.92e-19
C19 a_16203_12091# ringtest_0.x3.x2.GN3 0.048646f
C20 ringtest_0.x4._08_ a_24968_5308# 9.82e-20
C21 ringtest_0.x4._06_ ringtest_0.x4.net9 0.017291f
C22 a_16579_11759# ringtest_0.x3.x2.GN1 6.43e-20
C23 a_23809_4790# ringtest_0.x4._20_ 0.237238f
C24 ua[3] ui_in[4] 1.14709f
C25 ringtest_0.x4._11_ a_21395_6940# 0.055744f
C26 a_21509_4790# a_21948_5156# 0.273138f
C27 ringtest_0.x4._15_ a_22097_5334# 7.5e-20
C28 ringtest_0.x4.net6 a_24800_5334# 0.019975f
C29 ringtest_0.x4._03_ a_22116_4902# 0.006259f
C30 ringtest_0.x4._22_ a_27273_4220# 4.31e-19
C31 ringtest_0.x4._12_ a_22245_8054# 0.026119f
C32 muxtest_0.x1.x5.A muxtest_0.R7R8 4.52065f
C33 a_24527_5340# a_25168_5156# 7.62e-19
C34 a_24800_5334# a_24895_4790# 8.92e-19
C35 ringtest_0.x4._15_ ringtest_0.x4._16_ 0.656968f
C36 a_25393_5308# a_24729_4790# 0.002274f
C37 a_25977_4220# a_25975_3867# 0.01226f
C38 ringtest_0.x4.net7 ringtest_0.x4._06_ 0.141876f
C39 ringtest_0.x4.net7 a_24070_5852# 0.003377f
C40 ringtest_0.x4.clknet_0_clk a_25168_5156# 4.63e-19
C41 ringtest_0.x4._18_ a_23932_6128# 0.00112f
C42 ringtest_0.x4._17_ ringtest_0.x4._06_ 0.001225f
C43 muxtest_0.x1.x1.nSEL1 ui_in[1] 0.275603f
C44 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A 5.04e-19
C45 a_23879_6940# ringtest_0.x4._21_ 0.001038f
C46 ringtest_0.x4._16_ a_22541_5058# 1.37e-19
C47 a_26808_5308# a_26640_5334# 0.239923f
C48 a_26201_5340# a_27065_5334# 0.032244f
C49 a_23770_5308# a_23993_5654# 0.011458f
C50 a_26367_5340# a_27233_5308# 0.034054f
C51 ringtest_0.x4._17_ a_24070_5852# 0.062168f
C52 a_24968_5308# VDPWR 0.185172f
C53 ringtest_0.x4.net6 ringtest_0.x4._23_ 0.023006f
C54 a_24329_6640# a_24883_6800# 0.057611f
C55 a_24045_6654# a_24287_6422# 0.008508f
C56 ringtest_0.x4.net4 a_22457_5156# 8.77e-19
C57 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x5.GN 0.10521f
C58 muxtest_0.x2.x2.GP1 ua[2] 0.352897f
C59 a_24895_4790# a_26367_4790# 0.002814f
C60 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._03_ 0.00668f
C61 a_18662_32213# m2_18699_31802# 0.01297f
C62 muxtest_0.x2.x1.nSEL1 a_12977_24040# 4.08e-19
C63 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN2 0.209956f
C64 a_11845_23906# muxtest_0.x2.x2.GN1 0.12869f
C65 ringtest_0.x4.net10 ringtest_0.x4._09_ 0.081678f
C66 ringtest_0.counter7 ringtest_0.x4.net5 6.88e-20
C67 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR 0.636314f
C68 a_27233_5308# a_27065_5156# 7.04e-19
C69 a_22817_6146# ringtest_0.x4._06_ 1.81e-20
C70 a_25925_6788# VDPWR 0.455589f
C71 a_27065_5334# a_27233_5058# 7.04e-19
C72 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x1.nSEL1 0.352716f
C73 a_21395_6940# a_21785_5878# 5.49e-20
C74 a_21375_3867# ringtest_0.x4.counter[2] 4.98e-19
C75 a_22817_6146# a_24070_5852# 2.22e-20
C76 muxtest_0.x1.x5.A muxtest_0.R5R6 4.5214f
C77 uio_in[7] uio_in[6] 0.031023f
C78 ringtest_0.x4.net6 ringtest_0.x4._02_ 0.001309f
C79 ringtest_0.x4._11_ ringtest_0.x4._08_ 1.44e-20
C80 ringtest_0.x4.clknet_1_0__leaf_clk a_21939_8054# 3.8e-19
C81 a_15749_12123# VDPWR 9.25e-19
C82 ringtest_0.x4._22_ a_26201_4790# 4.68e-20
C83 muxtest_0.x2.x2.GN2 ua[0] 4.0283f
C84 a_19794_32347# muxtest_0.x1.x3.GP3 4.39e-19
C85 ringtest_0.x3.x2.GN3 m3_17036_9140# 0.001446f
C86 muxtest_0.x1.x5.A VDPWR 14.1646f
C87 ringtest_0.x4.net3 a_22021_4220# 0.002183f
C88 ringtest_0.x4.net7 a_26269_4612# 5.42e-19
C89 ringtest_0.x4._15_ a_26201_6788# 0.001194f
C90 ringtest_0.x4._11_ a_25336_4902# 0.039242f
C91 a_25925_6788# ringtest_0.x4._25_ 1.87e-19
C92 ringtest_0.x4._23_ a_27169_6641# 6.47e-19
C93 ringtest_0.x4.net11 a_27191_4790# 3e-19
C94 ringtest_0.x4._07_ a_25351_5712# 5.27e-19
C95 a_21675_9686# a_21465_9294# 3.08e-19
C96 a_19290_32287# muxtest_0.x1.x3.GN3 0.048646f
C97 ringtest_0.x4._02_ a_21055_5334# 0.01416f
C98 ringtest_0.counter7 a_21007_3867# 2.81e-20
C99 a_26749_6422# a_26808_4902# 1.02e-20
C100 a_26640_5156# a_26766_4790# 0.005525f
C101 a_19114_31955# VDPWR 0.164569f
C102 a_26555_4790# a_26735_5156# 0.001229f
C103 a_21233_5340# VDPWR 0.684183f
C104 a_21399_5340# a_22265_5308# 0.034054f
C105 a_21840_5308# a_21672_5334# 0.239923f
C106 ringtest_0.x4.net4 ringtest_0.x4._03_ 0.031989f
C107 ringtest_0.x4.net10 a_27659_4246# 0.003077f
C108 ringtest_0.ring_out ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.167117f
C109 muxtest_0.x2.x2.GN3 a_12977_24040# 0.001073f
C110 muxtest_0.x2.x2.GN2 a_13675_24012# 8.14e-21
C111 m2_11882_23495# VDPWR 0.139985f
C112 ringtest_0.x4.net8 a_24715_5334# 0.005878f
C113 ringtest_0.x4.net6 a_25593_5156# 4.38e-19
C114 ringtest_0.x4._15_ a_23467_4818# 7.85e-19
C115 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GN3 0.067465f
C116 ringtest_0.x4._11_ a_22223_5712# 6.78e-19
C117 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN4 0.001074f
C118 a_25364_5878# a_26808_5308# 0.006157f
C119 a_24045_6654# a_24329_6640# 0.030894f
C120 a_23949_6654# a_24336_6544# 0.034054f
C121 a_20492_32319# ui_in[0] 1.77e-19
C122 ringtest_0.x4._11_ VDPWR 5.18499f
C123 a_25336_4902# a_25761_5058# 1.28e-19
C124 a_24729_4790# a_25083_4790# 0.062224f
C125 a_24895_4790# a_25593_5156# 0.193199f
C126 a_19842_32287# ui_in[0] 0.279876f
C127 ringtest_0.x4.net4 a_23770_5308# 1.34e-19
C128 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN3 4.01e-20
C129 ringtest_0.x4.clknet_1_1__leaf_clk a_24895_5334# 0.002214f
C130 ringtest_0.x4._22_ a_27303_4246# 6.52e-20
C131 a_25975_3867# ringtest_0.x4.counter[9] 2.37e-20
C132 muxtest_0.R6R7 muxtest_0.R4R5 2.49e-19
C133 ringtest_0.x4._14_ a_22164_4362# 0.089653f
C134 a_25761_5058# VDPWR 0.400861f
C135 ringtest_0.x4.net8 a_25547_4612# 1.72e-20
C136 ringtest_0.x4._11_ a_23467_4584# 6.46e-19
C137 a_23879_6940# a_24968_5308# 8.05e-21
C138 ringtest_0.x4._11_ ringtest_0.x4._25_ 2.54e-20
C139 muxtest_0.x1.x3.GN1 muxtest_0.R2R3 2.55e-19
C140 a_25364_5878# a_26555_4790# 1.26e-19
C141 a_21675_4790# VDPWR 0.342267f
C142 ringtest_0.x4.net3 a_21561_8830# 0.006429f
C143 a_24536_6699# ringtest_0.x4._06_ 2.41e-19
C144 muxtest_0.x1.x3.GN1 ui_in[1] 0.312176f
C145 ringtest_0.x4.net1 ringtest_0.x4._11_ 0.002334f
C146 ringtest_0.x4.clknet_0_clk ringtest_0.x4._18_ 0.002702f
C147 a_24968_5308# a_25309_5334# 9.73e-19
C148 a_24800_5334# a_24895_5334# 0.007724f
C149 a_21561_9116# a_21852_8720# 1.53e-19
C150 a_21845_9116# a_21561_8830# 9.64e-20
C151 a_21852_9416# a_21845_8816# 3.36e-19
C152 a_24336_6544# a_24004_6128# 0.002652f
C153 a_24329_6640# a_24699_6200# 0.007926f
C154 ringtest_0.x4.net6 ringtest_0.x4._04_ 0.050232f
C155 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A 0.17253f
C156 a_23899_5654# VDPWR 5.6e-19
C157 a_26569_6422# ringtest_0.x4._24_ 0.095435f
C158 ringtest_0.x4.net2 a_21780_9142# 2.28e-19
C159 ringtest_0.x4._19_ a_24883_6800# 0.014678f
C160 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net6 6.56e-20
C161 ringtest_0.x3.nselect2 ui_in[3] 1.88e-19
C162 ringtest_0.ring_out ua[1] 4.51997f
C163 ringtest_0.x4.net2 a_21561_9116# 0.019416f
C164 ringtest_0.x4._09_ a_27191_4790# 0.001794f
C165 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN1 0.645006f
C166 muxtest_0.x1.x1.nSEL0 VDPWR 0.389106f
C167 ringtest_0.ring_out a_16755_12091# 2.55e-19
C168 a_24465_6800# ringtest_0.x4._15_ 2.35e-21
C169 ringtest_0.x4._09_ a_26808_4902# 0.039926f
C170 a_26201_4790# a_26640_5156# 0.273138f
C171 a_24763_6143# a_24527_5340# 0.003413f
C172 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP3 0.002437f
C173 a_21785_5878# VDPWR 0.6434f
C174 muxtest_0.x2.x1.nSEL0 a_13025_23980# 1.21e-20
C175 a_24045_6654# a_24317_4942# 5.98e-21
C176 ringtest_0.x4.clknet_0_clk a_24763_6143# 7.62e-19
C177 a_21951_5878# a_22265_5308# 0.003783f
C178 ringtest_0.x4.clknet_1_0__leaf_clk a_21055_5334# 1.21e-20
C179 a_24699_6200# a_24545_5878# 0.049785f
C180 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP1 1.16e-20
C181 a_22399_9142# VDPWR 0.080219f
C182 ringtest_0.x4.net9 a_26895_3867# 0.202772f
C183 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR 0.63819f
C184 ringtest_0.x4._11_ ringtest_0.x4._21_ 0.059807f
C185 muxtest_0.R7R8 ua[2] 4.51509f
C186 a_23949_6654# a_23899_5334# 2.76e-21
C187 ringtest_0.x4.clknet_1_1__leaf_clk a_24527_5340# 0.079788f
C188 muxtest_0.x1.x3.GN4 muxtest_0.R4R5 4.23588f
C189 muxtest_0.x2.x2.GP1 m3_13302_19985# 3.25e-21
C190 a_21852_8720# ringtest_0.x4._01_ 0.239739f
C191 ringtest_0.x4.net3 a_21049_8598# 0.042192f
C192 a_22052_8875# a_21981_8976# 0.239923f
C193 a_26367_5340# a_27149_5334# 6.32e-19
C194 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_1_1__leaf_clk 0.335671f
C195 muxtest_0.x1.x3.GN2 muxtest_0.R7R8 0.260757f
C196 a_25977_4220# a_26375_4612# 0.005781f
C197 ringtest_0.x4._14_ a_22373_5156# 0.002114f
C198 ringtest_0.x4.net6 ringtest_0.x4.net4 0.008308f
C199 a_21981_9142# ringtest_0.x4.clknet_1_0__leaf_clk 0.050329f
C200 a_12473_23980# ui_in[3] 0.143958f
C201 ringtest_0.x4.net2 ringtest_0.x4._01_ 9.85e-20
C202 ringtest_0.x4._11_ a_23349_6422# 0.001422f
C203 ringtest_0.x4.net7 a_24883_6800# 0.019182f
C204 ringtest_0.x4._11_ a_23879_6940# 4.59e-19
C205 ringtest_0.x4._17_ a_21951_5878# 9.29e-21
C206 ringtest_0.x4.net1 a_22399_9142# 5.53e-20
C207 a_24361_5340# a_25393_5308# 0.048748f
C208 a_24527_5340# a_24800_5334# 0.074815f
C209 a_18662_32213# a_18836_32319# 0.006584f
C210 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP2 0.043402f
C211 ringtest_0.x4._17_ a_24883_6800# 0.016586f
C212 ringtest_0.x4._15_ a_26201_4790# 0.02569f
C213 ringtest_0.x4._21_ a_23899_5654# 2.03e-19
C214 ringtest_0.ring_out ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C215 ringtest_0.x4.net9 a_26808_5308# 2.66e-21
C216 a_24045_6654# ringtest_0.x4._19_ 0.046625f
C217 a_24329_6640# a_25421_6641# 5.23e-20
C218 ringtest_0.x4.clknet_0_clk a_24800_5334# 4.59e-20
C219 ringtest_0.x4._08_ ringtest_0.x4.net10 0.001321f
C220 ringtest_0.counter3 VDPWR 2.51653f
C221 ringtest_0.x4._03_ a_22021_4220# 0.112166f
C222 a_21509_4790# a_22164_4362# 0.00127f
C223 a_24317_4942# a_24479_4790# 0.004009f
C224 muxtest_0.x2.x2.GN4 ua[3] 0.085877f
C225 ringtest_0.x4._15_ a_26555_5334# 0.007874f
C226 ringtest_0.x4.net8 ringtest_0.x4._07_ 0.001136f
C227 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x3.x2.GN3 7.01e-21
C228 ringtest_0.x4._24_ a_26640_5334# 0.010979f
C229 a_16579_11759# ui_in[4] 0.261734f
C230 ringtest_0.x3.x1.nSEL1 a_16755_12091# 1.59e-19
C231 a_23809_4790# a_24317_4942# 0.017774f
C232 a_22116_4902# ringtest_0.x4.net5 0.001073f
C233 a_21948_5156# a_22074_4790# 0.005525f
C234 ringtest_0.x4._00_ VDPWR 0.655201f
C235 a_27489_3702# a_27815_3867# 0.024477f
C236 ringtest_0.x4.net8 a_25055_3867# 3.76e-19
C237 muxtest_0.x1.x3.GP3 muxtest_0.R2R3 0.115101f
C238 a_22392_5990# a_22224_6244# 0.239923f
C239 a_21951_5878# a_22817_6146# 0.034054f
C240 ringtest_0.x4._16_ a_22765_4478# 0.01632f
C241 a_13501_23906# VDPWR 0.218058f
C242 VDPWR ua[2] 13.246901f
C243 a_21852_8720# a_21785_8054# 1.58e-19
C244 a_21981_8976# a_21803_8598# 9.73e-19
C245 a_22052_8875# a_22228_8598# 0.007724f
C246 ringtest_0.x4.net6 a_23837_5878# 4.02e-19
C247 a_21845_8816# ringtest_0.x4._10_ 0.011255f
C248 ringtest_0.x4._01_ a_22399_8976# 0.121379f
C249 muxtest_0.x1.x3.GP3 ui_in[1] 0.003199f
C250 ringtest_0.x4.clknet_0_clk ringtest_0.x4._23_ 2.29e-20
C251 ringtest_0.x4.net6 ringtest_0.x4._22_ 0.641715f
C252 ringtest_0.x4.net9 a_26555_4790# 0.016338f
C253 muxtest_0.x2.x2.GN4 m3_13316_18955# 0.084813f
C254 muxtest_0.x1.x3.GN2 muxtest_0.R5R6 0.122627f
C255 a_23949_6654# ringtest_0.x4._16_ 3.45e-20
C256 ringtest_0.x4._07_ a_24729_4790# 0.112051f
C257 ringtest_0.x4._19_ a_24699_6200# 1.87e-20
C258 ringtest_0.x4.net10 VDPWR 1.28398f
C259 ringtest_0.x4._22_ a_24895_4790# 0.02378f
C260 ringtest_0.x4.net2 a_21785_8054# 0.165774f
C261 ringtest_0.x4.net6 a_24135_3867# 0.195979f
C262 ringtest_0.x4.counter[0] ua[1] 3.21e-19
C263 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A 5.04e-19
C264 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP3 3.82e-20
C265 ringtest_0.drv_out ringtest_0.x4._05_ 0.0016f
C266 a_24729_4790# a_25055_3867# 1.63e-21
C267 muxtest_0.x1.x3.GN2 VDPWR 0.701394f
C268 ringtest_0.x4._00_ a_21803_9508# 3.7e-19
C269 ringtest_0.x4._24_ a_26735_5156# 7.21e-19
C270 ringtest_0.x4.net7 a_23381_4584# 2.04e-20
C271 ringtest_0.x4._04_ ringtest_0.x4.net5 0.003846f
C272 ua[1] ua[4] 0.001128f
C273 ringtest_0.x4.net7 a_26555_4790# 2.26e-19
C274 ringtest_0.x4.net1 ringtest_0.x4._00_ 0.056053f
C275 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net5 6.12e-20
C276 ringtest_0.x4._14_ a_21399_5340# 4.89e-20
C277 a_24045_6654# ringtest_0.x4.net7 0.037726f
C278 a_24627_6200# VDPWR 0.001301f
C279 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GP1 1.21e-19
C280 ringtest_0.x4.clknet_1_1__leaf_clk a_25168_5156# 0.042872f
C281 muxtest_0.x1.x3.GN4 ui_in[2] 5.71e-20
C282 ringtest_0.x4._06_ a_22765_5308# 1.6e-20
C283 ringtest_0.x4.counter[4] VDPWR 0.454642f
C284 ringtest_0.x4.net8 a_26201_5340# 0.001229f
C285 muxtest_0.R2R3 muxtest_0.R1R2 1.9897f
C286 ringtest_0.x3.x2.GN3 ua[1] 0.429944f
C287 ringtest_0.x4._11_ a_24968_5308# 7.26e-20
C288 ringtest_0.x4._17_ a_24045_6654# 0.036473f
C289 a_23399_3867# VDPWR 0.316408f
C290 a_16579_11759# ringtest_0.x3.x2.GP1 1.21e-20
C291 ui_in[3] ui_in[5] 0.13854f
C292 ringtest_0.x4._08_ a_25393_5308# 9.54e-19
C293 muxtest_0.x2.x1.nSEL1 a_12297_23648# 0.073392f
C294 a_16755_12091# ringtest_0.x3.x2.GN3 0.004288f
C295 a_24004_6128# ringtest_0.x4._16_ 0.029136f
C296 muxtest_0.x1.x1.nSEL1 ui_in[0] 0.169954f
C297 ringtest_0.x4.net9 ringtest_0.x4.counter[6] 3.69e-19
C298 a_24699_6200# ringtest_0.x4.net9 0.170073f
C299 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR 0.92605f
C300 ringtest_0.counter3 ringtest_0.x4.counter[2] 0.16993f
C301 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x3.x1.nSEL1 1.23e-19
C302 ringtest_0.x4.net6 a_25225_5334# 8.63e-19
C303 ringtest_0.x4._15_ a_23770_5308# 0.229149f
C304 a_21509_4790# a_22373_5156# 0.032244f
C305 a_23899_5334# ringtest_0.x4._20_ 1.05e-19
C306 ringtest_0.x4._03_ a_22541_5058# 3.08e-19
C307 a_25225_5334# a_24895_4790# 1.5e-19
C308 a_25393_5308# a_25336_4902# 6.84e-19
C309 ringtest_0.x4.net2 ringtest_0.x4._16_ 5.41e-20
C310 muxtest_0.x2.x2.GP1 ua[0] 0.128232f
C311 ringtest_0.x4._24_ a_25364_5878# 0.025563f
C312 a_26627_4246# a_26895_3867# 1.23e-19
C313 a_15575_12017# VDPWR 0.211635f
C314 ringtest_0.x4.net7 ringtest_0.x4.counter[6] 1.8e-19
C315 ringtest_0.x4._16_ a_23963_4790# 5.12e-19
C316 ringtest_0.x4._11_ a_25925_6788# 0.087773f
C317 a_22649_6244# a_22765_4478# 3.06e-22
C318 ringtest_0.x4.net7 a_24699_6200# 6.37e-20
C319 a_21840_5308# a_21863_4790# 6.87e-19
C320 ringtest_0.x4.net9 a_24479_4790# 8.5e-21
C321 a_22765_5308# a_22373_5156# 0.006202f
C322 a_19666_31955# muxtest_0.R7R8 7.47e-21
C323 ringtest_0.x4._16_ a_23381_4818# 0.113241f
C324 ringtest_0.x4.counter[2] ua[2] 1.11e-19
C325 a_26808_5308# a_27065_5334# 0.036838f
C326 a_22265_5308# a_22795_5334# 2.84e-19
C327 a_24361_5340# a_24715_5334# 0.057611f
C328 a_22097_5334# a_22181_5334# 0.008508f
C329 ringtest_0.x4._17_ a_24699_6200# 7.49e-19
C330 muxtest_0.x2.x1.nSEL0 ui_in[3] 0.32698f
C331 muxtest_0.R7R8 m3_13302_19985# 0.001045f
C332 a_25393_5308# VDPWR 0.406789f
C333 a_24336_6544# a_24287_6422# 4.04e-19
C334 a_24536_6699# a_24883_6800# 0.037333f
C335 a_24465_6800# a_24685_6788# 4.62e-19
C336 a_21425_9686# ringtest_0.x4._00_ 0.167554f
C337 ringtest_0.x4.net4 ringtest_0.x4.net5 0.483177f
C338 ringtest_0.x4.net7 a_24479_4790# 1.98e-19
C339 a_25421_6641# ringtest_0.x4._19_ 0.214472f
C340 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP1 0.001426f
C341 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.001676f
C342 a_12297_23648# muxtest_0.x2.x2.GN3 6.68e-19
C343 ringtest_0.x4.net7 a_23809_4790# 0.003261f
C344 a_12473_23980# muxtest_0.x2.x2.GN1 1.46e-19
C345 muxtest_0.R7R8 muxtest_0.x2.x2.GP2 1.13e-20
C346 a_23932_6128# a_23837_5878# 0.002032f
C347 ringtest_0.x4._11_ a_21233_5340# 0.00462f
C348 ringtest_0.x4._17_ a_23809_4790# 1e-20
C349 a_21951_5878# ringtest_0.x4._14_ 3.24e-22
C350 a_26749_6422# a_26201_5340# 6.06e-21
C351 ringtest_0.x4.net8 ringtest_0.x4._06_ 0.209874f
C352 a_27191_4790# VDPWR 4.71e-19
C353 ringtest_0.x4.net8 a_24070_5852# 0.028641f
C354 a_22392_5990# a_22139_5878# 3.39e-19
C355 a_26808_4902# VDPWR 0.186041f
C356 ringtest_0.counter3 a_21375_3867# 4.27e-20
C357 ringtest_0.x3.x2.GN4 VDPWR 1.23317f
C358 muxtest_0.x1.x4.A muxtest_0.R5R6 1.64e-20
C359 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_0_clk 0.004956f
C360 muxtest_0.x1.x3.GN3 ua[3] 0.014498f
C361 muxtest_0.x1.x5.GN muxtest_0.x2.nselect2 4.76e-21
C362 a_25421_6641# ringtest_0.x4.net9 3.61e-20
C363 ringtest_0.x3.x2.GP1 m3_17032_8096# 3.25e-21
C364 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._12_ 0.075464f
C365 ringtest_0.x3.x2.GN3 m3_17046_7066# 0.016026f
C366 ringtest_0.x4._24_ a_26913_4566# 0.002926f
C367 ringtest_0.x4._16_ ringtest_0.x4._20_ 0.011071f
C368 muxtest_0.x1.x4.A VDPWR 15.014299f
C369 a_21233_5340# a_21675_4790# 2.24e-19
C370 ringtest_0.x4._22_ ringtest_0.x4.net5 4.26e-20
C371 a_21399_5340# a_21509_4790# 0.010101f
C372 a_19794_32347# muxtest_0.x1.x3.GN4 3.22e-19
C373 ringtest_0.x4.net8 a_23891_4790# 4.38e-20
C374 muxtest_0.x1.x3.GN3 a_20492_32319# 1.07e-20
C375 a_22164_4362# a_22390_4566# 0.005961f
C376 ringtest_0.x4._11_ a_25761_5058# 0.028602f
C377 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A 0.17253f
C378 a_21465_9294# a_21780_9142# 7.84e-20
C379 a_27065_5156# a_27273_4220# 0.003595f
C380 a_19842_32287# muxtest_0.x1.x3.GN3 0.004289f
C381 a_21675_9686# a_21852_9416# 0.001655f
C382 a_21465_9294# a_21561_9116# 0.310858f
C383 ringtest_0.counter7 a_22295_3867# 2.81e-20
C384 ringtest_0.x4.net5 a_24135_3867# 0.001724f
C385 ringtest_0.x4._19_ ringtest_0.x4._24_ 8.27e-21
C386 a_19666_31955# VDPWR 0.171399f
C387 a_27233_5058# ringtest_0.x4.net11 0.092457f
C388 ringtest_0.x4._11_ a_21675_4790# 0.03376f
C389 ringtest_0.x4.net6 ringtest_0.x4._15_ 0.117386f
C390 a_21840_5308# a_22097_5334# 0.036838f
C391 a_25421_6641# ringtest_0.x4.net7 0.030401f
C392 muxtest_0.x1.x1.nSEL0 a_19114_31955# 0.03096f
C393 ringtest_0.x4._15_ a_24895_4790# 2.57e-20
C394 ringtest_0.x4._16_ a_21840_5308# 1.76e-20
C395 ringtest_0.x4._17_ a_25421_6641# 0.019971f
C396 a_23529_6422# ringtest_0.x4._05_ 4.91e-20
C397 a_23949_6654# a_24465_6800# 1.28e-19
C398 ringtest_0.x4._18_ ringtest_0.x4.clknet_1_1__leaf_clk 3.06e-19
C399 a_24329_6640# a_24336_6544# 0.961627f
C400 ringtest_0.x4._24_ a_26735_5334# 7.21e-19
C401 ringtest_0.x3.x2.GP2 ringtest_0.counter7 1.13e-20
C402 a_25336_4902# a_25083_4790# 3.39e-19
C403 ringtest_0.x3.x2.GP3 ui_in[4] 0.003259f
C404 muxtest_0.x1.x3.GN1 ui_in[0] 0.023343f
C405 a_21465_8830# VDPWR 0.399249f
C406 a_23381_4818# a_23467_4818# 0.006584f
C407 a_21785_5878# a_21233_5340# 0.002682f
C408 ringtest_0.x4._13_ a_21399_5340# 1.58e-19
C409 ringtest_0.x4.net6 a_24926_5712# 0.001426f
C410 a_27489_3702# ringtest_0.x4.counter[9] 0.109832f
C411 muxtest_0.x2.x2.GP2 VDPWR 1.81003f
C412 a_26201_5340# ringtest_0.x4._09_ 1.11e-19
C413 a_26367_5340# a_26201_4790# 2.64e-19
C414 ringtest_0.x4._14_ a_23381_4584# 9.06e-21
C415 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x1.nSEL1 2.53e-21
C416 ringtest_0.x4._11_ a_21785_5878# 0.205946f
C417 a_26721_4246# a_26895_3867# 2.21e-19
C418 a_25083_4790# VDPWR 0.079731f
C419 ringtest_0.x4._24_ ringtest_0.x4.net9 0.165357f
C420 muxtest_0.x1.x3.GP2 ua[3] 0.023177f
C421 a_25364_5878# a_25977_4220# 4.57e-20
C422 a_22399_9142# ringtest_0.x4._11_ 2.48e-19
C423 ringtest_0.x4.clknet_1_0__leaf_clk a_22245_8054# 0.00537f
C424 a_21948_5156# VDPWR 0.286549f
C425 ringtest_0.x4.net3 a_21852_8720# 0.005586f
C426 a_26367_5340# a_26555_5334# 0.097994f
C427 a_21852_9416# a_22052_8875# 1.26e-19
C428 a_21845_9116# a_21852_8720# 3.36e-19
C429 a_22052_9116# a_21845_8816# 6.88e-20
C430 a_24715_5334# VDPWR 0.084103f
C431 ringtest_0.x4._15_ a_22939_4584# 1.81e-19
C432 a_19842_32287# muxtest_0.x1.x3.GP2 2.95e-20
C433 ringtest_0.x4.net1 a_21465_8830# 0.081622f
C434 ringtest_0.x4.net2 ringtest_0.x4.net3 1.28152f
C435 ringtest_0.x4._15_ a_27169_6641# 8.98e-20
C436 muxtest_0.R7R8 ua[0] 2.33155f
C437 ringtest_0.x4.net7 ringtest_0.x4._24_ 2.68e-19
C438 ringtest_0.x4.net2 a_21845_9116# 4.59e-19
C439 ringtest_0.ring_out ringtest_0.x3.x2.GN1 4.6809f
C440 a_21951_5878# a_21509_4790# 1.21e-19
C441 a_21785_5878# a_21675_4790# 3.23e-21
C442 ringtest_0.x4._09_ a_27233_5058# 0.010518f
C443 a_26201_4790# a_27065_5156# 0.032244f
C444 ringtest_0.x4._07_ a_24361_5340# 0.022853f
C445 ringtest_0.x4._17_ ringtest_0.x4._24_ 0.004444f
C446 ringtest_0.counter7 ringtest_0.x4._23_ 0.004833f
C447 a_24763_6143# a_24800_5334# 1.41e-19
C448 ringtest_0.x4.net5 a_22021_4220# 0.006016f
C449 ringtest_0.x4._22_ a_24527_5340# 0.015364f
C450 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.025028f
C451 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP3 0.001226f
C452 ringtest_0.counter7 a_26367_4790# 5.88e-20
C453 muxtest_0.R1R2 ui_in[4] 8.73e-20
C454 ringtest_0.x4._04_ a_22983_5654# 0.002919f
C455 muxtest_0.x2.x1.nSEL0 a_12425_24040# 2.51e-19
C456 a_24361_5340# a_25055_3867# 1.7e-21
C457 a_21780_8964# VDPWR 3.44e-19
C458 a_22224_6244# a_22265_5308# 0.004197f
C459 a_22392_5990# a_22097_5334# 0.004484f
C460 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN1 0.004375f
C461 a_24336_6544# a_24317_4942# 2.42e-19
C462 ringtest_0.x4.clknet_1_0__leaf_clk a_22983_5654# 1.8e-20
C463 ringtest_0.x4.clknet_0_clk ringtest_0.x4._22_ 0.003156f
C464 muxtest_0.R7R8 muxtest_0.x2.x2.GN3 0.01204f
C465 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GP3 2.78e-20
C466 a_22392_5990# ringtest_0.x4._16_ 1.01e-19
C467 ringtest_0.ring_out ui_in[6] 0.550306f
C468 ringtest_0.x4._11_ ringtest_0.counter3 1.13e-19
C469 muxtest_0.x1.x4.A a_12849_23648# 1.34e-19
C470 uio_in[1] uio_in[0] 0.033505f
C471 ringtest_0.x4.clknet_1_1__leaf_clk a_24800_5334# 0.033626f
C472 ringtest_0.x4.clknet_0_clk a_23619_6788# 9.48e-20
C473 ringtest_0.x4._13_ a_21951_5878# 7.99e-20
C474 muxtest_0.x2.x1.nSEL1 VDPWR 0.649185f
C475 a_21981_8976# ringtest_0.x4._01_ 0.00226f
C476 ringtest_0.x4.net3 a_22399_8976# 4.27e-20
C477 ringtest_0.x4.clknet_1_0__leaf_clk a_21591_6128# 0.001585f
C478 ringtest_0.x4._00_ ringtest_0.x4._11_ 0.003231f
C479 a_26627_4246# a_26817_4566# 0.011458f
C480 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A 0.429373f
C481 a_27065_5156# a_27303_4246# 3.93e-20
C482 a_13025_23980# ui_in[3] 0.279858f
C483 ringtest_0.x4.net1 a_21780_8964# 1.42e-19
C484 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A 5.04e-19
C485 ringtest_0.x4.net7 a_26007_6788# 0.003849f
C486 a_24527_5340# a_25225_5334# 0.192206f
C487 a_21840_5308# a_21587_5334# 3.39e-19
C488 a_21399_5340# a_21798_5712# 8.12e-19
C489 a_24968_5308# a_25393_5308# 1.28e-19
C490 a_24361_5340# a_26201_5340# 0.002059f
C491 a_21948_5156# ringtest_0.x4.counter[2] 1.99e-20
C492 a_19114_31955# muxtest_0.x1.x3.GN2 0.106131f
C493 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._23_ 0.071442f
C494 ringtest_0.x4._11_ ringtest_0.x4.net10 0.36244f
C495 ringtest_0.x4.clknet_1_1__leaf_clk a_26367_4790# 0.031849f
C496 a_24336_6544# ringtest_0.x4._19_ 0.457296f
C497 VDPWR ua[0] 3.15952f
C498 a_12849_23648# muxtest_0.x2.x2.GP2 3.07e-19
C499 ringtest_0.x4.clknet_0_clk a_25225_5334# 0.013741f
C500 muxtest_0.x1.x3.GP3 ui_in[0] 2.74e-19
C501 ringtest_0.x4._15_ ringtest_0.x4.net5 0.016962f
C502 ringtest_0.x4._03_ a_22765_4478# 1.19e-19
C503 ringtest_0.x4.net4 a_22983_5654# 5.3e-19
C504 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2 2.14737f
C505 ringtest_0.drv_out VDPWR 16.4224f
C506 muxtest_0.x2.nselect2 ui_in[4] 0.001201f
C507 a_17231_12017# ui_in[4] 0.125445f
C508 ringtest_0.x4._11_ a_22775_5878# 8.02e-19
C509 ringtest_0.x4._24_ a_27065_5334# 0.013075f
C510 a_15575_12017# a_15749_12123# 0.006584f
C511 ringtest_0.x3.x1.nSEL1 a_16155_12151# 9.57e-19
C512 ringtest_0.x4._11_ a_24627_6200# 4.38e-19
C513 a_22541_5058# ringtest_0.x4.net5 0.13266f
C514 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN1 0.034862f
C515 ringtest_0.x4._08_ ringtest_0.x4._07_ 9.41e-21
C516 muxtest_0.R3R4 ua[3] 0.039417f
C517 ringtest_0.x4._11_ ringtest_0.x4.counter[4] 6.77e-20
C518 ringtest_0.x4._18_ a_23993_5654# 6.01e-19
C519 a_13675_24012# VDPWR 8.97e-19
C520 ringtest_0.x4.net8 a_26895_3867# 7.5e-19
C521 a_22392_5990# a_22649_6244# 0.036838f
C522 muxtest_0.x2.x2.GN3 VDPWR 0.650589f
C523 a_21951_5878# ringtest_0.x4.net8 0.001542f
C524 a_23879_6940# a_24715_5334# 2.19e-20
C525 ringtest_0.x4.net9 a_25977_4220# 9.8e-19
C526 a_22052_8875# ringtest_0.x4._10_ 2.11e-19
C527 a_23949_6654# a_23770_5308# 8.51e-20
C528 ringtest_0.x4._01_ a_22228_8598# 5.75e-19
C529 muxtest_0.x1.x3.GN4 muxtest_0.R2R3 0.127088f
C530 ringtest_0.x4.net9 a_25719_4790# 0.001933f
C531 muxtest_0.x1.x3.GN4 ui_in[1] 0.059771f
C532 a_24329_6640# ringtest_0.x4._16_ 1.49e-19
C533 ringtest_0.x4.net4 a_22486_4246# 0.003167f
C534 ringtest_0.x4._07_ a_25336_4902# 0.004454f
C535 a_24336_6544# ringtest_0.x4.net9 1.52e-20
C536 ringtest_0.x4._22_ a_25168_5156# 0.002895f
C537 ringtest_0.x3.x2.GP2 ui_in[3] 5.28e-19
C538 ringtest_0.x4._24_ a_26627_4246# 0.085832f
C539 muxtest_0.R3R4 m3_13316_18955# 1.46e-19
C540 ringtest_0.x4.net7 a_25977_4220# 0.023542f
C541 ringtest_0.x4._00_ a_22399_9142# 0.139872f
C542 ringtest_0.x4._18_ ringtest_0.x4._04_ 0.003255f
C543 ringtest_0.x4._24_ a_27149_5156# 8.56e-19
C544 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN4 9.02e-19
C545 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN3 0.012418f
C546 ringtest_0.x4._23_ a_26367_4790# 0.031117f
C547 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN2 0.154394f
C548 ringtest_0.x4._07_ VDPWR 0.322336f
C549 a_24336_6544# ringtest_0.x4.net7 0.027472f
C550 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.001676f
C551 ringtest_0.x4._06_ a_24361_5340# 0.091082f
C552 ringtest_0.x4.clknet_1_1__leaf_clk a_25593_5156# 0.044904f
C553 ringtest_0.x4.net8 a_26808_5308# 8.61e-20
C554 ringtest_0.x4._16_ a_24545_5878# 0.036674f
C555 ringtest_0.x4._11_ a_25393_5308# 1.18e-19
C556 ringtest_0.x4._17_ a_24336_6544# 0.050404f
C557 a_25055_3867# VDPWR 0.315151f
C558 a_16155_12151# ringtest_0.x3.x2.GN3 5.17e-20
C559 ringtest_0.x3.x2.GN2 a_16707_12151# 3.11e-20
C560 ringtest_0.x4.net2 ringtest_0.x4._03_ 5.34e-20
C561 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN3 0.002857f
C562 ringtest_0.x4._08_ a_26201_5340# 0.097891f
C563 muxtest_0.x2.x1.nSEL1 a_12849_23648# 7.84e-19
C564 a_25364_5878# ringtest_0.x4._16_ 0.001016f
C565 a_24264_6788# VDPWR 7.65e-20
C566 muxtest_0.x2.x1.nSEL0 ua[3] 7.05e-20
C567 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ui_in[6] 0.108977f
C568 ringtest_0.x4.net6 a_26367_5340# 1.27e-19
C569 ringtest_0.x4._03_ a_23381_4818# 2.2e-20
C570 ringtest_0.x4._15_ a_24527_5340# 0.027322f
C571 a_21509_4790# a_23809_4790# 1.62e-21
C572 a_21845_8816# a_21395_6940# 6.92e-20
C573 a_25225_5334# a_25168_5156# 7.26e-19
C574 a_27273_4220# a_27489_3702# 1.29e-21
C575 a_26817_4566# a_26721_4246# 1.26e-19
C576 muxtest_0.x1.x4.A muxtest_0.x1.x5.A 2.05508f
C577 ringtest_0.x4.clknet_0_clk ringtest_0.x4._15_ 4.05e-19
C578 a_16203_12091# VDPWR 0.192568f
C579 muxtest_0.x1.x3.GP1 muxtest_0.R7R8 4.13739f
C580 a_21561_8830# ringtest_0.x4._12_ 0.036321f
C581 ringtest_0.x4.net8 a_23381_4584# 9.57e-20
C582 ringtest_0.x4._11_ a_27191_4790# 9.67e-22
C583 ringtest_0.x4.net9 a_25677_5156# 8.89e-19
C584 ringtest_0.x4.net11 a_26895_3867# 3.2e-20
C585 ringtest_0.x4._11_ a_26808_4902# 8.51e-19
C586 ringtest_0.x4.counter[1] ua[1] 3.21e-19
C587 ringtest_0.x4._16_ a_24317_4942# 1.3e-19
C588 a_16707_12151# ui_in[3] 0.001558f
C589 a_24045_6654# ringtest_0.x4.net8 1.55e-19
C590 ringtest_0.x3.x2.GN2 ui_in[3] 0.114345f
C591 a_27233_5308# a_27065_5334# 0.310858f
C592 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._04_ 1.67e-21
C593 a_22265_5308# a_23899_5334# 2.67e-21
C594 a_22765_5308# a_22795_5334# 0.025037f
C595 a_24968_5308# a_24715_5334# 3.39e-19
C596 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A 0.159172f
C597 a_26201_5340# VDPWR 0.714632f
C598 ringtest_0.x4._05_ a_24883_6800# 0.114695f
C599 a_24465_6800# a_24287_6422# 9.73e-19
C600 ringtest_0.x4.net6 a_22765_4478# 5.34e-20
C601 ringtest_0.x4._16_ a_23151_5334# 0.010038f
C602 ringtest_0.x4._18_ ringtest_0.x4.net4 3.06e-19
C603 ringtest_0.counter7 ringtest_0.x4.net4 6.88e-20
C604 ringtest_0.drv_out a_23879_6940# 0.318051f
C605 ringtest_0.x4.net7 a_25677_5156# 0.002598f
C606 ringtest_0.x4._23_ a_25593_5156# 0.001187f
C607 a_25593_5156# a_26367_4790# 2.56e-19
C608 a_24729_4790# a_26555_4790# 4.76e-21
C609 a_23949_6654# ringtest_0.x4.net6 1.76e-19
C610 ringtest_0.x4.counter[5] VDPWR 0.450193f
C611 a_12849_23648# muxtest_0.x2.x2.GN3 0.104151f
C612 a_13025_23980# muxtest_0.x2.x2.GN1 3.78e-20
C613 ringtest_0.x4._21_ ringtest_0.x4._07_ 4.77e-20
C614 a_22224_6244# ringtest_0.x4._14_ 5.19e-22
C615 ringtest_0.x4.net7 a_23899_5334# 0.006434f
C616 ringtest_0.x4.net9 ringtest_0.x4.counter[9] 5.19e-19
C617 a_26749_6422# a_26808_5308# 2.48e-20
C618 ringtest_0.x4._25_ a_26201_5340# 1.01e-19
C619 m2_15612_11606# ui_in[3] 0.130999f
C620 ringtest_0.x3.nselect2 a_16579_11759# 1.29e-19
C621 a_22164_4362# VDPWR 0.108977f
C622 ringtest_0.counter3 ringtest_0.x4.counter[4] 0.07836f
C623 ringtest_0.x4.net8 ringtest_0.x4.counter[6] 0.079257f
C624 ringtest_0.x4.net8 a_24699_6200# 0.003186f
C625 ringtest_0.x4._17_ a_23899_5334# 9.12e-21
C626 a_27233_5058# VDPWR 0.462064f
C627 a_22224_6244# a_22319_6244# 0.007724f
C628 a_22392_5990# a_22733_6244# 9.73e-19
C629 ringtest_0.counter3 a_23399_3867# 0.110188f
C630 a_23529_6422# VDPWR 0.185924f
C631 ringtest_0.x4.net4 a_22295_3867# 0.202764f
C632 ringtest_0.x4._12_ a_21049_8598# 0.090947f
C633 ringtest_0.x4._19_ ringtest_0.x4._16_ 0.001191f
C634 muxtest_0.x1.x3.GP1 muxtest_0.R5R6 0.122287f
C635 a_23770_5308# ringtest_0.x4._20_ 3.36e-20
C636 ringtest_0.x4._18_ a_23837_5878# 0.002103f
C637 ringtest_0.x4.net6 a_24004_6128# 0.074355f
C638 ringtest_0.counter7 ringtest_0.x4._22_ 1.31e-20
C639 a_21672_5334# a_21509_4790# 4.57e-19
C640 a_21233_5340# a_21948_5156# 0.001041f
C641 a_21840_5308# ringtest_0.x4._03_ 0.009555f
C642 a_25977_4220# a_26627_4246# 0.010893f
C643 a_22765_4478# a_22939_4584# 0.006584f
C644 a_22021_4220# a_22486_4246# 0.005941f
C645 ringtest_0.x4.net8 a_24479_4790# 0.002158f
C646 ringtest_0.x4._11_ a_25083_4790# 0.016192f
C647 muxtest_0.x1.x3.GP1 VDPWR 3.2848f
C648 a_21465_9294# ringtest_0.x4.net3 9.98e-20
C649 a_24699_6200# a_24729_4790# 5.07e-21
C650 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN3 0.08518f
C651 ringtest_0.x4.net9 a_27149_5334# 1.06e-19
C652 a_21465_9294# a_21845_9116# 0.048748f
C653 a_21561_9116# a_21852_9416# 0.194892f
C654 ringtest_0.counter7 a_24135_3867# 2.81e-20
C655 ringtest_0.x4.net8 a_23809_4790# 7.44e-19
C656 a_20318_32213# VDPWR 0.217349f
C657 ringtest_0.x4._11_ a_21948_5156# 0.00274f
C658 a_22265_5308# a_22097_5334# 0.310858f
C659 ringtest_0.ring_out ui_in[4] 0.016625f
C660 muxtest_0.x1.x1.nSEL0 a_19666_31955# 1.91e-20
C661 ringtest_0.x4._16_ a_22265_5308# 7.03e-19
C662 ringtest_0.x4._06_ VDPWR 0.276236f
C663 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.025028f
C664 a_24336_6544# a_24536_6699# 0.074815f
C665 a_24329_6640# a_24465_6800# 0.136009f
C666 a_24045_6654# ringtest_0.x4._05_ 9.72e-20
C667 a_24070_5852# VDPWR 0.084816f
C668 a_25168_5156# a_25263_5156# 0.007724f
C669 a_21395_6940# a_21399_5340# 1.82e-21
C670 ringtest_0.x4.net6 a_23381_4818# 4.93e-21
C671 ringtest_0.x4.net9 ringtest_0.x4._16_ 0.243936f
C672 a_24763_6143# ringtest_0.x4._22_ 0.155189f
C673 a_21845_8816# VDPWR 0.446206f
C674 ringtest_0.x4._04_ ringtest_0.x4._02_ 1.6e-19
C675 a_23809_4790# a_24729_4790# 2.37e-21
C676 ringtest_0.x4._15_ a_22983_5654# 1.54e-19
C677 ringtest_0.x4.net2 a_21055_5334# 0.002977f
C678 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._02_ 0.254839f
C679 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ui_in[6] 6.29e-19
C680 a_21675_4790# a_21948_5156# 0.081834f
C681 a_23399_3867# ringtest_0.x4.counter[4] 0.001146f
C682 a_26640_5334# a_26201_4790# 1.73e-19
C683 a_23891_4790# VDPWR 2.86e-19
C684 ringtest_0.x4.net7 ringtest_0.x4._16_ 5.07e-19
C685 a_22164_4362# ringtest_0.x4.counter[2] 6.46e-19
C686 a_24465_6800# a_24545_5878# 1.71e-20
C687 a_22373_5156# VDPWR 0.183311f
C688 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._22_ 0.031888f
C689 ringtest_0.x3.x1.nSEL0 VDPWR 0.5228f
C690 ringtest_0.x4.net3 a_21981_8976# 2.06e-19
C691 a_26640_5334# a_26555_5334# 0.037333f
C692 a_26808_5308# a_26766_5712# 4.62e-19
C693 ringtest_0.x4._17_ ringtest_0.x4._16_ 0.048058f
C694 a_21845_9116# a_21981_8976# 5.28e-20
C695 a_21852_9416# ringtest_0.x4._01_ 8.68e-20
C696 a_22052_9116# a_22052_8875# 0.013851f
C697 ringtest_0.drv_out a_25925_6788# 1.34e-19
C698 ringtest_0.x4._05_ a_24699_6200# 3.16e-19
C699 muxtest_0.x2.x1.nSEL1 m2_11882_23495# 0.00815f
C700 ringtest_0.x3.x2.GN4 ringtest_0.counter3 0.237196f
C701 a_21767_5334# VDPWR 0.003619f
C702 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP2 0.068989f
C703 ringtest_0.x4.net1 a_21845_8816# 0.002755f
C704 ringtest_0.ring_out ringtest_0.x3.x2.GP1 4.09516f
C705 ringtest_0.x4.net2 a_21981_9142# 3.46e-19
C706 a_12977_24040# muxtest_0.x2.x2.GP3 4.39e-19
C707 a_22224_6244# a_21509_4790# 5.5e-20
C708 ringtest_0.x4._09_ a_26555_4790# 0.129132f
C709 a_26201_4790# a_26735_5156# 0.002698f
C710 a_21785_5878# a_21948_5156# 8.98e-19
C711 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP3 0.004298f
C712 ringtest_0.x4._07_ a_24968_5308# 0.011124f
C713 ringtest_0.x4._22_ a_24800_5334# 0.006172f
C714 ringtest_0.x4.net5 a_22765_4478# 0.081136f
C715 ringtest_0.x4.clknet_1_0__leaf_clk a_22116_4902# 0.001507f
C716 ringtest_0.x4.net6 ringtest_0.x4._20_ 0.00624f
C717 muxtest_0.x2.nselect2 muxtest_0.x2.x2.GN4 1.53e-20
C718 a_23349_6422# a_23529_6422# 0.185422f
C719 a_22201_8964# VDPWR 0.002269f
C720 ringtest_0.x4._20_ a_24895_4790# 0.003428f
C721 a_26269_4612# VDPWR 0.001259f
C722 ringtest_0.x4.net10 a_26808_4902# 1.26e-19
C723 a_13025_23980# ua[3] 9.59e-19
C724 ringtest_0.x4._21_ ringtest_0.x4._06_ 0.224771f
C725 ringtest_0.counter7 ua[3] 1.17e-19
C726 ringtest_0.x4.net4 ringtest_0.x4._02_ 1.19e-19
C727 a_22817_6146# ringtest_0.x4._16_ 0.001048f
C728 ringtest_0.x3.x1.nSEL1 ui_in[4] 0.272823f
C729 a_24070_5852# ringtest_0.x4._21_ 0.114705f
C730 a_22139_5878# a_22319_6244# 0.001229f
C731 a_27489_3702# ringtest_0.x4.counter[8] 0.006251f
C732 a_24004_6128# a_23932_6128# 0.005941f
C733 muxtest_0.x1.x4.A a_13501_23906# 0.001685f
C734 a_21395_6940# a_21951_5878# 1.63e-19
C735 ringtest_0.x4.clknet_1_1__leaf_clk a_25225_5334# 0.024694f
C736 ringtest_0.x4.net6 a_21840_5308# 6.4e-20
C737 ringtest_0.drv_out ringtest_0.x4._11_ 1.2e-19
C738 ringtest_0.x4.clknet_0_clk a_24685_6788# 4.62e-19
C739 ringtest_0.x4._23_ ringtest_0.x4._22_ 0.511385f
C740 ringtest_0.x4._13_ a_22224_6244# 5.02e-20
C741 a_22499_4790# VDPWR 4.65e-19
C742 ringtest_0.x4._22_ a_26367_4790# 3.15e-20
C743 a_27065_5334# a_27149_5334# 0.008508f
C744 ringtest_0.x4._24_ ringtest_0.x4.net8 1.23e-20
C745 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._04_ 0.005301f
C746 a_22021_4220# a_22295_3867# 4.71e-19
C747 a_25364_5878# a_26201_4790# 6.92e-20
C748 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A 0.429199f
C749 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 5.02073f
C750 muxtest_0.x2.x2.GN1 ui_in[3] 0.021261f
C751 a_23879_6940# ringtest_0.x4._06_ 1.96e-20
C752 ringtest_0.x4.net7 a_26201_6788# 5.71e-19
C753 ringtest_0.x4._17_ a_22649_6244# 1.03e-20
C754 a_23879_6940# a_24070_5852# 3.15e-19
C755 a_21672_5334# a_21798_5712# 0.005525f
C756 a_24527_5340# a_26367_5340# 0.001861f
C757 a_19666_31955# muxtest_0.x1.x3.GN2 1.61e-19
C758 ringtest_0.x4.net6 a_26569_6422# 2.84e-19
C759 ringtest_0.x4._17_ a_26201_6788# 3.01e-19
C760 a_21399_5340# VDPWR 0.341027f
C761 a_25364_5878# a_26555_5334# 9.53e-19
C762 muxtest_0.x1.x1.nSEL1 a_18662_32213# 0.193944f
C763 ringtest_0.x4.net4 a_22116_4902# 0.007782f
C764 ringtest_0.x4.clknet_1_1__leaf_clk a_26640_5156# 3.02e-19
C765 ringtest_0.x4._05_ a_25421_6641# 0.121098f
C766 muxtest_0.x2.x2.GP2 ua[2] 0.349855f
C767 a_24465_6800# ringtest_0.x4._19_ 0.040707f
C768 ringtest_0.x4._18_ ringtest_0.x4._15_ 0.045245f
C769 ringtest_0.counter7 ringtest_0.x4._15_ 0.003538f
C770 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.001676f
C771 a_24968_5308# ringtest_0.x4.counter[5] 2.7e-21
C772 ringtest_0.x4.net2 ringtest_0.x4.net5 7.09e-21
C773 muxtest_0.x1.x3.GN4 ui_in[0] 0.218694f
C774 muxtest_0.x1.x1.nSEL1 m2_18699_31802# 0.00815f
C775 ringtest_0.x4.net5 a_23963_4790# 1.04e-20
C776 a_17405_12123# ui_in[4] 8.84e-19
C777 ringtest_0.x4._15_ a_27191_5712# 6.51e-20
C778 ringtest_0.x3.x2.GN3 ui_in[4] 0.273713f
C779 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GP1 1.21e-19
C780 ringtest_0.x4._11_ ringtest_0.x4._07_ 0.161717f
C781 a_16027_11759# ringtest_0.x3.x2.GN2 0.106178f
C782 a_21863_4790# a_22043_5156# 0.001229f
C783 a_23381_4818# ringtest_0.x4.net5 4.5e-19
C784 muxtest_0.x1.x3.GN3 muxtest_0.R1R2 4.03753f
C785 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ui_in[6] 3.49e-19
C786 muxtest_0.R7R8 muxtest_0.R4R5 0.286971f
C787 a_22817_6146# a_22649_6244# 0.310858f
C788 a_22224_6244# ringtest_0.x4.net8 4.11e-20
C789 uio_in[6] uio_in[5] 0.031023f
C790 ringtest_0.x4.net9 a_27273_4220# 0.001158f
C791 ringtest_0.x4._01_ ringtest_0.x4._10_ 0.002197f
C792 a_24045_6654# a_24361_5340# 1.16e-21
C793 ringtest_0.x4.net4 ringtest_0.x4._04_ 0.689049f
C794 ringtest_0.x4.net9 a_26766_4790# 0.002793f
C795 ringtest_0.x4._15_ a_24763_6143# 1.57e-19
C796 muxtest_0.x1.x3.GN1 muxtest_0.R3R4 3.99705f
C797 a_24536_6699# ringtest_0.x4._16_ 1.35e-21
C798 ringtest_0.x4._07_ a_25761_5058# 3.3e-20
C799 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR 0.639695f
C800 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP3 0.09552f
C801 a_24465_6800# ringtest_0.x4.net9 0.004659f
C802 ringtest_0.x4._22_ a_25593_5156# 6.29e-19
C803 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net4 0.158995f
C804 ringtest_0.x4.clknet_0_clk a_23949_6654# 0.002548f
C805 ringtest_0.x4.net6 a_22392_5990# 3.85e-19
C806 ringtest_0.x4.net2 a_21007_3867# 0.223155f
C807 ringtest_0.x4._24_ a_26749_6422# 0.197975f
C808 ringtest_0.x4._24_ ringtest_0.x4.net11 0.002712f
C809 a_16027_11759# ui_in[3] 0.246189f
C810 ringtest_0.x4.net6 a_24287_6422# 1.73e-19
C811 ringtest_0.x4._23_ a_26640_5156# 0.011058f
C812 a_26808_4902# a_27191_4790# 4.67e-20
C813 ringtest_0.x4._05_ ringtest_0.x4._24_ 2.08e-20
C814 a_26367_4790# a_26640_5156# 0.078545f
C815 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._15_ 0.471647f
C816 ringtest_0.x4._14_ a_22097_5334# 2.97e-21
C817 a_24465_6800# ringtest_0.x4.net7 0.035198f
C818 ringtest_0.x4.clknet_1_1__leaf_clk a_25263_5156# 0.001835f
C819 ringtest_0.x4._06_ a_24968_5308# 0.001008f
C820 ringtest_0.x4._16_ ringtest_0.x4._14_ 0.202586f
C821 ringtest_0.x4.net8 a_27233_5308# 4.93e-20
C822 ringtest_0.x4._11_ a_26201_5340# 3.54e-20
C823 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP1 0.001426f
C824 a_24699_6200# a_24361_5340# 0.001396f
C825 ringtest_0.x4._17_ a_24465_6800# 0.016441f
C826 a_26895_3867# VDPWR 0.303091f
C827 a_21951_5878# VDPWR 0.304738f
C828 ringtest_0.x4._08_ a_26808_5308# 0.047112f
C829 ringtest_0.x4.net5 ringtest_0.x4._20_ 8.42e-21
C830 a_24883_6800# VDPWR 0.085296f
C831 muxtest_0.x1.x3.GP2 muxtest_0.R1R2 0.153531f
C832 ringtest_0.x4.clknet_0_clk a_24004_6128# 2.03e-19
C833 a_21509_4790# a_21863_4790# 0.062224f
C834 ringtest_0.x4._15_ a_24800_5334# 0.026278f
C835 muxtest_0.R5R6 muxtest_0.R4R5 2.29244f
C836 ringtest_0.x4._22_ a_25441_4612# 0.002353f
C837 a_21785_8054# ringtest_0.x4._10_ 0.107891f
C838 ringtest_0.x4._13_ a_22139_5878# 5.97e-20
C839 a_22052_8875# a_21395_6940# 2.84e-19
C840 VDPWR ua[1] 17.382101f
C841 ringtest_0.drv_out ringtest_0.counter3 1.91048f
C842 a_25225_5334# a_25593_5156# 3.78e-19
C843 a_26555_5334# a_26735_5334# 0.001229f
C844 a_16755_12091# VDPWR 0.26222f
C845 a_22224_6244# a_22390_4566# 4.44e-21
C846 ringtest_0.x4.net8 a_25977_4220# 0.004343f
C847 a_21852_8720# ringtest_0.x4._12_ 0.206007f
C848 ringtest_0.x4._11_ a_22164_4362# 1e-19
C849 muxtest_0.x1.x3.GP1 muxtest_0.x1.x5.A 0.353808f
C850 muxtest_0.R4R5 VDPWR 1.56678f
C851 ringtest_0.x4.net9 a_26201_4790# 0.11266f
C852 ringtest_0.x4.net11 a_27815_3867# 0.003661f
C853 ringtest_0.x4.net8 a_25719_4790# 5.67e-20
C854 ringtest_0.x4._11_ a_27233_5058# 5.38e-21
C855 ua[0] ua[2] 4.5205f
C856 a_24336_6544# ringtest_0.x4.net8 4.93e-19
C857 ringtest_0.x4.net2 ringtest_0.x4._12_ 0.10227f
C858 a_24800_5334# a_24926_5712# 0.005525f
C859 ringtest_0.x4._11_ a_23529_6422# 0.001495f
C860 a_19114_31955# muxtest_0.x1.x3.GP1 9.8e-19
C861 a_26808_5308# VDPWR 0.182123f
C862 ringtest_0.x4._15_ ringtest_0.x4._23_ 0.683594f
C863 ua[3] ui_in[3] 0.553118f
C864 a_24329_6640# a_24712_6422# 0.001632f
C865 ringtest_0.x4.net6 a_25149_4220# 0.211407f
C866 ringtest_0.x4._24_ ringtest_0.x4._09_ 0.151845f
C867 a_18662_32213# muxtest_0.x1.x3.GN1 0.128677f
C868 ringtest_0.x4._15_ a_26367_4790# 0.036316f
C869 muxtest_0.R7R8 ui_in[2] 0.054741f
C870 a_24895_4790# a_25149_4220# 0.002313f
C871 ringtest_0.x4.net7 a_26201_4790# 0.007864f
C872 a_24329_6640# ringtest_0.x4.net6 0.001597f
C873 a_13501_23906# a_13675_24012# 0.006584f
C874 muxtest_0.x1.x3.GN1 m2_18699_31802# 0.06935f
C875 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.025028f
C876 a_13501_23906# muxtest_0.x2.x2.GN3 1.07e-20
C877 muxtest_0.x2.x2.GN1 a_12425_24040# 1.22e-20
C878 a_12019_24012# muxtest_0.x2.x2.GN2 8.86e-19
C879 a_22116_4902# a_22021_4220# 1.66e-20
C880 muxtest_0.x2.x2.GN3 ua[2] 0.429994f
C881 a_21675_4790# a_22164_4362# 0.010312f
C882 a_24329_6640# a_24895_4790# 4.79e-20
C883 ringtest_0.x4._24_ a_26766_5712# 9.29e-19
C884 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP2 1.19e-20
C885 a_27065_5334# a_27273_4220# 9.49e-21
C886 ringtest_0.x4.net8 a_24986_5878# 1.76e-19
C887 ringtest_0.x3.nselect2 a_17231_12017# 9.77e-20
C888 a_23381_4584# VDPWR 0.2419f
C889 a_27233_5308# ringtest_0.x4.net11 1.16e-19
C890 ringtest_0.x4._11_ ringtest_0.x4._06_ 0.020042f
C891 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GN4 3.13e-20
C892 a_21675_9686# VDPWR 0.262851f
C893 a_22224_6244# a_22350_5878# 0.005525f
C894 a_21785_8054# a_21867_8054# 0.005167f
C895 a_21951_5878# ringtest_0.x4._21_ 2.75e-21
C896 a_26555_4790# VDPWR 0.079695f
C897 ringtest_0.x4.net9 a_27303_4246# 0.005829f
C898 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ui_in[6] 1.67e-19
C899 ringtest_0.x4._11_ a_24070_5852# 0.002559f
C900 ringtest_0.x4._19_ a_23770_5308# 8.51e-20
C901 muxtest_0.x1.x3.GP3 muxtest_0.R3R4 0.384927f
C902 a_24045_6654# VDPWR 0.175351f
C903 ringtest_0.x4.net6 a_24545_5878# 0.00514f
C904 a_21845_8816# ringtest_0.x4._11_ 9.54e-19
C905 ringtest_0.x4._12_ a_22399_8976# 0.023132f
C906 a_21852_8720# a_22245_8054# 0.011211f
C907 muxtest_0.x2.x2.GP2 m3_13302_19985# 0.005314f
C908 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR 0.637448f
C909 ringtest_0.x4.net6 a_25364_5878# 0.047825f
C910 ringtest_0.x4.net2 a_22245_8054# 3.45e-20
C911 ringtest_0.x4.counter[2] ua[1] 3.21e-19
C912 a_22097_5334# a_21509_4790# 0.002525f
C913 a_23381_4584# a_23467_4584# 0.006584f
C914 a_26627_4246# a_27273_4220# 0.016298f
C915 ringtest_0.x4._11_ a_23891_4790# 0.002312f
C916 a_25364_5878# a_24895_4790# 1.98e-20
C917 ringtest_0.x4.net11 a_25977_4220# 1.29e-21
C918 ringtest_0.x4._16_ a_21509_4790# 1.96e-20
C919 a_21233_5340# a_21767_5334# 0.002698f
C920 a_21852_9416# a_21845_9116# 0.966391f
C921 ringtest_0.counter7 a_25975_3867# 8.66e-19
C922 a_21465_9294# a_21981_9142# 1.28e-19
C923 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GP1 6.21e-20
C924 a_22392_5990# ringtest_0.x4.net5 1.47e-21
C925 ringtest_0.x4._11_ a_22373_5156# 0.045224f
C926 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP3 0.001226f
C927 muxtest_0.x1.x5.GN a_19242_32347# 1.08e-19
C928 muxtest_0.x1.x1.nSEL1 a_18836_32319# 0.00175f
C929 muxtest_0.R5R6 ui_in[2] 2.39e-19
C930 a_22265_5308# a_23770_5308# 1e-20
C931 ringtest_0.x4.net1 a_21675_9686# 0.073427f
C932 a_23879_6940# a_24883_6800# 8.9e-19
C933 ringtest_0.x4._15_ a_25593_5156# 1.98e-20
C934 ringtest_0.x4.net8 a_23899_5334# 2.79e-20
C935 ringtest_0.x4.net6 a_24551_4790# 7.29e-19
C936 ringtest_0.x4._11_ a_21767_5334# 3.45e-19
C937 ringtest_0.x4._16_ a_22765_5308# 0.243866f
C938 a_24336_6544# ringtest_0.x4._05_ 0.181338f
C939 ringtest_0.x4.counter[6] VDPWR 0.462317f
C940 a_24536_6699# a_24465_6800# 0.239923f
C941 a_24699_6200# VDPWR 0.2552f
C942 VDPWR ui_in[2] 4.46272f
C943 muxtest_0.R3R4 muxtest_0.R1R2 0.184502f
C944 a_21395_6940# a_21672_5334# 7.35e-19
C945 ringtest_0.x4.net6 a_24317_4942# 0.173962f
C946 muxtest_0.x2.x2.GN2 ui_in[4] 0.108808f
C947 ringtest_0.drv_out a_25393_5308# 1.4e-22
C948 a_22052_8875# VDPWR 0.271061f
C949 a_24317_4942# a_24895_4790# 0.00145f
C950 ringtest_0.x4.net9 ringtest_0.x4.counter[8] 2.39e-19
C951 ringtest_0.x4.net6 a_23151_5334# 7.79e-20
C952 ringtest_0.x4._15_ a_23993_5654# 0.004604f
C953 ringtest_0.x4.net8 ringtest_0.x4.counter[9] 1.68e-20
C954 ringtest_0.x4.net3 ringtest_0.x4._14_ 0.471315f
C955 a_27065_5334# a_26201_4790# 1.29e-19
C956 a_22116_4902# a_22541_5058# 1.28e-19
C957 a_27233_5308# ringtest_0.x4._09_ 5.87e-19
C958 a_21675_4790# a_22373_5156# 0.195152f
C959 ringtest_0.x4.net7 a_23770_5308# 0.142058f
C960 a_22399_8976# a_22245_8054# 6.31e-19
C961 a_21785_5878# a_24070_5852# 1.55e-21
C962 a_24479_4790# VDPWR 4.84e-19
C963 ringtest_0.x4._11_ a_26269_4612# 0.006396f
C964 ringtest_0.x4.clknet_0_clk a_26569_6422# 2.96e-20
C965 ringtest_0.x4._17_ a_23770_5308# 1.33e-19
C966 a_23809_4790# VDPWR 0.211123f
C967 a_21465_8830# a_21780_8964# 7.84e-20
C968 muxtest_0.x1.x3.GN3 muxtest_0.R6R7 0.260987f
C969 a_26201_5340# ringtest_0.x4.net10 4.73e-19
C970 ringtest_0.x4.net4 a_22021_4220# 0.021386f
C971 ringtest_0.x4.clknet_1_0__leaf_clk a_21561_8830# 0.044938f
C972 a_21981_9142# a_21981_8976# 0.013661f
C973 a_24045_6654# ringtest_0.x4._21_ 9.57e-19
C974 ringtest_0.x4._15_ ringtest_0.x4._04_ 3.75e-19
C975 a_22795_5334# VDPWR 0.261491f
C976 ringtest_0.x4._15_ a_25441_4612# 3.42e-21
C977 ringtest_0.x4.net1 a_22052_8875# 1.33e-19
C978 ringtest_0.x4._11_ a_22499_4790# 5.7e-19
C979 ringtest_0.drv_out ringtest_0.x3.x2.GN4 0.071598f
C980 a_26201_4790# a_26627_4246# 9.12e-19
C981 ringtest_0.x4._09_ a_25977_4220# 1.89e-19
C982 muxtest_0.x1.x4.A ua[0] 4.51511f
C983 a_21425_9686# a_21675_9686# 0.025037f
C984 a_21785_5878# a_22373_5156# 0.001131f
C985 ringtest_0.x4.net8 a_27149_5334# 2.29e-20
C986 ringtest_0.x4._04_ a_22541_5058# 7.11e-19
C987 ringtest_0.x4._07_ a_25393_5308# 0.008579f
C988 ringtest_0.x4._19_ ringtest_0.x4.net6 0.04173f
C989 a_21233_5340# a_21399_5340# 0.968904f
C990 ringtest_0.x4._22_ a_25225_5334# 1.1e-21
C991 ringtest_0.x4.net5 a_25149_4220# 1.18e-20
C992 ringtest_0.x4.clknet_1_0__leaf_clk a_22541_5058# 1.1e-19
C993 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.001676f
C994 ringtest_0.x4._18_ a_23949_6654# 0.006776f
C995 a_16579_11759# ringtest_0.x3.x2.GP2 3.07e-19
C996 a_21803_8598# VDPWR 0.004522f
C997 ringtest_0.x4._20_ a_25168_5156# 9.2e-20
C998 a_22649_6244# a_22765_5308# 0.001534f
C999 a_23879_6940# a_24045_6654# 0.017149f
C1000 m3_13302_19985# ua[0] 0.003764f
C1001 ringtest_0.x4._11_ a_21399_5340# 0.008371f
C1002 ringtest_0.x4.net10 a_27233_5058# 0.008159f
C1003 muxtest_0.x2.x2.GN1 ua[3] 4.69116f
C1004 muxtest_0.x1.x4.A a_13675_24012# 2.9e-19
C1005 ringtest_0.counter3 m3_17036_9140# 2.1e-20
C1006 ringtest_0.x4.net8 ringtest_0.x4._16_ 0.193029f
C1007 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN3 8.22e-19
C1008 a_24699_6200# ringtest_0.x4._21_ 0.001146f
C1009 ringtest_0.x4.counter[4] ringtest_0.x4.counter[5] 0.068962f
C1010 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[6] 5.64e-20
C1011 a_25421_6641# VDPWR 0.209324f
C1012 ringtest_0.x4.clknet_1_1__leaf_clk a_26367_5340# 0.026802f
C1013 ringtest_0.x4.net6 a_22265_5308# 6.37e-19
C1014 ringtest_0.x4.clknet_0_clk a_24287_6422# 2.01e-19
C1015 muxtest_0.x1.x3.GP2 muxtest_0.R6R7 4.11376f
C1016 muxtest_0.x2.x2.GP2 ua[0] 4.069f
C1017 ringtest_0.x4.net3 ringtest_0.x4._10_ 0.003052f
C1018 ringtest_0.x4.net11 ringtest_0.x4.counter[9] 0.066386f
C1019 ringtest_0.x4._22_ a_26640_5156# 0.004398f
C1020 a_21587_5334# a_21509_4790# 2.5e-19
C1021 ringtest_0.x4.net6 ringtest_0.x4.net9 0.566537f
C1022 ringtest_0.x4.clknet_1_0__leaf_clk a_21049_8598# 3.26e-19
C1023 ringtest_0.x4._23_ a_25975_3867# 2.99e-20
C1024 muxtest_0.x2.x2.GN3 m3_13302_19985# 0.087318f
C1025 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR 0.637284f
C1026 ringtest_0.x4._16_ a_24729_4790# 1.25e-20
C1027 a_21399_5340# a_21675_4790# 6.25e-19
C1028 ringtest_0.counter7 m3_17032_8096# 6.07e-21
C1029 ringtest_0.x4.net11 a_27491_4566# 0.001149f
C1030 ringtest_0.x4._24_ ringtest_0.x4._08_ 0.423487f
C1031 ringtest_0.x4.net9 a_24895_4790# 0.017191f
C1032 ringtest_0.x4._15_ ringtest_0.x4.net4 0.003757f
C1033 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP1 4.57902f
C1034 ringtest_0.x4._00_ a_21845_8816# 8.76e-20
C1035 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GN4 0.190572f
C1036 ringtest_0.x4._18_ a_24004_6128# 5.77e-19
C1037 a_23879_6940# a_24699_6200# 6.61e-19
C1038 ringtest_0.x4._21_ a_23809_4790# 0.087922f
C1039 a_19794_32347# VDPWR 0.001496f
C1040 a_25393_5308# a_26201_5340# 4.62e-19
C1041 a_20318_32213# muxtest_0.x1.x3.GN2 7.58e-21
C1042 muxtest_0.x1.x3.GN1 a_18836_32319# 0.001144f
C1043 a_25421_6641# ringtest_0.x4._25_ 6.03e-21
C1044 ringtest_0.x4._17_ a_24712_6422# 0.002153f
C1045 a_21672_5334# VDPWR 0.259474f
C1046 ringtest_0.x4.net6 ringtest_0.x4.net7 0.905861f
C1047 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP2 2.65608f
C1048 muxtest_0.x1.x1.nSEL1 a_19290_32287# 0.041068f
C1049 ringtest_0.x4.net4 a_22541_5058# 0.020834f
C1050 ringtest_0.x4.clknet_1_1__leaf_clk a_27065_5156# 2.2e-19
C1051 ringtest_0.ring_out ringtest_0.x3.nselect2 0.006614f
C1052 ringtest_0.x4.net7 a_24895_4790# 0.030766f
C1053 ringtest_0.x4.net3 a_21509_4790# 0.005671f
C1054 a_23949_6654# ringtest_0.x4.clknet_1_1__leaf_clk 1.77e-20
C1055 ringtest_0.x4._17_ ringtest_0.x4.net6 0.277113f
C1056 ringtest_0.x4.net2 ringtest_0.counter7 6.88e-20
C1057 muxtest_0.R7R8 muxtest_0.x2.x2.GP3 0.17349f
C1058 ringtest_0.x4._17_ a_24895_4790# 6.74e-21
C1059 a_16579_11759# a_16707_12151# 0.004764f
C1060 a_16579_11759# ringtest_0.x3.x2.GN2 1.63e-19
C1061 a_21785_5878# a_21399_5340# 1.36e-19
C1062 a_21951_5878# a_21233_5340# 9.16e-19
C1063 ringtest_0.x4._18_ a_23381_4818# 1.7e-19
C1064 ringtest_0.x4._23_ a_26367_5340# 0.031087f
C1065 a_22097_5334# a_22390_4566# 3.78e-21
C1066 ringtest_0.x4._24_ VDPWR 0.6956f
C1067 a_26367_5340# a_26367_4790# 0.027195f
C1068 a_26201_5340# a_26808_4902# 1.99e-20
C1069 ringtest_0.x4._16_ a_22390_4566# 3.76e-19
C1070 a_22649_6244# ringtest_0.x4.net8 3.5e-19
C1071 ringtest_0.x4._11_ a_21951_5878# 0.082924f
C1072 muxtest_0.x1.x5.A muxtest_0.R4R5 4.5151f
C1073 ringtest_0.x4.net3 a_21867_8054# 1.25e-19
C1074 a_24336_6544# a_24361_5340# 1.6e-20
C1075 a_24329_6640# a_24527_5340# 3.93e-19
C1076 ringtest_0.x4._15_ a_23837_5878# 9.44e-19
C1077 ringtest_0.x4._15_ ringtest_0.x4._22_ 0.422897f
C1078 ringtest_0.x4._11_ a_24883_6800# 7.39e-21
C1079 ringtest_0.x4._05_ ringtest_0.x4._16_ 0.001611f
C1080 ringtest_0.x4._07_ a_25083_4790# 0.128255f
C1081 ringtest_0.x4.net3 ringtest_0.x4._13_ 0.031667f
C1082 ringtest_0.x3.x2.GP2 m3_17032_8096# 0.005314f
C1083 ringtest_0.x4.clknet_0_clk a_24329_6640# 0.043419f
C1084 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP2 0.059353f
C1085 a_21465_9294# ringtest_0.x4._12_ 6.08e-20
C1086 ringtest_0.x4.net6 a_22817_6146# 0.129987f
C1087 ringtest_0.x4.clknet_1_1__leaf_clk a_24004_6128# 0.007927f
C1088 a_23891_4790# ringtest_0.x4.counter[4] 4.37e-20
C1089 ringtest_0.x4._14_ ringtest_0.x4._03_ 0.071143f
C1090 ringtest_0.x4._09_ a_27491_4566# 0.002954f
C1091 a_25083_4790# a_25055_3867# 7.39e-20
C1092 a_25593_5156# a_25975_3867# 3.85e-20
C1093 ringtest_0.x4._24_ ringtest_0.x4._25_ 0.095329f
C1094 a_16579_11759# ui_in[3] 0.086353f
C1095 ringtest_0.x4.net7 a_27169_6641# 2.85e-19
C1096 ringtest_0.x4._23_ a_27065_5156# 0.006274f
C1097 a_27233_5058# a_27191_4790# 7.84e-20
C1098 a_26808_4902# a_27233_5058# 1.28e-19
C1099 a_26367_4790# a_27065_5156# 0.194892f
C1100 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ui_in[4] 2.42e-19
C1101 ringtest_0.x4._06_ a_25393_5308# 1.75e-19
C1102 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.025028f
C1103 a_23879_6940# a_25421_6641# 1.59e-19
C1104 a_24699_6200# a_24968_5308# 1e-18
C1105 a_27815_3867# VDPWR 0.276039f
C1106 ringtest_0.x3.x2.GP3 ringtest_0.counter7 0.165274f
C1107 a_11845_23906# muxtest_0.x2.x2.GN2 0.039612f
C1108 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN3 0.012418f
C1109 a_22224_6244# VDPWR 0.255338f
C1110 ringtest_0.x4._08_ a_27233_5308# 0.004928f
C1111 ringtest_0.x4.clknet_1_1__leaf_clk a_23381_4818# 2.67e-20
C1112 a_22350_5878# ringtest_0.x4._16_ 2.63e-21
C1113 a_27149_5334# ringtest_0.x4._09_ 1.2e-19
C1114 a_26007_6788# VDPWR 0.001434f
C1115 ringtest_0.x4.clknet_0_clk a_25364_5878# 0.316676f
C1116 ringtest_0.x3.x1.nSEL0 a_15575_12017# 0.081627f
C1117 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.nselect2 0.047548f
C1118 muxtest_0.x2.x2.GP3 VDPWR 1.78328f
C1119 ringtest_0.x4._15_ a_25225_5334# 0.0351f
C1120 muxtest_0.R7R8 muxtest_0.R2R3 0.215077f
C1121 ringtest_0.x4._22_ a_26173_4612# 0.001961f
C1122 ringtest_0.x4._01_ a_21395_6940# 3.77e-19
C1123 muxtest_0.R7R8 ui_in[1] 4.98e-22
C1124 a_21785_5878# a_21951_5878# 0.966818f
C1125 a_16155_12151# VDPWR 2.96e-19
C1126 ringtest_0.x3.x2.GN1 VDPWR 1.47002f
C1127 a_21981_8976# ringtest_0.x4._12_ 0.039032f
C1128 ringtest_0.x4._11_ a_23381_4584# 0.002917f
C1129 a_22265_5308# ringtest_0.x4.net5 6.71e-21
C1130 muxtest_0.x1.x3.GP1 muxtest_0.x1.x4.A 0.354981f
C1131 muxtest_0.x2.x2.GN3 ua[0] 0.214839f
C1132 ringtest_0.x4._11_ a_26555_4790# 2.79e-20
C1133 ringtest_0.x3.x2.GN4 m3_17036_9140# 7.17e-19
C1134 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR 0.637855f
C1135 ringtest_0.x3.x2.GN2 m3_17032_8096# 0.016745f
C1136 ringtest_0.x4._17_ a_23932_6128# 0.002503f
C1137 a_24465_6800# ringtest_0.x4.net8 0.00192f
C1138 muxtest_0.x1.x5.GN muxtest_0.R7R8 0.558172f
C1139 ringtest_0.x4._11_ a_24045_6654# 1.82e-19
C1140 a_24361_5340# a_23899_5334# 1.44e-19
C1141 a_19666_31955# muxtest_0.x1.x3.GP1 1.19e-20
C1142 ringtest_0.x4.clknet_1_1__leaf_clk a_26375_4612# 5.67e-20
C1143 a_27233_5308# VDPWR 0.48745f
C1144 a_24536_6699# a_24712_6422# 0.007724f
C1145 ringtest_0.x4._15_ a_22021_4220# 3.5e-20
C1146 ringtest_0.x4.net6 a_26627_4246# 5.59e-20
C1147 a_19290_32287# muxtest_0.x1.x3.GN1 1.45e-19
C1148 ringtest_0.x4._15_ a_26640_5156# 0.001788f
C1149 a_25168_5156# a_25149_4220# 1.83e-19
C1150 VDPWR ui_in[6] 1.10022f
C1151 muxtest_0.x1.x5.A ui_in[2] 5.67943f
C1152 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x3.nselect2 2.88e-20
C1153 a_12977_24040# muxtest_0.x2.x2.GN4 3.22e-19
C1154 muxtest_0.x2.x2.GN3 a_13675_24012# 1.07e-20
C1155 a_24536_6699# ringtest_0.x4.net6 6.81e-19
C1156 a_25336_4902# a_25719_4790# 4.67e-20
C1157 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP3 0.031766f
C1158 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GN4 8.84e-19
C1159 a_21948_5156# a_22164_4362# 0.003601f
C1160 ua[3] ua[6] 0.008019f
C1161 muxtest_0.x2.x2.GP1 ui_in[4] 0.001143f
C1162 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._20_ 0.0051f
C1163 a_24329_6640# a_25168_5156# 7.91e-22
C1164 a_19114_31955# ui_in[2] 8.66e-20
C1165 a_12297_23648# ui_in[4] 0.03417f
C1166 ringtest_0.x3.nselect2 ringtest_0.x3.x2.GN3 7.39e-21
C1167 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN4 2.26e-20
C1168 a_21780_9142# VDPWR 4.59e-19
C1169 a_25977_4220# VDPWR 0.419035f
C1170 a_21785_8054# a_21395_6940# 5.68e-19
C1171 ringtest_0.x4._11_ ringtest_0.x4.counter[6] 0.002692f
C1172 ringtest_0.x4._10_ a_21939_8054# 5.49e-20
C1173 a_21561_9116# VDPWR 0.19379f
C1174 a_25719_4790# VDPWR 2.75e-19
C1175 ringtest_0.x4._11_ a_24699_6200# 0.042839f
C1176 uio_in[0] ui_in[7] 0.031023f
C1177 a_21509_4790# ringtest_0.x4._03_ 0.095111f
C1178 ringtest_0.x4._19_ a_24527_5340# 4.93e-21
C1179 a_24336_6544# VDPWR 0.321592f
C1180 ringtest_0.x4.net2 ringtest_0.x4._02_ 0.035742f
C1181 muxtest_0.x1.x3.GN4 muxtest_0.R3R4 0.237766f
C1182 ringtest_0.x4.net3 ringtest_0.x4.counter[1] 0.103986f
C1183 muxtest_0.R2R3 VDPWR 1.6072f
C1184 ringtest_0.x4.clknet_0_clk ringtest_0.x4._19_ 0.038005f
C1185 a_21465_8830# a_21845_8816# 0.048748f
C1186 VDPWR ui_in[1] 2.66846f
C1187 ringtest_0.x4._04_ a_22765_4478# 1.25e-20
C1188 ringtest_0.counter3 ua[1] 4.52195f
C1189 muxtest_0.x1.x5.GN muxtest_0.R5R6 7.03e-21
C1190 ringtest_0.x4.net3 a_22390_4566# 9.94e-20
C1191 a_25761_5058# ringtest_0.x4.counter[6] 4.54e-21
C1192 ringtest_0.x4.net8 a_26201_4790# 3.27e-19
C1193 ringtest_0.x4._23_ a_26375_4612# 1.08e-20
C1194 a_21981_9142# a_22201_9142# 4.62e-19
C1195 ringtest_0.x4._11_ a_24479_4790# 0.001677f
C1196 ringtest_0.x4.net11 a_27273_4220# 0.088145f
C1197 a_21845_9116# a_22052_9116# 0.273138f
C1198 a_21561_9116# a_21803_9508# 0.008508f
C1199 a_21852_9416# a_21981_9142# 0.110715f
C1200 ringtest_0.x4._18_ a_22392_5990# 1.41e-19
C1201 ringtest_0.counter7 a_27489_3702# 3.7e-19
C1202 a_21233_5340# a_22795_5334# 2.77e-19
C1203 ringtest_0.x4.net1 a_21780_9142# 2.14e-19
C1204 ringtest_0.x4._11_ a_23809_4790# 0.222369f
C1205 ringtest_0.x4._14_ a_21055_5334# 6.31e-19
C1206 ringtest_0.x4.clknet_1_1__leaf_clk a_26569_6422# 7.87e-19
C1207 muxtest_0.x1.x5.GN VDPWR 3.74211f
C1208 ringtest_0.x4.net1 a_21561_9116# 0.017118f
C1209 a_22111_10993# a_21852_9416# 4.65e-23
C1210 ringtest_0.x4._06_ a_24715_5334# 0.114717f
C1211 a_24986_5878# VDPWR 1.76e-19
C1212 ringtest_0.x4.net10 a_26895_3867# 2.65e-20
C1213 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[4] 8.27e-22
C1214 ringtest_0.x4._11_ a_22795_5334# 2.49e-20
C1215 ringtest_0.x4.net8 a_26555_5334# 1.28e-19
C1216 a_12849_23648# muxtest_0.x2.x2.GP3 0.00144f
C1217 ringtest_0.x4._16_ a_24361_5340# 1.57e-19
C1218 a_24465_6800# ringtest_0.x4._05_ 0.001005f
C1219 ringtest_0.x4.net9 a_24527_5340# 0.002182f
C1220 a_16707_12151# ringtest_0.x3.x2.GP3 4.39e-19
C1221 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.001676f
C1222 a_22139_5878# VDPWR 0.093135f
C1223 a_25336_4902# a_25677_5156# 9.73e-19
C1224 ua[2] ua[1] 1.12657f
C1225 a_24729_4790# a_26201_4790# 0.003146f
C1226 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP3 0.004296f
C1227 ringtest_0.x4._15_ a_22541_5058# 2.99e-20
C1228 muxtest_0.x2.nselect2 a_13025_23980# 6.01e-20
C1229 muxtest_0.x1.x1.nSEL0 ui_in[2] 0.131256f
C1230 ringtest_0.x4._01_ VDPWR 0.468919f
C1231 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net9 0.132797f
C1232 ringtest_0.x4._15_ a_24926_5712# 0.002542f
C1233 ringtest_0.x4._07_ a_25055_3867# 7.51e-19
C1234 ringtest_0.x4._22_ a_25975_3867# 2.78e-19
C1235 ringtest_0.x4._14_ a_22939_4584# 5.76e-19
C1236 ringtest_0.x4.net7 a_24527_5340# 0.456298f
C1237 ringtest_0.x4._04_ a_24004_6128# 3.15e-21
C1238 a_21007_3867# ringtest_0.x4.counter[0] 0.109791f
C1239 a_25677_5156# VDPWR 0.004788f
C1240 ringtest_0.x4._17_ a_24527_5340# 1.22e-20
C1241 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net7 0.043959f
C1242 a_21863_4790# VDPWR 0.083158f
C1243 muxtest_0.x1.x3.GN2 muxtest_0.R4R5 0.116214f
C1244 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR 0.637064f
C1245 a_26808_5308# ringtest_0.x4.net10 2.56e-19
C1246 ringtest_0.x4.clknet_1_0__leaf_clk a_21852_8720# 0.083453f
C1247 a_24336_6544# ringtest_0.x4._21_ 0.001538f
C1248 ringtest_0.x4.counter[4] ua[1] 3.21e-19
C1249 ringtest_0.x4._11_ a_25421_6641# 0.004334f
C1250 ringtest_0.x3.x2.GP3 ui_in[3] 2.82e-19
C1251 ringtest_0.x4.net4 a_22765_4478# 0.130038f
C1252 ringtest_0.x4.net2 ringtest_0.x4._04_ 4.09e-22
C1253 ringtest_0.x4.clknet_0_clk ringtest_0.x4._17_ 0.029087f
C1254 a_23899_5334# VDPWR 0.206364f
C1255 ringtest_0.x4.net6 a_26721_4246# 7.2e-20
C1256 ringtest_0.x4._15_ a_26173_4612# 0.006963f
C1257 ringtest_0.x4.net1 ringtest_0.x4._01_ 1.96e-19
C1258 a_25925_6788# ringtest_0.x4._24_ 4.18e-19
C1259 ringtest_0.x4._23_ a_26569_6422# 0.213625f
C1260 ringtest_0.x4.net2 ringtest_0.x4.clknet_1_0__leaf_clk 0.026712f
C1261 ringtest_0.x4._09_ a_27273_4220# 0.17213f
C1262 ringtest_0.x4._00_ a_21675_9686# 0.07841f
C1263 a_21425_9686# a_21561_9116# 7.31e-19
C1264 a_26749_6422# a_26201_4790# 3.35e-21
C1265 ringtest_0.x4._09_ a_26766_4790# 3.07e-19
C1266 a_26201_4790# ringtest_0.x4.net11 3.07e-19
C1267 ringtest_0.x4._02_ a_21840_5308# 4.65e-19
C1268 ringtest_0.x4._22_ a_26367_5340# 4.96e-21
C1269 a_21233_5340# a_21672_5334# 0.273138f
C1270 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x3.nselect2 5.69e-21
C1271 ringtest_0.x4._08_ a_27149_5334# 2.34e-19
C1272 ringtest_0.x4.counter[9] VDPWR 0.449609f
C1273 ringtest_0.x4._18_ a_24329_6640# 6.58e-19
C1274 a_23879_6940# a_24336_6544# 0.016444f
C1275 ringtest_0.x4.net8 a_23770_5308# 2.76e-19
C1276 a_21785_8054# VDPWR 0.266078f
C1277 ringtest_0.x4._20_ a_25593_5156# 1.2e-20
C1278 ringtest_0.x4.clknet_1_0__leaf_clk a_22181_5334# 3.7e-19
C1279 ringtest_0.x4._11_ a_21672_5334# 0.003174f
C1280 a_27491_4566# VDPWR 0.003335f
C1281 ringtest_0.x4._07_ ringtest_0.x4.counter[5] 1.62e-19
C1282 ringtest_0.counter3 m3_17046_7066# 8.01e-20
C1283 ringtest_0.x4.clknet_0_clk a_22817_6146# 3.43e-19
C1284 ringtest_0.drv_out m3_17036_9140# 0.132758f
C1285 muxtest_0.R7R8 ui_in[4] 0.104361f
C1286 a_25055_3867# ringtest_0.x4.counter[5] 0.1107f
C1287 ringtest_0.x4.clknet_1_1__leaf_clk a_26640_5334# 0.001015f
C1288 ringtest_0.x4.net6 a_22765_5308# 0.080758f
C1289 ringtest_0.x4.clknet_0_clk a_26095_6788# 9.17e-20
C1290 a_12019_24012# VDPWR 9.09e-19
C1291 ringtest_0.x4._11_ ringtest_0.x4._24_ 4.57e-19
C1292 ringtest_0.x4.clknet_1_0__leaf_clk a_22399_8976# 0.018091f
C1293 a_23949_6654# a_23837_5878# 2.76e-20
C1294 a_27273_4220# a_27659_4246# 0.006406f
C1295 ringtest_0.x4._23_ a_27489_3702# 9.55e-20
C1296 a_24329_6640# a_24763_6143# 0.00484f
C1297 ringtest_0.x4._14_ ringtest_0.x4.net5 0.258421f
C1298 ringtest_0.x4._16_ a_25336_4902# 8.82e-22
C1299 a_27149_5334# VDPWR 0.00533f
C1300 a_21399_5340# a_21948_5156# 0.002f
C1301 a_21672_5334# a_21675_4790# 0.004962f
C1302 ringtest_0.x4.net9 a_25168_5156# 0.003585f
C1303 ringtest_0.x4.net11 a_27303_4246# 0.01512f
C1304 a_26808_4902# a_26895_3867# 2.21e-20
C1305 ringtest_0.x4.net1 a_21785_8054# 0.232539f
C1306 ringtest_0.x4.net6 ringtest_0.x4._13_ 2.81e-21
C1307 a_25925_6788# a_26007_6788# 0.005781f
C1308 ringtest_0.x4.net2 ringtest_0.x4.net4 8.49e-21
C1309 a_22097_5334# a_22223_5712# 0.006169f
C1310 a_25225_5334# a_26367_5340# 8.68e-20
C1311 ringtest_0.x4.clknet_1_1__leaf_clk a_25149_4220# 1.84e-19
C1312 a_22097_5334# VDPWR 0.228175f
C1313 ringtest_0.x4.net4 a_23381_4818# 4.87e-19
C1314 muxtest_0.x1.x1.nSEL1 a_19842_32287# 1.59e-19
C1315 ringtest_0.x4._16_ VDPWR 2.17996f
C1316 a_26201_4790# ringtest_0.x4._09_ 0.098799f
C1317 ringtest_0.x4.net7 a_25168_5156# 0.005696f
C1318 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk 0.228247f
C1319 ringtest_0.x4._03_ a_22390_4566# 9.33e-19
C1320 a_22695_8304# VDPWR 0.006514f
C1321 ringtest_0.x3.x2.GN4 ua[1] 0.446629f
C1322 muxtest_0.x1.x3.GN2 ui_in[2] 0.001516f
C1323 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.025028f
C1324 a_24763_6143# a_24545_5878# 0.004465f
C1325 ringtest_0.x4._06_ ringtest_0.x4._07_ 5.11e-20
C1326 a_11845_23906# a_12297_23648# 0.002207f
C1327 a_16755_12091# ringtest_0.x3.x2.GN4 0.003699f
C1328 a_24004_6128# a_23837_5878# 0.046138f
C1329 a_17231_12017# ringtest_0.x3.x2.GN2 7.58e-21
C1330 a_21785_5878# a_21672_5334# 0.002054f
C1331 ringtest_0.x3.x2.GN1 a_15749_12123# 0.001144f
C1332 ringtest_0.x4._04_ a_21840_5308# 8.38e-20
C1333 ringtest_0.x4._14_ a_21007_3867# 0.001394f
C1334 ringtest_0.x4._23_ a_26640_5334# 0.012578f
C1335 ringtest_0.x4.clknet_1_0__leaf_clk a_21840_5308# 0.01796f
C1336 ringtest_0.x4._18_ a_23151_5334# 2.06e-20
C1337 a_26367_5340# a_26640_5156# 1.54e-19
C1338 a_26808_5308# a_26808_4902# 0.012451f
C1339 a_26640_5334# a_26367_4790# 1.54e-19
C1340 ringtest_0.x4._16_ a_23467_4584# 8.82e-20
C1341 ringtest_0.x4._11_ a_22224_6244# 0.054008f
C1342 a_21852_9416# ui_in[5] 4.56e-21
C1343 muxtest_0.x1.x4.A muxtest_0.R4R5 0.003925f
C1344 a_24465_6800# a_24361_5340# 5.48e-20
C1345 ringtest_0.x4.net3 a_21395_6940# 0.011213f
C1346 a_24536_6699# a_24527_5340# 8.21e-21
C1347 a_24329_6640# a_24800_5334# 8.34e-21
C1348 ringtest_0.x4._11_ a_26007_6788# 2.28e-19
C1349 ringtest_0.x4.clknet_1_1__leaf_clk a_24545_5878# 3.57e-20
C1350 ringtest_0.x4.net11 ringtest_0.x4.counter[8] 0.024563f
C1351 VDPWR ui_in[4] 9.60897f
C1352 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR 0.636224f
C1353 ringtest_0.x4.clknet_0_clk a_24536_6699# 0.004436f
C1354 ringtest_0.x4.clknet_1_1__leaf_clk a_25364_5878# 1.80017f
C1355 a_21425_9686# a_21785_8054# 2.44e-21
C1356 ringtest_0.x4.net6 ringtest_0.x4.net8 0.806426f
C1357 a_21852_9416# ringtest_0.x4._12_ 0.003541f
C1358 muxtest_0.x2.nselect2 ui_in[3] 1.88e-19
C1359 ringtest_0.x4._09_ a_27303_4246# 0.07143f
C1360 ringtest_0.x4.net8 a_24895_4790# 0.003497f
C1361 ringtest_0.x4._23_ a_25149_4220# 2.79e-19
C1362 a_17231_12017# ui_in[3] 0.220366f
C1363 a_23809_4790# ringtest_0.x4.counter[4] 2.6e-19
C1364 ringtest_0.x4._23_ a_26735_5156# 8.32e-19
C1365 a_26808_4902# a_26555_4790# 3.39e-19
C1366 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP1 8.08e-19
C1367 muxtest_0.R7R8 ui_in[0] 2.25e-21
C1368 ringtest_0.x4._06_ a_26201_5340# 4.19e-21
C1369 ringtest_0.x4.net10 a_26817_4566# 8.38e-19
C1370 ringtest_0.x4.net6 a_24729_4790# 0.083542f
C1371 ringtest_0.x4._18_ ringtest_0.x4._19_ 0.036736f
C1372 a_12473_23980# muxtest_0.x2.x2.GN2 0.017071f
C1373 a_22649_6244# VDPWR 0.169689f
C1374 a_24729_4790# a_24895_4790# 0.966391f
C1375 ringtest_0.x4.clknet_1_1__leaf_clk a_24317_4942# 0.050301f
C1376 ringtest_0.x4._21_ ringtest_0.x4._16_ 0.249175f
C1377 a_26201_6788# VDPWR 0.002272f
C1378 ringtest_0.x4._16_ ringtest_0.x4.counter[2] 3.86e-19
C1379 ringtest_0.x4.net4 a_21840_5308# 5.24e-19
C1380 ringtest_0.x4.clknet_1_1__leaf_clk a_23151_5334# 8.24e-20
C1381 ringtest_0.x3.x1.nSEL0 a_16203_12091# 0.001174f
C1382 ringtest_0.x4._15_ a_26367_5340# 0.058771f
C1383 a_21509_4790# ringtest_0.x4.net5 8.46e-19
C1384 ringtest_0.x4._03_ a_22074_4790# 0.001074f
C1385 ringtest_0.x4._22_ a_26375_4612# 2.76e-20
C1386 ringtest_0.x3.x2.GP1 VDPWR 1.86466f
C1387 ringtest_0.x4._04_ a_22392_5990# 0.04931f
C1388 a_21785_5878# a_22224_6244# 0.269567f
C1389 a_23467_4818# VDPWR 0.00273f
C1390 ringtest_0.x4._18_ a_22265_5308# 3.26e-20
C1391 ringtest_0.x4._11_ a_25977_4220# 0.19543f
C1392 a_22765_5308# ringtest_0.x4.net5 0.001034f
C1393 ringtest_0.x4._23_ a_25364_5878# 0.042503f
C1394 ringtest_0.x4.clknet_1_0__leaf_clk a_22392_5990# 5.16e-19
C1395 a_21852_9416# a_22245_8054# 6.42e-21
C1396 muxtest_0.x1.x3.GN1 ua[3] 4.34e-20
C1397 ringtest_0.x3.x2.GN4 m3_17046_7066# 0.084813f
C1398 ringtest_0.x4._11_ a_25719_4790# 2.44e-19
C1399 a_23837_5878# ringtest_0.x4._20_ 6.22e-20
C1400 a_25364_5878# a_26367_4790# 2.14e-19
C1401 a_19114_31955# ui_in[1] 0.03417f
C1402 a_23879_6940# ringtest_0.x4._16_ 4.51e-19
C1403 ringtest_0.x4._22_ ringtest_0.x4._20_ 2.69e-20
C1404 ringtest_0.counter7 ringtest_0.x4.net9 0.006102f
C1405 a_24361_5340# a_26555_5334# 2.33e-21
C1406 ringtest_0.x4._11_ a_24336_6544# 3.7e-19
C1407 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A 4.01025f
C1408 a_19242_32347# muxtest_0.x1.x3.GN3 5.17e-20
C1409 muxtest_0.x1.x3.GN2 a_19794_32347# 3.11e-20
C1410 a_21587_5334# VDPWR 0.075425f
C1411 ringtest_0.x4._15_ a_22765_4478# 1.84e-19
C1412 ringtest_0.ring_out ringtest_0.x3.x2.GP2 0.080385f
C1413 ringtest_0.x4.net6 a_26749_6422# 7.38e-20
C1414 a_19842_32287# muxtest_0.x1.x3.GN1 1.69e-20
C1415 a_25761_5058# a_25977_4220# 0.001105f
C1416 muxtest_0.x1.x5.GN a_19114_31955# 3.56e-19
C1417 muxtest_0.x1.x4.A ui_in[2] 4.96786f
C1418 ringtest_0.x4._05_ ringtest_0.x4.net6 0.03493f
C1419 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._19_ 0.060342f
C1420 a_23949_6654# ringtest_0.x4._15_ 1.78e-19
C1421 a_25761_5058# a_25719_4790# 7.84e-20
C1422 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ui_in[4] 4.96e-21
C1423 ringtest_0.x4._18_ ringtest_0.x4.net7 0.004371f
C1424 ringtest_0.counter7 ringtest_0.x4.net7 6.88e-20
C1425 a_22541_5058# a_22765_4478# 0.001036f
C1426 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.001676f
C1427 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 3.14e-21
C1428 ringtest_0.x4._24_ ringtest_0.x4.net10 0.13484f
C1429 a_19666_31955# ui_in[2] 0.009143f
C1430 VDPWR ui_in[0] 1.24711f
C1431 a_22139_5878# a_21233_5340# 3.23e-19
C1432 ringtest_0.x4._17_ ringtest_0.x4._18_ 0.181987f
C1433 muxtest_0.R3R4 muxtest_0.x2.x2.GN2 0.015374f
C1434 ringtest_0.x4.net9 a_24763_6143# 0.122363f
C1435 a_12849_23648# ui_in[4] 0.261734f
C1436 ringtest_0.x4.net3 VDPWR 2.1402f
C1437 a_27273_4220# VDPWR 0.230416f
C1438 a_24070_5852# ringtest_0.x4._06_ 0.004838f
C1439 a_21845_9116# VDPWR 0.721856f
C1440 a_22649_6244# ringtest_0.x4._21_ 8.88e-21
C1441 ringtest_0.x4.net8 a_23932_6128# 0.001644f
C1442 a_26766_4790# VDPWR -4.73e-35
C1443 ringtest_0.x4._11_ a_22139_5878# 0.020189f
C1444 a_27659_4246# ringtest_0.x4.counter[8] 1.28e-20
C1445 ringtest_0.x4._19_ a_24800_5334# 6.46e-21
C1446 a_24465_6800# VDPWR 0.191062f
C1447 ringtest_0.x4._01_ ringtest_0.x4._11_ 0.20957f
C1448 ringtest_0.x4._12_ ringtest_0.x4._10_ 0.002721f
C1449 ringtest_0.x4.net4 a_22392_5990# 0.034264f
C1450 ringtest_0.x4.net7 a_24763_6143# 1.85e-20
C1451 ringtest_0.x4._15_ a_24004_6128# 5.11e-20
C1452 a_21561_8830# a_21852_8720# 0.192341f
C1453 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net9 0.461828f
C1454 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR 0.636188f
C1455 ringtest_0.x4._23_ a_26913_4566# 2.44e-19
C1456 a_25149_4220# a_25441_4612# 0.001675f
C1457 ringtest_0.x4._17_ a_24763_6143# 2.72e-19
C1458 muxtest_0.x1.x1.nSEL0 ui_in[1] 0.137587f
C1459 a_25364_5878# a_25593_5156# 0.001605f
C1460 a_26749_6422# a_27169_6641# 0.017591f
C1461 ringtest_0.drv_out ua[1] 4.52048f
C1462 ringtest_0.x4.net2 a_21561_8830# 0.00144f
C1463 a_21465_9294# ringtest_0.x4.clknet_1_0__leaf_clk 0.007095f
C1464 ringtest_0.counter7 ringtest_0.x4.counter[0] 0.003899f
C1465 ringtest_0.x4._08_ a_26201_4790# 1.13e-19
C1466 a_22052_9116# a_21981_9142# 0.239923f
C1467 ringtest_0.x4._18_ a_22817_6146# 0.001543f
C1468 ringtest_0.x4.net1 ringtest_0.x4.net3 0.313425f
C1469 ringtest_0.x4.net8 ringtest_0.x4.net5 0.002187f
C1470 ringtest_0.x4._11_ a_21863_4790# 4.78e-19
C1471 ringtest_0.ring_out a_16707_12151# 2.99e-20
C1472 a_22111_10993# a_22052_9116# 2.02e-20
C1473 a_23770_5308# a_24361_5340# 0.044245f
C1474 ringtest_0.x4.net1 a_21845_9116# 0.003904f
C1475 ringtest_0.x4._19_ ringtest_0.x4._23_ 2.58e-20
C1476 ringtest_0.ring_out ringtest_0.x3.x2.GN2 0.23158f
C1477 ringtest_0.x4.net10 a_27815_3867# 0.219068f
C1478 ringtest_0.x4.net8 a_24895_5334# 4.84e-19
C1479 ringtest_0.x4.net6 ringtest_0.x4._09_ 1.5e-20
C1480 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net7 0.397702f
C1481 ringtest_0.x4._15_ a_23963_4790# 2.18e-19
C1482 ringtest_0.x4._11_ a_23899_5334# 0.07562f
C1483 muxtest_0.x2.x2.GP3 ua[2] 0.357853f
C1484 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x5.GN 0.043714f
C1485 ringtest_0.x4._16_ a_24968_5308# 0.001117f
C1486 ringtest_0.x4.net9 a_24800_5334# 6.38e-21
C1487 a_22733_6244# VDPWR 0.004177f
C1488 ringtest_0.x4._08_ a_26555_5334# 0.134213f
C1489 a_25168_5156# a_25294_4790# 0.005525f
C1490 ringtest_0.x4.clknet_0_clk a_22765_5308# 4.87e-21
C1491 ringtest_0.x4._15_ a_23381_4818# 0.22097f
C1492 ringtest_0.x4._17_ ringtest_0.x4.clknet_1_1__leaf_clk 0.044595f
C1493 ringtest_0.x4._23_ a_26735_5334# 8.32e-19
C1494 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN2 0.154394f
C1495 ringtest_0.x3.x2.GN3 ringtest_0.counter7 0.005062f
C1496 muxtest_0.R7R8 muxtest_0.x2.x2.GN4 3.97956f
C1497 a_22541_5058# a_23381_4818# 7.43e-20
C1498 a_21675_4790# a_21863_4790# 0.097994f
C1499 ringtest_0.x4._14_ a_22486_4246# 0.003598f
C1500 ringtest_0.x4.net7 a_24800_5334# 0.034093f
C1501 a_26201_4790# VDPWR 0.667506f
C1502 a_21785_5878# a_22139_5878# 0.062224f
C1503 ringtest_0.x4._10_ a_22245_8054# 0.423817f
C1504 a_21785_8054# ringtest_0.x4._11_ 0.005192f
C1505 uio_in[5] uio_in[4] 0.031023f
C1506 ringtest_0.ring_out ui_in[3] 3.69e-19
C1507 muxtest_0.x1.x3.GP3 ua[3] 0.023203f
C1508 ringtest_0.x4.net3 ringtest_0.x4.counter[2] 7.38e-19
C1509 a_11845_23906# VDPWR 0.211573f
C1510 ringtest_0.x4._23_ ringtest_0.x4.net9 0.065132f
C1511 ringtest_0.x4._17_ a_24800_5334# 9.6e-21
C1512 a_22457_5156# VDPWR 0.004797f
C1513 ringtest_0.x4.net9 a_26367_4790# 0.047741f
C1514 ua[3] ua[5] 0.008019f
C1515 a_23899_5654# a_23899_5334# 6.96e-20
C1516 a_27065_5334# a_27191_5712# 0.006169f
C1517 a_27233_5308# ringtest_0.x4.net10 0.084593f
C1518 ringtest_0.x4.clknet_1_0__leaf_clk a_21981_8976# 0.024273f
C1519 a_24465_6800# ringtest_0.x4._21_ 1.21e-19
C1520 a_26555_5334# VDPWR 0.078044f
C1521 ringtest_0.x4._15_ a_26375_4612# 0.002119f
C1522 ringtest_0.x4.net2 a_21049_8598# 0.07281f
C1523 a_19842_32287# muxtest_0.x1.x3.GP3 4.69e-19
C1524 muxtest_0.x2.x1.nSEL1 ui_in[2] 8.19e-21
C1525 a_19666_31955# a_19794_32347# 0.004764f
C1526 ringtest_0.x4.net7 ringtest_0.x4._23_ 0.074369f
C1527 a_21425_9686# a_21845_9116# 0.001828f
C1528 ringtest_0.x4._24_ a_26808_4902# 0.014122f
C1529 ringtest_0.x4._00_ a_21561_9116# 0.001635f
C1530 ringtest_0.x4.net7 a_26367_4790# 0.001362f
C1531 a_21233_5340# a_22097_5334# 0.032244f
C1532 ringtest_0.x4.net5 a_22390_4566# 0.075434f
C1533 ringtest_0.x4._02_ a_22265_5308# 1.8e-19
C1534 ringtest_0.counter7 a_26627_4246# 1.91e-19
C1535 ringtest_0.x4._17_ ringtest_0.x4._23_ 0.082072f
C1536 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ui_in[4] 4.96e-21
C1537 ringtest_0.x4._04_ a_23151_5334# 2.55e-19
C1538 ringtest_0.x4._15_ ringtest_0.x4._20_ 0.093509f
C1539 ringtest_0.x4._16_ a_21233_5340# 0.001516f
C1540 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP2 2.65608f
C1541 ringtest_0.x4._18_ a_24536_6699# 5.4e-20
C1542 ringtest_0.x4.net10 a_25977_4220# 0.158335f
C1543 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 7.08e-21
C1544 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.025028f
C1545 muxtest_0.R1R2 ua[3] 0.017912f
C1546 ringtest_0.x4.net8 a_24527_5340# 0.031957f
C1547 a_23879_6940# a_24465_6800# 0.013455f
C1548 ringtest_0.x4._11_ a_22097_5334# 0.017838f
C1549 a_27303_4246# VDPWR 0.283149f
C1550 ringtest_0.x3.x1.nSEL1 a_16707_12151# 4.08e-19
C1551 ringtest_0.x4._11_ ringtest_0.x4._16_ 0.223435f
C1552 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN2 0.209956f
C1553 a_22373_5156# a_22499_4790# 0.006169f
C1554 a_15575_12017# ringtest_0.x3.x2.GN1 0.12869f
C1555 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net8 8.45e-19
C1556 ringtest_0.x4._11_ a_22695_8304# 0.002858f
C1557 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A a_15575_12017# 6.58e-22
C1558 ringtest_0.x4.clknet_1_1__leaf_clk a_27065_5334# 1.84e-19
C1559 muxtest_0.x2.x2.GN4 VDPWR 1.23441f
C1560 ringtest_0.x4.net6 a_24361_5340# 0.0618f
C1561 a_21007_3867# ringtest_0.x4.counter[1] 0.057818f
C1562 ringtest_0.x4._22_ a_25149_4220# 0.106132f
C1563 a_24361_5340# a_24895_4790# 0.003047f
C1564 a_24527_5340# a_24729_4790# 0.003672f
C1565 muxtest_0.x1.x3.GN2 muxtest_0.R2R3 3.99837f
C1566 ringtest_0.x4.net3 a_21375_3867# 0.233128f
C1567 ringtest_0.x4.clknet_1_0__leaf_clk a_22228_8598# 0.002447f
C1568 a_24329_6640# ringtest_0.x4._22_ 1.01e-19
C1569 muxtest_0.x1.x3.GN2 ui_in[1] 0.108644f
C1570 ringtest_0.x4._03_ VDPWR 0.393273f
C1571 a_24536_6699# a_24763_6143# 3.7e-19
C1572 a_22265_5308# a_22116_4902# 0.001344f
C1573 ringtest_0.x4.net9 a_25593_5156# 0.031858f
C1574 a_22097_5334# a_21675_4790# 0.003824f
C1575 a_21672_5334# a_21948_5156# 4.47e-19
C1576 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR 0.638508f
C1577 ringtest_0.x4.counter[5] ua[1] 3.21e-19
C1578 ringtest_0.x4.clknet_0_clk a_24729_4790# 1.17e-21
C1579 ringtest_0.x4._00_ ringtest_0.x4._01_ 0.014628f
C1580 a_25925_6788# a_26201_6788# 0.00119f
C1581 m2_11882_23495# ui_in[4] 0.183786f
C1582 ringtest_0.x4._16_ a_21675_4790# 2.51e-21
C1583 ringtest_0.x3.x1.nSEL1 m2_15612_11606# 0.00815f
C1584 a_22765_5308# a_22983_5654# 0.007234f
C1585 a_26201_5340# a_26808_5308# 0.141453f
C1586 ringtest_0.x3.x1.nSEL1 ui_in[3] 0.168464f
C1587 ringtest_0.x4._15_ a_26569_6422# 0.001697f
C1588 a_23770_5308# VDPWR 0.17068f
C1589 a_24045_6654# a_24264_6788# 0.006169f
C1590 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN2 7.45e-19
C1591 ringtest_0.x4._16_ a_23899_5654# 0.001343f
C1592 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN1 0.034842f
C1593 ringtest_0.x4.net7 a_25593_5156# 0.040127f
C1594 ringtest_0.x4._03_ a_23467_4584# 5.07e-20
C1595 ringtest_0.x4.counter[8] VDPWR 0.228646f
C1596 a_12473_23980# muxtest_0.x2.x2.GP1 2.33e-21
C1597 a_24536_6699# ringtest_0.x4.clknet_1_1__leaf_clk 4.65e-20
C1598 a_21939_8054# VDPWR 3.14e-19
C1599 ringtest_0.x4.net4 a_23151_5334# 6.79e-19
C1600 ringtest_0.x4._22_ a_24545_5878# 9.75e-19
C1601 ringtest_0.x3.x2.GN3 a_16707_12151# 0.001073f
C1602 ringtest_0.x3.x2.GN2 a_17405_12123# 8.14e-21
C1603 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN4 0.001072f
C1604 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GN3 0.067463f
C1605 a_12297_23648# a_12473_23980# 0.185422f
C1606 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP3 0.005595f
C1607 a_21785_5878# a_22097_5334# 0.001393f
C1608 a_24699_6200# ringtest_0.x4._07_ 0.096566f
C1609 ringtest_0.x4._04_ a_22265_5308# 0.008333f
C1610 a_22074_4790# ringtest_0.x4.net5 3e-19
C1611 a_25364_5878# ringtest_0.x4._22_ 8.12e-19
C1612 ringtest_0.x4._14_ a_22295_3867# 4.42e-19
C1613 a_25225_5334# a_25149_4220# 3.32e-21
C1614 muxtest_0.x2.nselect2 ua[3] 0.005153f
C1615 a_21785_5878# ringtest_0.x4._16_ 6.86e-20
C1616 ringtest_0.x4.clknet_1_0__leaf_clk a_22265_5308# 0.002373f
C1617 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A a_16203_12091# 2.34e-20
C1618 a_26640_5334# a_26640_5156# 0.013839f
C1619 a_26367_5340# a_27065_5156# 1.3e-19
C1620 a_27065_5334# a_26367_4790# 1.3e-19
C1621 a_25055_3867# ringtest_0.x4.counter[6] 4.98e-19
C1622 ringtest_0.x4._11_ a_22649_6244# 0.043928f
C1623 ringtest_0.x4.net9 a_25441_4612# 6.97e-19
C1624 a_21951_5878# a_24070_5852# 8.39e-21
C1625 ringtest_0.x4._17_ a_23993_5654# 3.09e-20
C1626 a_22052_9116# ui_in[5] 1.46e-21
C1627 ringtest_0.x4._05_ a_24527_5340# 2.65e-21
C1628 ui_in[6] uio_in[0] 0.001316f
C1629 ringtest_0.x4._11_ a_26201_6788# 0.005861f
C1630 ringtest_0.x4.clknet_0_clk a_26749_6422# 1.5e-20
C1631 muxtest_0.x1.x3.GP1 muxtest_0.R4R5 0.123828f
C1632 muxtest_0.x2.x2.GP3 m3_13302_19985# 0.002824f
C1633 ringtest_0.x4._13_ a_21591_6128# 0.01129f
C1634 ringtest_0.ring_out a_17377_14114# 0.105448f
C1635 muxtest_0.x1.x3.GN3 muxtest_0.R7R8 0.129382f
C1636 ringtest_0.x4.net1 a_21939_8054# 0.002601f
C1637 ringtest_0.x4.clknet_0_clk ringtest_0.x4._05_ 0.067252f
C1638 a_22052_9116# ringtest_0.x4._12_ 5.69e-20
C1639 ringtest_0.x4._07_ a_23809_4790# 1.81e-20
C1640 a_17405_12123# ui_in[3] 1.4e-19
C1641 ringtest_0.x3.x2.GN3 ui_in[3] 0.254198f
C1642 ringtest_0.x4.net8 a_25168_5156# 0.001808f
C1643 ringtest_0.x4._23_ a_26627_4246# 0.04546f
C1644 ringtest_0.x4.net7 a_25441_4612# 0.006602f
C1645 ringtest_0.x4.net6 ringtest_0.x4._08_ 5.42e-20
C1646 ringtest_0.drv_out a_25421_6641# 0.012863f
C1647 ringtest_0.x4._11_ a_23467_4818# 0.003027f
C1648 ringtest_0.x4._17_ ringtest_0.x4._04_ 6.62e-21
C1649 a_26367_4790# a_26627_4246# 0.008374f
C1650 ringtest_0.x4.net10 ringtest_0.x4.counter[9] 0.092658f
C1651 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP3 0.031766f
C1652 a_21233_5340# a_21587_5334# 0.062224f
C1653 a_22392_5990# a_22541_5058# 8.5e-21
C1654 a_21951_5878# a_22373_5156# 0.001133f
C1655 a_26640_5156# a_26735_5156# 0.007724f
C1656 a_22224_6244# a_21948_5156# 9.19e-21
C1657 a_26367_4790# a_27149_5156# 6.32e-19
C1658 a_23899_5334# ringtest_0.x4.counter[4] 4.47e-20
C1659 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._17_ 3.38e-20
C1660 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ui_in[4] 4.1e-20
C1661 ringtest_0.x4.net10 a_27491_4566# 0.002502f
C1662 ringtest_0.x4.clknet_1_1__leaf_clk a_25294_4790# 4.82e-19
C1663 ringtest_0.x4.net6 a_25336_4902# 6.78e-21
C1664 ringtest_0.x4._11_ a_21587_5334# 2.52e-19
C1665 ringtest_0.x4._21_ a_23770_5308# 0.005326f
C1666 a_12849_23648# muxtest_0.x2.x2.GN4 6.84e-19
C1667 a_25364_5878# a_25225_5334# 5.73e-19
C1668 muxtest_0.R3R4 muxtest_0.x2.x2.GP1 0.011522f
C1669 a_13025_23980# muxtest_0.x2.x2.GN2 5.62e-20
C1670 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.001676f
C1671 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 1.11e-20
C1672 a_24895_4790# a_25336_4902# 0.110715f
C1673 a_24729_4790# a_25168_5156# 0.273138f
C1674 a_19114_31955# ui_in[0] 0.246193f
C1675 a_24712_6422# VDPWR 0.004407f
C1676 ringtest_0.counter3 ringtest_0.x4._16_ 1.05e-19
C1677 ringtest_0.x4.net4 a_22265_5308# 0.110738f
C1678 ringtest_0.x4.counter[5] ringtest_0.x4.counter[6] 0.070133f
C1679 ringtest_0.x4._15_ a_26640_5334# 0.001174f
C1680 ringtest_0.x3.x1.nSEL0 a_16755_12091# 1.21e-20
C1681 ringtest_0.x4.net3 a_21233_5340# 0.023332f
C1682 ringtest_0.x4._22_ a_26913_4566# 3.67e-19
C1683 ringtest_0.x4.net6 VDPWR 3.11824f
C1684 muxtest_0.x1.x4.A muxtest_0.R2R3 4.52053f
C1685 ringtest_0.x4._04_ a_22817_6146# 0.003723f
C1686 ringtest_0.x4.net10 a_27149_5334# 3.67e-19
C1687 a_21785_5878# a_22649_6244# 0.030894f
C1688 a_24895_4790# VDPWR 0.323392f
C1689 ringtest_0.x4.net3 ringtest_0.x4._11_ 0.005186f
C1690 ringtest_0.x4._18_ a_22765_5308# 0.002375f
C1691 ringtest_0.x4._11_ a_27273_4220# 2.01e-20
C1692 muxtest_0.x1.x3.GP2 muxtest_0.R7R8 0.131352f
C1693 a_23879_6940# a_23770_5308# 4.81e-21
C1694 ringtest_0.x4._19_ ringtest_0.x4._22_ 7e-20
C1695 ringtest_0.x4.clknet_1_0__leaf_clk a_22817_6146# 1.77e-20
C1696 muxtest_0.x1.x3.GN3 muxtest_0.R5R6 4.12612f
C1697 a_21845_9116# ringtest_0.x4._11_ 8.58e-21
C1698 ringtest_0.x4._11_ a_26766_4790# 4.03e-21
C1699 a_25364_5878# a_26640_5156# 6.58e-20
C1700 a_27169_6641# ringtest_0.x4._08_ 0.109717f
C1701 a_19666_31955# ui_in[1] 0.261734f
C1702 a_24361_5340# a_24895_5334# 0.001632f
C1703 ringtest_0.x4._11_ a_24465_6800# 5.19e-20
C1704 a_24045_6654# a_24070_5852# 0.006438f
C1705 a_21465_9294# a_21561_8830# 6.79e-19
C1706 a_21561_9116# a_21465_8830# 6.79e-19
C1707 a_23949_6654# a_24004_6128# 3.4e-19
C1708 muxtest_0.x1.x5.GN muxtest_0.x1.x4.A 4.14763f
C1709 a_21055_5334# VDPWR 0.006911f
C1710 muxtest_0.x1.x3.GN3 VDPWR 0.766397f
C1711 ringtest_0.x4._15_ a_25149_4220# 1.2e-20
C1712 ringtest_0.x4._19_ a_23619_6788# 8.17e-20
C1713 ringtest_0.x4.net6 ringtest_0.x4._25_ 2.22e-20
C1714 ringtest_0.x4._17_ ringtest_0.x4.net4 9.08e-20
C1715 ringtest_0.x4.net2 a_21507_9686# 0.00492f
C1716 muxtest_0.x1.x5.GN a_19666_31955# 3.51e-19
C1717 a_21509_4790# a_22295_3867# 8.97e-21
C1718 a_24329_6640# ringtest_0.x4._15_ 3.85e-20
C1719 ringtest_0.x4._14_ ringtest_0.x4._02_ 0.166596f
C1720 muxtest_0.x1.x3.GP1 ui_in[2] 5.64e-19
C1721 ringtest_0.x4.net3 a_21675_4790# 0.00115f
C1722 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GP1 6.21e-20
C1723 ringtest_0.x4._16_ a_22775_5878# 4.87e-20
C1724 a_16579_11759# ringtest_0.x3.x2.GP3 0.00144f
C1725 ringtest_0.x4.net9 ringtest_0.x4._22_ 0.369389f
C1726 a_13501_23906# ui_in[4] 0.125445f
C1727 ui_in[4] ua[2] 0.936267f
C1728 a_21951_5878# a_21399_5340# 5.5e-20
C1729 muxtest_0.x2.x1.nSEL0 a_12297_23648# 0.03096f
C1730 muxtest_0.x1.x1.nSEL0 ui_in[0] 0.325407f
C1731 a_22939_4584# VDPWR 3.83e-21
C1732 a_24699_6200# ringtest_0.x4._06_ 0.003245f
C1733 ringtest_0.x4._16_ a_23399_3867# 3.59e-21
C1734 a_27169_6641# VDPWR 0.28996f
C1735 a_21981_9142# VDPWR 0.211499f
C1736 ringtest_0.x4._11_ a_22733_6244# 0.002344f
C1737 a_22111_10993# VDPWR 0.305606f
C1738 ringtest_0.x4.clknet_1_1__leaf_clk a_22765_5308# 1.5e-19
C1739 ringtest_0.x4.net4 a_22817_6146# 7.5e-19
C1740 muxtest_0.x1.x3.GP2 muxtest_0.R5R6 0.312699f
C1741 muxtest_0.x2.x2.GP3 ua[0] 0.050476f
C1742 ringtest_0.x4.net7 ringtest_0.x4._22_ 0.179589f
C1743 ringtest_0.x4.net3 a_21785_5878# 1.48e-19
C1744 ringtest_0.x3.nselect2 VDPWR 1.23654f
C1745 ringtest_0.x4.net6 ringtest_0.x4._21_ 0.083542f
C1746 ringtest_0.x4._15_ a_25364_5878# 0.047247f
C1747 a_21561_8830# a_21981_8976# 0.036838f
C1748 a_21845_8816# a_22052_8875# 0.260055f
C1749 a_21465_8830# ringtest_0.x4._01_ 1.56e-19
C1750 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B a_17377_14114# 0.110771f
C1751 ringtest_0.x4._17_ a_23837_5878# 0.060488f
C1752 ringtest_0.x4._23_ a_26721_4246# 0.038842f
C1753 ringtest_0.x4._17_ ringtest_0.x4._22_ 1.76e-19
C1754 a_22390_4566# a_22486_4246# 0.002032f
C1755 ringtest_0.x4._11_ a_26201_4790# 0.012822f
C1756 a_11845_23906# m2_11882_23495# 0.01297f
C1757 ringtest_0.x4._14_ a_22116_4902# 1.1e-19
C1758 ringtest_0.x4.clknet_1_0__leaf_clk a_22201_9142# 0.002297f
C1759 ringtest_0.x3.x2.GP1 ringtest_0.counter3 5.62e-21
C1760 muxtest_0.x1.x3.GP2 VDPWR 3.26769f
C1761 a_27169_6641# ringtest_0.x4._25_ 0.227897f
C1762 a_26367_4790# a_26721_4246# 1.65e-19
C1763 a_21845_9116# a_22399_9142# 0.062224f
C1764 ringtest_0.x4.net2 a_21852_8720# 8.79e-19
C1765 ringtest_0.x4._18_ ringtest_0.x4.net8 0.01511f
C1766 a_22052_9116# a_22228_9508# 0.007724f
C1767 a_21852_9416# ringtest_0.x4.clknet_1_0__leaf_clk 0.470509f
C1768 a_21981_9142# a_21803_9508# 9.73e-19
C1769 ringtest_0.counter7 ringtest_0.x4.net8 6.32e-19
C1770 ringtest_0.x4.net7 a_23619_6788# 5.91e-19
C1771 ringtest_0.x4._11_ a_22457_5156# 0.002515f
C1772 a_24070_5852# a_23809_4790# 7.94e-19
C1773 ringtest_0.x4.net1 a_21981_9142# 0.002441f
C1774 a_24361_5340# a_24527_5340# 0.961627f
C1775 ringtest_0.drv_out ringtest_0.x3.x2.GN1 3.11e-19
C1776 ringtest_0.x4._17_ a_23619_6788# 7.93e-19
C1777 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 2.86851f
C1778 a_22111_10993# ringtest_0.x4.net1 0.10983f
C1779 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ui_in[4] 0.008686f
C1780 ringtest_0.x4.net9 a_25225_5334# 0.002503f
C1781 a_23932_6128# VDPWR 0.011634f
C1782 a_25761_5058# a_26201_4790# 0.001745f
C1783 ringtest_0.x4.clknet_0_clk a_24361_5340# 0.009291f
C1784 ringtest_0.x4._15_ a_24317_4942# 2.8e-19
C1785 a_23879_6940# ringtest_0.x4.net6 8.49e-19
C1786 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 1.99e-20
C1787 ua[0] ui_in[6] 0.619336f
C1788 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.025028f
C1789 a_23949_6654# ringtest_0.x4._20_ 1.63e-20
C1790 a_23809_4790# a_23891_4790# 0.005167f
C1791 a_22817_6146# a_23837_5878# 3.28e-20
C1792 ringtest_0.x4._04_ ringtest_0.x4._14_ 4.63e-22
C1793 a_22649_6244# a_22775_5878# 0.006169f
C1794 a_21395_6940# ringtest_0.x4.clknet_0_clk 0.317755f
C1795 a_15575_12017# ui_in[4] 0.02803f
C1796 ringtest_0.x4._24_ a_26201_5340# 0.031818f
C1797 ringtest_0.x4.net8 a_24763_6143# 0.003744f
C1798 a_21948_5156# a_21863_4790# 0.037333f
C1799 a_21675_4790# a_22457_5156# 3.14e-19
C1800 ringtest_0.x3.x1.nSEL1 a_16027_11759# 0.073392f
C1801 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A a_16755_12091# 9.97e-21
C1802 ringtest_0.x4.net7 a_25225_5334# 0.054488f
C1803 a_22265_5308# a_22021_4220# 2.52e-20
C1804 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._14_ 0.088295f
C1805 muxtest_0.R7R8 muxtest_0.R3R4 5.65992f
C1806 ringtest_0.x4._12_ a_21395_6940# 4.42e-19
C1807 a_12473_23980# VDPWR 0.193262f
C1808 ringtest_0.x4.net3 ringtest_0.counter3 6.21e-20
C1809 ringtest_0.x4._17_ a_25225_5334# 8.73e-21
C1810 ringtest_0.x4.clknet_1_0__leaf_clk a_22319_6244# 4.17e-19
C1811 muxtest_0.x1.x3.GN4 ua[3] 0.014367f
C1812 a_21132_8918# ringtest_0.x4._12_ 0.001776f
C1813 a_21852_8720# a_22399_8976# 0.099725f
C1814 a_21465_8830# a_21785_8054# 3.66e-19
C1815 a_22052_8875# a_22201_8964# 0.005525f
C1816 ringtest_0.x4.net5 VDPWR 0.923749f
C1817 ringtest_0.x4.net9 a_26640_5156# 0.023502f
C1818 ringtest_0.x3.x2.GP3 m3_17032_8096# 0.002824f
C1819 a_12977_24040# ui_in[3] 0.001558f
C1820 a_24895_5334# VDPWR 0.004219f
C1821 muxtest_0.x1.x3.GN4 a_20492_32319# 0.001562f
C1822 muxtest_0.x2.x2.GN2 ui_in[3] 0.11443f
C1823 ringtest_0.x4._02_ a_21509_4790# 3.71e-19
C1824 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net8 0.073766f
C1825 ringtest_0.x4.net2 a_22399_8976# 1.01e-21
C1826 a_21233_5340# ringtest_0.x4._03_ 0.001727f
C1827 ringtest_0.x4._15_ a_26913_4566# 0.001637f
C1828 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP3 0.075682f
C1829 muxtest_0.R2R3 ua[0] 2.39e-19
C1830 ringtest_0.counter7 ringtest_0.x4.counter[1] 0.003115f
C1831 a_24004_6128# ringtest_0.x4._20_ 4.3e-20
C1832 a_19842_32287# muxtest_0.x1.x3.GN4 0.003645f
C1833 ringtest_0.x4._24_ a_27233_5058# 0.009415f
C1834 ringtest_0.x4._00_ a_21845_9116# 0.118744f
C1835 ringtest_0.x4._11_ ringtest_0.x4._03_ 0.00174f
C1836 ringtest_0.x4._19_ ringtest_0.x4._15_ 6.2e-22
C1837 ringtest_0.x4.net7 a_26640_5156# 4.39e-19
C1838 ringtest_0.x4._02_ a_22765_5308# 7.66e-20
C1839 ringtest_0.x4.net5 a_23467_4584# 0.001706f
C1840 ringtest_0.x4.clknet_1_0__leaf_clk a_22043_5156# 5.04e-19
C1841 ringtest_0.counter7 ringtest_0.x4.net11 1.31e-19
C1842 ringtest_0.x4.clknet_1_1__leaf_clk a_24729_4790# 0.319108f
C1843 ringtest_0.x4.net10 a_27273_4220# 0.104575f
C1844 ringtest_0.x4._18_ ringtest_0.x4._05_ 1.11e-19
C1845 ringtest_0.x4.net8 a_24800_5334# 0.003635f
C1846 ringtest_0.x4._20_ a_23963_4790# 0.001506f
C1847 muxtest_0.x1.x3.GN2 ui_in[0] 0.114399f
C1848 ringtest_0.x4._11_ a_23770_5308# 0.058411f
C1849 a_21007_3867# VDPWR 0.25802f
C1850 ringtest_0.x3.x2.GN4 ui_in[4] 0.059808f
C1851 ringtest_0.x4._08_ a_24527_5340# 8.29e-20
C1852 a_16027_11759# ringtest_0.x3.x2.GN3 6.68e-19
C1853 a_16203_12091# ringtest_0.x3.x2.GN1 1.46e-19
C1854 ringtest_0.x4._13_ ringtest_0.x4._02_ 0.053355f
C1855 a_23381_4818# ringtest_0.x4._20_ 3.41e-19
C1856 ringtest_0.x4.net4 ringtest_0.x4._14_ 0.209869f
C1857 ringtest_0.x4._11_ a_21939_8054# 2.12e-19
C1858 ringtest_0.x4.net6 a_24968_5308# 0.012704f
C1859 ringtest_0.x4._03_ a_21675_4790# 0.260627f
C1860 a_21509_4790# a_22116_4902# 0.141453f
C1861 muxtest_0.x1.x4.A ui_in[4] 0.034362f
C1862 ringtest_0.x4._15_ a_22265_5308# 1.37e-19
C1863 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.173286f
C1864 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x1.nSEL0 1.14e-19
C1865 ringtest_0.x4._22_ a_26627_4246# 0.140356f
C1866 a_24968_5308# a_24895_4790# 0.001607f
C1867 a_24361_5340# a_25168_5156# 4.58e-19
C1868 a_24800_5334# a_24729_4790# 2.14e-19
C1869 a_24527_5340# a_25336_4902# 6.74e-19
C1870 ringtest_0.x4._15_ ringtest_0.x4.net9 0.08758f
C1871 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._10_ 0.006812f
C1872 muxtest_0.R3R4 VDPWR 3.2635f
C1873 ringtest_0.x4._16_ a_25083_4790# 1.98e-21
C1874 ringtest_0.x4._23_ ringtest_0.x4.net8 0.011201f
C1875 ringtest_0.x4._05_ a_24763_6143# 2.43e-19
C1876 a_22097_5334# a_21948_5156# 0.001152f
C1877 a_22265_5308# a_22541_5058# 0.007214f
C1878 ringtest_0.x4.net8 a_26367_4790# 1.04e-19
C1879 ringtest_0.x4.clknet_0_clk a_25336_4902# 8.09e-19
C1880 ringtest_0.x4._16_ a_21948_5156# 2.79e-19
C1881 ringtest_0.x4._21_ ringtest_0.x4.net5 2.83e-22
C1882 a_21672_5334# a_21767_5334# 0.007724f
C1883 a_23770_5308# a_23899_5654# 0.010132f
C1884 a_21840_5308# a_22181_5334# 9.73e-19
C1885 a_26201_5340# a_27233_5308# 0.048748f
C1886 a_26367_5340# a_26640_5334# 0.078545f
C1887 a_24527_5340# VDPWR 0.300379f
C1888 ringtest_0.x4.net7 ringtest_0.x4._15_ 0.590844f
C1889 ringtest_0.x4.clknet_1_1__leaf_clk a_26749_6422# 3.65e-19
C1890 ringtest_0.x4.net6 a_25925_6788# 0.157729f
C1891 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net11 1.82e-20
C1892 VDPWR ui_in[5] 0.255037f
C1893 ringtest_0.x4._04_ a_21509_4790# 2.08e-19
C1894 a_21785_5878# ringtest_0.x4._03_ 4.31e-20
C1895 ringtest_0.x4.net7 a_25263_5156# 5.23e-19
C1896 ringtest_0.x4._23_ a_24729_4790# 3.56e-21
C1897 a_13025_23980# muxtest_0.x2.x2.GP1 2.87e-20
C1898 ringtest_0.x4._17_ ringtest_0.x4._15_ 0.083602f
C1899 ringtest_0.x4._05_ ringtest_0.x4.clknet_1_1__leaf_clk 0.143201f
C1900 ringtest_0.x4.clknet_0_clk VDPWR 2.53166f
C1901 muxtest_0.x2.x2.GP2 ui_in[4] 4.34e-19
C1902 a_24729_4790# a_26367_4790# 8.05e-21
C1903 ringtest_0.x4.clknet_1_0__leaf_clk a_21509_4790# 0.293401f
C1904 ua[3] ua[4] 0.008019f
C1905 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP1 8.08e-19
C1906 ringtest_0.counter7 ringtest_0.x4._09_ 5.27e-21
C1907 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 5.48e-19
C1908 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y 0.001676f
C1909 muxtest_0.x2.x1.nSEL1 a_12019_24012# 0.00175f
C1910 a_12473_23980# a_12849_23648# 3.02e-19
C1911 ringtest_0.x4._12_ VDPWR 0.307826f
C1912 ringtest_0.x4._04_ a_22765_5308# 0.171873f
C1913 ringtest_0.x4.counter[9] ua[0] 0.004138f
C1914 ringtest_0.x4.net10 a_26201_4790# 0.001924f
C1915 a_27191_5712# ringtest_0.x4._09_ 1.66e-19
C1916 ringtest_0.x4.net7 a_24926_5712# 2.79e-19
C1917 ringtest_0.x4.clknet_1_0__leaf_clk a_22765_5308# 1.95e-19
C1918 a_27233_5308# a_27233_5058# 0.026048f
C1919 ringtest_0.x4._05_ a_24800_5334# 6.05e-21
C1920 ringtest_0.x4.net6 a_21233_5340# 1.88e-19
C1921 ringtest_0.x4._13_ ringtest_0.x4._04_ 1.41e-19
C1922 ringtest_0.x4.clknet_1_0__leaf_clk a_21867_8054# 2.61e-19
C1923 ringtest_0.x4.net1 ui_in[5] 0.067291f
C1924 a_26555_5334# ringtest_0.x4.net10 6.3e-20
C1925 muxtest_0.x2.x1.nSEL0 VDPWR 0.523833f
C1926 ringtest_0.x4._22_ a_25294_4790# 6.82e-19
C1927 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A 0.429924f
C1928 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._13_ 0.02176f
C1929 ringtest_0.x4.counter[6] ua[1] 3.21e-19
C1930 ringtest_0.x4._11_ ringtest_0.x4.net6 2.01574f
C1931 ringtest_0.x3.x2.GN1 m3_17036_9140# 6.03e-20
C1932 ringtest_0.x4.net1 ringtest_0.x4._12_ 0.312817f
C1933 ringtest_0.x4.net7 a_26173_4612# 6.49e-19
C1934 ringtest_0.x4.net8 a_25593_5156# 0.007067f
C1935 ringtest_0.x4._11_ a_24895_4790# 0.042209f
C1936 ringtest_0.x4._23_ a_26749_6422# 0.007723f
C1937 ringtest_0.x4._23_ ringtest_0.x4.net11 0.257634f
C1938 a_26640_5156# a_26627_4246# 2.47e-19
C1939 a_19114_31955# muxtest_0.x1.x3.GN3 6.68e-19
C1940 a_21233_5340# a_21055_5334# 5.87e-19
C1941 a_26749_6422# a_26367_4790# 3.03e-21
C1942 muxtest_0.R4R5 ui_in[2] 6.76e-20
C1943 a_26808_4902# a_26766_4790# 4.62e-19
C1944 a_22224_6244# a_22373_5156# 1.06e-19
C1945 a_26367_4790# ringtest_0.x4.net11 2.58e-19
C1946 a_18662_32213# VDPWR 0.213938f
C1947 ringtest_0.x4._05_ ringtest_0.x4._23_ 9.36e-20
C1948 a_21399_5340# a_21672_5334# 0.078737f
C1949 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._09_ 0.003413f
C1950 ringtest_0.x4.net4 a_21509_4790# 0.008383f
C1951 ringtest_0.x4.net10 a_27303_4246# 0.001384f
C1952 ringtest_0.x4.net6 a_25761_5058# 3.96e-21
C1953 m2_18699_31802# VDPWR 0.140918f
C1954 a_13501_23906# muxtest_0.x2.x2.GN4 0.134079f
C1955 muxtest_0.x2.x2.GN2 a_12425_24040# 0.002418f
C1956 muxtest_0.x2.x2.GN4 ua[2] 0.446579f
C1957 a_25364_5878# a_26367_5340# 0.008007f
C1958 ringtest_0.x4._21_ a_24527_5340# 0.002388f
C1959 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN2 0.065156f
C1960 a_23949_6654# a_24329_6640# 0.048635f
C1961 a_22245_8054# VDPWR 0.292813f
C1962 a_24895_4790# a_25761_5058# 0.034054f
C1963 a_24729_4790# a_25593_5156# 0.032244f
C1964 a_25336_4902# a_25168_5156# 0.239923f
C1965 a_19666_31955# ui_in[0] 0.086357f
C1966 ringtest_0.x4.net4 a_22765_5308# 0.005124f
C1967 muxtest_0.x2.x1.nSEL1 ui_in[4] 0.275874f
C1968 muxtest_0.x1.x3.GP3 muxtest_0.R1R2 4.25867f
C1969 ringtest_0.x3.x1.nSEL0 a_16155_12151# 2.51e-19
C1970 ringtest_0.x4.clknet_0_clk ringtest_0.x4._21_ 4.86e-19
C1971 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN1 0.004375f
C1972 ringtest_0.x4._15_ a_27065_5334# 2.78e-19
C1973 ringtest_0.x4._22_ a_26721_4246# 0.063386f
C1974 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 5.04e-19
C1975 ringtest_0.x4._14_ a_22021_4220# 0.134293f
C1976 ringtest_0.x4._04_ ringtest_0.x4.net8 7.52e-21
C1977 muxtest_0.x1.x3.GP1 muxtest_0.R2R3 0.127193f
C1978 a_25168_5156# VDPWR 0.256044f
C1979 a_21007_3867# a_21375_3867# 2.48e-19
C1980 ringtest_0.x4._18_ a_24361_5340# 5.99e-21
C1981 ringtest_0.x4.net8 a_25441_4612# 0.001229f
C1982 ringtest_0.x4._11_ a_22939_4584# 8.14e-19
C1983 a_23879_6940# a_24527_5340# 4.98e-20
C1984 ringtest_0.x4.net4 ringtest_0.x4._13_ 0.050083f
C1985 muxtest_0.x1.x3.GP1 ui_in[1] 8.43e-19
C1986 muxtest_0.x1.x3.GP2 muxtest_0.x1.x5.A 0.350698f
C1987 ringtest_0.x4.net3 a_21465_8830# 0.115857f
C1988 a_24336_6544# ringtest_0.x4._06_ 1.63e-21
C1989 a_20318_32213# ui_in[1] 0.125445f
C1990 a_25225_5334# a_25351_5712# 0.006169f
C1991 a_24527_5340# a_25309_5334# 3.14e-19
C1992 ringtest_0.x4.net1 a_22245_8054# 4.64e-19
C1993 ringtest_0.x4.clknet_0_clk a_23349_6422# 2.32e-20
C1994 a_21425_9686# ringtest_0.x4._12_ 1.27e-21
C1995 a_24329_6640# a_24004_6128# 0.001895f
C1996 ringtest_0.x4.net6 a_21785_5878# 0.006287f
C1997 a_21852_9416# a_21561_8830# 1.53e-19
C1998 a_21561_9116# a_21845_8816# 9.64e-20
C1999 ringtest_0.x4.clknet_0_clk a_23879_6940# 1.74729f
C2000 a_22983_5654# VDPWR 0.001324f
C2001 ringtest_0.x4._15_ a_26627_4246# 0.087822f
C2002 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP1 0.041018f
C2003 ringtest_0.x4._19_ a_24685_6788# 2.79e-19
C2004 ringtest_0.x4.net10 ringtest_0.x4.counter[8] 0.009948f
C2005 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN3 4.01e-20
C2006 ringtest_0.x4.net2 a_21465_9294# 0.092265f
C2007 ringtest_0.drv_out ui_in[4] 1.17e-19
C2008 ringtest_0.x4._23_ ringtest_0.x4._09_ 0.130147f
C2009 muxtest_0.x1.x5.GN a_20318_32213# 1.19e-19
C2010 ringtest_0.ring_out a_16579_11759# 5.47e-20
C2011 ringtest_0.x4._09_ a_26367_4790# 0.413296f
C2012 a_24536_6699# ringtest_0.x4._15_ 1.61e-21
C2013 a_26201_4790# a_26808_4902# 0.141453f
C2014 ui_in[6] ui_in[7] 0.03107f
C2015 ringtest_0.x4.net3 a_21948_5156# 3.32e-20
C2016 a_24763_6143# a_24361_5340# 0.004179f
C2017 a_13675_24012# ui_in[4] 8.84e-19
C2018 ringtest_0.x4._16_ ringtest_0.x4._07_ 0.003808f
C2019 ringtest_0.x4._06_ a_24986_5878# 6.53e-20
C2020 muxtest_0.x2.x2.GN3 ui_in[4] 0.273874f
C2021 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y 0.174714f
C2022 a_21591_6128# VDPWR 0.006535f
C2023 ringtest_0.x4._23_ a_26766_5712# 9.59e-19
C2024 muxtest_0.x2.x1.nSEL0 a_12849_23648# 1.91e-20
C2025 a_24004_6128# a_24545_5878# 4.72e-19
C2026 a_21951_5878# a_21672_5334# 0.001124f
C2027 ringtest_0.x4.clknet_1_0__leaf_clk a_21798_5712# 0.001807f
C2028 a_22486_4246# VDPWR 0.012117f
C2029 a_22228_9508# VDPWR 0.005789f
C2030 ringtest_0.x4.net9 a_25975_3867# 7.77e-19
C2031 ringtest_0.x4._11_ a_23932_6128# 0.002546f
C2032 ringtest_0.x4._15_ ringtest_0.x4._14_ 1.65e-19
C2033 ringtest_0.x4.clknet_1_1__leaf_clk a_24361_5340# 0.670964f
C2034 ringtest_0.x4.net4 ringtest_0.x4.net8 0.001699f
C2035 a_21852_8720# a_21981_8976# 0.124967f
C2036 a_21845_8816# ringtest_0.x4._01_ 0.092611f
C2037 ringtest_0.x4._24_ a_26895_3867# 0.00116f
C2038 muxtest_0.x2.x2.GP1 ui_in[3] 9.65e-19
C2039 muxtest_0.x1.x3.GN1 muxtest_0.R6R7 0.254376f
C2040 ringtest_0.counter3 ringtest_0.x4.net6 1.1e-21
C2041 ringtest_0.x4.net7 a_25975_3867# 4.41e-19
C2042 a_25977_4220# a_26269_4612# 0.001675f
C2043 ringtest_0.x4._23_ a_27659_4246# 0.009249f
C2044 ringtest_0.x4._14_ a_22541_5058# 1.14e-20
C2045 a_26640_5156# a_26721_4246# 7.6e-20
C2046 a_22052_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.040993f
C2047 a_12297_23648# ui_in[3] 0.246189f
C2048 ringtest_0.x4.net2 a_21981_8976# 8.2e-21
C2049 a_21981_9142# a_22399_9142# 3.39e-19
C2050 ringtest_0.drv_out ringtest_0.x3.x2.GP1 0.125793f
C2051 ringtest_0.x4.net7 a_24685_6788# 0.002551f
C2052 ringtest_0.x4._11_ ringtest_0.x4.net5 0.388184f
C2053 a_24004_6128# a_24317_4942# 2.49e-20
C2054 ringtest_0.x4.net1 a_22228_9508# 4.16e-19
C2055 a_24361_5340# a_24800_5334# 0.260055f
C2056 a_24527_5340# a_24968_5308# 0.110715f
C2057 ringtest_0.x4._06_ a_23899_5334# 2.02e-19
C2058 a_24070_5852# a_23899_5334# 1.06e-19
C2059 ringtest_0.x4.net9 a_26367_5340# 0.001054f
C2060 ringtest_0.counter3 a_21055_5334# 1.26e-20
C2061 a_23949_6654# ringtest_0.x4._19_ 0.065395f
C2062 ringtest_0.x4._08_ a_27191_5712# 7.43e-19
C2063 a_25593_5156# ringtest_0.x4._09_ 1.4e-19
C2064 ringtest_0.x4.clknet_0_clk a_24968_5308# 3.18e-19
C2065 a_21509_4790# a_22021_4220# 2.64e-19
C2066 ringtest_0.x4.net4 a_21798_5712# 1.81e-19
C2067 a_12977_24040# ua[3] 1.48e-19
C2068 ringtest_0.x4.net6 ringtest_0.x4.net10 1.08e-19
C2069 muxtest_0.x2.x2.GN2 ua[3] 0.234749f
C2070 ringtest_0.x4._15_ a_25351_5712# 0.00162f
C2071 ringtest_0.x4.net8 a_23837_5878# 0.057781f
C2072 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN4 0.011047f
C2073 a_16203_12091# ui_in[4] 0.254026f
C2074 ringtest_0.x4._24_ a_26808_5308# 0.015657f
C2075 ringtest_0.x4.net8 ringtest_0.x4._22_ 0.137056f
C2076 ringtest_0.x3.x1.nSEL1 a_16579_11759# 7.84e-19
C2077 a_21675_4790# ringtest_0.x4.net5 8.3e-19
C2078 a_22116_4902# a_22074_4790# 4.62e-19
C2079 ringtest_0.x4.net7 a_26367_5340# 2.99e-20
C2080 ringtest_0.x4._23_ a_24361_5340# 1.94e-21
C2081 a_21675_10006# VDPWR 5.43e-19
C2082 ringtest_0.x4._04_ a_22350_5878# 2.91e-19
C2083 muxtest_0.x1.x5.A muxtest_0.R3R4 4.07e-21
C2084 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.173286f
C2085 muxtest_0.x1.x3.GN3 a_13501_23906# 1.84e-20
C2086 ringtest_0.x4.net4 ringtest_0.x4.counter[1] 3.68e-19
C2087 a_21951_5878# a_22224_6244# 0.074434f
C2088 ringtest_0.x4._16_ a_22164_4362# 0.146025f
C2089 ringtest_0.x4._18_ VDPWR 0.686881f
C2090 a_13025_23980# VDPWR 0.261817f
C2091 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[3] 2.42e-19
C2092 ringtest_0.x4.clknet_1_0__leaf_clk a_22350_5878# 3.26e-19
C2093 a_21845_8816# a_21785_8054# 4.35e-19
C2094 a_21981_8976# a_22399_8976# 3.39e-19
C2095 ringtest_0.x4.net6 a_22775_5878# 5.88e-19
C2096 ringtest_0.counter7 VDPWR 2.42695f
C2097 ringtest_0.x4.clknet_0_clk a_25925_6788# 1.5e-19
C2098 ringtest_0.x4.net6 a_24627_6200# 4.57e-19
C2099 ringtest_0.x4.net9 a_27065_5156# 0.020729f
C2100 muxtest_0.x2.x2.GN4 m3_13302_19985# 7.07e-19
C2101 ringtest_0.x4.net6 ringtest_0.x4.counter[4] 0.003133f
C2102 a_23529_6422# ringtest_0.x4._16_ 1.86e-20
C2103 ringtest_0.x4.net4 a_22390_4566# 0.01239f
C2104 ringtest_0.x4._22_ a_24729_4790# 0.019806f
C2105 a_27191_5712# VDPWR 7.83e-19
C2106 ringtest_0.x4._15_ a_26721_4246# 0.038186f
C2107 ringtest_0.x4.net6 a_23399_3867# 3.58e-19
C2108 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN4 0.141966f
C2109 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GN3 0.175252f
C2110 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._08_ 0.00277f
C2111 ringtest_0.x4._00_ a_21981_9142# 0.005564f
C2112 ringtest_0.x4._24_ a_26555_4790# 3.3e-19
C2113 a_18836_32319# VDPWR 0.001273f
C2114 a_21785_5878# ringtest_0.x4.net5 1.51e-20
C2115 ringtest_0.x4.net7 a_27065_5156# 1.49e-19
C2116 a_22111_10993# ringtest_0.x4._00_ 4.57e-22
C2117 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP2 8.45e-19
C2118 ringtest_0.x4.net1 a_21675_10006# 0.003019f
C2119 a_23949_6654# ringtest_0.x4.net7 0.114197f
C2120 a_24763_6143# VDPWR 0.129866f
C2121 ringtest_0.x4.clknet_1_1__leaf_clk a_25336_4902# 0.046669f
C2122 ringtest_0.x4.net8 a_25225_5334# 0.00311f
C2123 ringtest_0.x4._11_ a_24527_5340# 8.46e-20
C2124 ringtest_0.x4._17_ a_23949_6654# 0.0702f
C2125 ringtest_0.x3.x2.GN1 ua[1] 0.430121f
C2126 a_22295_3867# VDPWR 0.317416f
C2127 a_22139_5878# a_21399_5340# 2.83e-19
C2128 a_16203_12091# ringtest_0.x3.x2.GP1 2.33e-21
C2129 ringtest_0.x4._06_ ringtest_0.x4._16_ 0.064563f
C2130 muxtest_0.x2.x1.nSEL1 a_11845_23906# 0.193944f
C2131 a_16579_11759# ringtest_0.x3.x2.GN3 0.104151f
C2132 ringtest_0.x4._08_ a_24800_5334# 1.22e-20
C2133 a_16755_12091# ringtest_0.x3.x2.GN1 3.78e-20
C2134 a_24070_5852# ringtest_0.x4._16_ 0.035189f
C2135 a_24317_4942# ringtest_0.x4._20_ 0.113204f
C2136 ringtest_0.x4._11_ ringtest_0.x4.clknet_0_clk 0.042991f
C2137 muxtest_0.x1.x3.GP2 a_13501_23906# 6.46e-20
C2138 ringtest_0.x4._15_ a_22765_5308# 8.84e-19
C2139 a_21509_4790# a_22541_5058# 0.048748f
C2140 ringtest_0.x4.net6 a_25393_5308# 0.002597f
C2141 ringtest_0.x4._03_ a_21948_5156# 0.010537f
C2142 ringtest_0.x4.clknet_1_1__leaf_clk VDPWR 3.34801f
C2143 ringtest_0.x4._12_ ringtest_0.x4._11_ 0.214271f
C2144 ringtest_0.x3.x2.GP2 VDPWR 1.81711f
C2145 a_22399_8976# a_22228_8598# 0.001229f
C2146 a_25393_5308# a_24895_4790# 0.002689f
C2147 ringtest_0.x4._22_ ringtest_0.x4.net11 1.96e-19
C2148 a_25225_5334# a_24729_4790# 0.004606f
C2149 muxtest_0.x1.x3.GP3 muxtest_0.R6R7 0.12263f
C2150 a_26569_6422# a_25364_5878# 0.010673f
C2151 ringtest_0.x4._16_ a_23891_4790# 0.00109f
C2152 ringtest_0.x4._05_ ringtest_0.x4._22_ 0.001519f
C2153 a_22765_5308# a_22541_5058# 0.002391f
C2154 a_22097_5334# a_22373_5156# 5.06e-19
C2155 ringtest_0.x4.net7 a_24004_6128# 3.79e-19
C2156 ringtest_0.x4._18_ ringtest_0.x4._21_ 0.005609f
C2157 ringtest_0.x4._23_ ringtest_0.x4._08_ 0.030554f
C2158 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2 3.78674f
C2159 muxtest_0.x2.x1.nSEL0 m2_11882_23495# 3.43e-19
C2160 ringtest_0.x4._16_ a_22373_5156# 6.21e-20
C2161 ringtest_0.x4._17_ a_24004_6128# 0.076419f
C2162 a_26808_5308# a_27233_5308# 1.28e-19
C2163 ringtest_0.x4._08_ a_26367_4790# 0.001269f
C2164 ringtest_0.counter7 ringtest_0.x4.counter[2] 0.003115f
C2165 a_26367_5340# a_27065_5334# 0.194892f
C2166 ringtest_0.counter3 ringtest_0.x4.net5 0.082815f
C2167 ringtest_0.ring_out ringtest_0.x3.x2.GP3 0.080819f
C2168 a_24800_5334# VDPWR 0.255475f
C2169 a_24465_6800# a_24264_6788# 4.67e-20
C2170 a_24336_6544# a_24883_6800# 0.095025f
C2171 a_24536_6699# a_24685_6788# 0.005525f
C2172 muxtest_0.R7R8 ui_in[3] 0.025566f
C2173 a_21425_9686# a_21675_10006# 0.007234f
C2174 ringtest_0.x4.net4 a_22074_4790# 6.57e-19
C2175 a_18662_32213# a_19114_31955# 0.002207f
C2176 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1 1.5157f
C2177 a_12297_23648# a_12425_24040# 0.004764f
C2178 a_12849_23648# a_13025_23980# 0.185422f
C2179 a_23349_6422# ringtest_0.x4._18_ 0.09549f
C2180 a_12297_23648# muxtest_0.x2.x2.GN1 0.012445f
C2181 ringtest_0.x4._21_ a_24763_6143# 1.69e-19
C2182 ringtest_0.x4._17_ a_23381_4818# 6.88e-22
C2183 ringtest_0.x3.x1.nSEL0 ui_in[4] 0.137394f
C2184 muxtest_0.R4R5 muxtest_0.R2R3 7.85e-20
C2185 a_27065_5334# a_27065_5156# 0.01464f
C2186 ringtest_0.x4._23_ VDPWR 1.70159f
C2187 a_21395_6940# ringtest_0.x4._04_ 0.00168f
C2188 a_21951_5878# a_22139_5878# 0.095025f
C2189 a_22817_6146# a_24004_6128# 1.25e-19
C2190 a_22245_8054# ringtest_0.x4._11_ 0.201886f
C2191 a_26367_4790# VDPWR 0.31984f
C2192 a_22295_3867# ringtest_0.x4.counter[2] 0.1107f
C2193 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C2194 ringtest_0.counter3 a_21007_3867# 2.11e-19
C2195 ringtest_0.x4.clknet_1_0__leaf_clk a_21395_6940# 1.67275f
C2196 a_16707_12151# VDPWR 0.001127f
C2197 ringtest_0.x3.x2.GN2 VDPWR 0.602894f
C2198 ringtest_0.x4._22_ ringtest_0.x4._09_ 0.009594f
C2199 muxtest_0.x2.x2.GN4 ua[0] 0.046938f
C2200 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._21_ 0.038033f
C2201 ringtest_0.x4._15_ ringtest_0.x4.net8 0.048599f
C2202 ringtest_0.x3.x2.GP1 m3_17036_9140# 5.81e-19
C2203 ringtest_0.x4.net2 ringtest_0.x4.counter[0] 0.010591f
C2204 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP3 5.60415f
C2205 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A 0.429865f
C2206 ringtest_0.x3.x2.GN3 m3_17032_8096# 0.087318f
C2207 ringtest_0.x4._24_ a_26817_4566# 9.33e-19
C2208 a_23879_6940# a_24763_6143# 1.03e-20
C2209 ringtest_0.x4.net9 ringtest_0.x4._20_ 1.35e-20
C2210 ringtest_0.x4.net3 a_22164_4362# 8.22e-19
C2211 ringtest_0.x4._11_ a_25168_5156# 0.026293f
C2212 ringtest_0.x4.net7 a_26375_4612# 6.33e-20
C2213 a_22021_4220# a_22390_4566# 0.046138f
C2214 ringtest_0.x4._23_ ringtest_0.x4._25_ 0.0063f
C2215 ringtest_0.x4.net5 ringtest_0.x4.counter[4] 0.001223f
C2216 a_27065_5156# a_26627_4246# 2.58e-19
C2217 a_27233_5058# a_27273_4220# 0.005283f
C2218 a_19666_31955# muxtest_0.x1.x3.GN3 0.104183f
C2219 a_21675_9686# a_21561_9116# 1.96e-19
C2220 ringtest_0.counter7 a_21375_3867# 2.81e-20
C2221 ringtest_0.x4.net5 a_23399_3867# 0.233889f
C2222 a_25421_6641# ringtest_0.x4._24_ 1.86e-20
C2223 a_19290_32287# VDPWR 0.194389f
C2224 a_27065_5156# a_27149_5156# 0.008508f
C2225 a_22649_6244# a_22373_5156# 2.6e-20
C2226 ringtest_0.x4._02_ VDPWR 0.325572f
C2227 a_21840_5308# a_22265_5308# 1.28e-19
C2228 a_21399_5340# a_22097_5334# 0.196846f
C2229 muxtest_0.x1.x1.nSEL0 a_18662_32213# 0.081627f
C2230 muxtest_0.x2.x2.GN4 a_13675_24012# 0.001562f
C2231 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GN4 0.071281f
C2232 ringtest_0.x4.net6 a_25083_4790# 0.00565f
C2233 ringtest_0.x4._15_ a_24729_4790# 4.49e-20
C2234 ringtest_0.x4.net8 a_24926_5712# 4.88e-19
C2235 m2_15612_11606# VDPWR 0.14037f
C2236 a_25364_5878# a_26640_5334# 0.01166f
C2237 ringtest_0.x4.net7 ringtest_0.x4._20_ 0.035834f
C2238 ringtest_0.x4._16_ a_21399_5340# 8.97e-20
C2239 muxtest_0.x1.x3.GP1 ui_in[0] 8.18e-19
C2240 VDPWR ui_in[3] 6.025721f
C2241 a_24045_6654# a_24336_6544# 0.192261f
C2242 a_23879_6940# ringtest_0.x4.clknet_1_1__leaf_clk 0.002451f
C2243 muxtest_0.x1.x1.nSEL0 m2_18699_31802# 3.43e-19
C2244 a_24895_4790# a_25083_4790# 0.095025f
C2245 a_25336_4902# a_25593_5156# 0.036838f
C2246 a_24729_4790# a_25263_5156# 0.002698f
C2247 a_20318_32213# ui_in[0] 0.220425f
C2248 ringtest_0.x4._17_ ringtest_0.x4._20_ 1.89e-19
C2249 ringtest_0.x3.nselect2 ringtest_0.x3.x2.GN4 1.53e-20
C2250 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GP1 6.21e-20
C2251 muxtest_0.R3R4 ua[2] 4.52137f
C2252 ui_in[2] ui_in[6] 0.264066f
C2253 ringtest_0.x4.clknet_1_1__leaf_clk a_25309_5334# 0.001538f
C2254 ringtest_0.x4.net6 a_24715_5334# 0.008614f
C2255 muxtest_0.x1.x3.GN4 muxtest_0.R1R2 0.628977f
C2256 a_26895_3867# ringtest_0.x4.counter[9] 2.34e-19
C2257 a_21395_6940# ringtest_0.x4.net4 4.87e-19
C2258 ringtest_0.x4._14_ a_22765_4478# 0.112679f
C2259 a_26201_5340# a_26201_4790# 0.037572f
C2260 uio_in[4] uio_in[3] 0.031023f
C2261 ringtest_0.x4._11_ a_21591_6128# 0.002118f
C2262 a_25593_5156# VDPWR 0.1878f
C2263 a_21375_3867# a_22295_3867# 1.37e-20
C2264 ringtest_0.x4._00_ ui_in[5] 2.67e-19
C2265 a_23879_6940# a_24800_5334# 5.07e-19
C2266 a_24329_6640# a_24545_5878# 2.84e-21
C2267 a_22399_9142# a_22245_8054# 9.03e-20
C2268 muxtest_0.x1.x3.GN2 muxtest_0.R3R4 0.271818f
C2269 muxtest_0.x1.x3.GP2 muxtest_0.x1.x4.A 0.350401f
C2270 a_22116_4902# VDPWR 0.219675f
C2271 ringtest_0.x4.net3 a_21845_8816# 0.008811f
C2272 a_24465_6800# ringtest_0.x4._06_ 4.29e-19
C2273 a_26201_5340# a_26555_5334# 0.062224f
C2274 a_21587_5334# a_21767_5334# 0.001229f
C2275 a_24336_6544# a_24699_6200# 6.47e-19
C2276 a_21845_9116# a_21845_8816# 0.040702f
C2277 ringtest_0.x4._00_ ringtest_0.x4._12_ 4.17e-19
C2278 a_21852_9416# a_21852_8720# 0.027204f
C2279 a_23993_5654# VDPWR 2.25e-21
C2280 a_19666_31955# muxtest_0.x1.x3.GP2 2.46e-19
C2281 ringtest_0.x4._15_ a_22390_4566# 8.81e-20
C2282 ringtest_0.x4._15_ a_26749_6422# 0.001357f
C2283 ringtest_0.x4._19_ a_24287_6422# 1.83e-19
C2284 ringtest_0.x4.net2 a_22201_9142# 1.37e-19
C2285 ringtest_0.x4._15_ ringtest_0.x4.net11 1.7e-19
C2286 ringtest_0.x4.net7 a_26569_6422# 6.19e-19
C2287 ringtest_0.x4.net2 a_21852_9416# 4.89e-19
C2288 ui_in[1] ui_in[2] 2.795f
C2289 ringtest_0.ring_out a_17231_12017# 0.001281f
C2290 ringtest_0.x4._05_ ringtest_0.x4._15_ 9.02e-20
C2291 a_26201_4790# a_27233_5058# 0.048748f
C2292 ringtest_0.x4._09_ a_26640_5156# 0.0221f
C2293 ringtest_0.x4._17_ a_26569_6422# 0.056144f
C2294 ringtest_0.x4.net3 a_22373_5156# 1.53e-21
C2295 ringtest_0.x4._22_ a_24361_5340# 0.016414f
C2296 a_24763_6143# a_24968_5308# 1.06e-19
C2297 a_22541_5058# a_22390_4566# 0.001062f
C2298 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 2.86851f
C2299 muxtest_0.x2.x2.GP1 ua[3] 4.09825f
C2300 ringtest_0.x4._04_ VDPWR 0.27578f
C2301 a_21951_5878# a_22097_5334# 3.42e-19
C2302 muxtest_0.x1.x5.GN ui_in[2] 3.98638f
C2303 a_24699_6200# a_24986_5878# 3.14e-19
C2304 a_22392_5990# a_22265_5308# 0.002135f
C2305 a_24329_6640# a_24317_4942# 8.37e-20
C2306 ringtest_0.x4.clknet_1_0__leaf_clk a_22223_5712# 4.11e-19
C2307 ringtest_0.x4.clknet_0_clk a_24627_6200# 2.68e-20
C2308 a_12297_23648# ua[3] 1.21e-19
C2309 ringtest_0.x4.clknet_1_0__leaf_clk VDPWR 3.74806f
C2310 a_21951_5878# ringtest_0.x4._16_ 1.01e-19
C2311 ringtest_0.x4.net9 a_27489_3702# 0.003439f
C2312 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ui_in[4] 9.08e-20
C2313 a_24045_6654# a_23899_5334# 4.21e-21
C2314 ringtest_0.x4.clknet_1_1__leaf_clk a_24968_5308# 0.01748f
C2315 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.173286f
C2316 ringtest_0.x4.net2 ringtest_0.x4._14_ 0.45134f
C2317 a_21591_6128# a_21785_5878# 5.05e-19
C2318 ringtest_0.x4._18_ a_21233_5340# 3.08e-21
C2319 a_22052_8875# ringtest_0.x4._01_ 0.004715f
C2320 a_26808_5308# a_27149_5334# 9.73e-19
C2321 a_26640_5334# a_26735_5334# 0.007724f
C2322 a_21852_9416# a_22399_8976# 4.5e-20
C2323 ringtest_0.x4._00_ a_22245_8054# 5.19e-20
C2324 a_27233_5058# a_27303_4246# 1.25e-19
C2325 a_21803_9508# ringtest_0.x4.clknet_1_0__leaf_clk 7.44e-19
C2326 a_12849_23648# ui_in[3] 0.086353f
C2327 a_22228_9508# a_22399_9142# 0.001229f
C2328 ringtest_0.drv_out ringtest_0.x4.net6 2.01e-20
C2329 ringtest_0.x4._11_ ringtest_0.x4._18_ 0.035586f
C2330 ringtest_0.x4.net7 a_24287_6422# 6.13e-20
C2331 ringtest_0.x4._11_ ringtest_0.counter7 2.85e-19
C2332 ringtest_0.x4._17_ a_22392_5990# 2.52e-22
C2333 a_24527_5340# a_25393_5308# 0.034054f
C2334 a_24361_5340# a_25225_5334# 0.030894f
C2335 ringtest_0.x4.net1 ringtest_0.x4.clknet_1_0__leaf_clk 0.561165f
C2336 a_21399_5340# a_21587_5334# 0.097818f
C2337 a_24968_5308# a_24800_5334# 0.239923f
C2338 a_18662_32213# muxtest_0.x1.x3.GN2 0.039612f
C2339 ringtest_0.x4._15_ ringtest_0.x4._09_ 0.030214f
C2340 ringtest_0.x4.clknet_1_1__leaf_clk a_25925_6788# 0.001522f
C2341 ringtest_0.x4._17_ a_24287_6422# 0.002375f
C2342 ringtest_0.x4._21_ a_23993_5654# 4.25e-19
C2343 muxtest_0.x1.x3.GN3 ua[0] 0.007815f
C2344 a_24329_6640# ringtest_0.x4._19_ 0.074331f
C2345 ringtest_0.x4.clknet_0_clk a_25393_5308# 0.01296f
C2346 ringtest_0.x4._03_ a_22164_4362# 0.005187f
C2347 ringtest_0.x4.net4 a_22223_5712# 3.33e-19
C2348 a_24317_4942# a_24551_4790# 0.005167f
C2349 ringtest_0.x4._15_ a_26766_5712# 4.15e-19
C2350 a_17377_14114# VDPWR 0.006305f
C2351 ringtest_0.x4.net4 VDPWR 1.18326f
C2352 a_16755_12091# ui_in[4] 0.127717f
C2353 ringtest_0.x4._24_ a_27233_5308# 0.009415f
C2354 ringtest_0.x4._11_ a_24763_6143# 0.004209f
C2355 a_21948_5156# ringtest_0.x4.net5 4.4e-19
C2356 a_22373_5156# a_22457_5156# 0.008508f
C2357 ringtest_0.x4.net3 a_21399_5340# 0.007798f
C2358 a_22765_5308# a_22765_4478# 8.07e-19
C2359 ringtest_0.x4._08_ ringtest_0.x4._22_ 1.19e-20
C2360 ringtest_0.x4.net8 a_25975_3867# 0.2272f
C2361 ringtest_0.x4._18_ a_23899_5654# 9.76e-19
C2362 ringtest_0.x4._11_ a_22295_3867# 3.83e-19
C2363 a_21951_5878# a_22649_6244# 0.194203f
C2364 a_22392_5990# a_22817_6146# 1.28e-19
C2365 ringtest_0.x4._16_ a_23381_4584# 0.039613f
C2366 a_12425_24040# VDPWR 4.32e-19
C2367 muxtest_0.x1.x4.A muxtest_0.R3R4 4.53278f
C2368 a_23899_5334# a_23809_4790# 8.68e-19
C2369 ringtest_0.x4.net9 a_25149_4220# 0.125008f
C2370 muxtest_0.x2.x2.GN1 VDPWR 1.60341f
C2371 ringtest_0.x4._01_ a_21803_8598# 2.39e-19
C2372 a_21852_8720# ringtest_0.x4._10_ 6.77e-19
C2373 ringtest_0.x4.net6 ringtest_0.x4._07_ 0.066033f
C2374 a_23529_6422# a_23770_5308# 6.83e-19
C2375 a_22052_8875# a_21785_8054# 0.0033f
C2376 a_24715_5334# a_24895_5334# 0.001229f
C2377 a_24045_6654# ringtest_0.x4._16_ 1.29e-20
C2378 ringtest_0.x4._07_ a_24895_4790# 0.195848f
C2379 a_24329_6640# ringtest_0.x4.net9 6.06e-20
C2380 ringtest_0.x4._22_ a_25336_4902# 0.001181f
C2381 ringtest_0.x4._19_ a_25364_5878# 6.04e-19
C2382 ringtest_0.x4.net2 ringtest_0.x4._10_ 0.006086f
C2383 ringtest_0.x4.net6 a_25055_3867# 0.013611f
C2384 ringtest_0.x4._11_ ringtest_0.x4.clknet_1_1__leaf_clk 0.367667f
C2385 muxtest_0.R3R4 m3_13302_19985# 0.136776f
C2386 a_24895_4790# a_25055_3867# 1.2e-20
C2387 ringtest_0.x4._00_ a_22228_9508# 8.32e-19
C2388 a_25925_6788# ringtest_0.x4._23_ 0.026998f
C2389 ringtest_0.x4._18_ a_21785_5878# 7.56e-20
C2390 ringtest_0.x4.net6 a_24264_6788# 1.91e-20
C2391 ringtest_0.x4.net7 a_25149_4220# 0.212284f
C2392 a_21425_9686# ringtest_0.x4.clknet_1_0__leaf_clk 3.24e-19
C2393 muxtest_0.x1.x5.GN a_19794_32347# 9.76e-20
C2394 muxtest_0.x1.x1.nSEL1 a_19242_32347# 9.57e-19
C2395 ringtest_0.x4.net7 a_26735_5156# 1.13e-19
C2396 muxtest_0.x1.x3.GP2 ua[0] 1.13e-20
C2397 a_21675_4790# a_22295_3867# 7.04e-21
C2398 a_23837_5878# VDPWR 0.004487f
C2399 a_24329_6640# ringtest_0.x4.net7 0.035144f
C2400 ringtest_0.x4._14_ a_21840_5308# 8.48e-21
C2401 ringtest_0.x4._22_ VDPWR 0.56354f
C2402 ringtest_0.x4._06_ a_23770_5308# 0.002127f
C2403 ringtest_0.x3.x2.GP1 ua[1] 0.352376f
C2404 ringtest_0.x4.clknet_1_1__leaf_clk a_25761_5058# 0.084941f
C2405 muxtest_0.R3R4 muxtest_0.x2.x2.GP2 0.171364f
C2406 ringtest_0.x4.net8 a_26367_5340# 5.19e-19
C2407 ringtest_0.x4._11_ a_24800_5334# 2.99e-20
C2408 ringtest_0.x4.net9 a_24545_5878# 0.063508f
C2409 ringtest_0.x4._19_ a_24317_4942# 4.85e-22
C2410 ringtest_0.x4._17_ a_24329_6640# 0.42661f
C2411 a_24070_5852# a_23770_5308# 8.74e-19
C2412 a_24135_3867# VDPWR 0.287214f
C2413 a_17231_12017# a_17405_12123# 0.006584f
C2414 a_16755_12091# ringtest_0.x3.x2.GP1 2.87e-20
C2415 ringtest_0.x4.net2 a_21509_4790# 5.19e-20
C2416 ringtest_0.x4._08_ a_25225_5334# 7.33e-20
C2417 muxtest_0.x2.x1.nSEL1 a_12473_23980# 0.041068f
C2418 a_15749_12123# ringtest_0.x3.x2.GN2 8.86e-19
C2419 a_17231_12017# ringtest_0.x3.x2.GN3 1.07e-20
C2420 ringtest_0.x3.x2.GN1 a_16155_12151# 1.22e-20
C2421 a_24699_6200# ringtest_0.x4._16_ 0.113309f
C2422 a_25364_5878# ringtest_0.x4.net9 0.111158f
C2423 a_23619_6788# VDPWR 0.002157f
C2424 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ui_in[4] 0.001652f
C2425 ringtest_0.x4.net6 a_26201_5340# 2.14e-19
C2426 a_21509_4790# a_23381_4818# 7.98e-21
C2427 ringtest_0.x4._03_ a_22373_5156# 0.001345f
C2428 ringtest_0.x4._15_ a_24361_5340# 0.034785f
C2429 muxtest_0.x1.x4.A muxtest_0.x2.x1.nSEL0 4.83e-20
C2430 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 5.04e-19
C2431 ringtest_0.x4.net4 ringtest_0.x4.counter[2] 0.006188f
C2432 ringtest_0.x4.net7 a_24545_5878# 2.13e-20
C2433 a_25225_5334# a_25336_4902# 0.001204f
C2434 a_25393_5308# a_25168_5156# 0.003655f
C2435 a_16027_11759# VDPWR 0.161536f
C2436 a_21465_8830# ringtest_0.x4._12_ 0.027335f
C2437 muxtest_0.x1.x3.GN4 muxtest_0.R6R7 0.156481f
C2438 ringtest_0.x4._16_ a_24479_4790# 7.06e-20
C2439 ringtest_0.x4._11_ ringtest_0.x4._23_ 0.090724f
C2440 ringtest_0.x4.net2 a_21867_8054# 6.45e-19
C2441 ringtest_0.x4.net7 a_25364_5878# 0.037674f
C2442 ringtest_0.x4.net6 ringtest_0.x4.counter[5] 0.080069f
C2443 ringtest_0.x4._11_ a_26367_4790# 7.13e-19
C2444 a_19842_32287# muxtest_0.R7R8 7.47e-21
C2445 ringtest_0.x4._16_ a_23809_4790# 0.105405f
C2446 ringtest_0.x4.net2 ringtest_0.x4._13_ 0.197255f
C2447 a_15749_12123# ui_in[3] 9.55e-19
C2448 a_23949_6654# ringtest_0.x4.net8 1.16e-19
C2449 a_24527_5340# a_24715_5334# 0.095025f
C2450 ringtest_0.x4._17_ a_25364_5878# 0.002308f
C2451 ringtest_0.x4.net9 a_24317_4942# 3.24e-20
C2452 ringtest_0.counter3 ringtest_0.counter7 3.44556f
C2453 a_25225_5334# VDPWR 0.182006f
C2454 ui_in[2] ui_in[4] 0.015983f
C2455 muxtest_0.R7R8 m3_13316_18955# 0.131878f
C2456 ringtest_0.x4._16_ a_22795_5334# 0.059496f
C2457 a_24465_6800# a_24883_6800# 3.39e-19
C2458 a_21675_10006# ringtest_0.x4._00_ 0.002065f
C2459 a_19114_31955# a_19290_32287# 0.185422f
C2460 ringtest_0.x4._23_ a_25761_5058# 1.37e-20
C2461 a_21233_5340# ringtest_0.x4._02_ 0.184941f
C2462 a_25761_5058# a_26367_4790# 8.52e-19
C2463 a_23529_6422# ringtest_0.x4.net6 1.5e-19
C2464 a_12473_23980# muxtest_0.x2.x2.GN3 0.048646f
C2465 ringtest_0.x4.net7 a_24317_4942# 0.084753f
C2466 a_12849_23648# muxtest_0.x2.x2.GN1 6.43e-20
C2467 ringtest_0.x4._21_ a_23837_5878# 0.002821f
C2468 ringtest_0.counter7 ua[2] 2.06e-19
C2469 ringtest_0.x4._11_ ringtest_0.x4._02_ 0.012298f
C2470 ringtest_0.x4._21_ ringtest_0.x4._22_ 2.96e-19
C2471 ringtest_0.x4._17_ a_24317_4942# 1.09e-21
C2472 a_26749_6422# a_26367_5340# 6.98e-21
C2473 m2_11882_23495# ui_in[3] 0.130999f
C2474 a_27169_6641# a_26201_5340# 7.7e-20
C2475 a_21509_4790# ringtest_0.x4._20_ 1.9e-21
C2476 ringtest_0.x4._03_ a_22499_4790# 9.96e-20
C2477 a_22021_4220# VDPWR 0.377321f
C2478 ringtest_0.counter7 ringtest_0.x4.net10 5.8e-20
C2479 ringtest_0.x4.net8 a_24004_6128# 0.063158f
C2480 a_21951_5878# a_22733_6244# 4.04e-19
C2481 a_22224_6244# a_22139_5878# 0.037333f
C2482 a_26640_5156# VDPWR 0.248502f
C2483 ringtest_0.counter3 a_22295_3867# 5.4e-19
C2484 ringtest_0.x4._12_ a_21780_8964# 0.001666f
C2485 a_21132_8918# a_21049_8598# 2.42e-19
C2486 ringtest_0.x4.net4 a_21375_3867# 7.77e-19
C2487 ringtest_0.x4.net6 ringtest_0.x4._06_ 0.037389f
C2488 ringtest_0.x4._19_ ringtest_0.x4.net9 4.58e-20
C2489 VDPWR ua[3] 11.3115f
C2490 a_23879_6940# a_23837_5878# 1.78e-20
C2491 ringtest_0.x4._24_ a_27491_4566# 5.3e-19
C2492 ringtest_0.x4.net6 a_24070_5852# 0.016498f
C2493 ringtest_0.x3.x2.GP2 ringtest_0.counter3 0.148166f
C2494 a_21399_5340# ringtest_0.x4._03_ 1.23e-19
C2495 a_21840_5308# a_21509_4790# 0.001425f
C2496 a_26201_4790# a_26895_3867# 4.75e-20
C2497 a_23879_6940# ringtest_0.x4._22_ 7.51e-19
C2498 a_21233_5340# a_22116_4902# 0.001786f
C2499 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP1 0.051787f
C2500 ringtest_0.x4.net8 a_23963_4790# 8.5e-20
C2501 ringtest_0.x4._15_ ringtest_0.x4._08_ 0.030258f
C2502 a_22765_4478# a_22390_4566# 4e-20
C2503 muxtest_0.R3R4 ua[0] 3.1523f
C2504 ringtest_0.x4._11_ a_25593_5156# 0.045045f
C2505 a_20492_32319# VDPWR 8.55e-19
C2506 ringtest_0.counter7 ringtest_0.x4.counter[4] 0.007159f
C2507 ui_in[1] ui_in[6] 0.239552f
C2508 a_21561_9116# a_21780_9142# 0.006169f
C2509 a_20318_32213# muxtest_0.x1.x3.GN3 1.07e-20
C2510 a_21675_9686# a_21845_9116# 5.23e-20
C2511 a_21465_9294# a_21852_9416# 0.034054f
C2512 muxtest_0.x1.x3.GN1 a_19242_32347# 1.22e-20
C2513 ringtest_0.counter7 a_23399_3867# 2.81e-20
C2514 a_18836_32319# muxtest_0.x1.x3.GN2 8.86e-19
C2515 a_19842_32287# VDPWR 0.261767f
C2516 a_27065_5156# ringtest_0.x4.net11 0.003417f
C2517 ringtest_0.x4._11_ a_22116_4902# 0.004479f
C2518 ringtest_0.x4._19_ ringtest_0.x4.net7 0.552257f
C2519 muxtest_0.x1.x1.nSEL0 a_19290_32287# 0.001174f
C2520 ringtest_0.x4._15_ a_25336_4902# 4.59e-21
C2521 a_22649_6244# a_22795_5334# 1.65e-19
C2522 ringtest_0.x4._11_ a_23993_5654# 5.64e-19
C2523 ringtest_0.x4._16_ a_21672_5334# 1.68e-20
C2524 a_24045_6654# a_24465_6800# 0.036838f
C2525 a_24329_6640# a_24536_6699# 0.260055f
C2526 a_23949_6654# ringtest_0.x4._05_ 1.85e-19
C2527 ringtest_0.x4._17_ ringtest_0.x4._19_ 0.214371f
C2528 ringtest_0.x4._24_ a_27149_5334# 8.56e-19
C2529 a_25168_5156# a_25083_4790# 0.037333f
C2530 a_25761_5058# a_25593_5156# 0.310858f
C2531 ua[0] ui_in[5] 0.483363f
C2532 muxtest_0.R3R4 muxtest_0.x2.x2.GN3 3.9625f
C2533 a_21561_8830# VDPWR 0.181976f
C2534 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net10 6.99e-20
C2535 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x1.nSEL1 0.352716f
C2536 ringtest_0.x4._04_ a_21233_5340# 0.001469f
C2537 ringtest_0.drv_out ui_in[5] 0.391919f
C2538 a_27815_3867# ringtest_0.x4.counter[9] 0.039377f
C2539 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ui_in[4] 1.79e-19
C2540 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x3.x2.GN1 2.09e-20
C2541 ringtest_0.x4._15_ VDPWR 1.72333f
C2542 ringtest_0.x4.clknet_1_0__leaf_clk a_21233_5340# 0.318658f
C2543 a_21675_4790# a_22116_4902# 0.127288f
C2544 a_26808_5308# a_26201_4790# 1.99e-20
C2545 ringtest_0.drv_out ringtest_0.x4.clknet_0_clk 0.00889f
C2546 ringtest_0.x4._11_ ringtest_0.x4._04_ 0.257603f
C2547 ui_in[0] ui_in[2] 0.450267f
C2548 a_25263_5156# VDPWR 0.003234f
C2549 a_22295_3867# a_23399_3867# 9e-21
C2550 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.173286f
C2551 a_25364_5878# a_26627_4246# 1.15e-20
C2552 a_24536_6699# a_24545_5878# 1.55e-20
C2553 ringtest_0.x4.net7 ringtest_0.x4.net9 0.742565f
C2554 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._11_ 0.317456f
C2555 a_22541_5058# VDPWR 0.391294f
C2556 ringtest_0.x4.net3 a_22052_8875# 3.02e-19
C2557 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.ring_out 0.083309f
C2558 ringtest_0.x4.net2 ringtest_0.x4.counter[1] 0.015257f
C2559 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP2 0.100463f
C2560 a_25225_5334# a_25309_5334# 0.008508f
C2561 a_26808_5308# a_26555_5334# 3.39e-19
C2562 ringtest_0.x4._17_ ringtest_0.x4.net9 7.02e-19
C2563 a_21845_9116# a_22052_8875# 6.88e-20
C2564 a_22052_9116# a_21852_8720# 1.26e-19
C2565 muxtest_0.x1.x5.GN ui_in[1] 0.141313f
C2566 a_24465_6800# a_24699_6200# 1.61e-19
C2567 a_21981_9142# a_21845_8816# 5.28e-20
C2568 a_24926_5712# VDPWR 0.001185f
C2569 ringtest_0.x3.x2.GN2 ringtest_0.counter3 0.004367f
C2570 ringtest_0.x4._15_ a_23467_4584# 0.001523f
C2571 ringtest_0.x4.net8 ringtest_0.x4._20_ 0.027217f
C2572 ringtest_0.x4._15_ ringtest_0.x4._25_ 0.003323f
C2573 ringtest_0.x4.net1 a_21561_8830# 0.030538f
C2574 ringtest_0.ring_out a_17405_12123# 1.86e-19
C2575 ringtest_0.x4.net2 a_22052_9116# 1.88e-19
C2576 ringtest_0.ring_out ringtest_0.x3.x2.GN3 0.080584f
C2577 a_26201_4790# a_26555_4790# 0.062224f
C2578 a_21951_5878# ringtest_0.x4._03_ 3.92e-19
C2579 ringtest_0.x4._09_ a_27065_5156# 0.024482f
C2580 ringtest_0.x4._07_ a_24527_5340# 0.029939f
C2581 ringtest_0.x4._22_ a_24968_5308# 0.01767f
C2582 ringtest_0.x4.net5 a_22164_4362# 3.95e-20
C2583 ringtest_0.x4._17_ ringtest_0.x4.net7 0.072785f
C2584 ringtest_0.x4.clknet_1_0__leaf_clk a_21675_4790# 0.021572f
C2585 ringtest_0.counter7 a_26808_4902# 1.4e-19
C2586 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN3 4.01e-20
C2587 a_24527_5340# a_25055_3867# 7.09e-22
C2588 ringtest_0.x4._23_ ringtest_0.x4.net10 0.188811f
C2589 ringtest_0.x4.clknet_0_clk ringtest_0.x4._07_ 0.114561f
C2590 a_21049_8598# VDPWR 0.229121f
C2591 ringtest_0.x3.x2.GN4 ringtest_0.counter7 3.94045f
C2592 ringtest_0.counter3 ringtest_0.x4._02_ 0.001266f
C2593 ringtest_0.x4._20_ a_24729_4790# 0.004564f
C2594 a_22224_6244# a_22097_5334# 0.002298f
C2595 ringtest_0.x4.net10 a_26367_4790# 0.003321f
C2596 a_26173_4612# VDPWR 0.001618f
C2597 a_12849_23648# ua[3] 0.001506f
C2598 ringtest_0.x4.net4 a_21233_5340# 0.007432f
C2599 a_22224_6244# ringtest_0.x4._16_ 1.81e-20
C2600 a_26895_3867# ringtest_0.x4.counter[8] 6.92e-19
C2601 muxtest_0.x1.x4.A a_13025_23980# 3.23e-19
C2602 ringtest_0.x4.clknet_1_1__leaf_clk a_25393_5308# 0.005058f
C2603 ringtest_0.x4.net6 a_21399_5340# 1.26e-19
C2604 ringtest_0.x4.clknet_0_clk a_24264_6788# 1.49e-19
C2605 ringtest_0.x4._11_ ringtest_0.x4.net4 0.952686f
C2606 a_21785_5878# ringtest_0.x4._04_ 0.09532f
C2607 ringtest_0.x4._15_ ringtest_0.x4._21_ 0.054317f
C2608 ringtest_0.x4.clknet_1_0__leaf_clk a_21785_5878# 0.245743f
C2609 a_26627_4246# a_26913_4566# 0.010132f
C2610 muxtest_0.x2.x2.GN1 m2_11882_23495# 0.06935f
C2611 a_13501_23906# ui_in[3] 0.220366f
C2612 a_22399_9142# ringtest_0.x4.clknet_1_0__leaf_clk 0.012004f
C2613 ui_in[3] ua[2] 1.63519f
C2614 ringtest_0.x4.net1 a_21049_8598# 0.060735f
C2615 a_21425_9686# a_21561_8830# 6.59e-20
C2616 ringtest_0.x4.net7 a_26095_6788# 0.00717f
C2617 ringtest_0.x4._21_ a_22541_5058# 1.79e-21
C2618 ringtest_0.x4._17_ a_22817_6146# 1.35e-20
C2619 a_21840_5308# a_21798_5712# 4.62e-19
C2620 a_21672_5334# a_21587_5334# 0.037333f
C2621 a_24527_5340# a_26201_5340# 1.33e-19
C2622 a_24968_5308# a_25225_5334# 0.036838f
C2623 a_24361_5340# a_26367_5340# 3.42e-21
C2624 a_19290_32287# muxtest_0.x1.x3.GN2 0.017048f
C2625 ringtest_0.x4.net9 a_27065_5334# 2.45e-19
C2626 ringtest_0.x4.clknet_1_1__leaf_clk a_26808_4902# 2.7e-19
C2627 ringtest_0.x4.net4 a_21675_4790# 0.019846f
C2628 a_13025_23980# muxtest_0.x2.x2.GP2 3.2e-20
C2629 a_24536_6699# ringtest_0.x4._19_ 0.034076f
C2630 muxtest_0.x2.x2.GP3 ui_in[4] 0.00356f
C2631 a_23879_6940# ringtest_0.x4._15_ 2.08e-20
C2632 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP2 8.45e-19
C2633 ringtest_0.x4._03_ a_23381_4584# 2.93e-20
C2634 a_19794_32347# ui_in[0] 0.001558f
C2635 ringtest_0.x4.net4 a_23899_5654# 7.88e-20
C2636 ringtest_0.x3.x2.GN1 ui_in[4] 0.312198f
C2637 ringtest_0.x4._11_ a_23837_5878# 3.73e-19
C2638 a_15575_12017# ringtest_0.x3.x2.GN2 0.039612f
C2639 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN3 0.012418f
C2640 ringtest_0.x4._11_ ringtest_0.x4._22_ 0.420712f
C2641 a_22373_5156# ringtest_0.x4.net5 0.019334f
C2642 ringtest_0.x4.net3 a_21672_5334# 8.21e-19
C2643 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ui_in[4] 1.03e-20
C2644 rst_n clk 0.031023f
C2645 a_22392_5990# ringtest_0.x4.net8 1.22e-20
C2646 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 5.04e-19
C2647 ringtest_0.x4.net9 a_26627_4246# 0.008597f
C2648 ringtest_0.x4._01_ a_21785_8054# 3.94e-19
C2649 a_21981_8976# ringtest_0.x4._10_ 6.67e-19
C2650 a_24045_6654# a_23770_5308# 7.28e-21
C2651 muxtest_0.x1.x3.GP1 muxtest_0.R3R4 4.16645f
C2652 ringtest_0.x4.net9 a_27149_5156# 1.5e-19
C2653 ringtest_0.x4.net4 a_21785_5878# 0.071607f
C2654 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ui_in[3] 1.18e-19
C2655 ringtest_0.x4._11_ a_23619_6788# 1.46e-19
C2656 ringtest_0.x4._07_ a_25168_5156# 0.008539f
C2657 a_24336_6544# ringtest_0.x4._16_ 6.29e-20
C2658 a_24883_6800# a_24712_6422# 0.001229f
C2659 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.ring_out 0.025177f
C2660 a_24536_6699# ringtest_0.x4.net9 4.56e-19
C2661 ringtest_0.x4._22_ a_25761_5058# 3.11e-19
C2662 ui_in[4] ui_in[6] 0.177925f
C2663 ui_in[0] rst_n 0.031023f
C2664 ringtest_0.x4.clknet_0_clk a_23529_6422# 8e-19
C2665 ringtest_0.x4.net6 a_21951_5878# 0.004467f
C2666 ringtest_0.x4._24_ a_27273_4220# 0.003347f
C2667 a_15575_12017# m2_15612_11606# 0.01297f
C2668 a_26569_6422# a_26749_6422# 0.185422f
C2669 a_15575_12017# ui_in[3] 0.048888f
C2670 ringtest_0.x4._24_ a_26766_4790# 6.57e-19
C2671 ringtest_0.x4.net6 a_24883_6800# 9.51e-20
C2672 ringtest_0.x4._00_ ringtest_0.x4.clknet_1_0__leaf_clk 0.144154f
C2673 ringtest_0.x4.net7 a_27149_5156# 3.05e-20
C2674 ringtest_0.x4._23_ a_26808_4902# 0.005759f
C2675 muxtest_0.x1.x1.nSEL1 VDPWR 0.475048f
C2676 a_24763_6143# a_24715_5334# 1.39e-19
C2677 ringtest_0.x4._05_ a_26569_6422# 6.38e-20
C2678 a_26367_4790# a_26808_4902# 0.118966f
C2679 a_24536_6699# ringtest_0.x4.net7 0.026259f
C2680 ringtest_0.x4._14_ a_22265_5308# 1.02e-20
C2681 ringtest_0.x4._06_ a_24527_5340# 0.183131f
C2682 ringtest_0.x4.clknet_1_1__leaf_clk a_25083_4790# 0.011819f
C2683 ringtest_0.x4._16_ a_24986_5878# 3.12e-19
C2684 ringtest_0.x4.net8 a_26640_5334# 2.79e-19
C2685 ringtest_0.x4._11_ a_25225_5334# 7.12e-21
C2686 ringtest_0.x4._17_ a_24536_6699# 0.032936f
C2687 a_24004_6128# a_24361_5340# 4.26e-19
C2688 a_16707_12151# ringtest_0.x3.x2.GN4 3.22e-19
C2689 a_25975_3867# VDPWR 0.309637f
C2690 ringtest_0.x3.x2.GN3 a_17405_12123# 1.07e-20
C2691 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1 1.51569f
C2692 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GN4 8.82e-19
C2693 muxtest_0.x2.x1.nSEL1 a_13025_23980# 1.59e-19
C2694 ringtest_0.x4._08_ a_26367_5340# 0.415957f
C2695 ringtest_0.x4.net5 a_22499_4790# 6.03e-19
C2696 ringtest_0.x4.clknet_0_clk ringtest_0.x4._06_ 2.8e-19
C2697 a_24685_6788# VDPWR 0.002269f
C2698 ringtest_0.x4._04_ a_22775_5878# 6.79e-19
C2699 a_21785_5878# a_23837_5878# 9.88e-21
C2700 ringtest_0.x4.clknet_0_clk a_24070_5852# 7.65e-20
C2701 ringtest_0.x4.clknet_1_1__leaf_clk a_24715_5334# 0.017223f
C2702 ui_in[1] ui_in[4] 4.85e-19
C2703 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x3.nselect2 1.41e-19
C2704 ringtest_0.x4._15_ a_24968_5308# 0.03519f
C2705 a_21233_5340# a_22021_4220# 3.4e-19
C2706 ringtest_0.x4._22_ a_25345_4612# 0.002279f
C2707 ringtest_0.x4._01_ a_22695_8304# 0.012244f
C2708 muxtest_0.x1.x5.A ua[3] 4.51865f
C2709 ringtest_0.counter3 ringtest_0.x4.net4 8.11e-19
C2710 a_25393_5308# a_25593_5156# 4.17e-19
C2711 a_24800_5334# a_25083_4790# 0.001307f
C2712 a_26913_4566# a_26721_4246# 6.96e-20
C2713 muxtest_0.x1.x3.GN3 muxtest_0.R4R5 0.123863f
C2714 a_16579_11759# VDPWR 0.179803f
C2715 ringtest_0.x4.net8 a_25149_4220# 0.1454f
C2716 a_21845_8816# ringtest_0.x4._12_ 0.062549f
C2717 ringtest_0.x4._11_ a_22021_4220# 7.66e-19
C2718 ringtest_0.x4.net9 a_25294_4790# 3.93e-19
C2719 a_23770_5308# a_23809_4790# 2.2e-19
C2720 muxtest_0.x1.x5.GN ui_in[4] 2.49e-19
C2721 ringtest_0.x4.net11 a_27489_3702# 0.250513f
C2722 ringtest_0.x4._11_ a_26640_5156# 5.04e-19
C2723 muxtest_0.x1.x3.GN1 muxtest_0.R7R8 4.45989f
C2724 ringtest_0.x3.x2.GN4 ui_in[3] 0.218716f
C2725 a_24800_5334# a_24715_5334# 0.037333f
C2726 a_24968_5308# a_24926_5712# 4.62e-19
C2727 ringtest_0.x4.net2 a_21132_8918# 0.010623f
C2728 a_22765_5308# a_23151_5334# 0.006406f
C2729 a_24329_6640# ringtest_0.x4.net8 0.001356f
C2730 ringtest_0.x4._08_ a_27065_5156# 3.02e-19
C2731 a_26367_5340# VDPWR 0.31297f
C2732 ringtest_0.x4.net6 a_23381_4584# 1.4e-20
C2733 ringtest_0.x4._16_ a_23899_5334# 0.008193f
C2734 ringtest_0.x4._15_ a_25925_6788# 0.142876f
C2735 ringtest_0.x4._24_ a_26201_4790# 0.03301f
C2736 ringtest_0.drv_out ringtest_0.counter7 2.39e-19
C2737 ringtest_0.x4.net9 a_25351_5712# 3.81e-19
C2738 a_19290_32287# a_19666_31955# 3.02e-19
C2739 muxtest_0.x1.x4.A ui_in[3] 0.00371f
C2740 a_24729_4790# a_25149_4220# 0.009169f
C2741 a_24045_6654# ringtest_0.x4.net6 8.38e-19
C2742 a_21675_4790# a_22021_4220# 0.010515f
C2743 a_13025_23980# muxtest_0.x2.x2.GN3 0.004288f
C2744 a_24329_6640# a_24729_4790# 2.6e-21
C2745 muxtest_0.x2.x2.GN1 ua[2] 0.430038f
C2746 ringtest_0.x4._24_ a_26555_5334# 4.8e-19
C2747 a_27233_5308# a_27273_4220# 1.35e-20
C2748 ringtest_0.x4.net7 a_25351_5712# 1.38e-19
C2749 ringtest_0.x4.net8 a_24545_5878# 0.009814f
C2750 ringtest_0.x4._25_ a_26367_5340# 1.11e-19
C2751 ui_in[0] ui_in[6] 0.281408f
C2752 a_22765_4478# VDPWR 0.201367f
C2753 ringtest_0.x3.nselect2 a_16755_12091# 6.01e-20
C2754 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ui_in[4] 7.73e-20
C2755 a_21507_9686# VDPWR 0.008578f
C2756 ringtest_0.x4.net9 a_26721_4246# 0.003753f
C2757 a_22392_5990# a_22350_5878# 4.62e-19
C2758 a_21951_5878# a_23932_6128# 1.01e-20
C2759 a_27065_5156# VDPWR 0.215619f
C2760 ringtest_0.x4.net8 a_25364_5878# 0.001798f
C2761 ringtest_0.x4._15_ a_21233_5340# 8.17e-21
C2762 a_23949_6654# VDPWR 0.376761f
C2763 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.173286f
C2764 muxtest_0.x1.x3.GP2 muxtest_0.R4R5 0.117653f
C2765 a_21845_8816# a_22245_8054# 4.04e-19
C2766 ringtest_0.x4._12_ a_22201_8964# 0.002771f
C2767 ringtest_0.x4.net4 a_23399_3867# 0.003224f
C2768 muxtest_0.x2.x2.GP2 ui_in[3] 6.63e-19
C2769 muxtest_0.x1.x3.GN1 muxtest_0.R5R6 0.250509f
C2770 ringtest_0.x4._11_ ringtest_0.x4._15_ 1.40124f
C2771 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B 0.163894f
C2772 ringtest_0.x4.net6 a_24699_6200# 0.09145f
C2773 a_21672_5334# ringtest_0.x4._03_ 0.001262f
C2774 a_22265_5308# a_21509_4790# 0.00142f
C2775 ringtest_0.x4.net8 a_24551_4790# 5.79e-19
C2776 a_25364_5878# a_24729_4790# 4.21e-21
C2777 a_24699_6200# a_24895_4790# 8.41e-19
C2778 ringtest_0.drv_out ringtest_0.x4.clknet_1_1__leaf_clk 0.008913f
C2779 ringtest_0.drv_out ringtest_0.x3.x2.GP2 4.09557f
C2780 ringtest_0.counter7 a_25055_3867# 2.81e-20
C2781 a_21561_9116# a_21845_9116# 0.032244f
C2782 ringtest_0.x4._22_ ringtest_0.x4.net10 0.074459f
C2783 a_21951_5878# ringtest_0.x4.net5 3.57e-21
C2784 muxtest_0.x1.x3.GN1 VDPWR 0.915833f
C2785 ringtest_0.x4.net8 a_24317_4942# 0.236033f
C2786 ringtest_0.x4._11_ a_22541_5058# 0.065594f
C2787 ringtest_0.x4.net1 a_21507_9686# 0.010028f
C2788 a_22265_5308# a_22765_5308# 0.016344f
C2789 muxtest_0.x1.x1.nSEL0 a_19842_32287# 1.21e-20
C2790 ui_in[0] ui_in[1] 4.44986f
C2791 ringtest_0.x4.net6 a_24479_4790# 1.78e-19
C2792 ringtest_0.x4._15_ a_25761_5058# 7.77e-19
C2793 ringtest_0.x4._16_ a_22097_5334# 1.35e-19
C2794 a_24329_6640# ringtest_0.x4._05_ 0.196756f
C2795 a_24336_6544# a_24465_6800# 0.110715f
C2796 muxtest_0.x1.x3.GN3 ui_in[2] 0.002225f
C2797 a_24004_6128# VDPWR 0.316019f
C2798 a_24729_4790# a_24551_4790# 1.43e-19
C2799 a_21395_6940# a_21840_5308# 3.17e-20
C2800 a_24763_6143# ringtest_0.x4._07_ 0.001092f
C2801 ringtest_0.x4.net6 a_23809_4790# 0.005791f
C2802 muxtest_0.x1.x5.GN ui_in[0] 0.149831f
C2803 a_21852_8720# VDPWR 0.309635f
C2804 a_24317_4942# a_24729_4790# 0.020429f
C2805 ringtest_0.x4._15_ a_23899_5654# 0.005043f
C2806 ringtest_0.x4.net6 a_22795_5334# 0.007899f
C2807 a_21675_4790# a_22541_5058# 0.034054f
C2808 a_24135_3867# ringtest_0.x4.counter[4] 0.110403f
C2809 a_22116_4902# a_21948_5156# 0.239923f
C2810 ringtest_0.x4.net2 VDPWR 2.41286f
C2811 a_23963_4790# VDPWR 3.08e-19
C2812 a_23399_3867# a_24135_3867# 2.31e-20
C2813 ringtest_0.x4._11_ a_26173_4612# 7.08e-19
C2814 muxtest_0.x1.x3.GP3 muxtest_0.R7R8 0.124327f
C2815 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._07_ 0.44529f
C2816 a_26749_6422# a_25364_5878# 0.006666f
C2817 a_23381_4818# VDPWR 0.254188f
C2818 ringtest_0.x4.net3 ringtest_0.x4._01_ 0.006403f
C2819 a_26640_5334# a_26766_5712# 0.005525f
C2820 ringtest_0.x4._19_ ringtest_0.x4.net8 2.14e-19
C2821 a_21845_9116# ringtest_0.x4._01_ 6.79e-20
C2822 ringtest_0.x4._05_ a_25364_5878# 0.003024f
C2823 a_23949_6654# ringtest_0.x4._21_ 0.001295f
C2824 a_21981_9142# a_22052_8875# 1.77e-19
C2825 a_22052_9116# a_21981_8976# 1.77e-19
C2826 ringtest_0.x4.clknet_1_0__leaf_clk a_21465_8830# 0.01132f
C2827 a_22181_5334# VDPWR 0.007439f
C2828 ringtest_0.x4.clknet_1_1__leaf_clk a_25055_3867# 4.13e-21
C2829 ringtest_0.x4._15_ a_25345_4612# 2.85e-21
C2830 ringtest_0.counter7 ringtest_0.x4.counter[5] 0.007023f
C2831 muxtest_0.x2.x1.nSEL1 ui_in[3] 0.168511f
C2832 ringtest_0.x4.net1 a_21852_8720# 0.00338f
C2833 a_26201_4790# a_25977_4220# 2.81e-20
C2834 ringtest_0.drv_out ringtest_0.x3.x2.GN2 3.92936f
C2835 a_21425_9686# a_21507_9686# 0.006406f
C2836 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP3 3.4436f
C2837 a_21785_5878# a_22541_5058# 3.85e-19
C2838 ringtest_0.x4.net8 a_26735_5334# 7.49e-20
C2839 ringtest_0.x4._04_ a_21948_5156# 3.52e-21
C2840 ringtest_0.x4._07_ a_24800_5334# 0.002926f
C2841 ringtest_0.x4.net1 ringtest_0.x4.net2 0.722672f
C2842 a_25421_6641# ringtest_0.x4.net6 0.019537f
C2843 ringtest_0.x4.net3 a_21863_4790# 7.76e-19
C2844 ringtest_0.x4.net5 a_23381_4584# 0.201023f
C2845 ringtest_0.x4._22_ a_25393_5308# 4.4e-21
C2846 muxtest_0.x1.x3.GP2 ui_in[2] 4.34e-19
C2847 ringtest_0.x4.clknet_1_0__leaf_clk a_21948_5156# 0.003461f
C2848 ringtest_0.x4._18_ a_23529_6422# 0.190808f
C2849 a_24800_5334# a_25055_3867# 3e-19
C2850 a_22399_8976# VDPWR 0.074934f
C2851 ringtest_0.x4._20_ a_25336_4902# 6.25e-20
C2852 a_23879_6940# a_23949_6654# 0.022122f
C2853 a_22817_6146# a_22765_5308# 0.004132f
C2854 muxtest_0.R7R8 muxtest_0.R1R2 0.216753f
C2855 ringtest_0.x4.net10 a_26640_5156# 5.45e-19
C2856 a_26375_4612# VDPWR 1.16e-19
C2857 a_13501_23906# ua[3] 0.003273f
C2858 ua[3] ua[2] 8.93455f
C2859 a_24883_6800# a_24527_5340# 1.11e-20
C2860 a_22649_6244# ringtest_0.x4._16_ 0.003542f
C2861 a_27815_3867# ringtest_0.x4.counter[8] 0.111116f
C2862 ringtest_0.x4.net8 ringtest_0.x4.net9 0.748324f
C2863 a_24004_6128# ringtest_0.x4._21_ 0.128337f
C2864 a_15575_12017# a_16027_11759# 0.002207f
C2865 muxtest_0.R4R5 muxtest_0.R3R4 1.39313f
C2866 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN1 1.38e-21
C2867 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ui_in[4] 1.2e-19
C2868 ringtest_0.x4.clknet_1_1__leaf_clk a_26201_5340# 0.285659f
C2869 ringtest_0.x3.x2.GP3 VDPWR 1.79155f
C2870 ringtest_0.x4._13_ ringtest_0.x4.counter[0] 3.39e-20
C2871 ringtest_0.x4.net6 a_21672_5334# 6.57e-20
C2872 ringtest_0.x4.clknet_0_clk a_24883_6800# 0.004448f
C2873 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 5.04e-19
C2874 muxtest_0.x1.x3.GP3 muxtest_0.R5R6 4.11451f
C2875 ringtest_0.x4._20_ VDPWR 0.175404f
C2876 ringtest_0.x4.net3 a_21785_8054# 0.079675f
C2877 ringtest_0.x4._22_ a_26808_4902# 8.71e-19
C2878 muxtest_0.x1.x3.GN2 ua[3] 0.01442f
C2879 a_22164_4362# a_22295_3867# 0.002548f
C2880 a_26627_4246# a_26721_4246# 0.062574f
C2881 a_27273_4220# a_27491_4566# 0.007234f
C2882 ringtest_0.x4.clknet_1_0__leaf_clk a_21780_8964# 0.001172f
C2883 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B 5.04e-19
C2884 a_13675_24012# ui_in[3] 1.4e-19
C2885 ringtest_0.x4._16_ a_23467_4818# 5.76e-19
C2886 ringtest_0.x4.net7 ringtest_0.x4.net8 1.22349f
C2887 a_25364_5878# ringtest_0.x4._09_ 3.55e-20
C2888 muxtest_0.x2.x2.GN3 ui_in[3] 0.254283f
C2889 ringtest_0.x4.net9 a_24729_4790# 0.006834f
C2890 ringtest_0.x4._18_ ringtest_0.x4._06_ 3.12e-20
C2891 ringtest_0.x4.net1 a_22399_8976# 6.38e-20
C2892 muxtest_0.x1.x3.GP3 VDPWR 3.24635f
C2893 muxtest_0.x1.x3.GN2 a_20492_32319# 8.14e-21
C2894 muxtest_0.x1.x3.GN3 a_19794_32347# 0.001073f
C2895 ringtest_0.x4.net7 a_26839_6788# 1.83e-19
C2896 ringtest_0.x4._18_ a_24070_5852# 7.58e-19
C2897 a_23879_6940# a_24004_6128# 1.01e-19
C2898 ringtest_0.x4._17_ ringtest_0.x4.net8 0.172731f
C2899 a_21840_5308# a_22223_5712# 4.67e-20
C2900 a_25393_5308# a_25225_5334# 0.310858f
C2901 a_19842_32287# muxtest_0.x1.x3.GN2 9.62e-20
C2902 ringtest_0.x4.net6 ringtest_0.x4._24_ 0.002355f
C2903 a_21840_5308# VDPWR 0.200136f
C2904 ringtest_0.x4._16_ a_21587_5334# 4.26e-21
C2905 ringtest_0.x4.net2 a_21425_9686# 0.107098f
C2906 muxtest_0.x1.x1.nSEL1 a_19114_31955# 0.073392f
C2907 ringtest_0.x4.net4 a_21948_5156# 0.004091f
C2908 ringtest_0.x4.clknet_1_1__leaf_clk a_27233_5058# 1.1e-19
C2909 ua[2] ua[6] 0.001584f
C2910 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP2 0.005194f
C2911 ringtest_0.x4._05_ ringtest_0.x4._19_ 0.284135f
C2912 ringtest_0.x4.net7 a_24729_4790# 0.003956f
C2913 a_23529_6422# ringtest_0.x4.clknet_1_1__leaf_clk 1.19e-21
C2914 ringtest_0.x3.x2.GP1 ui_in[4] 8.45e-19
C2915 ringtest_0.x4._17_ a_24729_4790# 1.69e-21
C2916 ringtest_0.x4._15_ ringtest_0.x4.net10 0.289356f
C2917 ringtest_0.x4._06_ a_24763_6143# 9.69e-19
C2918 a_16203_12091# ringtest_0.x3.x2.GN2 0.017071f
C2919 a_23809_4790# ringtest_0.x4.net5 5.06e-20
C2920 ringtest_0.x4._23_ a_26201_5340# 0.029216f
C2921 a_26569_6422# VDPWR 0.206381f
C2922 a_26201_5340# a_26367_4790# 2.64e-19
C2923 muxtest_0.R1R2 VDPWR 1.61319f
C2924 ringtest_0.x4.net3 ringtest_0.x4._16_ 6.72e-19
C2925 ringtest_0.x4._11_ a_25975_3867# 2.18e-19
C2926 a_22817_6146# ringtest_0.x4.net8 5.45e-19
C2927 a_26749_6422# ringtest_0.x4.net9 7.48e-22
C2928 a_24329_6640# a_24361_5340# 0.001493f
C2929 ringtest_0.x4.net9 ringtest_0.x4.net11 0.055197f
C2930 ringtest_0.x4._15_ ringtest_0.x4.counter[4] 9.07e-20
C2931 a_24465_6800# ringtest_0.x4._16_ 2.16e-20
C2932 ringtest_0.x4._07_ a_25593_5156# 5.62e-20
C2933 ringtest_0.x3.x2.GP2 m3_17036_9140# 0.004119f
C2934 ringtest_0.x4._05_ ringtest_0.x4.net9 1.93e-19
C2935 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._06_ 0.005269f
C2936 ringtest_0.x4._22_ a_25083_4790# 0.012798f
C2937 ringtest_0.x4.clknet_0_clk a_24045_6654# 0.00222f
C2938 ringtest_0.x4.net6 a_22224_6244# 3.12e-19
C2939 ringtest_0.x4.net2 a_21375_3867# 0.016821f
C2940 ringtest_0.x4._21_ ringtest_0.x4._20_ 0.296715f
C2941 ringtest_0.x4._14_ a_21509_4790# 0.008544f
C2942 a_25761_5058# a_25975_3867# 2.93e-21
C2943 a_26569_6422# ringtest_0.x4._25_ 0.001476f
C2944 ringtest_0.x4._24_ a_27169_6641# 0.006166f
C2945 a_16203_12091# ui_in[3] 0.143958f
C2946 ringtest_0.x4.net7 a_26749_6422# 5.4e-19
C2947 muxtest_0.R3R4 ui_in[2] 2.94e-19
C2948 ringtest_0.x4._23_ a_27233_5058# 2.3e-19
C2949 ringtest_0.x4.net7 ringtest_0.x4.net11 2.47e-20
C2950 a_26367_4790# a_27233_5058# 0.034054f
C2951 a_26808_4902# a_26640_5156# 0.239923f
C2952 ringtest_0.x4._14_ a_22765_5308# 1.74e-20
C2953 ringtest_0.x4._05_ ringtest_0.x4.net7 0.232588f
C2954 ringtest_0.x4._17_ a_26749_6422# 8.24e-19
C2955 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x1.nSEL1 0.352716f
C2956 ringtest_0.x4._06_ a_24800_5334# 3.32e-19
C2957 ringtest_0.x4.net8 a_27065_5334# 1.1e-19
C2958 ringtest_0.x4._11_ a_26367_5340# 2.03e-20
C2959 a_27489_3702# VDPWR 0.293517f
C2960 ringtest_0.x4._17_ ringtest_0.x4._05_ 0.0576f
C2961 a_24699_6200# a_24527_5340# 1.08e-19
C2962 muxtest_0.x2.x1.nSEL1 a_12425_24040# 9.57e-19
C2963 a_11845_23906# a_12019_24012# 0.006584f
C2964 a_22392_5990# VDPWR 0.177502f
C2965 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN1 0.034862f
C2966 ringtest_0.x4._08_ a_26640_5334# 0.030723f
C2967 ui_in[2] ui_in[5] 0.211146f
C2968 a_24287_6422# VDPWR 0.004852f
C2969 ringtest_0.x4._13_ ringtest_0.x4._14_ 0.074354f
C2970 ringtest_0.x4.clknet_0_clk a_24699_6200# 0.034583f
C2971 a_21509_4790# a_22043_5156# 0.002698f
C2972 ringtest_0.x4._15_ a_25393_5308# 0.031321f
C2973 ringtest_0.x4.counter[0] ringtest_0.x4.counter[1] 0.079742f
C2974 ringtest_0.x4._03_ a_21863_4790# 0.13856f
C2975 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ui_in[4] 1.2e-19
C2976 ringtest_0.x4._22_ a_25547_4612# 0.002069f
C2977 uio_in[3] uio_in[2] 0.031023f
C2978 a_21981_8976# a_21395_6940# 1.29e-20
C2979 muxtest_0.x1.x4.A ua[3] 6.48818f
C2980 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.173286f
C2981 muxtest_0.x2.nselect2 VDPWR 1.22451f
C2982 a_17231_12017# VDPWR 0.217593f
C2983 a_22052_8875# ringtest_0.x4._12_ 0.032034f
C2984 ringtest_0.x4.net8 a_26627_4246# 4.33e-20
C2985 ringtest_0.x4._11_ a_22765_4478# 0.159397f
C2986 a_24361_5340# a_24317_4942# 1.28e-19
C2987 ringtest_0.x4.net9 ringtest_0.x4._09_ 0.571636f
C2988 muxtest_0.x2.x2.GN1 ua[0] 2.35e-19
C2989 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A 0.17253f
C2990 ringtest_0.x4._11_ a_27065_5156# 3.81e-21
C2991 ringtest_0.x3.x2.GN2 m3_17036_9140# 0.099332f
C2992 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A 0.4308f
C2993 a_23770_5308# a_23899_5334# 0.062574f
C2994 a_24536_6699# ringtest_0.x4.net8 5.83e-19
C2995 ringtest_0.x4._11_ a_23949_6654# 8.65e-19
C2996 ringtest_0.x4.clknet_1_1__leaf_clk a_26269_4612# 3.29e-19
C2997 a_26640_5334# VDPWR 0.247111f
C2998 ringtest_0.x4.net6 a_25977_4220# 0.009771f
C2999 a_19114_31955# muxtest_0.x1.x3.GN1 0.012335f
C3000 a_19666_31955# a_19842_32287# 0.185422f
C3001 ringtest_0.x4._15_ a_26808_4902# 0.002208f
C3002 ringtest_0.x4.net7 ringtest_0.x4._09_ 2.46e-19
C3003 a_25336_4902# a_25149_4220# 3.07e-19
C3004 a_24336_6544# ringtest_0.x4.net6 0.001918f
C3005 a_12425_24040# muxtest_0.x2.x2.GN3 5.17e-20
C3006 muxtest_0.x2.x2.GN2 a_12977_24040# 3.11e-20
C3007 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN3 0.002859f
C3008 a_21948_5156# a_22021_4220# 3.53e-19
C3009 a_22116_4902# a_22164_4362# 5.83e-19
C3010 muxtest_0.x2.x2.GP2 ua[3] 0.085048f
C3011 a_18662_32213# ui_in[2] 4.33e-19
C3012 m3_13302_19985# m3_13316_18955# 0.003741f
C3013 ringtest_0.x4.net3 a_21587_5334# 0.003111f
C3014 a_11845_23906# ui_in[4] 0.02803f
C3015 ringtest_0.x4.counter[9] ringtest_0.x4.counter[8] 0.299988f
C3016 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN2 0.154394f
C3017 a_25149_4220# VDPWR 0.405792f
C3018 m2_18699_31802# ui_in[2] 4.4e-19
C3019 a_21465_9294# VDPWR 0.415615f
C3020 ringtest_0.x4._10_ a_21867_8054# 4.63e-20
C3021 a_21785_8054# a_21939_8054# 0.004009f
C3022 ringtest_0.x4.net9 a_27659_4246# 3.29e-19
C3023 a_26735_5156# VDPWR 0.002923f
C3024 a_22649_6244# a_22733_6244# 0.008508f
C3025 ringtest_0.x4._11_ a_24004_6128# 0.043142f
C3026 ringtest_0.x4._19_ a_24361_5340# 9.86e-21
C3027 muxtest_0.R7R8 muxtest_0.R6R7 2.27687f
C3028 a_24287_6422# ringtest_0.x4._21_ 1.26e-19
C3029 ringtest_0.x4._08_ a_25364_5878# 0.011527f
C3030 a_24329_6640# VDPWR 0.438492f
C3031 a_22052_8875# a_22245_8054# 2.48e-20
C3032 ringtest_0.x4._12_ a_21803_8598# 1.13e-19
C3033 ringtest_0.x4.net2 a_21233_5340# 3.28e-19
C3034 a_21852_8720# ringtest_0.x4._11_ 4.06e-19
C3035 ringtest_0.x4.net6 a_24986_5878# 0.001357f
C3036 muxtest_0.x1.x3.GN3 muxtest_0.R2R3 0.27459f
C3037 muxtest_0.x2.x2.GP2 m3_13316_18955# 2.65e-20
C3038 muxtest_0.x1.x3.GN3 ui_in[1] 0.273672f
C3039 a_21465_8830# a_21561_8830# 0.310858f
C3040 ringtest_0.x4.clknet_0_clk a_25421_6641# 0.012442f
C3041 ringtest_0.x4.net6 a_22139_5878# 5.63e-21
C3042 ringtest_0.x4.net2 ringtest_0.x4._11_ 0.001125f
C3043 a_22052_9116# a_22201_9142# 0.005525f
C3044 a_21981_9142# a_21780_9142# 4.67e-20
C3045 ringtest_0.x4._11_ a_23963_4790# 0.001879f
C3046 a_24699_6200# a_25168_5156# 5.18e-21
C3047 a_25364_5878# a_25336_4902# 2.72e-20
C3048 ringtest_0.x4.net11 a_26627_4246# 2.78e-19
C3049 ringtest_0.x4._16_ ringtest_0.x4._03_ 0.005745f
C3050 a_21561_9116# a_21981_9142# 0.036838f
C3051 a_21852_9416# a_22052_9116# 0.074815f
C3052 ringtest_0.x3.x1.nSEL0 m2_15612_11606# 3.43e-19
C3053 ringtest_0.counter7 a_26895_3867# 0.110188f
C3054 ringtest_0.x4._18_ a_21951_5878# 8.49e-20
C3055 ringtest_0.x3.x1.nSEL0 ui_in[3] 0.324822f
C3056 a_22224_6244# ringtest_0.x4.net5 1.47e-19
C3057 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN3 1.7e-19
C3058 ringtest_0.x4._11_ a_23381_4818# 0.163973f
C3059 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN2 0.209954f
C3060 ringtest_0.x4.net1 a_21465_9294# 0.045364f
C3061 ringtest_0.x4._18_ a_24883_6800# 2.19e-20
C3062 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN1 0.002605f
C3063 a_24545_5878# VDPWR 0.011033f
C3064 ringtest_0.x4._06_ a_23993_5654# 6.56e-20
C3065 ringtest_0.x4._15_ a_25083_4790# 7.24e-21
C3066 ringtest_0.x4._13_ a_21509_4790# 6.65e-20
C3067 ringtest_0.x4._11_ a_22181_5334# 7.61e-19
C3068 ringtest_0.x4._16_ a_23770_5308# 0.01721f
C3069 a_24536_6699# ringtest_0.x4._05_ 3.36e-19
C3070 ringtest_0.x4.net9 a_24361_5340# 5.55e-19
C3071 a_24895_4790# a_25677_5156# 3.14e-19
C3072 a_25083_4790# a_25263_5156# 0.001229f
C3073 a_25364_5878# VDPWR 1.3575f
C3074 ringtest_0.counter7 ua[1] 5.26868f
C3075 muxtest_0.x2.x2.GN4 ui_in[4] 0.063283f
C3076 ringtest_0.x4._22_ ringtest_0.x4._07_ 0.503878f
C3077 ringtest_0.x4.net2 a_21675_4790# 3.95e-20
C3078 muxtest_0.x2.nselect2 a_12849_23648# 1.29e-19
C3079 ringtest_0.drv_out a_25225_5334# 2.32e-21
C3080 ringtest_0.x4._14_ ringtest_0.x4.counter[1] 1.03e-21
C3081 a_21981_8976# VDPWR 0.211083f
C3082 ringtest_0.x4.net6 a_23899_5334# 0.044713f
C3083 ringtest_0.x4._15_ a_24715_5334# 0.019231f
C3084 ringtest_0.x4._22_ a_25055_3867# 8.8e-19
C3085 ringtest_0.x4._14_ a_22390_4566# 0.122283f
C3086 a_22116_4902# a_22373_5156# 0.036838f
C3087 a_27065_5334# ringtest_0.x4._09_ 0.001217f
C3088 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ui_in[4] 2.29e-19
C3089 ringtest_0.x4.net7 a_24361_5340# 0.088061f
C3090 a_22399_8976# ringtest_0.x4._11_ 0.001319f
C3091 muxtest_0.R6R7 muxtest_0.R5R6 2.03637f
C3092 a_21785_5878# a_24004_6128# 1.89e-21
C3093 a_24135_3867# a_25055_3867# 1.37e-20
C3094 ringtest_0.x4._04_ a_24070_5852# 8.65e-21
C3095 a_24551_4790# VDPWR 9.47e-20
C3096 muxtest_0.x1.x3.GP2 muxtest_0.R2R3 4.15159f
C3097 ringtest_0.x4.net8 a_26721_4246# 6.89e-20
C3098 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 5.04e-19
C3099 ringtest_0.x4._11_ a_26375_4612# 0.001561f
C3100 muxtest_0.x1.x3.GP2 ui_in[1] 3.1e-20
C3101 ringtest_0.x4._17_ a_24361_5340# 1.12e-20
C3102 a_21465_8830# a_21049_8598# 5.03e-19
C3103 ringtest_0.counter3 a_22765_4478# 8.56e-20
C3104 muxtest_0.x1.x3.GP3 muxtest_0.x1.x5.A 0.358703f
C3105 a_21561_8830# a_21780_8964# 0.006169f
C3106 a_24317_4942# VDPWR 0.226919f
C3107 muxtest_0.x1.x3.GN4 muxtest_0.R7R8 0.13848f
C3108 a_26808_5308# a_27191_5712# 4.67e-20
C3109 muxtest_0.R6R7 VDPWR 1.6078f
C3110 a_26367_5340# ringtest_0.x4.net10 5.04e-19
C3111 a_22399_9142# a_21852_8720# 4.5e-20
C3112 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A 5.04e-19
C3113 ringtest_0.x4.clknet_1_0__leaf_clk a_21845_8816# 0.683552f
C3114 a_24329_6640# ringtest_0.x4._21_ 8.19e-20
C3115 ringtest_0.x4.net4 a_22164_4362# 0.007901f
C3116 ringtest_0.x4.net2 a_21785_5878# 2.26e-20
C3117 a_23151_5334# VDPWR 0.009139f
C3118 ringtest_0.x4._15_ a_25547_4612# 5.62e-21
C3119 ua[3] ua[0] 1.8361f
C3120 ringtest_0.x4.net1 a_21981_8976# 0.001727f
C3121 ringtest_0.x4._11_ ringtest_0.x4._20_ 0.174111f
C3122 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP2 1.7e-20
C3123 ringtest_0.x4.net2 a_22399_9142# 1.04e-19
C3124 ringtest_0.x4._09_ a_26627_4246# 0.001692f
C3125 ringtest_0.x4.clknet_1_1__leaf_clk a_24883_6800# 3.41e-20
C3126 a_21425_9686# a_21465_9294# 1.32e-19
C3127 ringtest_0.x4._00_ a_21507_9686# 6.18e-19
C3128 ringtest_0.x4._09_ a_27149_5156# 6.12e-19
C3129 ringtest_0.x4._04_ a_22373_5156# 0.001409f
C3130 ringtest_0.x4._07_ a_25225_5334# 0.009837f
C3131 ringtest_0.x4._22_ a_26201_5340# 5.82e-21
C3132 ringtest_0.x4._02_ a_21399_5340# 0.275992f
C3133 a_21233_5340# a_21840_5308# 0.141453f
C3134 ringtest_0.x3.x2.GP2 ua[1] 0.349381f
C3135 ringtest_0.x4.clknet_1_0__leaf_clk a_22373_5156# 6.12e-19
C3136 ringtest_0.counter7 a_26555_4790# 2.77e-20
C3137 muxtest_0.R3R4 muxtest_0.x2.x2.GP3 4.09931f
C3138 ringtest_0.x4._18_ a_24045_6654# 2.33e-19
C3139 a_23349_6422# a_24329_6640# 6.46e-21
C3140 a_22228_8598# VDPWR 0.004407f
C3141 a_16755_12091# ringtest_0.x3.x2.GP2 3.2e-20
C3142 a_23879_6940# a_24329_6640# 0.022305f
C3143 ringtest_0.x4._21_ a_24545_5878# 0.053333f
C3144 a_13675_24012# ua[3] 3.17e-19
C3145 ringtest_0.x4._20_ a_25761_5058# 3.47e-20
C3146 ringtest_0.x4.clknet_1_0__leaf_clk a_21767_5334# 0.001355f
C3147 ringtest_0.x4._11_ a_21840_5308# 0.005658f
C3148 a_26913_4566# VDPWR 4.51e-19
C3149 ringtest_0.x4.net10 a_27065_5156# 0.003817f
C3150 muxtest_0.x2.x2.GN3 ua[3] 0.087947f
C3151 ringtest_0.ring_out VDPWR 4.36398f
C3152 ringtest_0.counter3 m3_17032_8096# 0.119717f
C3153 a_16027_11759# a_16203_12091# 0.185422f
C3154 a_25364_5878# ringtest_0.x4._21_ 3.33e-20
C3155 a_22116_4902# a_22499_4790# 4.67e-20
C3156 a_24135_3867# ringtest_0.x4.counter[5] 4.98e-19
C3157 ringtest_0.x4._19_ VDPWR 0.197759f
C3158 ringtest_0.x4.clknet_1_1__leaf_clk a_26808_5308# 5.16e-19
C3159 ringtest_0.x4._08_ ringtest_0.x4.net9 0.003243f
C3160 ringtest_0.x4.clknet_0_clk a_26007_6788# 5.18e-20
C3161 ringtest_0.x4.net6 a_22097_5334# 5.09e-19
C3162 ringtest_0.x4.net6 ringtest_0.x4._16_ 0.291584f
C3163 muxtest_0.x1.x3.GN4 muxtest_0.R5R6 0.304696f
C3164 ringtest_0.x4.clknet_1_0__leaf_clk a_22201_8964# 4.64e-19
C3165 muxtest_0.x2.x2.GN3 m3_13316_18955# 0.016026f
C3166 ringtest_0.x4._23_ a_26895_3867# 7.52e-20
C3167 a_27273_4220# a_27303_4246# 0.025037f
C3168 ringtest_0.x4.net2 ringtest_0.counter3 0.003151f
C3169 a_23879_6940# a_24545_5878# 2.81e-20
C3170 ringtest_0.x4._16_ a_24895_4790# 4.88e-21
C3171 a_26735_5334# VDPWR 0.002923f
C3172 ringtest_0.x4.net9 a_25336_4902# 0.007121f
C3173 a_21840_5308# a_21675_4790# 3.46e-19
C3174 a_21399_5340# a_22116_4902# 0.001879f
C3175 ringtest_0.counter7 m3_17046_7066# 0.117708f
C3176 ringtest_0.drv_out ringtest_0.x4._15_ 0.005511f
C3177 ringtest_0.x4.net7 ringtest_0.x4._08_ 1.97e-19
C3178 ringtest_0.x4._00_ a_21852_8720# 4.06e-19
C3179 ringtest_0.counter7 ringtest_0.x4.counter[6] 0.087745f
C3180 muxtest_0.x1.x3.GN4 VDPWR 1.35388f
C3181 ringtest_0.x4._21_ a_24317_4942# 0.011629f
C3182 a_22265_5308# a_22223_5712# 7.84e-20
C3183 a_25393_5308# a_26367_5340# 2.73e-19
C3184 a_25225_5334# a_26201_5340# 1.07e-19
C3185 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN2 0.142718f
C3186 ringtest_0.x4._19_ ringtest_0.x4._25_ 9.05e-21
C3187 a_22265_5308# VDPWR 0.421579f
C3188 ringtest_0.x4.net2 ringtest_0.x4._00_ 0.002662f
C3189 a_23529_6422# a_23619_6788# 0.004764f
C3190 muxtest_0.x1.x1.nSEL1 a_19666_31955# 7.84e-19
C3191 ringtest_0.x4.clknet_1_1__leaf_clk a_26555_4790# 6.27e-19
C3192 ringtest_0.x4.net4 a_22373_5156# 0.022715f
C3193 ringtest_0.x4.net7 a_25336_4902# 0.005145f
C3194 ringtest_0.x4.net3 ringtest_0.x4._03_ 0.019455f
C3195 ringtest_0.x4.net9 VDPWR 0.964697f
C3196 a_24045_6654# ringtest_0.x4.clknet_1_1__leaf_clk 1.54e-20
C3197 ui_in[6] ui_in[5] 6.50488f
C3198 a_21509_4790# a_22390_4566# 3.11e-19
C3199 ringtest_0.x3.x2.GN2 ua[1] 0.42933f
C3200 ringtest_0.x4._06_ a_23837_5878# 4.79e-19
C3201 a_16579_11759# ringtest_0.x3.x2.GN4 6.84e-19
C3202 ringtest_0.x4._06_ ringtest_0.x4._22_ 0.004416f
C3203 a_16755_12091# ringtest_0.x3.x2.GN2 5.62e-20
C3204 ringtest_0.x4._04_ a_21399_5340# 0.011144f
C3205 a_24070_5852# a_23837_5878# 0.005961f
C3206 a_21785_5878# a_21840_5308# 0.002941f
C3207 a_24699_6200# a_24763_6143# 0.266837f
C3208 a_21863_4790# ringtest_0.x4.net5 2.02e-19
C3209 muxtest_0.R3R4 muxtest_0.R2R3 2.48395f
C3210 ringtest_0.x4._23_ a_26808_5308# 0.006211f
C3211 ringtest_0.x4.clknet_1_0__leaf_clk a_21399_5340# 0.158653f
C3212 ringtest_0.x4._18_ a_22795_5334# 4.57e-20
C3213 a_26808_5308# a_26367_4790# 2.96e-21
C3214 ringtest_0.x4.net7 VDPWR 1.83862f
C3215 a_26367_5340# a_26808_4902# 2.96e-21
C3216 a_26201_5340# a_26640_5156# 1.73e-19
C3217 ringtest_0.x4._11_ a_22392_5990# 0.032361f
C3218 a_21561_9116# ui_in[5] 2.06e-20
C3219 a_24336_6544# a_24527_5340# 6.46e-19
C3220 ringtest_0.x4.net3 a_21939_8054# 8.45e-20
C3221 a_24329_6640# a_24968_5308# 2.9e-20
C3222 ringtest_0.x4._15_ ringtest_0.x4._07_ 0.022092f
C3223 a_24536_6699# a_24361_5340# 2.08e-22
C3224 a_27273_4220# ringtest_0.x4.counter[8] 0.001844f
C3225 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.173286f
C3226 muxtest_0.x1.x3.GN3 ui_in[4] 7.93e-20
C3227 ringtest_0.x4._17_ VDPWR 2.38225f
C3228 ringtest_0.x4._07_ a_25263_5156# 2.91e-19
C3229 ringtest_0.x3.x2.GP2 m3_17046_7066# 2.65e-20
C3230 ringtest_0.x3.x1.nSEL1 VDPWR 0.646724f
C3231 ringtest_0.x4._19_ ringtest_0.x4._21_ 7.87e-20
C3232 ringtest_0.x4.clknet_0_clk a_24336_6544# 0.025079f
C3233 ringtest_0.x4.net6 a_22649_6244# 0.021756f
C3234 ui_in[3] ua[1] 4.1e-22
C3235 ringtest_0.x3.x2.GP3 ringtest_0.counter3 4.0653f
C3236 ringtest_0.x4.clknet_1_1__leaf_clk a_24699_6200# 7.2e-19
C3237 ringtest_0.x4._00_ a_22399_8976# 0.001531f
C3238 a_21561_9116# ringtest_0.x4._12_ 1.23e-19
C3239 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y 0.17253f
C3240 a_23963_4790# ringtest_0.x4.counter[4] 4.17e-20
C3241 ui_in[1] ui_in[5] 0.187526f
C3242 ringtest_0.x4._09_ a_26721_4246# 2.04e-21
C3243 a_16755_12091# ui_in[3] 0.279858f
C3244 a_22021_4220# a_22164_4362# 0.221119f
C3245 ringtest_0.x4.net8 a_24729_4790# 0.009204f
C3246 ringtest_0.x4.net7 ringtest_0.x4._25_ 3.01e-19
C3247 a_27065_5156# a_27191_4790# 0.006169f
C3248 ringtest_0.x4._23_ a_26555_4790# 0.012973f
C3249 ringtest_0.x4.net4 a_22499_4790# 0.00133f
C3250 a_26367_4790# a_26555_4790# 0.097994f
C3251 a_26808_4902# a_27065_5156# 0.036838f
C3252 a_24329_6640# a_25925_6788# 2.69e-21
C3253 ringtest_0.x4._17_ ringtest_0.x4._25_ 1.89e-19
C3254 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP1 2.55932f
C3255 ringtest_0.x4._06_ a_25225_5334# 9.38e-20
C3256 a_23349_6422# ringtest_0.x4._19_ 0.001413f
C3257 ringtest_0.x4._11_ a_26640_5334# 6.96e-20
C3258 a_24699_6200# a_24800_5334# 0.001605f
C3259 a_23879_6940# ringtest_0.x4._19_ 5.98e-19
C3260 ringtest_0.x4.counter[0] VDPWR 0.661077f
C3261 a_12297_23648# muxtest_0.x2.x2.GN2 0.106178f
C3262 a_22817_6146# VDPWR 0.386139f
C3263 ringtest_0.x4.clknet_1_1__leaf_clk a_23809_4790# 2.42e-19
C3264 ringtest_0.x4._08_ a_27065_5334# 0.013878f
C3265 ringtest_0.x4._21_ ringtest_0.x4.net9 0.170283f
C3266 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR 0.787508f
C3267 a_26095_6788# VDPWR 0.002069f
C3268 ringtest_0.x4.net4 a_21399_5340# 0.002039f
C3269 ringtest_0.x3.nselect2 ui_in[4] 0.001177f
C3270 ringtest_0.x4.clknet_1_1__leaf_clk a_22795_5334# 7.11e-20
C3271 ringtest_0.x4._15_ a_26201_5340# 0.069151f
C3272 ringtest_0.x4.net6 a_21587_5334# 1.35e-20
C3273 ringtest_0.x3.x1.nSEL0 a_16027_11759# 0.03096f
C3274 ringtest_0.x4._22_ a_26269_4612# 6.12e-20
C3275 ringtest_0.x4._13_ a_22350_5878# 2.65e-20
C3276 a_17405_12123# VDPWR 7.45e-19
C3277 ua[2] ua[5] 0.002786f
C3278 ringtest_0.x4._04_ a_21951_5878# 0.215918f
C3279 a_21785_5878# a_22392_5990# 0.136461f
C3280 ringtest_0.x3.x2.GN3 VDPWR 0.649844f
C3281 muxtest_0.x1.x3.GP1 ua[3] 0.0076f
C3282 ringtest_0.x4._01_ ringtest_0.x4._12_ 0.353697f
C3283 ringtest_0.x4._11_ a_25149_4220# 2.67e-19
C3284 a_25925_6788# a_25364_5878# 0.010774f
C3285 ringtest_0.x4.net7 ringtest_0.x4._21_ 0.326643f
C3286 ringtest_0.x4.clknet_1_0__leaf_clk a_21951_5878# 0.020113f
C3287 ringtest_0.x3.x2.GN4 m3_17032_8096# 7.07e-19
C3288 a_26749_6422# a_26839_6788# 0.004764f
C3289 a_18662_32213# ui_in[1] 0.02803f
C3290 ringtest_0.x4._16_ ringtest_0.x4.net5 0.096932f
C3291 ringtest_0.x4._17_ ringtest_0.x4._21_ 0.019243f
C3292 a_23879_6940# ringtest_0.x4.net9 1.97e-19
C3293 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A 0.428132f
C3294 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP3 0.060268f
C3295 ringtest_0.x4._08_ a_27149_5156# 1.22e-19
C3296 ringtest_0.x4._11_ a_24329_6640# 2.33e-19
C3297 a_20318_32213# a_20492_32319# 0.006584f
C3298 a_27065_5334# VDPWR 0.233266f
C3299 ringtest_0.x4._15_ a_22164_4362# 4.86e-20
C3300 ringtest_0.x4.net6 a_27273_4220# 4.97e-21
C3301 m2_18699_31802# ui_in[1] 0.183786f
C3302 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ui_in[3] 1.1e-22
C3303 a_19666_31955# muxtest_0.x1.x3.GN1 7.37e-20
C3304 muxtest_0.x1.x5.GN a_18662_32213# 0.001336f
C3305 a_24465_6800# ringtest_0.x4.net6 0.001158f
C3306 ringtest_0.x4.clknet_1_1__leaf_clk a_25421_6641# 0.035969f
C3307 a_23529_6422# ringtest_0.x4._15_ 2e-21
C3308 a_13501_23906# muxtest_0.R1R2 5.05e-21
C3309 a_23349_6422# ringtest_0.x4.net7 2.88e-19
C3310 a_23879_6940# ringtest_0.x4.net7 0.002812f
C3311 muxtest_0.x1.x5.GN m2_18699_31802# 4e-19
C3312 muxtest_0.x1.x3.GN3 ui_in[0] 0.254198f
C3313 a_19290_32287# ui_in[2] 1.22e-19
C3314 ringtest_0.x4._17_ a_23349_6422# 0.250762f
C3315 a_23879_6940# ringtest_0.x4._17_ 7.15e-19
C3316 ringtest_0.x4.net7 a_25309_5334# 0.001255f
C3317 a_12473_23980# ui_in[4] 0.254026f
C3318 ringtest_0.x4._11_ a_24545_5878# 1.22e-19
C3319 a_22201_9142# VDPWR 0.003202f
C3320 a_26627_4246# VDPWR 0.152186f
C3321 a_21852_9416# VDPWR 0.335402f
C3322 a_22817_6146# ringtest_0.x4._21_ 1.76e-19
C3323 a_27149_5156# VDPWR 0.005629f
C3324 ui_in[2] ui_in[3] 0.170107f
C3325 ringtest_0.x4._11_ a_25364_5878# 0.049204f
C3326 muxtest_0.x1.x3.GN2 muxtest_0.R1R2 0.006936f
C3327 a_24536_6699# VDPWR 0.266088f
C3328 muxtest_0.x1.x5.A muxtest_0.R6R7 4.52052f
C3329 ringtest_0.x4._01_ a_22245_8054# 0.014882f
C3330 ringtest_0.x4._12_ a_21785_8054# 0.001375f
C3331 ringtest_0.x4.net4 a_21951_5878# 0.34974f
C3332 ringtest_0.x4._15_ ringtest_0.x4._06_ 0.139237f
C3333 a_21561_8830# a_21845_8816# 0.030894f
C3334 ringtest_0.x4._15_ a_24070_5852# 6.77e-20
C3335 a_21465_8830# a_21852_8720# 0.034054f
C3336 ringtest_0.x4.net8 ringtest_0.x4._09_ 2.1e-20
C3337 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y 5.04e-19
C3338 ringtest_0.x4._23_ a_26817_4566# 4.18e-19
C3339 a_25149_4220# a_25345_4612# 0.00119f
C3340 ringtest_0.x4._11_ a_24551_4790# 0.001398f
C3341 a_25593_5156# ringtest_0.x4.counter[6] 2e-19
C3342 a_25364_5878# a_25761_5058# 0.001883f
C3343 a_21845_9116# a_21981_9142# 0.141453f
C3344 a_21233_5340# a_23151_5334# 4.04e-20
C3345 a_21852_9416# a_21803_9508# 6.32e-19
C3346 a_21675_9686# ringtest_0.x4.clknet_1_0__leaf_clk 2.59e-19
C3347 ringtest_0.x4.net2 a_21465_8830# 0.004306f
C3348 ringtest_0.x4._18_ a_22224_6244# 5.13e-20
C3349 a_22649_6244# ringtest_0.x4.net5 4.89e-20
C3350 ringtest_0.x4._11_ a_24317_4942# 0.046716f
C3351 a_25421_6641# ringtest_0.x4._23_ 1.03e-19
C3352 ringtest_0.x4._05_ a_26749_6422# 4.21e-20
C3353 ringtest_0.x4.net1 a_21852_9416# 0.006588f
C3354 a_22111_10993# a_21845_9116# 6.9e-23
C3355 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._24_ 0.041474f
C3356 ringtest_0.x4.net10 a_27489_3702# 1.3e-21
C3357 ringtest_0.x4._14_ VDPWR 0.685574f
C3358 ringtest_0.x4.net6 a_26201_4790# 5.6e-22
C3359 ringtest_0.x4._15_ a_23891_4790# 1.25e-19
C3360 ringtest_0.x4._11_ a_23151_5334# 0.00137f
C3361 ringtest_0.x4._16_ a_24527_5340# 9.89e-20
C3362 a_13025_23980# muxtest_0.x2.x2.GP3 5.21e-19
C3363 ringtest_0.x4.net9 a_24968_5308# 2.05e-20
C3364 muxtest_0.x1.x3.GP2 ui_in[0] 4.71e-19
C3365 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP3 3.4436f
C3366 a_22319_6244# VDPWR 0.003961f
C3367 a_25336_4902# a_25294_4790# 4.62e-19
C3368 a_24895_4790# a_26201_4790# 3.23e-19
C3369 ringtest_0.x4._15_ a_22373_5156# 1.6e-20
C3370 muxtest_0.x2.nselect2 a_13501_23906# 9.77e-20
C3371 ringtest_0.x4.clknet_0_clk ringtest_0.x4._16_ 0.019509f
C3372 ringtest_0.x4.net5 a_23467_4818# 2.72e-19
C3373 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR 0.639974f
C3374 ringtest_0.x4.net6 a_26555_5334# 3.93e-20
C3375 muxtest_0.R7R8 muxtest_0.x2.x2.GN2 1.22e-19
C3376 ringtest_0.x4._22_ a_26895_3867# 1.85e-19
C3377 a_22392_5990# a_22775_5878# 4.67e-20
C3378 muxtest_0.R3R4 ui_in[4] 3.8e-21
C3379 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x2.GN2 3.88e-22
C3380 a_22541_5058# a_22373_5156# 0.310858f
C3381 clk ena 0.031023f
C3382 ringtest_0.x4.net7 a_24968_5308# 0.040813f
C3383 a_24883_6800# ringtest_0.x4._22_ 0.001069f
C3384 a_21785_8054# a_22245_8054# 0.001479f
C3385 ringtest_0.x4._12_ a_22695_8304# 0.001754f
C3386 a_25055_3867# a_25975_3867# 1.37e-20
C3387 a_25294_4790# VDPWR 1.42e-19
C3388 ringtest_0.x4._17_ a_24968_5308# 1.03e-20
C3389 a_22043_5156# VDPWR 0.005794f
C3390 muxtest_0.x1.x3.GP3 muxtest_0.x1.x4.A 0.358376f
C3391 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A 0.446595f
C3392 a_26640_5334# ringtest_0.x4.net10 3.33e-19
C3393 a_27233_5308# a_27191_5712# 7.84e-20
C3394 ringtest_0.x4.clknet_1_0__leaf_clk a_22052_8875# 0.037641f
C3395 ringtest_0.x4.net4 a_23381_4584# 0.083888f
C3396 a_24536_6699# ringtest_0.x4._21_ 0.0043f
C3397 ui_in[4] ui_in[5] 0.278355f
C3398 ringtest_0.x4._11_ ringtest_0.x4._19_ 0.032711f
C3399 ringtest_0.x4._15_ a_26269_4612# 0.00403f
C3400 a_19666_31955# muxtest_0.x1.x3.GP3 0.001353f
C3401 ringtest_0.x4._23_ ringtest_0.x4._24_ 0.206353f
C3402 ringtest_0.x4.net7 a_25925_6788# 0.168744f
C3403 ringtest_0.x4._24_ a_26367_4790# 0.03707f
C3404 ringtest_0.x4._00_ a_21465_9294# 0.001095f
C3405 a_21425_9686# a_21852_9416# 0.00324f
C3406 a_26749_6422# ringtest_0.x4._09_ 2.51e-21
C3407 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ui_in[3] 0.001551f
C3408 ringtest_0.x4._09_ ringtest_0.x4.net11 0.071633f
C3409 ringtest_0.x4.net3 ringtest_0.x4.net5 9.15e-21
C3410 ringtest_0.x4._02_ a_21672_5334# 8.22e-19
C3411 a_21233_5340# a_22265_5308# 0.048748f
C3412 ringtest_0.x4._22_ a_26808_5308# 9.3e-20
C3413 ringtest_0.x4._17_ a_25925_6788# 0.139841f
C3414 ringtest_0.x4._04_ a_22795_5334# 0.072162f
C3415 ringtest_0.x4._18_ a_24336_6544# 1.59e-19
C3416 ringtest_0.x4._10_ VDPWR 0.249351f
C3417 ringtest_0.x4._20_ a_25083_4790# 5.09e-20
C3418 ringtest_0.x4.net8 a_24361_5340# 0.036074f
C3419 a_23879_6940# a_24536_6699# 0.007109f
C3420 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP2 0.005192f
C3421 ringtest_0.x4._11_ a_22265_5308# 0.033019f
C3422 a_26721_4246# VDPWR 0.191262f
C3423 muxtest_0.x1.x4.A muxtest_0.R1R2 4.5214f
C3424 muxtest_0.x2.x1.nSEL0 ui_in[4] 0.13767f
C3425 a_16203_12091# a_16579_11759# 3.02e-19
C3426 ringtest_0.x3.x1.nSEL1 a_15749_12123# 0.00175f
C3427 a_22541_5058# a_22499_4790# 7.84e-20
C3428 ringtest_0.x4._11_ ringtest_0.x4.net9 0.233741f
C3429 ringtest_0.x4.clknet_1_1__leaf_clk a_27233_5308# 9.45e-20
C3430 muxtest_0.x1.x3.GN3 muxtest_0.x2.x2.GN4 8.02e-21
C3431 a_12977_24040# VDPWR 0.001496f
C3432 ringtest_0.x4.net6 a_23770_5308# 0.050235f
C3433 ringtest_0.x4.clknet_0_clk a_26201_6788# 6.75e-20
C3434 muxtest_0.x2.x2.GN2 VDPWR 0.601936f
C3435 a_24361_5340# a_24729_4790# 0.012779f
C3436 ringtest_0.x4.net3 a_21007_3867# 0.006292f
C3437 ringtest_0.x4.clknet_1_0__leaf_clk a_21803_8598# 0.002574f
C3438 a_24045_6654# a_23837_5878# 9.42e-20
C3439 ringtest_0.x4._16_ a_25168_5156# 7.37e-22
C3440 a_24336_6544# a_24763_6143# 0.003687f
C3441 ringtest_0.x4._11_ ringtest_0.x4.net7 0.966176f
C3442 a_21509_4790# VDPWR 0.741952f
C3443 ringtest_0.x4.net9 a_25761_5058# 0.115737f
C3444 a_22265_5308# a_21675_4790# 0.00183f
C3445 a_26640_5156# a_26895_3867# 6.36e-19
C3446 ringtest_0.x4.net11 a_27659_4246# 0.004987f
C3447 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A 0.17253f
C3448 ringtest_0.x4.net1 ringtest_0.x4._10_ 0.033245f
C3449 a_25925_6788# a_26095_6788# 0.001675f
C3450 ringtest_0.x4._11_ ringtest_0.x4._17_ 0.113734f
C3451 a_26201_5340# a_26367_5340# 0.970499f
C3452 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GP1 1.17e-19
C3453 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN4 2.26e-20
C3454 a_22765_5308# VDPWR 0.252112f
C3455 ringtest_0.x4.clknet_1_1__leaf_clk a_25977_4220# 3.39e-19
C3456 a_23949_6654# a_24264_6788# 7.84e-20
C3457 ringtest_0.x4._16_ a_22983_5654# 3.98e-19
C3458 a_25364_5878# ringtest_0.x4.net10 3.58e-19
C3459 muxtest_0.x1.x5.GN a_18836_32319# 1.95e-19
C3460 ringtest_0.x4.net7 a_25761_5058# 0.064911f
C3461 ringtest_0.x4._03_ a_22939_4584# 1.17e-19
C3462 a_24336_6544# ringtest_0.x4.clknet_1_1__leaf_clk 0.013843f
C3463 a_12297_23648# muxtest_0.x2.x2.GP1 9.92e-19
C3464 a_21867_8054# VDPWR 2.01e-19
C3465 ringtest_0.x4.net4 a_22795_5334# 0.005199f
C3466 a_24627_6200# a_24545_5878# 2.78e-19
C3467 a_24763_6143# a_24986_5878# 3.74e-19
C3468 ringtest_0.x4._13_ VDPWR 0.524973f
C3469 a_17231_12017# ringtest_0.x3.x2.GN4 0.134079f
C3470 ringtest_0.x3.x2.GN2 a_16155_12151# 0.002418f
C3471 ua[3] ua[1] 0.003505f
C3472 a_21785_5878# a_22265_5308# 4.12e-19
C3473 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN2 0.065153f
C3474 ringtest_0.x4._04_ a_21672_5334# 3.3e-20
C3475 ringtest_0.x4._22_ ringtest_0.x4.counter[6] 9.35e-22
C3476 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR 0.636657f
C3477 a_24699_6200# ringtest_0.x4._22_ 0.019192f
C3478 ui_in[0] ui_in[5] 0.21609f
C3479 ringtest_0.x4._23_ a_27233_5308# 1.75e-20
C3480 ringtest_0.x4.clknet_1_0__leaf_clk a_21672_5334# 0.032164f
C3481 a_26201_5340# a_27065_5156# 1.29e-19
C3482 a_26640_5334# a_26808_4902# 3.15e-19
C3483 a_26808_5308# a_26640_5156# 3.15e-19
C3484 ringtest_0.x4._18_ a_23899_5334# 3.94e-20
C3485 ringtest_0.x4._16_ a_22486_4246# 0.00427f
C3486 muxtest_0.x1.x4.A muxtest_0.x2.nselect2 0.01287f
C3487 ringtest_0.x4._11_ a_22817_6146# 0.052724f
C3488 a_21845_9116# ui_in[5] 1.25e-19
C3489 ringtest_0.x4.net9 a_25345_4612# 0.001755f
C3490 a_24336_6544# a_24800_5334# 9.47e-20
C3491 ringtest_0.x4._08_ ringtest_0.x4.net8 2.38e-19
C3492 ringtest_0.x4._11_ a_26095_6788# 0.001703f
C3493 muxtest_0.x2.x2.GP3 ui_in[3] 4.18e-19
C3494 ringtest_0.x4.net3 ringtest_0.x4._12_ 0.271994f
C3495 ringtest_0.x4._15_ a_26895_3867# 0.006207f
C3496 muxtest_0.x1.x3.GN2 muxtest_0.R6R7 4.03742f
C3497 ringtest_0.x4.net1 a_21867_8054# 0.00162f
C3498 ringtest_0.x4.clknet_0_clk a_24465_6800# 0.003343f
C3499 a_21845_9116# ringtest_0.x4._12_ 2.52e-19
C3500 ringtest_0.x4._07_ a_23381_4818# 2.73e-21
C3501 ringtest_0.x3.x2.GN1 m2_15612_11606# 0.06935f
C3502 ringtest_0.x4._09_ a_27659_4246# 2.25e-19
C3503 ringtest_0.counter7 ringtest_0.x4.counter[9] 2.14e-19
C3504 ringtest_0.x4._23_ a_25977_4220# 0.130093f
C3505 ringtest_0.x3.x2.GN1 ui_in[3] 0.021168f
C3506 ringtest_0.x4.net8 a_25336_4902# 0.00264f
C3507 ringtest_0.drv_out ringtest_0.x3.x2.GP3 0.077808f
C3508 ringtest_0.x4._17_ a_21785_5878# 1.5e-21
C3509 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ui_in[3] 1.61e-19
C3510 muxtest_0.x1.x3.GP3 ua[0] 0.17111f
C3511 a_26640_5156# a_26555_4790# 0.037333f
C3512 a_21951_5878# a_22541_5058# 8.13e-20
C3513 a_27233_5058# a_27065_5156# 0.310858f
C3514 ringtest_0.x4.net10 a_26913_4566# 0.002966f
C3515 ringtest_0.x4.clknet_1_1__leaf_clk a_25677_5156# 1.62e-19
C3516 ringtest_0.x4.net6 a_24895_4790# 0.045685f
C3517 a_12849_23648# a_12977_24040# 0.004764f
C3518 a_25364_5878# a_25393_5308# 0.009572f
C3519 a_23529_6422# a_23949_6654# 0.017007f
C3520 ringtest_0.x4.net8 VDPWR 1.78891f
C3521 a_12849_23648# muxtest_0.x2.x2.GN2 1.63e-19
C3522 a_24729_4790# a_25336_4902# 0.141453f
C3523 ui_in[3] ui_in[6] 0.153563f
C3524 a_18662_32213# ui_in[0] 0.048888f
C3525 a_26839_6788# VDPWR 6.35e-19
C3526 ringtest_0.x4.net4 a_21672_5334# 4.27e-19
C3527 ringtest_0.x4.clknet_1_1__leaf_clk a_23899_5334# 0.001857f
C3528 ringtest_0.x4._03_ ringtest_0.x4.net5 3.86e-19
C3529 ringtest_0.x3.x1.nSEL0 a_16579_11759# 1.91e-20
C3530 ringtest_0.x4._15_ a_26808_5308# 4.57e-19
C3531 m2_18699_31802# ui_in[0] 0.130999f
C3532 ringtest_0.x4._22_ a_26817_4566# 1.37e-20
C3533 ringtest_0.x4.net10 a_26735_5334# 8.52e-20
C3534 a_21785_5878# a_22817_6146# 0.048608f
C3535 ringtest_0.x4._04_ a_22224_6244# 0.01404f
C3536 a_24729_4790# VDPWR 0.727748f
C3537 ringtest_0.x4.net3 a_22245_8054# 0.001478f
C3538 ringtest_0.x4._11_ a_26627_4246# 0.054652f
C3539 muxtest_0.R1R2 ua[0] 2.31469f
C3540 ringtest_0.x4.clknet_1_0__leaf_clk a_22224_6244# 0.002436f
C3541 a_21845_9116# a_22245_8054# 4.52e-21
C3542 ringtest_0.x4._18_ ringtest_0.x4._16_ 0.283975f
C3543 ringtest_0.x4._07_ ringtest_0.x4._20_ 1.72e-19
C3544 a_25364_5878# a_26808_4902# 7.13e-20
C3545 a_26749_6422# ringtest_0.x4._08_ 0.001905f
C3546 a_19290_32287# ui_in[1] 0.254026f
C3547 ringtest_0.x4._25_ a_26839_6788# 8.17e-20
C3548 a_24968_5308# a_25351_5712# 4.67e-20
C3549 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A 5.04e-19
C3550 ringtest_0.x4._11_ a_24536_6699# 3.53e-20
C3551 a_23949_6654# a_24070_5852# 0.002561f
C3552 a_21465_9294# a_21465_8830# 0.025128f
C3553 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GN4 0.057602f
C3554 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1 2.99928f
C3555 a_21798_5712# VDPWR 4.21e-19
C3556 a_19242_32347# VDPWR 5.13e-19
C3557 ringtest_0.x4._15_ a_23381_4584# 0.110742f
C3558 ringtest_0.x4.net9 ringtest_0.x4.net10 0.022804f
C3559 ringtest_0.x4.net6 a_27169_6641# 1.17e-21
C3560 ui_in[1] ui_in[3] 0.006066f
C3561 ui_in[2] ua[3] 0.781024f
C3562 ringtest_0.x4._15_ a_26555_4790# 0.005742f
C3563 a_25593_5156# a_25977_4220# 0.009905f
C3564 muxtest_0.x1.x5.GN a_19290_32287# 3.26e-19
C3565 a_25593_5156# a_25719_4790# 0.006169f
C3566 a_24045_6654# ringtest_0.x4._15_ 1.09e-20
C3567 ringtest_0.x4._14_ a_21233_5340# 0.001276f
C3568 a_22373_5156# a_22765_4478# 0.001309f
C3569 ringtest_0.x4.counter[1] VDPWR 0.349593f
C3570 a_24763_6143# ringtest_0.x4._16_ 0.060109f
C3571 m3_17036_9140# m3_17032_8096# 0.003764f
C3572 muxtest_0.R3R4 muxtest_0.x2.x2.GN4 0.269437f
C3573 ringtest_0.x4.net9 a_24627_6200# 0.004319f
C3574 ringtest_0.x4.net7 ringtest_0.x4.net10 6.54e-19
C3575 a_13025_23980# ui_in[4] 0.127717f
C3576 ringtest_0.x4._11_ ringtest_0.x4._14_ 0.007676f
C3577 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.nselect2 0.047548f
C3578 muxtest_0.x2.x1.nSEL0 a_11845_23906# 0.081627f
C3579 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR 0.636415f
C3580 a_22390_4566# VDPWR 0.007674f
C3581 ringtest_0.x4._16_ a_22295_3867# 4.24e-19
C3582 a_24004_6128# ringtest_0.x4._06_ 0.111795f
C3583 a_26749_6422# VDPWR 0.178246f
C3584 a_22052_9116# VDPWR 0.286747f
C3585 ringtest_0.x4.net11 VDPWR 0.794015f
C3586 ringtest_0.x4.net8 ringtest_0.x4._21_ 0.333812f
C3587 ringtest_0.x4._11_ a_22319_6244# 0.00121f
C3588 ringtest_0.counter3 ringtest_0.x4.counter[0] 0.117902f
C3589 a_24070_5852# a_24004_6128# 0.221119f
C3590 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A a_16027_11759# 2.51e-19
C3591 a_24329_6640# a_24715_5334# 6.17e-21
C3592 ringtest_0.x4._05_ VDPWR 0.240335f
C3593 ringtest_0.x4._24_ ringtest_0.x4._22_ 0.01067f
C3594 ringtest_0.x4.net4 a_22224_6244# 0.034877f
C3595 ringtest_0.x4._23_ ringtest_0.x4.counter[9] 7.62e-19
C3596 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._16_ 0.001692f
C3597 ringtest_0.x4.net3 a_21591_6128# 0.001185f
C3598 a_21465_8830# a_21981_8976# 1.28e-19
C3599 ringtest_0.x4._15_ a_24699_6200# 2.91e-20
C3600 a_21845_8816# a_21852_8720# 0.969092f
C3601 ringtest_0.x4.net6 a_23932_6128# 0.002624f
C3602 ringtest_0.x4.net3 a_22486_4246# 1.66e-19
C3603 ringtest_0.x4._17_ a_24627_6200# 4.44e-20
C3604 ringtest_0.x4._23_ a_27491_4566# 3.52e-19
C3605 a_25149_4220# a_25547_4612# 0.005781f
C3606 ringtest_0.x4._11_ a_25294_4790# 0.002651f
C3607 ringtest_0.x4._14_ a_21675_4790# 5.98e-19
C3608 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP2 4.55678f
C3609 ringtest_0.x4._21_ a_24729_4790# 5.62e-21
C3610 ringtest_0.x4.clknet_1_0__leaf_clk a_21780_9142# 0.001704f
C3611 a_26749_6422# ringtest_0.x4._25_ 0.082413f
C3612 ringtest_0.x3.x2.GN3 ringtest_0.counter3 3.89796f
C3613 ringtest_0.x4.counter[0] ua[2] 1.11e-19
C3614 a_21852_9416# a_22399_9142# 0.095025f
C3615 ringtest_0.x4._08_ ringtest_0.x4._09_ 0.013938f
C3616 a_21561_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.038899f
C3617 ringtest_0.x4.net2 a_21845_8816# 3.07e-19
C3618 a_21845_9116# a_22228_9508# 0.002698f
C3619 ringtest_0.x4._18_ a_22649_6244# 3.43e-19
C3620 a_23879_6940# ringtest_0.x4.net8 0.001938f
C3621 ringtest_0.x4._11_ a_22043_5156# 6.67e-19
C3622 ringtest_0.ring_out ringtest_0.x3.x2.GN4 0.080391f
C3623 ringtest_0.x4._05_ ringtest_0.x4._25_ 4.6e-21
C3624 ringtest_0.x4.net1 a_22052_9116# 0.002893f
C3625 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ui_in[3] 5.64e-20
C3626 ringtest_0.drv_out a_17231_12017# 3.86e-20
C3627 ringtest_0.x4.net8 a_25309_5334# 9.28e-20
C3628 ua[2] ua[4] 0.002786f
C3629 ringtest_0.x4._16_ a_24800_5334# 0.00213f
C3630 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP3 0.002439f
C3631 ringtest_0.x4.net9 a_25393_5308# 0.007609f
C3632 ringtest_0.x4._08_ a_26766_5712# 0.001882f
C3633 a_22350_5878# VDPWR 3.37e-19
C3634 a_25593_5156# a_25677_5156# 0.008508f
C3635 ringtest_0.x4.clknet_0_clk a_23770_5308# 8.98e-21
C3636 ringtest_0.x4.net6 ringtest_0.x4.net5 0.003368f
C3637 ringtest_0.x4._15_ a_23809_4790# 0.080244f
C3638 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN4 2.26e-20
C3639 muxtest_0.x2.nselect2 muxtest_0.x2.x2.GN3 7.39e-21
C3640 ringtest_0.x3.x2.GP2 ui_in[4] 1.37e-19
C3641 ringtest_0.x4.net6 a_24895_5334# 0.001259f
C3642 a_22817_6146# a_22775_5878# 7.84e-20
C3643 a_17377_14114# ui_in[6] 0.040112f
C3644 ringtest_0.x4.counter[1] ringtest_0.x4.counter[2] 0.070133f
C3645 a_22116_4902# a_21863_4790# 3.39e-19
C3646 a_22541_5058# a_23809_4790# 3.71e-21
C3647 ringtest_0.x3.x1.nSEL1 a_15575_12017# 0.193944f
C3648 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A a_16579_11759# 2.51e-19
C3649 ringtest_0.x4.net7 a_25393_5308# 0.08513f
C3650 muxtest_0.x2.x2.GP1 VDPWR 1.85798f
C3651 a_25975_3867# a_26895_3867# 1.37e-20
C3652 a_21785_5878# a_22319_6244# 0.002698f
C3653 ringtest_0.x4._09_ VDPWR 0.262387f
C3654 ringtest_0.x4._04_ a_22139_5878# 0.126198f
C3655 ringtest_0.x4._10_ ringtest_0.x4._11_ 0.033565f
C3656 ringtest_0.x4._11_ a_26721_4246# 0.039972f
C3657 a_22795_5334# a_22541_5058# 0.001352f
C3658 ringtest_0.x4._23_ ringtest_0.x4._16_ 3.32e-22
C3659 ringtest_0.x4.net9 a_27191_4790# 6.87e-19
C3660 a_12297_23648# VDPWR 0.161892f
C3661 ringtest_0.x4._17_ a_25393_5308# 4.35e-22
C3662 ringtest_0.x4.clknet_1_0__leaf_clk a_22139_5878# 0.003123f
C3663 a_21852_8720# a_22201_8964# 2.36e-19
C3664 a_21981_8976# a_21780_8964# 4.67e-20
C3665 a_21845_8816# a_22399_8976# 0.057611f
C3666 a_21561_8830# a_21803_8598# 0.008508f
C3667 a_22074_4790# VDPWR 0.003212f
C3668 ringtest_0.x4.net9 a_26808_4902# 0.022365f
C3669 ringtest_0.x3.x2.GP3 m3_17036_9140# 9.67e-19
C3670 a_27065_5334# ringtest_0.x4.net10 0.00375f
C3671 a_23993_5654# a_23899_5334# 1.26e-19
C3672 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._01_ 0.05158f
C3673 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A 0.446529f
C3674 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP3 0.061475f
C3675 a_12019_24012# ui_in[3] 9.55e-19
C3676 a_21233_5340# a_21509_4790# 0.001876f
C3677 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A 0.17253f
C3678 ringtest_0.x4._15_ a_26817_4566# 0.004129f
C3679 a_19666_31955# muxtest_0.x1.x3.GN4 6.84e-19
C3680 ringtest_0.drv_out a_24329_6640# 4.16e-19
C3681 ringtest_0.x4._24_ a_26640_5156# 0.010089f
C3682 ringtest_0.x4._00_ a_21852_9416# 0.208988f
C3683 ringtest_0.x4._11_ a_21509_4790# 0.005486f
C3684 ringtest_0.x4.net7 a_26808_4902# 1.23e-19
C3685 ringtest_0.x4.net3 ringtest_0.counter7 4.2e-20
C3686 a_21233_5340# a_22765_5308# 1.05e-19
C3687 ringtest_0.x4._02_ a_22097_5334# 3.18e-19
C3688 ringtest_0.x4.net5 a_22939_4584# 0.002311f
C3689 ringtest_0.x4.clknet_1_0__leaf_clk a_21863_4790# 0.003207f
C3690 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP2 0.043302f
C3691 ringtest_0.x4._16_ ringtest_0.x4._02_ 3.22e-20
C3692 ringtest_0.x4._18_ a_24465_6800# 7.52e-20
C3693 ringtest_0.x4.net10 a_26627_4246# 0.27342f
C3694 a_23349_6422# ringtest_0.x4._05_ 4.45e-20
C3695 a_23879_6940# ringtest_0.x4._05_ 0.005813f
C3696 ringtest_0.x4.net8 a_24968_5308# 0.001066f
C3697 a_18836_32319# ui_in[0] 9.55e-19
C3698 ringtest_0.x4._11_ a_22765_5308# 0.001227f
C3699 a_27659_4246# VDPWR 0.009314f
C3700 ringtest_0.x4.net10 a_27149_5156# 3.08e-19
C3701 ringtest_0.x3.x2.GN2 ui_in[4] 0.108649f
C3702 a_16027_11759# a_16155_12151# 0.004764f
C3703 ringtest_0.x4._08_ a_24361_5340# 3.42e-20
C3704 a_16027_11759# ringtest_0.x3.x2.GN1 0.012445f
C3705 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR 0.636415f
C3706 a_16579_11759# a_16755_12091# 0.185422f
C3707 ringtest_0.x4._13_ a_21233_5340# 3.88e-19
C3708 muxtest_0.x1.x3.GP1 muxtest_0.R1R2 2.46e-21
C3709 ringtest_0.x4._11_ a_21867_8054# 1.17e-19
C3710 ringtest_0.x4._07_ a_25149_4220# 9.24e-19
C3711 uio_in[2] uio_in[1] 0.031023f
C3712 a_21509_4790# a_21675_4790# 0.970278f
C3713 ringtest_0.x4.net6 a_24527_5340# 0.048602f
C3714 a_21375_3867# ringtest_0.x4.counter[1] 0.1107f
C3715 ringtest_0.x4.clknet_0_clk a_24712_6422# 4.01e-19
C3716 ringtest_0.drv_out a_25364_5878# 1.27e-19
C3717 ringtest_0.x4._22_ a_25977_4220# 0.191159f
C3718 ringtest_0.x4.net4 a_22139_5878# 0.011292f
C3719 ringtest_0.x4._11_ ringtest_0.x4._13_ 0.217373f
C3720 a_24361_5340# a_25336_4902# 3.92e-19
C3721 ringtest_0.x4._22_ a_25719_4790# 7.63e-20
C3722 a_24968_5308# a_24729_4790# 1.62e-19
C3723 a_24527_5340# a_24895_4790# 1.17e-19
C3724 muxtest_0.x1.x3.GN3 muxtest_0.R3R4 0.377005f
C3725 ringtest_0.x4.net3 a_22295_3867# 0.001252f
C3726 ringtest_0.x4.clknet_1_0__leaf_clk a_21785_8054# 0.024338f
C3727 a_25149_4220# a_25055_3867# 3.27e-19
C3728 a_24329_6640# ringtest_0.x4._07_ 5.99e-19
C3729 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net6 0.087511f
C3730 a_24336_6544# ringtest_0.x4._22_ 8.56e-19
C3731 ringtest_0.x4.net9 a_25083_4790# 1.61e-19
C3732 a_27233_5058# a_27489_3702# 3.35e-20
C3733 a_22265_5308# a_21948_5156# 0.005602f
C3734 a_22097_5334# a_22116_4902# 3.73e-19
C3735 ringtest_0.x4.clknet_0_clk a_24895_4790# 3.43e-21
C3736 ringtest_0.x4._18_ a_22733_6244# 1.72e-19
C3737 m2_15612_11606# ui_in[4] 0.183786f
C3738 ringtest_0.x4._16_ a_22116_4902# 0.005579f
C3739 a_26367_5340# a_26808_5308# 0.118966f
C3740 a_26201_5340# a_26640_5334# 0.273138f
C3741 a_21399_5340# a_22181_5334# 6.32e-19
C3742 ui_in[3] ui_in[4] 13.523f
C3743 ringtest_0.x4._15_ ringtest_0.x4._24_ 0.032103f
C3744 a_24361_5340# VDPWR 0.421866f
C3745 ringtest_0.x4._16_ a_23993_5654# 3.31e-19
C3746 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ui_in[3] 9.57e-20
C3747 ringtest_0.x4.net4 a_21863_4790# 4.45e-19
C3748 ringtest_0.x4.net9 a_24715_5334# 1.41e-19
C3749 a_21785_5878# a_21509_4790# 2.82e-20
C3750 ringtest_0.x4.net7 a_25083_4790# 4.68e-19
C3751 a_12849_23648# muxtest_0.x2.x2.GP1 1.21e-20
C3752 a_24465_6800# ringtest_0.x4.clknet_1_1__leaf_clk 1.17e-20
C3753 a_21395_6940# VDPWR 1.52032f
C3754 ringtest_0.counter7 a_26201_4790# 2.09e-20
C3755 ringtest_0.x3.x2.GN4 a_17405_12123# 0.001562f
C3756 ringtest_0.x4._22_ a_24986_5878# 0.006962f
C3757 muxtest_0.x2.x2.GP3 ua[3] 0.084041f
C3758 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP1 2.56189f
C3759 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GN4 0.071282f
C3760 a_21132_8918# VDPWR 4.93e-19
C3761 muxtest_0.x1.x1.nSEL1 ui_in[2] 0.164995f
C3762 ringtest_0.x4._04_ a_22097_5334# 0.001211f
C3763 a_21785_5878# a_22765_5308# 0.002539f
C3764 a_25364_5878# ringtest_0.x4._07_ 0.022424f
C3765 ringtest_0.x4.net7 a_24715_5334# 0.014734f
C3766 ringtest_0.x4._04_ ringtest_0.x4._16_ 0.025302f
C3767 ringtest_0.x4.clknet_1_0__leaf_clk a_22097_5334# 0.004501f
C3768 a_25975_3867# ringtest_0.x4.counter[6] 0.1107f
C3769 a_26367_5340# a_26555_4790# 1.41e-20
C3770 ringtest_0.x4._11_ ringtest_0.x4.net8 0.418201f
C3771 ringtest_0.x4.net9 a_25547_4612# 6.77e-19
C3772 a_21951_5878# a_24004_6128# 1.23e-20
C3773 a_21981_9142# ui_in[5] 2.79e-20
C3774 muxtest_0.R7R8 muxtest_0.R5R6 0.318606f
C3775 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._16_ 4.14e-20
C3776 ringtest_0.x4._05_ a_24968_5308# 8.7e-19
C3777 muxtest_0.x1.x3.GP2 muxtest_0.R3R4 0.170487f
C3778 ringtest_0.x4._13_ a_21785_5878# 0.002226f
C3779 muxtest_0.x2.x2.GP3 m3_13316_18955# 0.006132f
C3780 a_22111_10993# ui_in[5] 0.231636f
C3781 ringtest_0.ring_out ringtest_0.drv_out 2.13841f
C3782 muxtest_0.x1.x3.GN1 muxtest_0.R4R5 0.334962f
C3783 ringtest_0.x4.net1 a_21395_6940# 0.001584f
C3784 muxtest_0.R7R8 VDPWR 3.21675f
C3785 a_21981_9142# ringtest_0.x4._12_ 7.61e-20
C3786 ringtest_0.x4._07_ a_24317_4942# 1.81e-19
C3787 ringtest_0.x3.x2.GP1 ui_in[3] 8.3e-19
C3788 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A 5.04e-19
C3789 ringtest_0.x4._23_ a_27273_4220# 0.220841f
C3790 ringtest_0.x4.net1 a_21132_8918# 0.001512f
C3791 ringtest_0.x4.net7 a_25547_4612# 0.001525f
C3792 a_22765_4478# a_23381_4584# 0.013543f
C3793 ringtest_0.drv_out ringtest_0.x4._19_ 0.013619f
C3794 ringtest_0.x4.net8 a_25761_5058# 0.020836f
C3795 ringtest_0.x4._11_ a_24729_4790# 0.029022f
C3796 a_26808_4902# a_26627_4246# 3.15e-19
C3797 ringtest_0.x4._23_ a_26766_4790# 6.82e-19
C3798 a_19114_31955# a_19242_32347# 0.004764f
C3799 ringtest_0.x4._02_ a_21587_5334# 0.114994f
C3800 a_26808_4902# a_27149_5156# 9.73e-19
C3801 a_22224_6244# a_22541_5058# 2.18e-19
C3802 ringtest_0.x4._05_ a_25925_6788# 1.27e-19
C3803 muxtest_0.x1.x3.GN4 ua[0] 4.10932f
C3804 a_21399_5340# a_21840_5308# 0.127288f
C3805 ringtest_0.x4.clknet_1_1__leaf_clk a_26201_4790# 0.306202f
C3806 ringtest_0.x4.net10 a_26721_4246# 0.007482f
C3807 ringtest_0.x4.net6 a_25168_5156# 6.05e-21
C3808 a_13025_23980# muxtest_0.x2.x2.GN4 0.003699f
C3809 ringtest_0.x4._11_ a_21798_5712# 4.01e-19
C3810 ringtest_0.x4._21_ a_24361_5340# 0.016583f
C3811 a_25364_5878# a_26201_5340# 0.016172f
C3812 a_13501_23906# muxtest_0.x2.x2.GN2 7.58e-21
C3813 muxtest_0.x2.x2.GN1 a_12019_24012# 0.001144f
C3814 a_23949_6654# a_24045_6654# 0.310858f
C3815 a_23529_6422# a_24329_6640# 2.3e-20
C3816 muxtest_0.x2.x2.GN2 ua[2] 0.429379f
C3817 a_24895_4790# a_25168_5156# 0.074022f
C3818 a_24729_4790# a_25761_5058# 0.048748f
C3819 a_19290_32287# ui_in[0] 0.143958f
C3820 ringtest_0.x4._08_ VDPWR 0.467036f
C3821 ringtest_0.x4.net4 a_22097_5334# 0.006897f
C3822 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR 0.636362f
C3823 ringtest_0.x4.clknet_1_1__leaf_clk a_26555_5334# 3.58e-19
C3824 muxtest_0.R2R3 ua[3] 0.017699f
C3825 ringtest_0.x4._15_ a_27233_5308# 1.61e-19
C3826 ringtest_0.x4.net6 a_22983_5654# 0.001315f
C3827 ringtest_0.x4.net3 ringtest_0.x4._02_ 0.031079f
C3828 ringtest_0.x4._22_ a_27491_4566# 3.34e-21
C3829 ringtest_0.x4.net4 ringtest_0.x4._16_ 0.442589f
C3830 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GN3 1.1e-19
C3831 ringtest_0.drv_out ringtest_0.x4.net9 4.05e-20
C3832 ui_in[0] ui_in[3] 0.001641f
C3833 ringtest_0.counter3 ringtest_0.x4._13_ 0.003357f
C3834 ringtest_0.x4._04_ a_22649_6244# 0.006456f
C3835 a_21785_5878# ringtest_0.x4.net8 9.67e-20
C3836 a_25336_4902# VDPWR 0.183641f
C3837 ringtest_0.x4.net8 a_25345_4612# 0.005557f
C3838 ringtest_0.x4._18_ a_23770_5308# 0.079699f
C3839 ringtest_0.x4._11_ a_22390_4566# 9.44e-19
C3840 a_23879_6940# a_24361_5340# 3.84e-19
C3841 a_20492_32319# ui_in[1] 8.84e-19
C3842 ringtest_0.x4.clknet_1_0__leaf_clk a_22649_6244# 6.75e-21
C3843 ringtest_0.x4._11_ ringtest_0.x4.net11 2.31e-19
C3844 muxtest_0.R5R6 VDPWR 1.61253f
C3845 muxtest_0.x1.x5.GN ua[3] 0.820663f
C3846 a_24329_6640# ringtest_0.x4._06_ 0.002324f
C3847 ringtest_0.x4._25_ ringtest_0.x4._08_ 0.208467f
C3848 a_19842_32287# ui_in[1] 0.127717f
C3849 a_25393_5308# a_25351_5712# 7.84e-20
C3850 ringtest_0.x4._11_ ringtest_0.x4._05_ 0.023537f
C3851 a_24045_6654# a_24004_6128# 0.001715f
C3852 ringtest_0.x4.net6 a_21591_6128# 4.71e-21
C3853 a_21561_9116# a_21561_8830# 0.015931f
C3854 ringtest_0.counter7 ringtest_0.x4.counter[8] 0.068429f
C3855 ringtest_0.drv_out ringtest_0.x4.net7 6.87e-19
C3856 a_22223_5712# VDPWR 0.002609f
C3857 ringtest_0.x4._15_ a_25977_4220# 0.086673f
C3858 ringtest_0.x4._19_ a_24264_6788# 1.38e-19
C3859 muxtest_0.x1.x1.nSEL1 a_19794_32347# 4.08e-19
C3860 ringtest_0.drv_out ringtest_0.x4._17_ 1.68e-19
C3861 muxtest_0.x1.x1.nSEL0 a_19242_32347# 2.51e-19
C3862 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ui_in[3] 9.57e-20
C3863 ringtest_0.x4.net2 a_21675_9686# 0.008042f
C3864 ringtest_0.x4._23_ a_26201_4790# 0.029061f
C3865 muxtest_0.x1.x5.GN a_19842_32287# 2.26e-19
C3866 a_26201_4790# a_26367_4790# 0.970499f
C3867 a_24336_6544# ringtest_0.x4._15_ 1.53e-20
C3868 ringtest_0.x4.net3 a_22116_4902# 3.22e-20
C3869 ringtest_0.x3.x2.GP3 ua[1] 0.357364f
C3870 a_21675_4790# a_22390_4566# 4.63e-19
C3871 a_23381_4818# a_23381_4584# 0.012876f
C3872 ringtest_0.x4._16_ a_23837_5878# 0.061172f
C3873 ringtest_0.x4._04_ a_21587_5334# 3.27e-21
C3874 muxtest_0.x1.x3.GN1 ui_in[2] 0.054229f
C3875 m3_17032_8096# m3_17046_7066# 0.003741f
C3876 ringtest_0.x4._06_ a_24545_5878# 0.046896f
C3877 ringtest_0.x4.net9 ringtest_0.x4._07_ 0.03749f
C3878 ringtest_0.x4._22_ ringtest_0.x4._16_ 0.135659f
C3879 a_16755_12091# ringtest_0.x3.x2.GP3 5.21e-19
C3880 muxtest_0.x2.x2.GN1 ui_in[4] 0.312374f
C3881 ringtest_0.x4._23_ a_26555_5334# 0.014354f
C3882 a_22795_5334# a_22765_4478# 6.77e-20
C3883 muxtest_0.x2.x1.nSEL0 a_12473_23980# 0.001174f
C3884 ringtest_0.x4.clknet_1_0__leaf_clk a_21587_5334# 0.03291f
C3885 a_23467_4584# VDPWR 0.002731f
C3886 a_26555_5334# a_26367_4790# 1.41e-20
C3887 ringtest_0.x4._25_ VDPWR 0.22908f
C3888 a_21803_9508# VDPWR 0.005315f
C3889 ringtest_0.x4._11_ a_22350_5878# 0.003523f
C3890 a_24004_6128# a_24699_6200# 5.89e-19
C3891 ringtest_0.x4.net1 VDPWR 1.47718f
C3892 ringtest_0.x4.clknet_1_1__leaf_clk a_23770_5308# 0.048773f
C3893 muxtest_0.x1.x3.GP3 muxtest_0.R4R5 0.346864f
C3894 ringtest_0.x4.net4 a_22649_6244# 0.002624f
C3895 ringtest_0.x4.net7 ringtest_0.x4._07_ 0.047771f
C3896 muxtest_0.x1.x3.GP1 muxtest_0.R6R7 0.271251f
C3897 ringtest_0.x4.net3 ringtest_0.x4._04_ 5.28e-22
C3898 a_21852_8720# a_22052_8875# 0.080195f
C3899 a_21785_5878# a_22390_4566# 4.07e-21
C3900 a_21561_8830# ringtest_0.x4._01_ 8.93e-19
C3901 a_21845_8816# a_21981_8976# 0.136009f
C3902 a_26201_5340# a_26735_5334# 0.002698f
C3903 ringtest_0.x4._17_ ringtest_0.x4._07_ 3.97e-20
C3904 ringtest_0.x4._23_ a_27303_4246# 0.113094f
C3905 ringtest_0.x4.net7 a_25055_3867# 0.201574f
C3906 a_25977_4220# a_26173_4612# 0.00119f
C3907 ringtest_0.x4._11_ ringtest_0.x4._09_ 0.004259f
C3908 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net3 0.373279f
C3909 ringtest_0.x4._14_ a_21948_5156# 9.43e-20
C3910 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A 0.17253f
C3911 a_26808_4902# a_26721_4246# 5.71e-20
C3912 a_11845_23906# ui_in[3] 0.048888f
C3913 ringtest_0.x4._06_ a_24317_4942# 2.49e-19
C3914 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.308902f
C3915 ringtest_0.x4.net2 a_22052_8875# 3.35e-21
C3916 a_22052_9116# a_22399_9142# 0.037333f
C3917 ringtest_0.x4.net7 a_24264_6788# 0.001683f
C3918 ringtest_0.drv_out ringtest_0.x3.x2.GN3 0.243642f
C3919 a_24004_6128# a_23809_4790# 5.65e-20
C3920 a_24361_5340# a_24968_5308# 0.136009f
C3921 ringtest_0.x4.net1 a_21803_9508# 8.57e-19
C3922 ringtest_0.x4.net8 ringtest_0.x4.net10 1.02e-19
C3923 ringtest_0.x4.net9 a_26201_5340# 8.34e-19
C3924 a_25593_5156# a_26201_4790# 3.54e-19
C3925 a_23529_6422# ringtest_0.x4._19_ 0.082191f
C3926 ringtest_0.x4._18_ ringtest_0.x4.net6 0.081404f
C3927 a_25761_5058# ringtest_0.x4._09_ 0.001669f
C3928 ringtest_0.x4._21_ VDPWR 0.492491f
C3929 ringtest_0.x4.clknet_0_clk a_24527_5340# 5.94e-19
C3930 ringtest_0.x4.counter[2] VDPWR 0.494938f
C3931 ringtest_0.counter7 ringtest_0.x4.net6 6.88e-20
C3932 a_24045_6654# ringtest_0.x4._20_ 1.76e-19
C3933 ringtest_0.x4.net4 a_21587_5334# 1.97e-19
C3934 a_23809_4790# a_23963_4790# 0.004009f
C3935 ringtest_0.x4._15_ a_23899_5334# 0.046541f
C3936 a_16027_11759# ui_in[4] 0.03417f
C3937 muxtest_0.x1.x4.A a_12977_24040# 3.86e-20
C3938 ringtest_0.x4._24_ a_26367_5340# 0.035946f
C3939 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR 0.636314f
C3940 ringtest_0.x3.x1.nSEL1 a_16203_12091# 0.041068f
C3941 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN2 1.03e-20
C3942 a_21675_4790# a_22074_4790# 0.001351f
C3943 a_22116_4902# a_22457_5156# 9.73e-19
C3944 a_23381_4818# a_23809_4790# 0.00155f
C3945 a_21948_5156# a_22043_5156# 0.007724f
C3946 ringtest_0.counter3 ringtest_0.x4.counter[1] 0.099026f
C3947 ringtest_0.x4.net7 a_26201_5340# 8.61e-20
C3948 a_22265_5308# a_22164_4362# 6.81e-19
C3949 a_21425_9686# VDPWR 0.260172f
C3950 ringtest_0.x4._16_ a_22021_4220# 0.184103f
C3951 a_21951_5878# a_22392_5990# 0.111047f
C3952 a_23349_6422# VDPWR 0.252612f
C3953 a_12849_23648# VDPWR 0.180589f
C3954 ringtest_0.x4._23_ ringtest_0.x4.counter[8] 9.18e-19
C3955 a_21845_8816# a_22228_8598# 0.001632f
C3956 a_21852_8720# a_21803_8598# 4.04e-19
C3957 a_23879_6940# VDPWR 1.29479f
C3958 a_22052_8875# a_22399_8976# 0.037333f
C3959 a_21981_8976# a_22201_8964# 4.62e-19
C3960 ringtest_0.x4.net6 a_24763_6143# 0.027058f
C3961 ringtest_0.x4.net9 a_27233_5058# 0.001937f
C3962 ringtest_0.x3.x2.GP3 m3_17046_7066# 0.006132f
C3963 ringtest_0.x4._19_ ringtest_0.x4._06_ 7.42e-21
C3964 ringtest_0.x4.net7 ringtest_0.x4.counter[5] 0.002945f
C3965 ringtest_0.x4.net3 ringtest_0.x4.net4 0.0313f
C3966 muxtest_0.x2.x2.GN2 m3_13302_19985# 0.016745f
C3967 muxtest_0.x2.x2.GN4 ui_in[3] 0.218988f
C3968 a_25309_5334# VDPWR 0.004428f
C3969 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP1 0.062377f
C3970 ringtest_0.x4.counter[1] ua[2] 1.11e-19
C3971 ua[4] VGND 0.139799f
C3972 ua[5] VGND 0.141076f
C3973 ua[6] VGND 0.141964f
C3974 ua[7] VGND 0.146962f
C3975 ena VGND 0.072324f
C3976 clk VGND 0.044814f
C3977 rst_n VGND 0.044814f
C3978 ui_in[7] VGND 0.044814f
C3979 uio_in[0] VGND 0.047326f
C3980 uio_in[1] VGND 0.048926f
C3981 uio_in[2] VGND 0.044814f
C3982 uio_in[3] VGND 0.044814f
C3983 uio_in[4] VGND 0.044814f
C3984 uio_in[5] VGND 0.044814f
C3985 uio_in[6] VGND 0.044814f
C3986 uio_in[7] VGND 0.075838f
C3987 ua[1] VGND 28.486887f
C3988 ui_in[5] VGND 17.64489f
C3989 ui_in[6] VGND 24.291725f
C3990 ua[2] VGND 34.46381f
C3991 ua[0] VGND 51.530293f
C3992 ui_in[4] VGND 31.64427f
C3993 ui_in[3] VGND 32.74676f
C3994 ua[3] VGND 54.146942f
C3995 ui_in[2] VGND 26.529623f
C3996 ui_in[1] VGND 10.570298f
C3997 ui_in[0] VGND 10.700917f
C3998 VDPWR VGND 0.699931p
C3999 m3_17046_7066# VGND 0.075151f $ **FLOATING
C4000 m3_17032_8096# VGND 0.073094f $ **FLOATING
C4001 m3_17036_9140# VGND 0.148749f $ **FLOATING
C4002 m3_13316_18955# VGND 0.066786f $ **FLOATING
C4003 m3_13302_19985# VGND 0.064102f $ **FLOATING
C4004 m2_15612_11606# VGND 0.070212f $ **FLOATING
C4005 m2_11882_23495# VGND 0.065655f $ **FLOATING
C4006 m2_18699_31802# VGND 0.065655f $ **FLOATING
C4007 ringtest_0.x4.counter[8] VGND 0.58641f
C4008 ringtest_0.x4.counter[9] VGND 0.88818f
C4009 ringtest_0.x4.counter[6] VGND 0.659827f
C4010 ringtest_0.x4.counter[5] VGND 0.636589f
C4011 ringtest_0.x4.counter[4] VGND 0.791173f
C4012 ringtest_0.x4.counter[2] VGND 0.606277f
C4013 ringtest_0.x4.counter[1] VGND 0.591348f
C4014 ringtest_0.x4.counter[0] VGND 0.938564f
C4015 a_27815_3867# VGND 0.270206f
C4016 a_27489_3702# VGND 0.257101f
C4017 a_26895_3867# VGND 0.296141f
C4018 a_25975_3867# VGND 0.269288f
C4019 a_25055_3867# VGND 0.278393f
C4020 a_24135_3867# VGND 0.327843f
C4021 a_23399_3867# VGND 0.269041f
C4022 a_22295_3867# VGND 0.276333f
C4023 a_21375_3867# VGND 0.316834f
C4024 a_21007_3867# VGND 0.25238f
C4025 a_27659_4246# VGND 8.84e-19
C4026 a_27303_4246# VGND 0.004608f
C4027 a_26721_4246# VGND 0.01879f
C4028 a_27491_4566# VGND 0.00589f
C4029 a_26913_4566# VGND 0.010025f
C4030 a_26817_4566# VGND 0.006433f
C4031 a_26375_4612# VGND 0.001566f
C4032 a_26269_4612# VGND 0.003693f
C4033 a_26173_4612# VGND 0.003656f
C4034 a_25547_4612# VGND 0.003203f
C4035 a_25441_4612# VGND 0.005457f
C4036 a_25345_4612# VGND 0.005167f
C4037 a_22486_4246# VGND 0.001114f
C4038 a_23467_4584# VGND 0.004685f
C4039 a_22939_4584# VGND 0.007506f
C4040 a_22390_4566# VGND 0.183329f
C4041 a_27273_4220# VGND 0.369297f
C4042 a_26627_4246# VGND 0.344415f
C4043 a_25977_4220# VGND 0.261046f
C4044 a_25149_4220# VGND 0.294745f
C4045 a_23381_4584# VGND 0.255389f
C4046 a_22765_4478# VGND 0.284107f
C4047 a_22164_4362# VGND 0.207092f
C4048 a_22021_4220# VGND 0.20644f
C4049 a_27191_4790# VGND 0.004938f
C4050 ringtest_0.x4.net11 VGND 0.763831f
C4051 a_26766_4790# VGND 0.009249f
C4052 a_27149_5156# VGND 3.75e-19
C4053 a_25719_4790# VGND 0.004164f
C4054 a_26735_5156# VGND 0.002645f
C4055 a_26555_4790# VGND 0.063923f
C4056 a_27065_5156# VGND 0.26998f
C4057 a_27233_5058# VGND 0.379784f
C4058 a_26640_5156# VGND 0.228155f
C4059 a_26808_4902# VGND 0.258239f
C4060 a_26367_4790# VGND 0.335157f
C4061 ringtest_0.x4._09_ VGND 0.545207f
C4062 a_26201_4790# VGND 0.497148f
C4063 a_25294_4790# VGND 0.008691f
C4064 a_25677_5156# VGND 2.5e-19
C4065 a_24551_4790# VGND 7.68e-19
C4066 a_24479_4790# VGND 0.002515f
C4067 a_23963_4790# VGND 0.002664f
C4068 a_23891_4790# VGND 7.95e-19
C4069 a_25263_5156# VGND 7.5e-19
C4070 a_25083_4790# VGND 0.062716f
C4071 a_25593_5156# VGND 0.275541f
C4072 a_25761_5058# VGND 0.356576f
C4073 a_25168_5156# VGND 0.218254f
C4074 a_25336_4902# VGND 0.278138f
C4075 a_24895_4790# VGND 0.323857f
C4076 a_24729_4790# VGND 0.485385f
C4077 a_23467_4818# VGND 0.004685f
C4078 ringtest_0.x4._20_ VGND 0.296302f
C4079 a_22499_4790# VGND 0.004794f
C4080 ringtest_0.x4.net5 VGND 1.52232f
C4081 a_22074_4790# VGND 0.007478f
C4082 a_22457_5156# VGND 3.28e-19
C4083 a_21863_4790# VGND 0.069011f
C4084 a_24317_4942# VGND 0.233023f
C4085 a_23809_4790# VGND 0.25233f
C4086 a_23381_4818# VGND 0.250617f
C4087 a_22373_5156# VGND 0.29125f
C4088 a_22541_5058# VGND 0.405228f
C4089 a_21948_5156# VGND 0.210325f
C4090 a_22116_4902# VGND 0.255348f
C4091 a_21675_4790# VGND 0.417108f
C4092 ringtest_0.x4._03_ VGND 0.578555f
C4093 a_21509_4790# VGND 0.557931f
C4094 a_27149_5334# VGND 0.001033f
C4095 a_26735_5334# VGND 0.002645f
C4096 ringtest_0.x4.net10 VGND 1.58326f
C4097 a_27191_5712# VGND 0.005282f
C4098 a_25309_5334# VGND 0.002002f
C4099 a_26766_5712# VGND 0.010952f
C4100 a_26555_5334# VGND 0.070151f
C4101 a_25351_5712# VGND 0.005844f
C4102 a_23899_5334# VGND 0.014804f
C4103 a_23151_5334# VGND 0.001519f
C4104 a_22795_5334# VGND 0.026188f
C4105 a_22181_5334# VGND 4.07e-19
C4106 a_21767_5334# VGND 6.93e-19
C4107 a_24926_5712# VGND 0.006941f
C4108 a_24715_5334# VGND 0.060618f
C4109 a_23993_5654# VGND 0.006538f
C4110 a_23899_5654# VGND 0.008165f
C4111 a_22983_5654# VGND 0.007253f
C4112 a_22223_5712# VGND 0.004473f
C4113 a_21055_5334# VGND 4.64e-19
C4114 a_21798_5712# VGND 0.008558f
C4115 a_21587_5334# VGND 0.080622f
C4116 a_27065_5334# VGND 0.275172f
C4117 a_27233_5308# VGND 0.371259f
C4118 a_26640_5334# VGND 0.237292f
C4119 a_26808_5308# VGND 0.266551f
C4120 a_26367_5340# VGND 0.344626f
C4121 a_26201_5340# VGND 0.532322f
C4122 a_25225_5334# VGND 0.288597f
C4123 a_25393_5308# VGND 0.391747f
C4124 a_24800_5334# VGND 0.200127f
C4125 a_24968_5308# VGND 0.247676f
C4126 a_24527_5340# VGND 0.312142f
C4127 a_24361_5340# VGND 0.480598f
C4128 a_23770_5308# VGND 0.352433f
C4129 a_22765_5308# VGND 0.430766f
C4130 a_22097_5334# VGND 0.280567f
C4131 a_22265_5308# VGND 0.367396f
C4132 a_21672_5334# VGND 0.214988f
C4133 a_21840_5308# VGND 0.263107f
C4134 a_21399_5340# VGND 0.41156f
C4135 ringtest_0.x4._02_ VGND 0.384112f
C4136 a_21233_5340# VGND 0.551857f
C4137 ringtest_0.x4._14_ VGND 1.2474f
C4138 a_24986_5878# VGND 0.004249f
C4139 a_24545_5878# VGND 0.154917f
C4140 ringtest_0.x4._07_ VGND 0.467795f
C4141 a_23837_5878# VGND 0.204157f
C4142 a_22775_5878# VGND 0.00681f
C4143 ringtest_0.x4._16_ VGND 2.102403f
C4144 ringtest_0.x4._22_ VGND 1.57042f
C4145 a_24627_6200# VGND 8.25e-20
C4146 a_24763_6143# VGND 0.189132f
C4147 ringtest_0.x4.net9 VGND 1.9761f
C4148 ringtest_0.x4._06_ VGND 0.355082f
C4149 ringtest_0.x4._21_ VGND 0.491639f
C4150 a_23932_6128# VGND 9.9e-19
C4151 a_22350_5878# VGND 0.007439f
C4152 a_22733_6244# VGND 0.002478f
C4153 a_22319_6244# VGND 5.31e-19
C4154 a_22139_5878# VGND 0.062654f
C4155 a_25364_5878# VGND 2.07482f
C4156 a_24699_6200# VGND 0.166512f
C4157 a_24004_6128# VGND 0.208373f
C4158 a_24070_5852# VGND 0.228425f
C4159 ringtest_0.x4.net8 VGND 1.78641f
C4160 a_22649_6244# VGND 0.331871f
C4161 a_22817_6146# VGND 0.427232f
C4162 a_22224_6244# VGND 0.220057f
C4163 a_22392_5990# VGND 0.267836f
C4164 a_21951_5878# VGND 0.384412f
C4165 ringtest_0.x4._04_ VGND 0.647447f
C4166 a_21785_5878# VGND 0.561386f
C4167 a_21591_6128# VGND 0.005123f
C4168 ringtest_0.x4._13_ VGND 1.13412f
C4169 ringtest_0.x4.net4 VGND 1.31635f
C4170 ringtest_0.x4._08_ VGND 0.728198f
C4171 a_26839_6788# VGND 0.008414f
C4172 a_26201_6788# VGND 0.003851f
C4173 a_26095_6788# VGND 0.003674f
C4174 a_26007_6788# VGND 0.001688f
C4175 a_24287_6422# VGND 7.93e-19
C4176 a_24883_6800# VGND 0.060853f
C4177 a_24685_6788# VGND 0.006624f
C4178 a_24264_6788# VGND 0.005539f
C4179 a_23619_6788# VGND 0.005238f
C4180 ringtest_0.x4._25_ VGND 0.368024f
C4181 a_27169_6641# VGND 0.273817f
C4182 a_26749_6422# VGND 0.263282f
C4183 ringtest_0.x4._24_ VGND 0.69832f
C4184 a_26569_6422# VGND 0.271803f
C4185 ringtest_0.x4._23_ VGND 0.976575f
C4186 a_25925_6788# VGND 0.264561f
C4187 ringtest_0.x4._15_ VGND 3.54948f
C4188 ringtest_0.x4.net7 VGND 2.72071f
C4189 ringtest_0.x4.net6 VGND 3.218643f
C4190 ringtest_0.x4._19_ VGND 0.32708f
C4191 a_25421_6641# VGND 0.252712f
C4192 ringtest_0.x4.clknet_1_1__leaf_clk VGND 3.414301f
C4193 ringtest_0.x4._05_ VGND 0.318608f
C4194 a_24465_6800# VGND 0.241882f
C4195 a_24536_6699# VGND 0.198121f
C4196 a_24336_6544# VGND 0.303545f
C4197 a_24329_6640# VGND 0.46613f
C4198 a_24045_6654# VGND 0.281525f
C4199 a_23949_6654# VGND 0.378965f
C4200 a_23529_6422# VGND 0.234926f
C4201 ringtest_0.x4._18_ VGND 0.468402f
C4202 a_23349_6422# VGND 0.254342f
C4203 ringtest_0.x4._17_ VGND 0.622485f
C4204 ringtest_0.counter7 VGND 17.349024f
C4205 a_23879_6940# VGND 2.29287f
C4206 ringtest_0.x4.clknet_0_clk VGND 4.193551f
C4207 a_21395_6940# VGND 2.29289f
C4208 a_21939_8054# VGND 0.002457f
C4209 a_21867_8054# VGND 0.001303f
C4210 a_22695_8304# VGND 0.005104f
C4211 ringtest_0.counter3 VGND 14.338387f
C4212 ringtest_0.x4._11_ VGND 5.669866f
C4213 a_22245_8054# VGND 0.298451f
C4214 ringtest_0.x4._10_ VGND 0.339714f
C4215 a_21785_8054# VGND 0.252154f
C4216 a_21803_8598# VGND 6.89e-19
C4217 a_22399_8976# VGND 0.064411f
C4218 a_22201_8964# VGND 0.006624f
C4219 a_21049_8598# VGND 0.017559f
C4220 a_21780_8964# VGND 0.004183f
C4221 ringtest_0.x4._12_ VGND 1.2616f
C4222 a_21132_8918# VGND 0.004429f
C4223 ringtest_0.x4._01_ VGND 0.405148f
C4224 a_21981_8976# VGND 0.238144f
C4225 a_22052_8875# VGND 0.195482f
C4226 a_21852_8720# VGND 0.31379f
C4227 a_21845_8816# VGND 0.552106f
C4228 a_21561_8830# VGND 0.279727f
C4229 a_21465_8830# VGND 0.390267f
C4230 ringtest_0.x4.net3 VGND 2.298238f
C4231 a_22201_9142# VGND 0.007478f
C4232 a_21780_9142# VGND 0.004654f
C4233 ringtest_0.x4.clknet_1_0__leaf_clk VGND 4.010709f
C4234 a_22399_9142# VGND 0.069779f
C4235 a_21803_9508# VGND 6.84e-19
C4236 a_21981_9142# VGND 0.264386f
C4237 a_22052_9116# VGND 0.210923f
C4238 a_21845_9116# VGND 0.580201f
C4239 a_21852_9416# VGND 0.340144f
C4240 a_21561_9116# VGND 0.287469f
C4241 a_21465_9294# VGND 0.412387f
C4242 a_21675_9686# VGND 0.013142f
C4243 a_21507_9686# VGND 0.006974f
C4244 ringtest_0.x4._00_ VGND 0.757573f
C4245 a_21675_10006# VGND 0.006222f
C4246 a_21425_9686# VGND 0.393994f
C4247 ringtest_0.x4.net2 VGND 3.500251f
C4248 ringtest_0.x4.net1 VGND 1.81106f
C4249 a_22111_10993# VGND 0.293097f
C4250 ringtest_0.x3.x2.GP3 VGND 1.64575f
C4251 ringtest_0.x3.x2.GP2 VGND 5.54164f
C4252 ringtest_0.x3.x2.GP1 VGND 4.63625f
C4253 a_17405_12123# VGND 0.006782f
C4254 ringtest_0.x3.x2.GN4 VGND 3.79271f
C4255 a_16707_12151# VGND 0.007327f
C4256 ringtest_0.x3.x2.GN3 VGND 3.64172f
C4257 a_16155_12151# VGND 0.004704f
C4258 ringtest_0.x3.x2.GN2 VGND 3.91967f
C4259 a_15749_12123# VGND 0.006793f
C4260 ringtest_0.x3.x2.GN1 VGND 4.84443f
C4261 a_17231_12017# VGND 0.3167f
C4262 a_16755_12091# VGND 0.251626f
C4263 a_16579_11759# VGND 0.236732f
C4264 a_16203_12091# VGND 0.236633f
C4265 a_16027_11759# VGND 0.222621f
C4266 a_15575_12017# VGND 0.270062f
C4267 ringtest_0.x3.nselect2 VGND 0.455447f
C4268 ringtest_0.x3.x1.nSEL1 VGND 0.740163f
C4269 ringtest_0.x3.x1.nSEL0 VGND 0.685116f
C4270 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VGND 0.505562f
C4271 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VGND 0.498424f
C4272 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VGND 0.498285f
C4273 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VGND 0.499488f
C4274 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VGND 0.500758f
C4275 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VGND 0.50136f
C4276 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VGND 0.501617f
C4277 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VGND 0.52312f
C4278 ringtest_0.drv_out VGND 29.368195f
C4279 a_17377_14114# VGND 0.332619f
C4280 ringtest_0.ring_out VGND 16.289782f
C4281 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VGND 0.632983f
C4282 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VGND 0.508122f
C4283 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VGND 0.498331f
C4284 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VGND 0.498331f
C4285 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VGND 0.498339f
C4286 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VGND 0.498632f
C4287 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VGND 0.498682f
C4288 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VGND 0.498707f
C4289 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VGND 0.507755f
C4290 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VGND 0.971227f
C4291 muxtest_0.x2.x2.GP3 VGND 1.68554f
C4292 muxtest_0.x2.x2.GP2 VGND 5.5641f
C4293 muxtest_0.x2.x2.GP1 VGND 4.625069f
C4294 muxtest_0.R1R2 VGND 6.645505f
C4295 a_13675_24012# VGND 0.006439f
C4296 muxtest_0.x2.x2.GN4 VGND 3.796f
C4297 a_12977_24040# VGND 0.006801f
C4298 muxtest_0.x2.x2.GN3 VGND 3.65554f
C4299 a_12425_24040# VGND 0.004461f
C4300 muxtest_0.x2.x2.GN2 VGND 3.88834f
C4301 a_12019_24012# VGND 0.006505f
C4302 muxtest_0.x2.x2.GN1 VGND 4.79625f
C4303 a_13501_23906# VGND 0.306555f
C4304 a_13025_23980# VGND 0.249538f
C4305 a_12849_23648# VGND 0.232764f
C4306 a_12473_23980# VGND 0.23458f
C4307 a_12297_23648# VGND 0.220868f
C4308 a_11845_23906# VGND 0.267622f
C4309 muxtest_0.x2.nselect2 VGND 0.451665f
C4310 muxtest_0.x2.x1.nSEL1 VGND 0.686441f
C4311 muxtest_0.x2.x1.nSEL0 VGND 0.647345f
C4312 muxtest_0.R2R3 VGND 7.982832f
C4313 muxtest_0.R3R4 VGND 15.859409f
C4314 muxtest_0.R4R5 VGND 7.656276f
C4315 muxtest_0.R5R6 VGND 7.957228f
C4316 muxtest_0.R6R7 VGND 7.795067f
C4317 muxtest_0.R7R8 VGND 29.82938f
C4318 muxtest_0.x1.x5.A VGND 13.867701f
C4319 muxtest_0.x1.x4.A VGND 16.1317f
C4320 muxtest_0.x1.x3.GP3 VGND 3.18231f
C4321 muxtest_0.x1.x3.GP2 VGND 10.304811f
C4322 muxtest_0.x1.x3.GP1 VGND 10.781407f
C4323 a_20492_32319# VGND 0.006616f
C4324 muxtest_0.x1.x3.GN4 VGND 7.04004f
C4325 a_19794_32347# VGND 0.006984f
C4326 muxtest_0.x1.x3.GN3 VGND 6.77674f
C4327 a_19242_32347# VGND 0.004523f
C4328 muxtest_0.x1.x3.GN2 VGND 7.175951f
C4329 a_18836_32319# VGND 0.006515f
C4330 muxtest_0.x1.x3.GN1 VGND 8.91731f
C4331 a_20318_32213# VGND 0.311491f
C4332 a_19842_32287# VGND 0.24978f
C4333 a_19666_31955# VGND 0.233122f
C4334 a_19290_32287# VGND 0.234813f
C4335 a_19114_31955# VGND 0.221018f
C4336 a_18662_32213# VGND 0.267639f
C4337 muxtest_0.x1.x5.GN VGND 5.73587f
C4338 muxtest_0.x1.x1.nSEL1 VGND 0.683011f
C4339 muxtest_0.x1.x1.nSEL0 VGND 0.650421f
C4340 ui_in[5].t1 VGND 0.0025f
C4341 ui_in[5].t0 VGND 0.004008f
C4342 ui_in[5].n0 VGND 0.008077f
C4343 ui_in[5].n1 VGND 0.003407f
C4344 ui_in[5].n2 VGND 0.33124f
C4345 ui_in[5].n3 VGND 3.27797f
C4346 ui_in[6].t0 VGND 0.00254f
C4347 ui_in[6].t2 VGND 0.001497f
C4348 ui_in[6].n0 VGND 0.003424f
C4349 ui_in[6].t1 VGND 0.00254f
C4350 ui_in[6].t3 VGND 0.001497f
C4351 ui_in[6].n1 VGND 0.003424f
C4352 ui_in[6].n2 VGND 0.001687f
C4353 ui_in[6].n3 VGND 0.224459f
C4354 muxtest_0.R2R3.t0 VGND 0.626391f
C4355 muxtest_0.R2R3.t1 VGND 0.443113f
C4356 muxtest_0.R2R3.n0 VGND 3.43546f
C4357 muxtest_0.R2R3.t2 VGND 0.347912f
C4358 muxtest_0.R2R3.t3 VGND 0.638083f
C4359 muxtest_0.R2R3.n1 VGND 3.5698f
C4360 muxtest_0.R2R3.n2 VGND 0.568983f
C4361 muxtest_0.R2R3.n3 VGND 0.116677f
C4362 muxtest_0.R2R3.t4 VGND 0.210663f
C4363 muxtest_0.R2R3.t5 VGND 0.170342f
C4364 muxtest_0.R2R3.n4 VGND 3.38019f
C4365 muxtest_0.R4R5.t1 VGND 0.627578f
C4366 muxtest_0.R4R5.t2 VGND 0.443953f
C4367 muxtest_0.R4R5.n0 VGND 3.44197f
C4368 muxtest_0.R4R5.t4 VGND 0.348571f
C4369 muxtest_0.R4R5.t5 VGND 0.639293f
C4370 muxtest_0.R4R5.n1 VGND 3.57657f
C4371 muxtest_0.R4R5.n2 VGND 0.570061f
C4372 muxtest_0.R4R5.n3 VGND 0.119407f
C4373 muxtest_0.R4R5.t0 VGND 0.212944f
C4374 muxtest_0.R4R5.t3 VGND 0.170665f
C4375 muxtest_0.R4R5.n4 VGND 3.47489f
C4376 muxtest_0.x2.x2.x4.GP VGND 2.57727f
C4377 muxtest_0.x2.x1.gpo3 VGND 1.20603f
C4378 muxtest_0.x2.x2.GP4.t1 VGND 0.012374f
C4379 muxtest_0.x2.x2.GP4.t0 VGND 0.012374f
C4380 muxtest_0.x2.x2.GP4.n0 VGND 0.027184f
C4381 muxtest_0.x2.x1.x14.Y VGND 0.076955f
C4382 muxtest_0.x2.x2.GP4.n1 VGND 0.01052f
C4383 muxtest_0.x2.x2.GP4.t5 VGND 0.626223f
C4384 muxtest_0.x2.x2.GP4.t4 VGND 0.643686f
C4385 muxtest_0.x2.x2.GP4.n2 VGND 2.28835f
C4386 muxtest_0.x2.x2.GP4.n3 VGND 0.048401f
C4387 muxtest_0.x2.x2.GP4.t3 VGND 0.019037f
C4388 muxtest_0.x2.x2.GP4.t2 VGND 0.019037f
C4389 muxtest_0.x2.x2.GP4.n4 VGND 0.043773f
C4390 muxtest_0.x2.x2.GP4.n5 VGND 0.088779f
C4391 ringtest_0.x3.x2.GP2.t1 VGND 0.016198f
C4392 ringtest_0.x3.x2.GP2.t0 VGND 0.016198f
C4393 ringtest_0.x3.x2.GP2.n0 VGND 0.035585f
C4394 ringtest_0.x3.x2.GP2.n1 VGND 0.023f
C4395 ringtest_0.x3.x2.GP2.t5 VGND 0.819754f
C4396 ringtest_0.x3.x2.GP2.t4 VGND 0.842614f
C4397 ringtest_0.x3.x2.GP2.n2 VGND 2.98946f
C4398 ringtest_0.x3.x2.GP2.t3 VGND 0.02492f
C4399 ringtest_0.x3.x2.GP2.t2 VGND 0.02492f
C4400 ringtest_0.x3.x2.GP2.n3 VGND 0.051391f
C4401 ringtest_0.x3.x2.GP2.n4 VGND 0.120168f
C4402 ringtest_0.x3.x2.GP2.n5 VGND 0.027176f
C4403 ringtest_0.ring_out.t13 VGND 0.143976f
C4404 ringtest_0.ring_out.t12 VGND 0.066482f
C4405 ringtest_0.ring_out.n0 VGND 1.43742f
C4406 ringtest_0.ring_out.t2 VGND 0.011895f
C4407 ringtest_0.ring_out.t1 VGND 0.011895f
C4408 ringtest_0.ring_out.n1 VGND 0.036116f
C4409 ringtest_0.ring_out.t7 VGND 0.011895f
C4410 ringtest_0.ring_out.t8 VGND 0.011895f
C4411 ringtest_0.ring_out.n2 VGND 0.026441f
C4412 ringtest_0.ring_out.n3 VGND 0.119642f
C4413 ringtest_0.ring_out.t9 VGND 0.007732f
C4414 ringtest_0.ring_out.t0 VGND 0.007732f
C4415 ringtest_0.ring_out.n4 VGND 0.017154f
C4416 ringtest_0.ring_out.n5 VGND 0.032249f
C4417 ringtest_0.ring_out.n6 VGND 0.009203f
C4418 ringtest_0.ring_out.t14 VGND 0.010903f
C4419 ringtest_0.ring_out.t10 VGND 0.018503f
C4420 ringtest_0.ring_out.t15 VGND 0.010903f
C4421 ringtest_0.ring_out.t11 VGND 0.018503f
C4422 ringtest_0.ring_out.n7 VGND 0.031045f
C4423 ringtest_0.ring_out.n8 VGND 0.04596f
C4424 ringtest_0.ring_out.n9 VGND 0.181049f
C4425 ringtest_0.ring_out.n10 VGND 0.421446f
C4426 ringtest_0.ring_out.t5 VGND 0.673389f
C4427 ringtest_0.ring_out.t6 VGND 0.47636f
C4428 ringtest_0.ring_out.n11 VGND 3.69323f
C4429 ringtest_0.ring_out.t3 VGND 0.374016f
C4430 ringtest_0.ring_out.t4 VGND 0.685959f
C4431 ringtest_0.ring_out.n12 VGND 3.83764f
C4432 ringtest_0.ring_out.n13 VGND 0.611674f
C4433 ringtest_0.x3.x2.GP1.t1 VGND 0.012908f
C4434 ringtest_0.x3.x2.GP1.t0 VGND 0.012908f
C4435 ringtest_0.x3.x2.GP1.n0 VGND 0.028358f
C4436 ringtest_0.x3.x2.GP1.n1 VGND 0.018329f
C4437 ringtest_0.x3.x2.GP1.t4 VGND 0.653268f
C4438 ringtest_0.x3.x2.GP1.t5 VGND 0.671486f
C4439 ringtest_0.x3.x2.GP1.n2 VGND 2.37213f
C4440 ringtest_0.x3.x2.GP1.t3 VGND 0.019859f
C4441 ringtest_0.x3.x2.GP1.t2 VGND 0.019859f
C4442 ringtest_0.x3.x2.GP1.n3 VGND 0.04092f
C4443 ringtest_0.x3.x2.GP1.n4 VGND 0.100085f
C4444 ringtest_0.x3.x2.GP1.n5 VGND 0.021877f
C4445 ui_in[3].t3 VGND 0.007332f
C4446 ui_in[3].t12 VGND 0.00432f
C4447 ui_in[3].t18 VGND 0.007332f
C4448 ui_in[3].t2 VGND 0.00432f
C4449 ui_in[3].n0 VGND 0.012301f
C4450 ui_in[3].n1 VGND 0.018181f
C4451 ui_in[3].n2 VGND 0.005713f
C4452 ui_in[3].t6 VGND 0.003611f
C4453 ui_in[3].t10 VGND 0.005245f
C4454 ui_in[3].n3 VGND 0.012493f
C4455 ui_in[3].n4 VGND 0.006939f
C4456 ui_in[3].t9 VGND 0.004276f
C4457 ui_in[3].t19 VGND 0.006297f
C4458 ui_in[3].n5 VGND 0.014878f
C4459 ui_in[3].n6 VGND 0.00309f
C4460 ui_in[3].n7 VGND 0.001204f
C4461 ui_in[3].n8 VGND 0.110032f
C4462 ui_in[3].t17 VGND 0.007155f
C4463 ui_in[3].t15 VGND 0.003393f
C4464 ui_in[3].n9 VGND 0.025691f
C4465 ui_in[3].n10 VGND 0.004978f
C4466 ui_in[3].n11 VGND 0.126236f
C4467 ui_in[3].n12 VGND 0.082029f
C4468 ui_in[3].t8 VGND 0.007332f
C4469 ui_in[3].t16 VGND 0.00432f
C4470 ui_in[3].t5 VGND 0.007332f
C4471 ui_in[3].t13 VGND 0.00432f
C4472 ui_in[3].n13 VGND 0.012301f
C4473 ui_in[3].n14 VGND 0.018181f
C4474 ui_in[3].n15 VGND 0.005713f
C4475 ui_in[3].t7 VGND 0.003611f
C4476 ui_in[3].t11 VGND 0.005245f
C4477 ui_in[3].n16 VGND 0.012493f
C4478 ui_in[3].n17 VGND 0.006939f
C4479 ui_in[3].t14 VGND 0.004276f
C4480 ui_in[3].t0 VGND 0.006297f
C4481 ui_in[3].n18 VGND 0.014878f
C4482 ui_in[3].n19 VGND 0.00309f
C4483 ui_in[3].n20 VGND 0.001204f
C4484 ui_in[3].n21 VGND 0.110032f
C4485 ui_in[3].t4 VGND 0.007155f
C4486 ui_in[3].t1 VGND 0.003393f
C4487 ui_in[3].n22 VGND 0.025691f
C4488 ui_in[3].n23 VGND 0.004978f
C4489 ui_in[3].n24 VGND 0.126236f
C4490 ui_in[3].n25 VGND 0.082029f
C4491 ui_in[3].n26 VGND 10.0315f
C4492 muxtest_0.R7R8.t4 VGND 0.570638f
C4493 muxtest_0.R7R8.t3 VGND 0.403673f
C4494 muxtest_0.R7R8.n0 VGND 3.12968f
C4495 muxtest_0.R7R8.t0 VGND 0.316945f
C4496 muxtest_0.R7R8.t1 VGND 0.58129f
C4497 muxtest_0.R7R8.n1 VGND 3.25206f
C4498 muxtest_0.R7R8.n2 VGND 0.51834f
C4499 muxtest_0.R7R8.n3 VGND 0.107649f
C4500 muxtest_0.R7R8.t9 VGND 0.157299f
C4501 muxtest_0.R7R8.t2 VGND 0.858788f
C4502 muxtest_0.R7R8.n4 VGND 1.55412f
C4503 muxtest_0.R7R8.t5 VGND 0.570638f
C4504 muxtest_0.R7R8.t6 VGND 0.403673f
C4505 muxtest_0.R7R8.n5 VGND 3.12968f
C4506 muxtest_0.R7R8.t7 VGND 0.316945f
C4507 muxtest_0.R7R8.t8 VGND 0.58129f
C4508 muxtest_0.R7R8.n6 VGND 3.25206f
C4509 muxtest_0.R7R8.n7 VGND 0.51834f
C4510 muxtest_0.R7R8.n8 VGND 0.108573f
C4511 muxtest_0.R7R8.n9 VGND 9.50513f
C4512 ua[0].t5 VGND 0.319126f
C4513 ua[0].t6 VGND 0.225752f
C4514 ua[0].n0 VGND 1.75026f
C4515 ua[0].t8 VGND 0.17725f
C4516 ua[0].t7 VGND 0.325083f
C4517 ua[0].n1 VGND 1.8187f
C4518 ua[0].n2 VGND 0.289879f
C4519 ua[0].n3 VGND 0.060719f
C4520 ua[0].t4 VGND 0.086784f
C4521 ua[0].n4 VGND 1.50131f
C4522 ua[0].n5 VGND 11.5833f
C4523 ua[0].t3 VGND 0.319126f
C4524 ua[0].t2 VGND 0.225752f
C4525 ua[0].n6 VGND 1.75026f
C4526 ua[0].t1 VGND 0.17725f
C4527 ua[0].t0 VGND 0.325083f
C4528 ua[0].n7 VGND 1.8187f
C4529 ua[0].n8 VGND 0.289879f
C4530 ua[0].n9 VGND 0.059443f
C4531 muxtest_0.R6R7.t1 VGND 0.693927f
C4532 muxtest_0.R6R7.t0 VGND 0.490889f
C4533 muxtest_0.R6R7.n0 VGND 3.80587f
C4534 muxtest_0.R6R7.t2 VGND 0.385423f
C4535 muxtest_0.R6R7.t3 VGND 0.706881f
C4536 muxtest_0.R6R7.n1 VGND 3.95469f
C4537 muxtest_0.R6R7.n2 VGND 0.63033f
C4538 muxtest_0.R6R7.n3 VGND 0.129257f
C4539 muxtest_0.R6R7.t4 VGND 0.920517f
C4540 muxtest_0.R6R7.t5 VGND 0.188708f
C4541 muxtest_0.R6R7.n4 VGND 2.80582f
C4542 muxtest_0.R6R7.n5 VGND 1.24461f
C4543 muxtest_0.x2.x2.GP2.t0 VGND 0.016198f
C4544 muxtest_0.x2.x2.GP2.t1 VGND 0.016198f
C4545 muxtest_0.x2.x2.GP2.n0 VGND 0.035585f
C4546 muxtest_0.x2.x2.GP2.n1 VGND 0.023f
C4547 muxtest_0.x2.x2.GP2.t5 VGND 0.819754f
C4548 muxtest_0.x2.x2.GP2.t4 VGND 0.842614f
C4549 muxtest_0.x2.x2.GP2.n2 VGND 2.98946f
C4550 muxtest_0.x2.x2.GP2.t3 VGND 0.02492f
C4551 muxtest_0.x2.x2.GP2.t2 VGND 0.02492f
C4552 muxtest_0.x2.x2.GP2.n3 VGND 0.051391f
C4553 muxtest_0.x2.x2.GP2.n4 VGND 0.120168f
C4554 muxtest_0.x2.x2.GP2.n5 VGND 0.027176f
C4555 ringtest_0.x4._16_.t0 VGND 0.046376f
C4556 ringtest_0.x4._16_.n0 VGND 0.026397f
C4557 ringtest_0.x4._16_.t7 VGND 0.021164f
C4558 ringtest_0.x4._16_.t2 VGND 0.017507f
C4559 ringtest_0.x4._16_.n1 VGND 0.047954f
C4560 ringtest_0.x4._16_.n2 VGND 0.154756f
C4561 ringtest_0.x4._16_.t9 VGND 0.020065f
C4562 ringtest_0.x4._16_.t3 VGND 0.031953f
C4563 ringtest_0.x4._16_.n3 VGND 0.045672f
C4564 ringtest_0.x4._16_.n4 VGND 0.0375f
C4565 ringtest_0.x4._16_.t4 VGND 0.020065f
C4566 ringtest_0.x4._16_.t8 VGND 0.031953f
C4567 ringtest_0.x4._16_.n5 VGND 0.058943f
C4568 ringtest_0.x4._16_.n6 VGND 0.063595f
C4569 ringtest_0.x4._16_.n7 VGND 0.426096f
C4570 ringtest_0.x4._16_.t5 VGND 0.012893f
C4571 ringtest_0.x4._16_.t6 VGND 0.013824f
C4572 ringtest_0.x4._16_.n8 VGND 0.03796f
C4573 ringtest_0.x4._16_.n9 VGND 0.022428f
C4574 ringtest_0.x4._16_.n10 VGND 0.327394f
C4575 ringtest_0.x4._16_.n11 VGND 0.020414f
C4576 ringtest_0.x4._16_.t1 VGND 0.119992f
C4577 ringtest_0.x4._16_.n12 VGND 0.021583f
C4578 ringtest_0.x4._16_.n13 VGND 0.021194f
C4579 muxtest_0.R5R6.t0 VGND 0.695132f
C4580 muxtest_0.R5R6.t1 VGND 0.491742f
C4581 muxtest_0.R5R6.n0 VGND 3.81248f
C4582 muxtest_0.R5R6.t5 VGND 0.386092f
C4583 muxtest_0.R5R6.t4 VGND 0.708108f
C4584 muxtest_0.R5R6.n1 VGND 3.96156f
C4585 muxtest_0.R5R6.n2 VGND 0.631424f
C4586 muxtest_0.R5R6.n3 VGND 0.129973f
C4587 muxtest_0.R5R6.t3 VGND 0.191095f
C4588 muxtest_0.R5R6.t2 VGND 1.13104f
C4589 muxtest_0.R5R6.n4 VGND 2.8297f
C4590 muxtest_0.x1.x3.GP2.t0 VGND 0.018287f
C4591 muxtest_0.x1.x3.GP2.t1 VGND 0.018287f
C4592 muxtest_0.x1.x3.GP2.n0 VGND 0.040174f
C4593 muxtest_0.x1.x3.GP2.n1 VGND 0.025967f
C4594 muxtest_0.x1.x3.GP2.t6 VGND 0.925483f
C4595 muxtest_0.x1.x3.GP2.t7 VGND 0.951291f
C4596 muxtest_0.x1.x3.GP2.n2 VGND 3.37503f
C4597 muxtest_0.x1.x3.GP2.t5 VGND 0.925483f
C4598 muxtest_0.x1.x3.GP2.t4 VGND 0.951291f
C4599 muxtest_0.x1.x3.GP2.n3 VGND 3.37503f
C4600 muxtest_0.x1.x3.GP2.n4 VGND 1.97357f
C4601 muxtest_0.x1.x3.GP2.t2 VGND 0.028134f
C4602 muxtest_0.x1.x3.GP2.t3 VGND 0.028134f
C4603 muxtest_0.x1.x3.GP2.n5 VGND 0.058019f
C4604 muxtest_0.x1.x3.GP2.n6 VGND 0.132927f
C4605 muxtest_0.x1.x3.GP2.n7 VGND 0.030681f
C4606 ringtest_0.counter3.t3 VGND 0.033829f
C4607 ringtest_0.counter3.n0 VGND 0.005886f
C4608 ringtest_0.counter3.t2 VGND 0.023398f
C4609 ringtest_0.counter3.n1 VGND 0.028682f
C4610 ringtest_0.counter3.n2 VGND 0.036901f
C4611 ringtest_0.counter3.n3 VGND 0.371589f
C4612 ringtest_0.counter3.t1 VGND 0.740343f
C4613 ringtest_0.counter3.t0 VGND 0.523724f
C4614 ringtest_0.counter3.n4 VGND 4.06044f
C4615 ringtest_0.counter3.t4 VGND 0.410954f
C4616 ringtest_0.counter3.t5 VGND 0.761665f
C4617 ringtest_0.counter3.n5 VGND 4.29752f
C4618 ringtest_0.counter3.n6 VGND 0.672491f
C4619 ringtest_0.x4.clknet_1_0__leaf_clk.t38 VGND 0.022262f
C4620 ringtest_0.x4.clknet_1_0__leaf_clk.t41 VGND 0.014894f
C4621 ringtest_0.x4.clknet_1_0__leaf_clk.n0 VGND 0.04068f
C4622 ringtest_0.x4.clknet_1_0__leaf_clk.n1 VGND 0.107083f
C4623 ringtest_0.x4.clknet_1_0__leaf_clk.t37 VGND 0.014894f
C4624 ringtest_0.x4.clknet_1_0__leaf_clk.t32 VGND 0.022262f
C4625 ringtest_0.x4.clknet_1_0__leaf_clk.n2 VGND 0.041145f
C4626 ringtest_0.x4.clknet_1_0__leaf_clk.n3 VGND 0.437523f
C4627 ringtest_0.x4.clknet_1_0__leaf_clk.t30 VGND 0.014222f
C4628 ringtest_0.x4.clknet_1_0__leaf_clk.t16 VGND 0.014222f
C4629 ringtest_0.x4.clknet_1_0__leaf_clk.n4 VGND 0.029978f
C4630 ringtest_0.x4.clknet_1_0__leaf_clk.t27 VGND 0.014222f
C4631 ringtest_0.x4.clknet_1_0__leaf_clk.t29 VGND 0.014222f
C4632 ringtest_0.x4.clknet_1_0__leaf_clk.n5 VGND 0.029589f
C4633 ringtest_0.x4.clknet_1_0__leaf_clk.t8 VGND 0.005973f
C4634 ringtest_0.x4.clknet_1_0__leaf_clk.t11 VGND 0.005973f
C4635 ringtest_0.x4.clknet_1_0__leaf_clk.n6 VGND 0.021211f
C4636 ringtest_0.x4.clknet_1_0__leaf_clk.t13 VGND 0.005973f
C4637 ringtest_0.x4.clknet_1_0__leaf_clk.t15 VGND 0.005973f
C4638 ringtest_0.x4.clknet_1_0__leaf_clk.n7 VGND 0.013636f
C4639 ringtest_0.x4.clknet_1_0__leaf_clk.n8 VGND 0.086164f
C4640 ringtest_0.x4.clknet_1_0__leaf_clk.t10 VGND 0.005973f
C4641 ringtest_0.x4.clknet_1_0__leaf_clk.t12 VGND 0.005973f
C4642 ringtest_0.x4.clknet_1_0__leaf_clk.n9 VGND 0.013636f
C4643 ringtest_0.x4.clknet_1_0__leaf_clk.n10 VGND 0.051791f
C4644 ringtest_0.x4.clknet_1_0__leaf_clk.t14 VGND 0.005973f
C4645 ringtest_0.x4.clknet_1_0__leaf_clk.t9 VGND 0.005973f
C4646 ringtest_0.x4.clknet_1_0__leaf_clk.n11 VGND 0.013644f
C4647 ringtest_0.x4.clknet_1_0__leaf_clk.n12 VGND 0.053424f
C4648 ringtest_0.x4.clknet_1_0__leaf_clk.t1 VGND 0.005973f
C4649 ringtest_0.x4.clknet_1_0__leaf_clk.t4 VGND 0.005973f
C4650 ringtest_0.x4.clknet_1_0__leaf_clk.n13 VGND 0.013636f
C4651 ringtest_0.x4.clknet_1_0__leaf_clk.n14 VGND 0.051791f
C4652 ringtest_0.x4.clknet_1_0__leaf_clk.t6 VGND 0.005973f
C4653 ringtest_0.x4.clknet_1_0__leaf_clk.t7 VGND 0.005973f
C4654 ringtest_0.x4.clknet_1_0__leaf_clk.n15 VGND 0.013636f
C4655 ringtest_0.x4.clknet_1_0__leaf_clk.n16 VGND 0.05205f
C4656 ringtest_0.x4.clknet_1_0__leaf_clk.t3 VGND 0.005973f
C4657 ringtest_0.x4.clknet_1_0__leaf_clk.t5 VGND 0.005973f
C4658 ringtest_0.x4.clknet_1_0__leaf_clk.n17 VGND 0.013636f
C4659 ringtest_0.x4.clknet_1_0__leaf_clk.n18 VGND 0.04471f
C4660 ringtest_0.x4.clknet_1_0__leaf_clk.t0 VGND 0.005973f
C4661 ringtest_0.x4.clknet_1_0__leaf_clk.t2 VGND 0.005973f
C4662 ringtest_0.x4.clknet_1_0__leaf_clk.n19 VGND 0.013163f
C4663 ringtest_0.x4.clknet_1_0__leaf_clk.n20 VGND 0.043256f
C4664 ringtest_0.x4.clknet_1_0__leaf_clk.n21 VGND 0.09308f
C4665 ringtest_0.x4.clknet_1_0__leaf_clk.n22 VGND 0.067594f
C4666 ringtest_0.x4.clknet_1_0__leaf_clk.t19 VGND 0.014222f
C4667 ringtest_0.x4.clknet_1_0__leaf_clk.t22 VGND 0.014222f
C4668 ringtest_0.x4.clknet_1_0__leaf_clk.n23 VGND 0.036128f
C4669 ringtest_0.x4.clknet_1_0__leaf_clk.t24 VGND 0.014222f
C4670 ringtest_0.x4.clknet_1_0__leaf_clk.t26 VGND 0.014222f
C4671 ringtest_0.x4.clknet_1_0__leaf_clk.n24 VGND 0.029978f
C4672 ringtest_0.x4.clknet_1_0__leaf_clk.n25 VGND 0.136621f
C4673 ringtest_0.x4.clknet_1_0__leaf_clk.t21 VGND 0.014222f
C4674 ringtest_0.x4.clknet_1_0__leaf_clk.t23 VGND 0.014222f
C4675 ringtest_0.x4.clknet_1_0__leaf_clk.n26 VGND 0.029978f
C4676 ringtest_0.x4.clknet_1_0__leaf_clk.n27 VGND 0.0787f
C4677 ringtest_0.x4.clknet_1_0__leaf_clk.t25 VGND 0.014222f
C4678 ringtest_0.x4.clknet_1_0__leaf_clk.t20 VGND 0.014222f
C4679 ringtest_0.x4.clknet_1_0__leaf_clk.n28 VGND 0.029978f
C4680 ringtest_0.x4.clknet_1_0__leaf_clk.n29 VGND 0.078334f
C4681 ringtest_0.x4.clknet_1_0__leaf_clk.t28 VGND 0.014222f
C4682 ringtest_0.x4.clknet_1_0__leaf_clk.t31 VGND 0.014222f
C4683 ringtest_0.x4.clknet_1_0__leaf_clk.n30 VGND 0.029978f
C4684 ringtest_0.x4.clknet_1_0__leaf_clk.n31 VGND 0.078334f
C4685 ringtest_0.x4.clknet_1_0__leaf_clk.n32 VGND 0.04742f
C4686 ringtest_0.x4.clknet_1_0__leaf_clk.t17 VGND 0.014222f
C4687 ringtest_0.x4.clknet_1_0__leaf_clk.t18 VGND 0.014222f
C4688 ringtest_0.x4.clknet_1_0__leaf_clk.n33 VGND 0.028445f
C4689 ringtest_0.x4.clknet_1_0__leaf_clk.n34 VGND 0.022411f
C4690 ringtest_0.x4.clknet_1_0__leaf_clk.n35 VGND 0.171468f
C4691 ringtest_0.x4.clknet_1_0__leaf_clk.t39 VGND 0.014894f
C4692 ringtest_0.x4.clknet_1_0__leaf_clk.t36 VGND 0.022262f
C4693 ringtest_0.x4.clknet_1_0__leaf_clk.n36 VGND 0.040782f
C4694 ringtest_0.x4.clknet_1_0__leaf_clk.n37 VGND 0.024896f
C4695 ringtest_0.x4.clknet_1_0__leaf_clk.t33 VGND 0.022262f
C4696 ringtest_0.x4.clknet_1_0__leaf_clk.t40 VGND 0.014894f
C4697 ringtest_0.x4.clknet_1_0__leaf_clk.n38 VGND 0.040732f
C4698 ringtest_0.x4.clknet_1_0__leaf_clk.n39 VGND 0.086433f
C4699 ringtest_0.x4.clknet_1_0__leaf_clk.n40 VGND 0.225449f
C4700 ringtest_0.x4.clknet_1_0__leaf_clk.t35 VGND 0.022262f
C4701 ringtest_0.x4.clknet_1_0__leaf_clk.t34 VGND 0.014894f
C4702 ringtest_0.x4.clknet_1_0__leaf_clk.n41 VGND 0.04068f
C4703 ringtest_0.x4.clknet_1_0__leaf_clk.n42 VGND 0.027948f
C4704 ringtest_0.x4.clknet_1_0__leaf_clk.n43 VGND 0.145937f
C4705 ua[1].t0 VGND 0.322568f
C4706 ua[1].n0 VGND 0.401178f
C4707 ua[1].t5 VGND 0.24977f
C4708 ua[1].t1 VGND 0.33145f
C4709 ua[1].n1 VGND 1.6726f
C4710 ua[1].n2 VGND 0.565936f
C4711 ua[1].t6 VGND 0.244855f
C4712 ua[1].n3 VGND 0.365612f
C4713 ua[1].n4 VGND 0.509787f
C4714 ua[1].t4 VGND 0.322568f
C4715 ua[1].n5 VGND 0.401178f
C4716 ua[1].t8 VGND 0.24977f
C4717 ua[1].t12 VGND 0.33145f
C4718 ua[1].n6 VGND 1.6726f
C4719 ua[1].n7 VGND 0.565936f
C4720 ua[1].t9 VGND 0.244855f
C4721 ua[1].n8 VGND 0.365612f
C4722 ua[1].n9 VGND 0.495416f
C4723 ua[1].n10 VGND 0.270615f
C4724 ua[1].t13 VGND 0.322568f
C4725 ua[1].n11 VGND 0.401178f
C4726 ua[1].t11 VGND 0.24977f
C4727 ua[1].t7 VGND 0.33145f
C4728 ua[1].n12 VGND 1.6726f
C4729 ua[1].n13 VGND 0.565936f
C4730 ua[1].t10 VGND 0.244855f
C4731 ua[1].n14 VGND 0.365612f
C4732 ua[1].n15 VGND 0.495991f
C4733 ua[1].n16 VGND 0.268745f
C4734 ua[1].n17 VGND 0.801201f
C4735 ua[1].t3 VGND 0.322568f
C4736 ua[1].n18 VGND 0.401178f
C4737 ua[1].t15 VGND 0.24977f
C4738 ua[1].t2 VGND 0.33145f
C4739 ua[1].n19 VGND 1.6726f
C4740 ua[1].n20 VGND 0.565936f
C4741 ua[1].t14 VGND 0.244855f
C4742 ua[1].n21 VGND 0.365612f
C4743 ua[1].n22 VGND 0.500412f
C4744 ua[1].n23 VGND 0.264233f
C4745 ua[1].n24 VGND 0.382993f
C4746 ua[1].n25 VGND 7.827061f
C4747 ringtest_0.counter7.t5 VGND 0.031678f
C4748 ringtest_0.counter7.n0 VGND 0.005512f
C4749 ringtest_0.counter7.t4 VGND 0.021911f
C4750 ringtest_0.counter7.n1 VGND 0.026858f
C4751 ringtest_0.counter7.n2 VGND 0.039564f
C4752 ringtest_0.counter7.n3 VGND 0.38767f
C4753 ringtest_0.counter7.t0 VGND 0.693272f
C4754 ringtest_0.counter7.t1 VGND 0.490426f
C4755 ringtest_0.counter7.n4 VGND 3.80227f
C4756 ringtest_0.counter7.t2 VGND 0.385059f
C4757 ringtest_0.counter7.t3 VGND 0.706213f
C4758 ringtest_0.counter7.n5 VGND 3.95096f
C4759 ringtest_0.counter7.n6 VGND 0.629734f
C4760 ringtest_0.x3.x2.x4.GP VGND 2.5438f
C4761 ringtest_0.x3.x1.gpo3 VGND 1.19037f
C4762 ringtest_0.x3.x2.GP4.t1 VGND 0.012213f
C4763 ringtest_0.x3.x2.GP4.t0 VGND 0.012213f
C4764 ringtest_0.x3.x2.GP4.n0 VGND 0.026831f
C4765 ringtest_0.x3.x1.x14.Y VGND 0.075955f
C4766 ringtest_0.x3.x2.GP4.n1 VGND 0.010383f
C4767 ringtest_0.x3.x2.GP4.t4 VGND 0.618091f
C4768 ringtest_0.x3.x2.GP4.t5 VGND 0.635327f
C4769 ringtest_0.x3.x2.GP4.n2 VGND 2.25863f
C4770 ringtest_0.x3.x2.GP4.n3 VGND 0.047772f
C4771 ringtest_0.x3.x2.GP4.t3 VGND 0.01879f
C4772 ringtest_0.x3.x2.GP4.t2 VGND 0.01879f
C4773 ringtest_0.x3.x2.GP4.n4 VGND 0.043205f
C4774 ringtest_0.x3.x2.GP4.n5 VGND 0.087626f
C4775 ui_in[2].t7 VGND 0.320078f
C4776 ui_in[2].t1 VGND 0.312355f
C4777 ui_in[2].n0 VGND 1.40142f
C4778 ui_in[2].n1 VGND 0.46615f
C4779 ui_in[2].t6 VGND 0.375993f
C4780 ui_in[2].t0 VGND 0.386477f
C4781 ui_in[2].n2 VGND 1.40813f
C4782 ui_in[2].n3 VGND 0.945344f
C4783 ui_in[2].n4 VGND 2.4766f
C4784 ui_in[2].t3 VGND 0.01778f
C4785 ui_in[2].t5 VGND 0.010478f
C4786 ui_in[2].t2 VGND 0.01778f
C4787 ui_in[2].t4 VGND 0.010478f
C4788 ui_in[2].n5 VGND 0.029832f
C4789 ui_in[2].n6 VGND 0.044104f
C4790 ui_in[2].n7 VGND 0.043804f
C4791 ui_in[2].n8 VGND 0.708274f
C4792 ringtest_0.x4.net3.t1 VGND 0.067779f
C4793 ringtest_0.x4.net3.t2 VGND 0.019614f
C4794 ringtest_0.x4.net3.t7 VGND 0.031428f
C4795 ringtest_0.x4.net3.n0 VGND 0.061838f
C4796 ringtest_0.x4.net3.n1 VGND 0.008618f
C4797 ringtest_0.x4.net3.n2 VGND 0.005246f
C4798 ringtest_0.x4.net3.t6 VGND 0.029572f
C4799 ringtest_0.x4.net3.t5 VGND 0.018443f
C4800 ringtest_0.x4.net3.n3 VGND 0.059457f
C4801 ringtest_0.x4.net3.n4 VGND 0.019056f
C4802 ringtest_0.x4.net3.t4 VGND 0.030361f
C4803 ringtest_0.x4.net3.t3 VGND 0.055573f
C4804 ringtest_0.x4.net3.n5 VGND 0.744487f
C4805 ringtest_0.x4.net3.n6 VGND 0.124162f
C4806 ringtest_0.x4.net3.n7 VGND 0.092279f
C4807 ringtest_0.x4.net3.t0 VGND 0.037792f
C4808 ringtest_0.x4.net3.n8 VGND 0.040884f
C4809 ringtest_0.drv_out.t19 VGND 0.591341f
C4810 ringtest_0.drv_out.t0 VGND 0.418319f
C4811 ringtest_0.drv_out.n0 VGND 3.24323f
C4812 ringtest_0.drv_out.t2 VGND 0.328444f
C4813 ringtest_0.drv_out.t1 VGND 0.602379f
C4814 ringtest_0.drv_out.n1 VGND 3.37005f
C4815 ringtest_0.drv_out.n2 VGND 0.537145f
C4816 ringtest_0.drv_out.n3 VGND 0.110148f
C4817 ringtest_0.drv_out.t21 VGND 0.015262f
C4818 ringtest_0.drv_out.t25 VGND 0.007138f
C4819 ringtest_0.drv_out.t20 VGND 0.015262f
C4820 ringtest_0.drv_out.t24 VGND 0.007138f
C4821 ringtest_0.drv_out.t23 VGND 0.015262f
C4822 ringtest_0.drv_out.t27 VGND 0.007138f
C4823 ringtest_0.drv_out.t22 VGND 0.015262f
C4824 ringtest_0.drv_out.t26 VGND 0.007138f
C4825 ringtest_0.drv_out.n4 VGND 0.034841f
C4826 ringtest_0.drv_out.n5 VGND 0.04589f
C4827 ringtest_0.drv_out.n6 VGND 0.04589f
C4828 ringtest_0.drv_out.n7 VGND 0.055736f
C4829 ringtest_0.drv_out.n8 VGND 0.015444f
C4830 ringtest_0.drv_out.n9 VGND 0.346765f
C4831 ringtest_0.drv_out.n10 VGND 0.764086f
C4832 ringtest_0.drv_out.n11 VGND 5.53733f
C4833 ringtest_0.drv_out.t17 VGND 0.1149f
C4834 ringtest_0.drv_out.t12 VGND 0.1149f
C4835 ringtest_0.drv_out.n12 VGND 0.273611f
C4836 ringtest_0.drv_out.t14 VGND 0.1149f
C4837 ringtest_0.drv_out.t16 VGND 0.1149f
C4838 ringtest_0.drv_out.n13 VGND 0.273611f
C4839 ringtest_0.drv_out.t13 VGND 0.1149f
C4840 ringtest_0.drv_out.t15 VGND 0.1149f
C4841 ringtest_0.drv_out.n14 VGND 0.273611f
C4842 ringtest_0.drv_out.t18 VGND 0.1149f
C4843 ringtest_0.drv_out.t11 VGND 0.1149f
C4844 ringtest_0.drv_out.n15 VGND 0.273611f
C4845 ringtest_0.drv_out.n16 VGND 4.32f
C4846 ringtest_0.drv_out.t6 VGND 0.0383f
C4847 ringtest_0.drv_out.t8 VGND 0.0383f
C4848 ringtest_0.drv_out.n17 VGND 0.093269f
C4849 ringtest_0.drv_out.t7 VGND 0.0383f
C4850 ringtest_0.drv_out.t9 VGND 0.0383f
C4851 ringtest_0.drv_out.n18 VGND 0.093269f
C4852 ringtest_0.drv_out.t3 VGND 0.0383f
C4853 ringtest_0.drv_out.t4 VGND 0.0383f
C4854 ringtest_0.drv_out.n19 VGND 0.093269f
C4855 ringtest_0.drv_out.t10 VGND 0.0383f
C4856 ringtest_0.drv_out.t5 VGND 0.0383f
C4857 ringtest_0.drv_out.n20 VGND 0.093269f
C4858 ringtest_0.drv_out.n21 VGND 1.9949f
C4859 ringtest_0.drv_out.n22 VGND 2.14485f
C4860 a_19289_13081.t12 VGND 0.136375f
C4861 a_19289_13081.t2 VGND 0.13635f
C4862 a_19289_13081.n0 VGND 0.157675f
C4863 a_19289_13081.t13 VGND 0.13635f
C4864 a_19289_13081.n1 VGND 0.086028f
C4865 a_19289_13081.t7 VGND 0.13635f
C4866 a_19289_13081.n2 VGND 0.160734f
C4867 a_19289_13081.t4 VGND 0.049796f
C4868 a_19289_13081.t15 VGND 0.049764f
C4869 a_19289_13081.n3 VGND 0.09498f
C4870 a_19289_13081.t5 VGND 0.049764f
C4871 a_19289_13081.n4 VGND 0.055718f
C4872 a_19289_13081.t11 VGND 0.049764f
C4873 a_19289_13081.n5 VGND 0.086134f
C4874 a_19289_13081.t0 VGND 0.098833f
C4875 a_19289_13081.n6 VGND 0.831842f
C4876 a_19289_13081.t6 VGND 0.049771f
C4877 a_19289_13081.t9 VGND 0.13635f
C4878 a_19289_13081.n7 VGND 0.503671f
C4879 a_19289_13081.t16 VGND 0.049764f
C4880 a_19289_13081.n8 VGND 0.212248f
C4881 a_19289_13081.t17 VGND 0.13635f
C4882 a_19289_13081.n9 VGND 0.242932f
C4883 a_19289_13081.t8 VGND 0.049764f
C4884 a_19289_13081.n10 VGND 0.212248f
C4885 a_19289_13081.t10 VGND 0.13635f
C4886 a_19289_13081.n11 VGND 0.242932f
C4887 a_19289_13081.t3 VGND 0.049764f
C4888 a_19289_13081.n12 VGND 0.212248f
C4889 a_19289_13081.t14 VGND 0.13635f
C4890 a_19289_13081.n13 VGND 0.494157f
C4891 a_19289_13081.n14 VGND 1.47337f
C4892 a_19289_13081.n15 VGND 2.33573f
C4893 a_19289_13081.t1 VGND 0.309542f
C4894 muxtest_0.R1R2.t1 VGND 0.625209f
C4895 muxtest_0.R1R2.t0 VGND 0.442278f
C4896 muxtest_0.R1R2.n0 VGND 3.42898f
C4897 muxtest_0.R1R2.t4 VGND 0.347255f
C4898 muxtest_0.R1R2.t5 VGND 0.63688f
C4899 muxtest_0.R1R2.n1 VGND 3.56307f
C4900 muxtest_0.R1R2.n2 VGND 0.56791f
C4901 muxtest_0.R1R2.n3 VGND 0.116899f
C4902 muxtest_0.R1R2.t3 VGND 0.207548f
C4903 muxtest_0.R1R2.t2 VGND 0.169702f
C4904 muxtest_0.R1R2.n4 VGND 3.13805f
C4905 muxtest_0.R1R2.n5 VGND 1.09366f
C4906 ui_in[4].t4 VGND 0.008207f
C4907 ui_in[4].t10 VGND 0.004836f
C4908 ui_in[4].t6 VGND 0.008207f
C4909 ui_in[4].t16 VGND 0.004836f
C4910 ui_in[4].n0 VGND 0.01377f
C4911 ui_in[4].n1 VGND 0.020344f
C4912 ui_in[4].n2 VGND 0.012412f
C4913 ui_in[4].t19 VGND 0.008009f
C4914 ui_in[4].t13 VGND 0.003797f
C4915 ui_in[4].n3 VGND 0.028758f
C4916 ui_in[4].n4 VGND 0.005576f
C4917 ui_in[4].n5 VGND 0.00476f
C4918 ui_in[4].t7 VGND 0.003976f
C4919 ui_in[4].t12 VGND 0.005786f
C4920 ui_in[4].n6 VGND 0.016813f
C4921 ui_in[4].n7 VGND 0.003873f
C4922 ui_in[4].n8 VGND 0.027736f
C4923 ui_in[4].n9 VGND 0.100485f
C4924 ui_in[4].t5 VGND 0.004786f
C4925 ui_in[4].t0 VGND 0.007049f
C4926 ui_in[4].n10 VGND 0.016654f
C4927 ui_in[4].n11 VGND 0.002169f
C4928 ui_in[4].n12 VGND 0.024508f
C4929 ui_in[4].n13 VGND 0.115979f
C4930 ui_in[4].n14 VGND 0.151491f
C4931 ui_in[4].n15 VGND 0.034981f
C4932 ui_in[4].t15 VGND 0.008207f
C4933 ui_in[4].t2 VGND 0.004836f
C4934 ui_in[4].t9 VGND 0.008207f
C4935 ui_in[4].t18 VGND 0.004836f
C4936 ui_in[4].n16 VGND 0.01377f
C4937 ui_in[4].n17 VGND 0.020344f
C4938 ui_in[4].n18 VGND 0.012412f
C4939 ui_in[4].t1 VGND 0.008009f
C4940 ui_in[4].t17 VGND 0.003797f
C4941 ui_in[4].n19 VGND 0.028758f
C4942 ui_in[4].n20 VGND 0.005576f
C4943 ui_in[4].n21 VGND 0.00476f
C4944 ui_in[4].t11 VGND 0.003976f
C4945 ui_in[4].t14 VGND 0.005786f
C4946 ui_in[4].n22 VGND 0.016813f
C4947 ui_in[4].n23 VGND 0.003873f
C4948 ui_in[4].n24 VGND 0.027736f
C4949 ui_in[4].n25 VGND 0.100485f
C4950 ui_in[4].t8 VGND 0.004786f
C4951 ui_in[4].t3 VGND 0.007049f
C4952 ui_in[4].n26 VGND 0.016654f
C4953 ui_in[4].n27 VGND 0.002169f
C4954 ui_in[4].n28 VGND 0.024508f
C4955 ui_in[4].n29 VGND 0.115979f
C4956 ui_in[4].n30 VGND 0.151491f
C4957 ui_in[4].n31 VGND 12.0273f
C4958 muxtest_0.R3R4.t6 VGND 0.65338f
C4959 muxtest_0.R3R4.t5 VGND 0.462206f
C4960 muxtest_0.R3R4.n0 VGND 3.58348f
C4961 muxtest_0.R3R4.t1 VGND 0.362902f
C4962 muxtest_0.R3R4.t0 VGND 0.665576f
C4963 muxtest_0.R3R4.n1 VGND 3.72361f
C4964 muxtest_0.R3R4.n2 VGND 0.593498f
C4965 muxtest_0.R3R4.n3 VGND 0.123258f
C4966 muxtest_0.R3R4.t4 VGND 1.02738f
C4967 muxtest_0.R3R4.t7 VGND 0.177328f
C4968 muxtest_0.R3R4.n4 VGND 2.29699f
C4969 muxtest_0.R3R4.t3 VGND 0.65338f
C4970 muxtest_0.R3R4.t2 VGND 0.462206f
C4971 muxtest_0.R3R4.n5 VGND 3.58348f
C4972 muxtest_0.R3R4.t8 VGND 0.362902f
C4973 muxtest_0.R3R4.t9 VGND 0.665576f
C4974 muxtest_0.R3R4.n6 VGND 3.72361f
C4975 muxtest_0.R3R4.n7 VGND 0.593498f
C4976 muxtest_0.R3R4.n8 VGND 0.122166f
C4977 muxtest_0.R3R4.n9 VGND 0.05979f
C4978 muxtest_0.R3R4.n10 VGND 6.98972f
C4979 muxtest_0.R3R4.n11 VGND 7.31123f
C4980 muxtest_0.R3R4.n12 VGND 1.03011f
C4981 ui_in[0].t6 VGND 0.006125f
C4982 ui_in[0].t0 VGND 0.003609f
C4983 ui_in[0].t8 VGND 0.006125f
C4984 ui_in[0].t3 VGND 0.003609f
C4985 ui_in[0].n0 VGND 0.010276f
C4986 ui_in[0].n1 VGND 0.015187f
C4987 ui_in[0].n2 VGND 0.004773f
C4988 ui_in[0].t9 VGND 0.003016f
C4989 ui_in[0].t5 VGND 0.004381f
C4990 ui_in[0].n3 VGND 0.010436f
C4991 ui_in[0].n4 VGND 0.005796f
C4992 ui_in[0].t1 VGND 0.003572f
C4993 ui_in[0].t7 VGND 0.00526f
C4994 ui_in[0].n5 VGND 0.012428f
C4995 ui_in[0].n6 VGND 0.002581f
C4996 ui_in[0].n7 VGND 0.001006f
C4997 ui_in[0].n8 VGND 0.091917f
C4998 ui_in[0].t4 VGND 0.005977f
C4999 ui_in[0].t2 VGND 0.002834f
C5000 ui_in[0].n9 VGND 0.021461f
C5001 ui_in[0].n10 VGND 0.004159f
C5002 ui_in[0].n11 VGND 0.105454f
C5003 ui_in[0].n12 VGND 0.068524f
C5004 ui_in[0].n13 VGND 2.54475f
C5005 ringtest_0.x4._11_.t3 VGND 0.02558f
C5006 ringtest_0.x4._11_.t2 VGND 0.02558f
C5007 ringtest_0.x4._11_.n0 VGND 0.053419f
C5008 ringtest_0.x4._11_.t12 VGND 0.042601f
C5009 ringtest_0.x4._11_.t9 VGND 0.026392f
C5010 ringtest_0.x4._11_.n1 VGND 0.086305f
C5011 ringtest_0.x4._11_.n2 VGND 0.024278f
C5012 ringtest_0.x4._11_.t7 VGND 0.027069f
C5013 ringtest_0.x4._11_.t13 VGND 0.043108f
C5014 ringtest_0.x4._11_.n3 VGND 0.058737f
C5015 ringtest_0.x4._11_.n4 VGND 0.032841f
C5016 ringtest_0.x4._11_.t17 VGND 0.023619f
C5017 ringtest_0.x4._11_.t5 VGND 0.034667f
C5018 ringtest_0.x4._11_.n5 VGND 0.06984f
C5019 ringtest_0.x4._11_.n6 VGND 0.034707f
C5020 ringtest_0.x4._11_.n7 VGND 0.494881f
C5021 ringtest_0.x4._11_.t21 VGND 0.027069f
C5022 ringtest_0.x4._11_.t10 VGND 0.043108f
C5023 ringtest_0.x4._11_.n8 VGND 0.058739f
C5024 ringtest_0.x4._11_.n9 VGND 0.133927f
C5025 ringtest_0.x4._11_.n10 VGND 0.765831f
C5026 ringtest_0.x4._11_.t11 VGND 0.021102f
C5027 ringtest_0.x4._11_.t18 VGND 0.017461f
C5028 ringtest_0.x4._11_.n11 VGND 0.092223f
C5029 ringtest_0.x4._11_.n12 VGND 0.043963f
C5030 ringtest_0.x4._11_.n13 VGND 0.150035f
C5031 ringtest_0.x4._11_.t14 VGND 0.028052f
C5032 ringtest_0.x4._11_.t4 VGND 0.019277f
C5033 ringtest_0.x4._11_.n14 VGND 0.081517f
C5034 ringtest_0.x4._11_.n15 VGND 0.011369f
C5035 ringtest_0.x4._11_.n16 VGND 0.03744f
C5036 ringtest_0.x4._11_.n17 VGND 0.156255f
C5037 ringtest_0.x4._11_.t15 VGND 0.019598f
C5038 ringtest_0.x4._11_.t19 VGND 0.028465f
C5039 ringtest_0.x4._11_.n18 VGND 0.067767f
C5040 ringtest_0.x4._11_.n19 VGND 0.143997f
C5041 ringtest_0.x4._11_.n20 VGND 0.492685f
C5042 ringtest_0.x4._11_.t8 VGND 0.042359f
C5043 ringtest_0.x4._11_.t16 VGND 0.026451f
C5044 ringtest_0.x4._11_.n21 VGND 0.080165f
C5045 ringtest_0.x4._11_.n22 VGND 0.023455f
C5046 ringtest_0.x4._11_.n23 VGND 0.356691f
C5047 ringtest_0.x4._11_.t20 VGND 0.023619f
C5048 ringtest_0.x4._11_.t6 VGND 0.034667f
C5049 ringtest_0.x4._11_.n24 VGND 0.06984f
C5050 ringtest_0.x4._11_.n25 VGND 0.014495f
C5051 ringtest_0.x4._11_.n26 VGND 0.490885f
C5052 ringtest_0.x4._11_.n27 VGND 1.19049f
C5053 ringtest_0.x4._11_.n28 VGND 0.353781f
C5054 ringtest_0.x4._11_.n29 VGND 0.021904f
C5055 ringtest_0.x4._11_.t0 VGND 0.010743f
C5056 ringtest_0.x4._11_.t1 VGND 0.010743f
C5057 ringtest_0.x4._11_.n30 VGND 0.02648f
C5058 muxtest_0.x1.x3.x4.GP VGND 2.932f
C5059 muxtest_0.x1.x2.x4.GP VGND 2.29581f
C5060 muxtest_0.x1.x1.gpo3 VGND 1.43031f
C5061 muxtest_0.x1.x3.GP4.t1 VGND 0.01297f
C5062 muxtest_0.x1.x3.GP4.t0 VGND 0.01297f
C5063 muxtest_0.x1.x3.GP4.n0 VGND 0.028494f
C5064 muxtest_0.x1.x1.x14.Y VGND 0.080663f
C5065 muxtest_0.x1.x3.GP4.n1 VGND 0.011026f
C5066 muxtest_0.x1.x3.GP4.t6 VGND 0.656398f
C5067 muxtest_0.x1.x3.GP4.t7 VGND 0.674702f
C5068 muxtest_0.x1.x3.GP4.n2 VGND 2.39862f
C5069 muxtest_0.x1.x3.GP4.t4 VGND 0.656398f
C5070 muxtest_0.x1.x3.GP4.t5 VGND 0.674702f
C5071 muxtest_0.x1.x3.GP4.n3 VGND 2.39862f
C5072 muxtest_0.x1.x3.GP4.n4 VGND 2.8073f
C5073 muxtest_0.x1.x3.GP4.n5 VGND 0.050183f
C5074 muxtest_0.x1.x3.GP4.t2 VGND 0.019954f
C5075 muxtest_0.x1.x3.GP4.t3 VGND 0.019954f
C5076 muxtest_0.x1.x3.GP4.n6 VGND 0.045883f
C5077 muxtest_0.x1.x3.GP4.n7 VGND 0.093057f
C5078 muxtest_0.x1.x3.GP1.t1 VGND 0.018021f
C5079 muxtest_0.x1.x3.GP1.t0 VGND 0.018021f
C5080 muxtest_0.x1.x3.GP1.n0 VGND 0.039591f
C5081 muxtest_0.x1.x3.GP1.n1 VGND 0.02559f
C5082 muxtest_0.x1.x3.GP1.t7 VGND 0.912037f
C5083 muxtest_0.x1.x3.GP1.t6 VGND 0.937471f
C5084 muxtest_0.x1.x3.GP1.n2 VGND 3.31176f
C5085 muxtest_0.x1.x3.GP1.t5 VGND 0.912037f
C5086 muxtest_0.x1.x3.GP1.t4 VGND 0.937471f
C5087 muxtest_0.x1.x3.GP1.n3 VGND 3.31176f
C5088 muxtest_0.x1.x3.GP1.n4 VGND 1.73806f
C5089 muxtest_0.x1.x3.GP1.t2 VGND 0.027725f
C5090 muxtest_0.x1.x3.GP1.t3 VGND 0.027725f
C5091 muxtest_0.x1.x3.GP1.n5 VGND 0.057129f
C5092 muxtest_0.x1.x3.GP1.n6 VGND 0.132634f
C5093 muxtest_0.x1.x3.GP1.n7 VGND 0.030542f
C5094 ui_in[1].t2 VGND 0.013664f
C5095 ui_in[1].t6 VGND 0.008052f
C5096 ui_in[1].t0 VGND 0.013664f
C5097 ui_in[1].t5 VGND 0.008052f
C5098 ui_in[1].n0 VGND 0.022926f
C5099 ui_in[1].n1 VGND 0.033873f
C5100 ui_in[1].n2 VGND 0.020666f
C5101 ui_in[1].t1 VGND 0.013334f
C5102 ui_in[1].t4 VGND 0.006323f
C5103 ui_in[1].n3 VGND 0.047881f
C5104 ui_in[1].n4 VGND 0.009284f
C5105 ui_in[1].n5 VGND 0.007925f
C5106 ui_in[1].t3 VGND 0.00662f
C5107 ui_in[1].t7 VGND 0.009633f
C5108 ui_in[1].n6 VGND 0.027992f
C5109 ui_in[1].n7 VGND 0.006448f
C5110 ui_in[1].n8 VGND 0.04618f
C5111 ui_in[1].n9 VGND 0.167305f
C5112 ui_in[1].t9 VGND 0.007969f
C5113 ui_in[1].t8 VGND 0.011736f
C5114 ui_in[1].n10 VGND 0.027728f
C5115 ui_in[1].n11 VGND 0.003611f
C5116 ui_in[1].n12 VGND 0.040805f
C5117 ui_in[1].n13 VGND 0.193102f
C5118 ui_in[1].n14 VGND 0.252228f
C5119 ui_in[1].n15 VGND 0.051098f
C5120 ui_in[1].n16 VGND 5.24829f
C5121 ringtest_0.x4.clknet_1_1__leaf_clk.t13 VGND 0.005541f
C5122 ringtest_0.x4.clknet_1_1__leaf_clk.t14 VGND 0.005541f
C5123 ringtest_0.x4.clknet_1_1__leaf_clk.n0 VGND 0.019676f
C5124 ringtest_0.x4.clknet_1_1__leaf_clk.t15 VGND 0.005541f
C5125 ringtest_0.x4.clknet_1_1__leaf_clk.t12 VGND 0.005541f
C5126 ringtest_0.x4.clknet_1_1__leaf_clk.n1 VGND 0.01265f
C5127 ringtest_0.x4.clknet_1_1__leaf_clk.n2 VGND 0.07993f
C5128 ringtest_0.x4.clknet_1_1__leaf_clk.t11 VGND 0.005541f
C5129 ringtest_0.x4.clknet_1_1__leaf_clk.t10 VGND 0.005541f
C5130 ringtest_0.x4.clknet_1_1__leaf_clk.n3 VGND 0.01265f
C5131 ringtest_0.x4.clknet_1_1__leaf_clk.n4 VGND 0.048044f
C5132 ringtest_0.x4.clknet_1_1__leaf_clk.t6 VGND 0.005541f
C5133 ringtest_0.x4.clknet_1_1__leaf_clk.t8 VGND 0.005541f
C5134 ringtest_0.x4.clknet_1_1__leaf_clk.n5 VGND 0.012657f
C5135 ringtest_0.x4.clknet_1_1__leaf_clk.n6 VGND 0.049559f
C5136 ringtest_0.x4.clknet_1_1__leaf_clk.t2 VGND 0.005541f
C5137 ringtest_0.x4.clknet_1_1__leaf_clk.t4 VGND 0.005541f
C5138 ringtest_0.x4.clknet_1_1__leaf_clk.n7 VGND 0.01265f
C5139 ringtest_0.x4.clknet_1_1__leaf_clk.n8 VGND 0.048044f
C5140 ringtest_0.x4.clknet_1_1__leaf_clk.t5 VGND 0.005541f
C5141 ringtest_0.x4.clknet_1_1__leaf_clk.t7 VGND 0.005541f
C5142 ringtest_0.x4.clknet_1_1__leaf_clk.n9 VGND 0.011247f
C5143 ringtest_0.x4.clknet_1_1__leaf_clk.t37 VGND 0.013817f
C5144 ringtest_0.x4.clknet_1_1__leaf_clk.t32 VGND 0.020651f
C5145 ringtest_0.x4.clknet_1_1__leaf_clk.n10 VGND 0.038168f
C5146 ringtest_0.x4.clknet_1_1__leaf_clk.t41 VGND 0.020651f
C5147 ringtest_0.x4.clknet_1_1__leaf_clk.t35 VGND 0.013817f
C5148 ringtest_0.x4.clknet_1_1__leaf_clk.n11 VGND 0.037785f
C5149 ringtest_0.x4.clknet_1_1__leaf_clk.n12 VGND 0.039947f
C5150 ringtest_0.x4.clknet_1_1__leaf_clk.t38 VGND 0.013817f
C5151 ringtest_0.x4.clknet_1_1__leaf_clk.t34 VGND 0.020651f
C5152 ringtest_0.x4.clknet_1_1__leaf_clk.n13 VGND 0.038168f
C5153 ringtest_0.x4.clknet_1_1__leaf_clk.n14 VGND 0.30833f
C5154 ringtest_0.x4.clknet_1_1__leaf_clk.t33 VGND 0.020651f
C5155 ringtest_0.x4.clknet_1_1__leaf_clk.t40 VGND 0.013817f
C5156 ringtest_0.x4.clknet_1_1__leaf_clk.n15 VGND 0.037785f
C5157 ringtest_0.x4.clknet_1_1__leaf_clk.n16 VGND 0.030886f
C5158 ringtest_0.x4.clknet_1_1__leaf_clk.n17 VGND 0.118422f
C5159 ringtest_0.x4.clknet_1_1__leaf_clk.t39 VGND 0.013817f
C5160 ringtest_0.x4.clknet_1_1__leaf_clk.t36 VGND 0.020651f
C5161 ringtest_0.x4.clknet_1_1__leaf_clk.n18 VGND 0.037832f
C5162 ringtest_0.x4.clknet_1_1__leaf_clk.n19 VGND 0.022005f
C5163 ringtest_0.x4.clknet_1_1__leaf_clk.n20 VGND 0.128874f
C5164 ringtest_0.x4.clknet_1_1__leaf_clk.n21 VGND 0.280206f
C5165 ringtest_0.x4.clknet_1_1__leaf_clk.n22 VGND 0.023331f
C5166 ringtest_0.x4.clknet_1_1__leaf_clk.n23 VGND 0.030986f
C5167 ringtest_0.x4.clknet_1_1__leaf_clk.t1 VGND 0.005541f
C5168 ringtest_0.x4.clknet_1_1__leaf_clk.t9 VGND 0.005541f
C5169 ringtest_0.x4.clknet_1_1__leaf_clk.n24 VGND 0.01265f
C5170 ringtest_0.x4.clknet_1_1__leaf_clk.n25 VGND 0.041476f
C5171 ringtest_0.x4.clknet_1_1__leaf_clk.t25 VGND 0.013193f
C5172 ringtest_0.x4.clknet_1_1__leaf_clk.t22 VGND 0.013193f
C5173 ringtest_0.x4.clknet_1_1__leaf_clk.n26 VGND 0.027449f
C5174 ringtest_0.x4.clknet_1_1__leaf_clk.t19 VGND 0.013193f
C5175 ringtest_0.x4.clknet_1_1__leaf_clk.t20 VGND 0.013193f
C5176 ringtest_0.x4.clknet_1_1__leaf_clk.n27 VGND 0.033515f
C5177 ringtest_0.x4.clknet_1_1__leaf_clk.t21 VGND 0.013193f
C5178 ringtest_0.x4.clknet_1_1__leaf_clk.t18 VGND 0.013193f
C5179 ringtest_0.x4.clknet_1_1__leaf_clk.n28 VGND 0.02781f
C5180 ringtest_0.x4.clknet_1_1__leaf_clk.n29 VGND 0.126738f
C5181 ringtest_0.x4.clknet_1_1__leaf_clk.t17 VGND 0.013193f
C5182 ringtest_0.x4.clknet_1_1__leaf_clk.t16 VGND 0.013193f
C5183 ringtest_0.x4.clknet_1_1__leaf_clk.n30 VGND 0.02781f
C5184 ringtest_0.x4.clknet_1_1__leaf_clk.n31 VGND 0.073006f
C5185 ringtest_0.x4.clknet_1_1__leaf_clk.t28 VGND 0.013193f
C5186 ringtest_0.x4.clknet_1_1__leaf_clk.t30 VGND 0.013193f
C5187 ringtest_0.x4.clknet_1_1__leaf_clk.n32 VGND 0.02781f
C5188 ringtest_0.x4.clknet_1_1__leaf_clk.n33 VGND 0.072667f
C5189 ringtest_0.x4.clknet_1_1__leaf_clk.t24 VGND 0.013193f
C5190 ringtest_0.x4.clknet_1_1__leaf_clk.t26 VGND 0.013193f
C5191 ringtest_0.x4.clknet_1_1__leaf_clk.n34 VGND 0.02781f
C5192 ringtest_0.x4.clknet_1_1__leaf_clk.n35 VGND 0.072667f
C5193 ringtest_0.x4.clknet_1_1__leaf_clk.t27 VGND 0.013193f
C5194 ringtest_0.x4.clknet_1_1__leaf_clk.t29 VGND 0.013193f
C5195 ringtest_0.x4.clknet_1_1__leaf_clk.n36 VGND 0.02781f
C5196 ringtest_0.x4.clknet_1_1__leaf_clk.n37 VGND 0.073006f
C5197 ringtest_0.x4.clknet_1_1__leaf_clk.t23 VGND 0.013193f
C5198 ringtest_0.x4.clknet_1_1__leaf_clk.t31 VGND 0.013193f
C5199 ringtest_0.x4.clknet_1_1__leaf_clk.n38 VGND 0.02781f
C5200 ringtest_0.x4.clknet_1_1__leaf_clk.n39 VGND 0.062704f
C5201 ringtest_0.x4.clknet_1_1__leaf_clk.n40 VGND 0.086346f
C5202 ringtest_0.x4.clknet_1_1__leaf_clk.n41 VGND 0.040127f
C5203 ringtest_0.x4.clknet_1_1__leaf_clk.t3 VGND 0.005541f
C5204 ringtest_0.x4.clknet_1_1__leaf_clk.t0 VGND 0.005541f
C5205 ringtest_0.x4.clknet_1_1__leaf_clk.n42 VGND 0.012211f
C5206 ringtest_0.x4.net6.t8 VGND 0.023291f
C5207 ringtest_0.x4.net6.t4 VGND 0.034395f
C5208 ringtest_0.x4.net6.n0 VGND 0.095831f
C5209 ringtest_0.x4.net6.t2 VGND 0.040459f
C5210 ringtest_0.x4.net6.t12 VGND 0.025233f
C5211 ringtest_0.x4.net6.n1 VGND 0.081347f
C5212 ringtest_0.x4.net6.n2 VGND 0.124436f
C5213 ringtest_0.x4.net6.t6 VGND 0.023291f
C5214 ringtest_0.x4.net6.t13 VGND 0.034395f
C5215 ringtest_0.x4.net6.n3 VGND 0.095831f
C5216 ringtest_0.x4.net6.n4 VGND 0.41789f
C5217 ringtest_0.x4.net6.t10 VGND 0.021456f
C5218 ringtest_0.x4.net6.t3 VGND 0.017754f
C5219 ringtest_0.x4.net6.n5 VGND 0.093771f
C5220 ringtest_0.x4.net6.n6 VGND 0.080526f
C5221 ringtest_0.x4.net6.n7 VGND 0.286209f
C5222 ringtest_0.x4.net6.t11 VGND 0.027524f
C5223 ringtest_0.x4.net6.t5 VGND 0.043832f
C5224 ringtest_0.x4.net6.n8 VGND 0.059723f
C5225 ringtest_0.x4.net6.n9 VGND 0.146037f
C5226 ringtest_0.x4.net6.n10 VGND 0.772479f
C5227 ringtest_0.x4.net6.n11 VGND 0.732404f
C5228 ringtest_0.x4.net6.t9 VGND 0.023842f
C5229 ringtest_0.x4.net6.t14 VGND 0.040459f
C5230 ringtest_0.x4.net6.n12 VGND 0.051672f
C5231 ringtest_0.x4.net6.t15 VGND 0.023842f
C5232 ringtest_0.x4.net6.t7 VGND 0.040459f
C5233 ringtest_0.x4.net6.n13 VGND 0.057394f
C5234 ringtest_0.x4.net6.n14 VGND 0.027196f
C5235 ringtest_0.x4.net6.n15 VGND 0.1061f
C5236 ringtest_0.x4.net6.n16 VGND 0.491563f
C5237 ringtest_0.x4.net6.t1 VGND 0.092732f
C5238 ringtest_0.x4.net6.n17 VGND 0.127274f
C5239 ringtest_0.x4.net6.t0 VGND 0.050895f
C5240 ringtest_0.x4.net6.n18 VGND 0.064268f
C5241 ringtest_0.x4.clknet_0_clk.t2 VGND 0.004717f
C5242 ringtest_0.x4.clknet_0_clk.t15 VGND 0.004717f
C5243 ringtest_0.x4.clknet_0_clk.n0 VGND 0.016749f
C5244 ringtest_0.x4.clknet_0_clk.t4 VGND 0.004717f
C5245 ringtest_0.x4.clknet_0_clk.t6 VGND 0.004717f
C5246 ringtest_0.x4.clknet_0_clk.n1 VGND 0.010767f
C5247 ringtest_0.x4.clknet_0_clk.n2 VGND 0.068037f
C5248 ringtest_0.x4.clknet_0_clk.t8 VGND 0.004717f
C5249 ringtest_0.x4.clknet_0_clk.t10 VGND 0.004717f
C5250 ringtest_0.x4.clknet_0_clk.n3 VGND 0.010767f
C5251 ringtest_0.x4.clknet_0_clk.n4 VGND 0.040895f
C5252 ringtest_0.x4.clknet_0_clk.t5 VGND 0.004717f
C5253 ringtest_0.x4.clknet_0_clk.t7 VGND 0.004717f
C5254 ringtest_0.x4.clknet_0_clk.n5 VGND 0.010774f
C5255 ringtest_0.x4.clknet_0_clk.n6 VGND 0.042184f
C5256 ringtest_0.x4.clknet_0_clk.t9 VGND 0.004717f
C5257 ringtest_0.x4.clknet_0_clk.t11 VGND 0.004717f
C5258 ringtest_0.x4.clknet_0_clk.n7 VGND 0.010767f
C5259 ringtest_0.x4.clknet_0_clk.n8 VGND 0.040895f
C5260 ringtest_0.x4.clknet_0_clk.t0 VGND 0.004717f
C5261 ringtest_0.x4.clknet_0_clk.t13 VGND 0.004717f
C5262 ringtest_0.x4.clknet_0_clk.n9 VGND 0.009573f
C5263 ringtest_0.x4.clknet_0_clk.t39 VGND 0.015823f
C5264 ringtest_0.x4.clknet_0_clk.t47 VGND 0.0074f
C5265 ringtest_0.x4.clknet_0_clk.t40 VGND 0.015823f
C5266 ringtest_0.x4.clknet_0_clk.t32 VGND 0.0074f
C5267 ringtest_0.x4.clknet_0_clk.t37 VGND 0.015823f
C5268 ringtest_0.x4.clknet_0_clk.t44 VGND 0.0074f
C5269 ringtest_0.x4.clknet_0_clk.t41 VGND 0.015823f
C5270 ringtest_0.x4.clknet_0_clk.t33 VGND 0.0074f
C5271 ringtest_0.x4.clknet_0_clk.n10 VGND 0.036121f
C5272 ringtest_0.x4.clknet_0_clk.n11 VGND 0.047576f
C5273 ringtest_0.x4.clknet_0_clk.n12 VGND 0.047576f
C5274 ringtest_0.x4.clknet_0_clk.n13 VGND 0.057784f
C5275 ringtest_0.x4.clknet_0_clk.n14 VGND 0.075138f
C5276 ringtest_0.x4.clknet_0_clk.t46 VGND 0.015823f
C5277 ringtest_0.x4.clknet_0_clk.t38 VGND 0.0074f
C5278 ringtest_0.x4.clknet_0_clk.t43 VGND 0.015823f
C5279 ringtest_0.x4.clknet_0_clk.t35 VGND 0.0074f
C5280 ringtest_0.x4.clknet_0_clk.t42 VGND 0.015823f
C5281 ringtest_0.x4.clknet_0_clk.t34 VGND 0.0074f
C5282 ringtest_0.x4.clknet_0_clk.t45 VGND 0.015823f
C5283 ringtest_0.x4.clknet_0_clk.t36 VGND 0.0074f
C5284 ringtest_0.x4.clknet_0_clk.n15 VGND 0.036121f
C5285 ringtest_0.x4.clknet_0_clk.n16 VGND 0.047576f
C5286 ringtest_0.x4.clknet_0_clk.n17 VGND 0.047576f
C5287 ringtest_0.x4.clknet_0_clk.n18 VGND 0.057941f
C5288 ringtest_0.x4.clknet_0_clk.n19 VGND 0.038186f
C5289 ringtest_0.x4.clknet_0_clk.n20 VGND 0.145873f
C5290 ringtest_0.x4.clknet_0_clk.n21 VGND 0.015919f
C5291 ringtest_0.x4.clknet_0_clk.n22 VGND 0.026375f
C5292 ringtest_0.x4.clknet_0_clk.t14 VGND 0.004717f
C5293 ringtest_0.x4.clknet_0_clk.t12 VGND 0.004717f
C5294 ringtest_0.x4.clknet_0_clk.n23 VGND 0.010767f
C5295 ringtest_0.x4.clknet_0_clk.n24 VGND 0.035304f
C5296 ringtest_0.x4.clknet_0_clk.t26 VGND 0.01123f
C5297 ringtest_0.x4.clknet_0_clk.t28 VGND 0.01123f
C5298 ringtest_0.x4.clknet_0_clk.n25 VGND 0.023364f
C5299 ringtest_0.x4.clknet_0_clk.t23 VGND 0.01123f
C5300 ringtest_0.x4.clknet_0_clk.t21 VGND 0.01123f
C5301 ringtest_0.x4.clknet_0_clk.n26 VGND 0.023672f
C5302 ringtest_0.x4.clknet_0_clk.t25 VGND 0.01123f
C5303 ringtest_0.x4.clknet_0_clk.t22 VGND 0.01123f
C5304 ringtest_0.x4.clknet_0_clk.n27 VGND 0.023672f
C5305 ringtest_0.x4.clknet_0_clk.t18 VGND 0.01123f
C5306 ringtest_0.x4.clknet_0_clk.t20 VGND 0.01123f
C5307 ringtest_0.x4.clknet_0_clk.n28 VGND 0.023672f
C5308 ringtest_0.x4.clknet_0_clk.t30 VGND 0.01123f
C5309 ringtest_0.x4.clknet_0_clk.t16 VGND 0.01123f
C5310 ringtest_0.x4.clknet_0_clk.n29 VGND 0.023672f
C5311 ringtest_0.x4.clknet_0_clk.t17 VGND 0.01123f
C5312 ringtest_0.x4.clknet_0_clk.t19 VGND 0.01123f
C5313 ringtest_0.x4.clknet_0_clk.n30 VGND 0.023672f
C5314 ringtest_0.x4.clknet_0_clk.t27 VGND 0.01123f
C5315 ringtest_0.x4.clknet_0_clk.t24 VGND 0.01123f
C5316 ringtest_0.x4.clknet_0_clk.n31 VGND 0.028528f
C5317 ringtest_0.x4.clknet_0_clk.t29 VGND 0.01123f
C5318 ringtest_0.x4.clknet_0_clk.t31 VGND 0.01123f
C5319 ringtest_0.x4.clknet_0_clk.n32 VGND 0.023672f
C5320 ringtest_0.x4.clknet_0_clk.n33 VGND 0.107879f
C5321 ringtest_0.x4.clknet_0_clk.n34 VGND 0.062143f
C5322 ringtest_0.x4.clknet_0_clk.n35 VGND 0.061854f
C5323 ringtest_0.x4.clknet_0_clk.n36 VGND 0.061854f
C5324 ringtest_0.x4.clknet_0_clk.n37 VGND 0.062143f
C5325 ringtest_0.x4.clknet_0_clk.n38 VGND 0.053374f
C5326 ringtest_0.x4.clknet_0_clk.n39 VGND 0.073498f
C5327 ringtest_0.x4.clknet_0_clk.n40 VGND 0.034156f
C5328 ringtest_0.x4.clknet_0_clk.t1 VGND 0.004717f
C5329 ringtest_0.x4.clknet_0_clk.t3 VGND 0.004717f
C5330 ringtest_0.x4.clknet_0_clk.n41 VGND 0.010394f
C5331 ua[2].t8 VGND 0.247385f
C5332 ua[2].n0 VGND 0.307673f
C5333 ua[2].t12 VGND 0.191554f
C5334 ua[2].t9 VGND 0.254197f
C5335 ua[2].n1 VGND 1.28275f
C5336 ua[2].n2 VGND 0.434029f
C5337 ua[2].t13 VGND 0.187785f
C5338 ua[2].n3 VGND 0.280396f
C5339 ua[2].n4 VGND 0.390968f
C5340 ua[2].t3 VGND 0.247385f
C5341 ua[2].n5 VGND 0.307673f
C5342 ua[2].t15 VGND 0.191554f
C5343 ua[2].t2 VGND 0.254197f
C5344 ua[2].n6 VGND 1.28275f
C5345 ua[2].n7 VGND 0.434029f
C5346 ua[2].t14 VGND 0.187785f
C5347 ua[2].n8 VGND 0.280396f
C5348 ua[2].n9 VGND 0.385643f
C5349 ua[2].n10 VGND 0.201153f
C5350 ua[2].n11 VGND 0.0295f
C5351 ua[2].n12 VGND 0.068599f
C5352 ua[2].n13 VGND 0.274656f
C5353 ua[2].t7 VGND 0.247385f
C5354 ua[2].n14 VGND 0.307673f
C5355 ua[2].t1 VGND 0.191554f
C5356 ua[2].t6 VGND 0.254197f
C5357 ua[2].n15 VGND 1.28275f
C5358 ua[2].n16 VGND 0.434029f
C5359 ua[2].t0 VGND 0.187785f
C5360 ua[2].n17 VGND 0.280396f
C5361 ua[2].n18 VGND 0.380387f
C5362 ua[2].n19 VGND 0.206106f
C5363 ua[2].n20 VGND 0.522334f
C5364 ua[2].t5 VGND 0.247385f
C5365 ua[2].n21 VGND 0.307673f
C5366 ua[2].t10 VGND 0.191554f
C5367 ua[2].t4 VGND 0.254197f
C5368 ua[2].n22 VGND 1.28275f
C5369 ua[2].n23 VGND 0.434029f
C5370 ua[2].t11 VGND 0.187785f
C5371 ua[2].n24 VGND 0.280396f
C5372 ua[2].n25 VGND 0.383777f
C5373 ua[2].n26 VGND 0.202647f
C5374 ua[2].n27 VGND 0.509311f
C5375 ua[2].n28 VGND 9.99833f
C5376 ua[3].t7 VGND 0.195583f
C5377 ua[3].n0 VGND 0.292041f
C5378 ua[3].t9 VGND 0.199509f
C5379 ua[3].t3 VGND 0.264753f
C5380 ua[3].n1 VGND 1.33602f
C5381 ua[3].n2 VGND 0.452054f
C5382 ua[3].t2 VGND 0.257658f
C5383 ua[3].n3 VGND 0.32045f
C5384 ua[3].n4 VGND 0.405279f
C5385 ua[3].t0 VGND 0.195583f
C5386 ua[3].n5 VGND 0.292041f
C5387 ua[3].t1 VGND 0.199509f
C5388 ua[3].t6 VGND 0.264753f
C5389 ua[3].n6 VGND 1.33602f
C5390 ua[3].n7 VGND 0.452054f
C5391 ua[3].t8 VGND 0.257658f
C5392 ua[3].n8 VGND 0.32045f
C5393 ua[3].n9 VGND 0.407204f
C5394 ua[3].t4 VGND 0.370241f
C5395 ua[3].t5 VGND 0.261912f
C5396 ua[3].n10 VGND 2.0306f
C5397 ua[3].t11 VGND 0.205641f
C5398 ua[3].t10 VGND 0.377153f
C5399 ua[3].n11 VGND 2.11001f
C5400 ua[3].n12 VGND 0.336309f
C5401 ua[3].n13 VGND 0.069845f
C5402 ua[3].n14 VGND 0.028001f
C5403 ua[3].n15 VGND 1.71586f
C5404 ua[3].n16 VGND 0.514233f
C5405 ua[3].n17 VGND 0.337655f
C5406 muxtest_0.x2.x2.GP1.t1 VGND 0.012908f
C5407 muxtest_0.x2.x2.GP1.t0 VGND 0.012908f
C5408 muxtest_0.x2.x2.GP1.n0 VGND 0.028358f
C5409 muxtest_0.x2.x2.GP1.n1 VGND 0.018329f
C5410 muxtest_0.x2.x2.GP1.t5 VGND 0.653268f
C5411 muxtest_0.x2.x2.GP1.t4 VGND 0.671486f
C5412 muxtest_0.x2.x2.GP1.n2 VGND 2.37213f
C5413 muxtest_0.x2.x2.GP1.t3 VGND 0.019859f
C5414 muxtest_0.x2.x2.GP1.t2 VGND 0.019859f
C5415 muxtest_0.x2.x2.GP1.n3 VGND 0.04092f
C5416 muxtest_0.x2.x2.GP1.n4 VGND 0.100085f
C5417 muxtest_0.x2.x2.GP1.n5 VGND 0.021877f
C5418 VDPWR.n0 VGND 0.003488f
C5419 VDPWR.t881 VGND 0.007172f
C5420 VDPWR.n1 VGND 0.007983f
C5421 VDPWR.t113 VGND 7.56e-19
C5422 VDPWR.t197 VGND 0.001148f
C5423 VDPWR.n2 VGND 0.001983f
C5424 VDPWR.t879 VGND 0.007175f
C5425 VDPWR.t307 VGND 0.00704f
C5426 VDPWR.n3 VGND 0.006705f
C5427 VDPWR.n4 VGND 0.003488f
C5428 VDPWR.n5 VGND 0.003158f
C5429 VDPWR.t56 VGND 0.001036f
C5430 VDPWR.n6 VGND 0.00294f
C5431 VDPWR.t217 VGND 0.004259f
C5432 VDPWR.n7 VGND 0.00392f
C5433 VDPWR.n8 VGND 0.003499f
C5434 VDPWR.t305 VGND 0.007175f
C5435 VDPWR.n9 VGND 5.76e-19
C5436 VDPWR.t988 VGND 0.003015f
C5437 VDPWR.t662 VGND 0.004984f
C5438 VDPWR.n10 VGND 0.004913f
C5439 VDPWR.n11 VGND 0.005888f
C5440 VDPWR.t1217 VGND 0.020799f
C5441 VDPWR.n12 VGND 0.018812f
C5442 VDPWR.t261 VGND 5.64e-19
C5443 VDPWR.t793 VGND 0.001513f
C5444 VDPWR.n13 VGND 0.006904f
C5445 VDPWR.n14 VGND 0.003647f
C5446 VDPWR.t663 VGND 0.004984f
C5447 VDPWR.n15 VGND 0.01361f
C5448 VDPWR.n16 VGND 0.010753f
C5449 VDPWR.n17 VGND 0.013967f
C5450 VDPWR.n18 VGND 0.008065f
C5451 VDPWR.n19 VGND 0.005888f
C5452 VDPWR.n20 VGND 0.004416f
C5453 VDPWR.n21 VGND 0.005354f
C5454 VDPWR.n22 VGND 0.006068f
C5455 VDPWR.n23 VGND 0.013691f
C5456 VDPWR.t1038 VGND 0.014151f
C5457 VDPWR.n24 VGND 7.37e-19
C5458 VDPWR.n25 VGND 0.004416f
C5459 VDPWR.n26 VGND 0.00136f
C5460 VDPWR.t131 VGND 7.56e-19
C5461 VDPWR.t961 VGND 0.001148f
C5462 VDPWR.n27 VGND 0.001983f
C5463 VDPWR.n28 VGND 0.005856f
C5464 VDPWR.n29 VGND 0.003488f
C5465 VDPWR.t1282 VGND 0.020799f
C5466 VDPWR.n30 VGND 0.005184f
C5467 VDPWR.n31 VGND 0.003488f
C5468 VDPWR.t207 VGND 5.64e-19
C5469 VDPWR.t909 VGND 0.001513f
C5470 VDPWR.n32 VGND 0.006904f
C5471 VDPWR.t1268 VGND 0.020799f
C5472 VDPWR.t927 VGND 0.003047f
C5473 VDPWR.n33 VGND 0.009651f
C5474 VDPWR.n34 VGND 0.005344f
C5475 VDPWR.n35 VGND 0.002933f
C5476 VDPWR.t529 VGND 0.004984f
C5477 VDPWR.n36 VGND 0.004913f
C5478 VDPWR.n37 VGND 0.018812f
C5479 VDPWR.n38 VGND 0.008065f
C5480 VDPWR.n39 VGND 0.013967f
C5481 VDPWR.t926 VGND 0.02849f
C5482 VDPWR.t908 VGND 0.027547f
C5483 VDPWR.t528 VGND 0.020377f
C5484 VDPWR.t206 VGND 0.029245f
C5485 VDPWR.t1136 VGND 0.02849f
C5486 VDPWR.t930 VGND 0.032453f
C5487 VDPWR.t960 VGND 0.023585f
C5488 VDPWR.t130 VGND 0.012641f
C5489 VDPWR.t208 VGND 0.005849f
C5490 VDPWR.t210 VGND 0.020566f
C5491 VDPWR.n40 VGND 0.026837f
C5492 VDPWR.t211 VGND 0.007137f
C5493 VDPWR.n41 VGND 0.002016f
C5494 VDPWR.n42 VGND 0.0024f
C5495 VDPWR.n43 VGND 0.018611f
C5496 VDPWR.n44 VGND 0.005471f
C5497 VDPWR.t530 VGND 0.004984f
C5498 VDPWR.n45 VGND 0.008777f
C5499 VDPWR.n46 VGND 0.010753f
C5500 VDPWR.n47 VGND 0.003648f
C5501 VDPWR.n48 VGND 0.02906f
C5502 VDPWR.n49 VGND 0.039529f
C5503 VDPWR.t712 VGND 0.004984f
C5504 VDPWR.n50 VGND 0.009746f
C5505 VDPWR.n51 VGND 0.018812f
C5506 VDPWR.n52 VGND 0.011593f
C5507 VDPWR.t950 VGND 0.007172f
C5508 VDPWR.n53 VGND 0.00838f
C5509 VDPWR.n54 VGND 0.003488f
C5510 VDPWR.n55 VGND 0.001519f
C5511 VDPWR.n56 VGND 0.001519f
C5512 VDPWR.n57 VGND 0.1025f
C5513 VDPWR.t569 VGND 0.004984f
C5514 VDPWR.n58 VGND 0.004913f
C5515 VDPWR.n59 VGND 0.005888f
C5516 VDPWR.t1215 VGND 0.020799f
C5517 VDPWR.n60 VGND 0.018812f
C5518 VDPWR.n61 VGND 0.003647f
C5519 VDPWR.t570 VGND 0.004984f
C5520 VDPWR.n62 VGND 0.01361f
C5521 VDPWR.n63 VGND 0.014953f
C5522 VDPWR.n64 VGND 0.011593f
C5523 VDPWR.n65 VGND 0.005888f
C5524 VDPWR.n66 VGND 0.004416f
C5525 VDPWR.n67 VGND 0.005604f
C5526 VDPWR.t1032 VGND 0.007175f
C5527 VDPWR.n68 VGND 0.009278f
C5528 VDPWR.n69 VGND 0.003488f
C5529 VDPWR.n70 VGND 0.005888f
C5530 VDPWR.n71 VGND 0.004416f
C5531 VDPWR.t60 VGND 0.007172f
C5532 VDPWR.n72 VGND 0.00847f
C5533 VDPWR.t929 VGND 0.007175f
C5534 VDPWR.n73 VGND 0.009165f
C5535 VDPWR.n74 VGND 0.003488f
C5536 VDPWR.n75 VGND 0.005888f
C5537 VDPWR.n76 VGND 0.004416f
C5538 VDPWR.t1022 VGND 0.007172f
C5539 VDPWR.n77 VGND 0.00847f
C5540 VDPWR.t947 VGND 0.007175f
C5541 VDPWR.n78 VGND 0.009165f
C5542 VDPWR.n79 VGND 0.001519f
C5543 VDPWR.n80 VGND 0.005888f
C5544 VDPWR.n81 VGND 0.004416f
C5545 VDPWR.n82 VGND 0.00224f
C5546 VDPWR.t711 VGND 0.064097f
C5547 VDPWR.t568 VGND 0.039378f
C5548 VDPWR.t1031 VGND 0.016158f
C5549 VDPWR.t59 VGND 0.022364f
C5550 VDPWR.t928 VGND 0.016158f
C5551 VDPWR.t1021 VGND 0.022364f
C5552 VDPWR.t946 VGND 0.016158f
C5553 VDPWR.t949 VGND 0.024184f
C5554 VDPWR.n83 VGND 0.026472f
C5555 VDPWR.n84 VGND 0.012237f
C5556 VDPWR.n85 VGND 0.005471f
C5557 VDPWR.t713 VGND 0.004984f
C5558 VDPWR.n86 VGND 0.008777f
C5559 VDPWR.n87 VGND 0.014953f
C5560 VDPWR.n88 VGND 0.002976f
C5561 VDPWR.n89 VGND 0.027044f
C5562 VDPWR.n90 VGND 0.026223f
C5563 VDPWR.n91 VGND 6.08e-19
C5564 VDPWR.t209 VGND 0.007136f
C5565 VDPWR.n92 VGND 0.013312f
C5566 VDPWR.t1138 VGND 0.007172f
C5567 VDPWR.n93 VGND 0.008357f
C5568 VDPWR.t931 VGND 0.002363f
C5569 VDPWR.t1039 VGND 0.006281f
C5570 VDPWR.n94 VGND 0.003563f
C5571 VDPWR.t1137 VGND 0.007041f
C5572 VDPWR.n95 VGND 0.007429f
C5573 VDPWR.n96 VGND 0.009555f
C5574 VDPWR.n97 VGND 0.001258f
C5575 VDPWR.n98 VGND 0.005888f
C5576 VDPWR.n99 VGND 0.003488f
C5577 VDPWR.n100 VGND 0.002016f
C5578 VDPWR.n101 VGND 0.00224f
C5579 VDPWR.n102 VGND 0.012275f
C5580 VDPWR.n103 VGND 0.032875f
C5581 VDPWR.t112 VGND 0.006226f
C5582 VDPWR.t880 VGND 0.016226f
C5583 VDPWR.t878 VGND 0.018113f
C5584 VDPWR.t196 VGND 0.012641f
C5585 VDPWR.t55 VGND 0.023585f
C5586 VDPWR.t306 VGND 0.033207f
C5587 VDPWR.t304 VGND 0.016226f
C5588 VDPWR.t216 VGND 0.012641f
C5589 VDPWR.t260 VGND 0.029245f
C5590 VDPWR.t661 VGND 0.020377f
C5591 VDPWR.t792 VGND 0.027547f
C5592 VDPWR.t987 VGND 0.02849f
C5593 VDPWR.n104 VGND 0.019402f
C5594 VDPWR.n105 VGND 0.005637f
C5595 VDPWR.n106 VGND 0.003862f
C5596 VDPWR.n107 VGND 0.009272f
C5597 VDPWR.n108 VGND 0.002696f
C5598 VDPWR.n109 VGND 0.005888f
C5599 VDPWR.n110 VGND 0.004416f
C5600 VDPWR.n111 VGND 0.002625f
C5601 VDPWR.n112 VGND 0.008924f
C5602 VDPWR.n113 VGND 0.006148f
C5603 VDPWR.n114 VGND 0.004064f
C5604 VDPWR.n115 VGND 0.011493f
C5605 VDPWR.n116 VGND 0.0731f
C5606 VDPWR.n117 VGND 7.840919f
C5607 VDPWR.n118 VGND 0.489074f
C5608 VDPWR.t893 VGND 0.007172f
C5609 VDPWR.n119 VGND 0.00838f
C5610 VDPWR.t369 VGND 0.007175f
C5611 VDPWR.n120 VGND 0.009029f
C5612 VDPWR.n121 VGND 0.023921f
C5613 VDPWR.t371 VGND 0.007172f
C5614 VDPWR.t75 VGND 0.007175f
C5615 VDPWR.n122 VGND 0.010921f
C5616 VDPWR.t77 VGND 0.007172f
C5617 VDPWR.n123 VGND 0.00847f
C5618 VDPWR.t245 VGND 0.007175f
C5619 VDPWR.t247 VGND 0.007172f
C5620 VDPWR.n124 VGND 0.00847f
C5621 VDPWR.t87 VGND 0.007175f
C5622 VDPWR.t85 VGND 0.007172f
C5623 VDPWR.n125 VGND 0.00847f
C5624 VDPWR.t89 VGND 0.007175f
C5625 VDPWR.t91 VGND 0.007172f
C5626 VDPWR.n126 VGND 0.00847f
C5627 VDPWR.n127 VGND 0.014476f
C5628 VDPWR.n128 VGND 0.013372f
C5629 VDPWR.t885 VGND 0.007172f
C5630 VDPWR.n129 VGND 0.00847f
C5631 VDPWR.n130 VGND 0.001519f
C5632 VDPWR.n131 VGND 0.001519f
C5633 VDPWR.n132 VGND 0.001519f
C5634 VDPWR.n133 VGND 0.001519f
C5635 VDPWR.n134 VGND 0.022941f
C5636 VDPWR.t905 VGND 0.007172f
C5637 VDPWR.n135 VGND 0.00838f
C5638 VDPWR.n136 VGND 0.01181f
C5639 VDPWR.n137 VGND 0.008587f
C5640 VDPWR.n138 VGND 0.013249f
C5641 VDPWR.t241 VGND 0.007179f
C5642 VDPWR.t861 VGND 0.0018f
C5643 VDPWR.t243 VGND 0.0018f
C5644 VDPWR.n139 VGND 0.003864f
C5645 VDPWR.n140 VGND 0.005287f
C5646 VDPWR.t859 VGND 0.006979f
C5647 VDPWR.n141 VGND 0.009924f
C5648 VDPWR.n142 VGND 0.04768f
C5649 VDPWR.n143 VGND 0.001711f
C5650 VDPWR.n144 VGND 0.010005f
C5651 VDPWR.n145 VGND 0.01181f
C5652 VDPWR.t858 VGND 0.041519f
C5653 VDPWR.t860 VGND 0.017977f
C5654 VDPWR.t242 VGND 0.017977f
C5655 VDPWR.t240 VGND 0.015837f
C5656 VDPWR.n146 VGND 0.021229f
C5657 VDPWR.n147 VGND 0.022941f
C5658 VDPWR.n148 VGND 0.01181f
C5659 VDPWR.n149 VGND 0.008587f
C5660 VDPWR.n150 VGND 0.008587f
C5661 VDPWR.n151 VGND 0.013372f
C5662 VDPWR.n152 VGND 0.001519f
C5663 VDPWR.n153 VGND 0.001519f
C5664 VDPWR.n154 VGND 0.001519f
C5665 VDPWR.t887 VGND 0.007175f
C5666 VDPWR.n155 VGND 0.009165f
C5667 VDPWR.n156 VGND 0.013372f
C5668 VDPWR.n157 VGND 0.022572f
C5669 VDPWR.n158 VGND 0.016929f
C5670 VDPWR.t889 VGND 0.007172f
C5671 VDPWR.n159 VGND 0.00847f
C5672 VDPWR.t181 VGND 0.007175f
C5673 VDPWR.n160 VGND 0.009165f
C5674 VDPWR.n161 VGND 0.013372f
C5675 VDPWR.n162 VGND 0.022572f
C5676 VDPWR.n163 VGND 0.016929f
C5677 VDPWR.t183 VGND 0.007172f
C5678 VDPWR.n164 VGND 0.00847f
C5679 VDPWR.t171 VGND 0.007175f
C5680 VDPWR.n165 VGND 0.009165f
C5681 VDPWR.n166 VGND 0.013372f
C5682 VDPWR.n167 VGND 0.022572f
C5683 VDPWR.n168 VGND 0.016929f
C5684 VDPWR.t173 VGND 0.007172f
C5685 VDPWR.n169 VGND 0.00847f
C5686 VDPWR.t903 VGND 0.007175f
C5687 VDPWR.n170 VGND 0.009165f
C5688 VDPWR.n171 VGND 0.001519f
C5689 VDPWR.n172 VGND 0.022572f
C5690 VDPWR.n173 VGND 0.016929f
C5691 VDPWR.n174 VGND 0.008587f
C5692 VDPWR.n175 VGND 0.011946f
C5693 VDPWR.n176 VGND 0.028292f
C5694 VDPWR.t904 VGND 0.024184f
C5695 VDPWR.t902 VGND 0.015813f
C5696 VDPWR.t172 VGND 0.022364f
C5697 VDPWR.t170 VGND 0.016158f
C5698 VDPWR.t182 VGND 0.022364f
C5699 VDPWR.t180 VGND 0.016158f
C5700 VDPWR.t888 VGND 0.022364f
C5701 VDPWR.t886 VGND 0.016158f
C5702 VDPWR.t884 VGND 0.022364f
C5703 VDPWR.t882 VGND 0.016158f
C5704 VDPWR.t291 VGND 0.022364f
C5705 VDPWR.t289 VGND 0.016158f
C5706 VDPWR.t842 VGND 0.022364f
C5707 VDPWR.t844 VGND 0.016158f
C5708 VDPWR.t840 VGND 0.022364f
C5709 VDPWR.t838 VGND 0.016158f
C5710 VDPWR.t898 VGND 0.022364f
C5711 VDPWR.t896 VGND 0.016158f
C5712 VDPWR.n177 VGND 0.008587f
C5713 VDPWR.n178 VGND 0.026055f
C5714 VDPWR.t897 VGND 0.007175f
C5715 VDPWR.n179 VGND 0.009029f
C5716 VDPWR.n180 VGND 0.013372f
C5717 VDPWR.n181 VGND 0.022572f
C5718 VDPWR.n182 VGND 0.016929f
C5719 VDPWR.t899 VGND 0.007172f
C5720 VDPWR.n183 VGND 0.00847f
C5721 VDPWR.t839 VGND 0.007175f
C5722 VDPWR.n184 VGND 0.009165f
C5723 VDPWR.n185 VGND 0.013372f
C5724 VDPWR.n186 VGND 0.022572f
C5725 VDPWR.n187 VGND 0.016929f
C5726 VDPWR.t841 VGND 0.007172f
C5727 VDPWR.n188 VGND 0.00847f
C5728 VDPWR.t845 VGND 0.007175f
C5729 VDPWR.n189 VGND 0.009165f
C5730 VDPWR.n190 VGND 0.013372f
C5731 VDPWR.n191 VGND 0.022572f
C5732 VDPWR.n192 VGND 0.016929f
C5733 VDPWR.t843 VGND 0.007172f
C5734 VDPWR.n193 VGND 0.00847f
C5735 VDPWR.t290 VGND 0.007175f
C5736 VDPWR.n194 VGND 0.009165f
C5737 VDPWR.n195 VGND 0.013372f
C5738 VDPWR.n196 VGND 0.022572f
C5739 VDPWR.n197 VGND 0.016929f
C5740 VDPWR.t292 VGND 0.007172f
C5741 VDPWR.n198 VGND 0.00847f
C5742 VDPWR.t883 VGND 0.007175f
C5743 VDPWR.n199 VGND 0.009165f
C5744 VDPWR.n200 VGND 0.001519f
C5745 VDPWR.n201 VGND 0.01374f
C5746 VDPWR.n202 VGND 1.62819f
C5747 VDPWR.n203 VGND 1.62991f
C5748 VDPWR.t313 VGND 0.007175f
C5749 VDPWR.t311 VGND 0.007172f
C5750 VDPWR.n204 VGND 0.00847f
C5751 VDPWR.t276 VGND 0.007175f
C5752 VDPWR.t274 VGND 0.007172f
C5753 VDPWR.n205 VGND 0.00847f
C5754 VDPWR.t278 VGND 0.007175f
C5755 VDPWR.t280 VGND 0.007172f
C5756 VDPWR.n206 VGND 0.00847f
C5757 VDPWR.t895 VGND 0.007175f
C5758 VDPWR.n207 VGND 0.023921f
C5759 VDPWR.n208 VGND 0.028948f
C5760 VDPWR.n209 VGND 0.001519f
C5761 VDPWR.n210 VGND 0.009165f
C5762 VDPWR.n211 VGND 0.010921f
C5763 VDPWR.n212 VGND 0.023921f
C5764 VDPWR.n213 VGND 0.028948f
C5765 VDPWR.n214 VGND 0.001519f
C5766 VDPWR.n215 VGND 0.009165f
C5767 VDPWR.n216 VGND 0.010921f
C5768 VDPWR.n217 VGND 0.023921f
C5769 VDPWR.n218 VGND 0.028948f
C5770 VDPWR.n219 VGND 0.001519f
C5771 VDPWR.n220 VGND 0.009165f
C5772 VDPWR.n221 VGND 0.010921f
C5773 VDPWR.n222 VGND 0.023921f
C5774 VDPWR.n223 VGND 0.028948f
C5775 VDPWR.n224 VGND 0.001519f
C5776 VDPWR.n225 VGND 0.009165f
C5777 VDPWR.n226 VGND 0.010921f
C5778 VDPWR.n227 VGND 0.023921f
C5779 VDPWR.n228 VGND 0.019415f
C5780 VDPWR.n229 VGND 0.001519f
C5781 VDPWR.n230 VGND 0.009165f
C5782 VDPWR.n231 VGND 0.010921f
C5783 VDPWR.n232 VGND 0.023921f
C5784 VDPWR.n233 VGND 0.028948f
C5785 VDPWR.n234 VGND 0.001519f
C5786 VDPWR.n235 VGND 0.009165f
C5787 VDPWR.n236 VGND 0.010921f
C5788 VDPWR.n237 VGND 0.023921f
C5789 VDPWR.n238 VGND 0.028948f
C5790 VDPWR.n239 VGND 0.001519f
C5791 VDPWR.n240 VGND 0.009165f
C5792 VDPWR.n241 VGND 0.010921f
C5793 VDPWR.n242 VGND 0.023921f
C5794 VDPWR.n243 VGND 0.028948f
C5795 VDPWR.n244 VGND 0.001519f
C5796 VDPWR.n245 VGND 0.009165f
C5797 VDPWR.n246 VGND 0.00847f
C5798 VDPWR.n247 VGND 0.001519f
C5799 VDPWR.n248 VGND 0.028948f
C5800 VDPWR.n249 VGND 0.010921f
C5801 VDPWR.n250 VGND 0.031124f
C5802 VDPWR.t368 VGND 0.01252f
C5803 VDPWR.t370 VGND 0.026002f
C5804 VDPWR.t74 VGND 0.01252f
C5805 VDPWR.t76 VGND 0.026002f
C5806 VDPWR.t244 VGND 0.01252f
C5807 VDPWR.t246 VGND 0.026002f
C5808 VDPWR.t86 VGND 0.01252f
C5809 VDPWR.t84 VGND 0.026002f
C5810 VDPWR.t88 VGND 0.01252f
C5811 VDPWR.t90 VGND 0.026002f
C5812 VDPWR.t312 VGND 0.01252f
C5813 VDPWR.t310 VGND 0.026002f
C5814 VDPWR.t275 VGND 0.01252f
C5815 VDPWR.t273 VGND 0.026002f
C5816 VDPWR.t277 VGND 0.01252f
C5817 VDPWR.t279 VGND 0.026002f
C5818 VDPWR.t894 VGND 0.01252f
C5819 VDPWR.t892 VGND 0.03644f
C5820 VDPWR.n251 VGND 0.035343f
C5821 VDPWR.n252 VGND 0.012134f
C5822 VDPWR.n253 VGND 3.92216f
C5823 VDPWR.n254 VGND 0.058044f
C5824 VDPWR.n255 VGND 0.105387f
C5825 VDPWR.n256 VGND 4.47053f
C5826 VDPWR.n257 VGND 2.12953f
C5827 VDPWR.n258 VGND 0.003488f
C5828 VDPWR.t177 VGND 0.007172f
C5829 VDPWR.n259 VGND 0.007983f
C5830 VDPWR.t109 VGND 7.56e-19
C5831 VDPWR.t990 VGND 0.001148f
C5832 VDPWR.n260 VGND 0.001983f
C5833 VDPWR.t179 VGND 0.007175f
C5834 VDPWR.t71 VGND 0.00704f
C5835 VDPWR.n261 VGND 0.006705f
C5836 VDPWR.n262 VGND 0.003488f
C5837 VDPWR.n263 VGND 0.003158f
C5838 VDPWR.t1090 VGND 0.001036f
C5839 VDPWR.n264 VGND 0.00294f
C5840 VDPWR.t189 VGND 0.004259f
C5841 VDPWR.n265 VGND 0.00392f
C5842 VDPWR.n266 VGND 0.003499f
C5843 VDPWR.t73 VGND 0.007175f
C5844 VDPWR.n267 VGND 5.76e-19
C5845 VDPWR.t765 VGND 0.003015f
C5846 VDPWR.t540 VGND 0.004984f
C5847 VDPWR.n268 VGND 0.004913f
C5848 VDPWR.n269 VGND 0.005888f
C5849 VDPWR.t1228 VGND 0.020799f
C5850 VDPWR.n270 VGND 0.018812f
C5851 VDPWR.t286 VGND 5.64e-19
C5852 VDPWR.t62 VGND 0.001513f
C5853 VDPWR.n271 VGND 0.006904f
C5854 VDPWR.n272 VGND 0.003647f
C5855 VDPWR.t541 VGND 0.004984f
C5856 VDPWR.n273 VGND 0.01361f
C5857 VDPWR.n274 VGND 0.010753f
C5858 VDPWR.n275 VGND 0.013967f
C5859 VDPWR.n276 VGND 0.008065f
C5860 VDPWR.n277 VGND 0.005888f
C5861 VDPWR.n278 VGND 0.004416f
C5862 VDPWR.n279 VGND 0.005354f
C5863 VDPWR.n280 VGND 0.006068f
C5864 VDPWR.n281 VGND 0.013691f
C5865 VDPWR.t110 VGND 0.014151f
C5866 VDPWR.n282 VGND 7.37e-19
C5867 VDPWR.n283 VGND 0.004416f
C5868 VDPWR.n284 VGND 0.00136f
C5869 VDPWR.t236 VGND 7.56e-19
C5870 VDPWR.t849 VGND 0.001148f
C5871 VDPWR.n285 VGND 0.001983f
C5872 VDPWR.n286 VGND 0.005856f
C5873 VDPWR.n287 VGND 0.003488f
C5874 VDPWR.t1201 VGND 0.020799f
C5875 VDPWR.n288 VGND 0.005184f
C5876 VDPWR.n289 VGND 0.003488f
C5877 VDPWR.t303 VGND 5.64e-19
C5878 VDPWR.t1092 VGND 0.001513f
C5879 VDPWR.n290 VGND 0.006904f
C5880 VDPWR.t1200 VGND 0.020799f
C5881 VDPWR.t107 VGND 0.003047f
C5882 VDPWR.n291 VGND 0.009651f
C5883 VDPWR.n292 VGND 0.005344f
C5884 VDPWR.n293 VGND 0.002933f
C5885 VDPWR.t600 VGND 0.004984f
C5886 VDPWR.n294 VGND 0.004913f
C5887 VDPWR.n295 VGND 0.018812f
C5888 VDPWR.n296 VGND 0.008065f
C5889 VDPWR.n297 VGND 0.013967f
C5890 VDPWR.t106 VGND 0.02849f
C5891 VDPWR.t1091 VGND 0.027547f
C5892 VDPWR.t599 VGND 0.020377f
C5893 VDPWR.t302 VGND 0.029245f
C5894 VDPWR.t851 VGND 0.02849f
C5895 VDPWR.t104 VGND 0.032453f
C5896 VDPWR.t848 VGND 0.023585f
C5897 VDPWR.t235 VGND 0.012641f
C5898 VDPWR.t1010 VGND 0.005849f
C5899 VDPWR.t1008 VGND 0.020566f
C5900 VDPWR.n298 VGND 0.026837f
C5901 VDPWR.t1009 VGND 0.007137f
C5902 VDPWR.n299 VGND 0.002016f
C5903 VDPWR.n300 VGND 0.0024f
C5904 VDPWR.n301 VGND 0.018611f
C5905 VDPWR.n302 VGND 0.005471f
C5906 VDPWR.t601 VGND 0.004984f
C5907 VDPWR.n303 VGND 0.008777f
C5908 VDPWR.n304 VGND 0.010753f
C5909 VDPWR.n305 VGND 0.003648f
C5910 VDPWR.n306 VGND 0.02906f
C5911 VDPWR.n307 VGND 0.039529f
C5912 VDPWR.t597 VGND 0.004984f
C5913 VDPWR.n308 VGND 0.009746f
C5914 VDPWR.n309 VGND 0.018812f
C5915 VDPWR.n310 VGND 0.011593f
C5916 VDPWR.t1097 VGND 0.007172f
C5917 VDPWR.n311 VGND 0.00838f
C5918 VDPWR.n312 VGND 0.003488f
C5919 VDPWR.n313 VGND 0.001519f
C5920 VDPWR.n314 VGND 0.001519f
C5921 VDPWR.n315 VGND 0.1025f
C5922 VDPWR.t436 VGND 0.004984f
C5923 VDPWR.n316 VGND 0.004913f
C5924 VDPWR.n317 VGND 0.005888f
C5925 VDPWR.t1263 VGND 0.020799f
C5926 VDPWR.n318 VGND 0.018812f
C5927 VDPWR.t437 VGND 0.004984f
C5928 VDPWR.n319 VGND 0.003647f
C5929 VDPWR.n320 VGND 0.01361f
C5930 VDPWR.n321 VGND 0.014953f
C5931 VDPWR.n322 VGND 0.011593f
C5932 VDPWR.n323 VGND 0.005888f
C5933 VDPWR.n324 VGND 0.004416f
C5934 VDPWR.n325 VGND 0.005604f
C5935 VDPWR.t234 VGND 0.007175f
C5936 VDPWR.n326 VGND 0.009278f
C5937 VDPWR.n327 VGND 0.003488f
C5938 VDPWR.n328 VGND 0.005888f
C5939 VDPWR.n329 VGND 0.004416f
C5940 VDPWR.t238 VGND 0.007172f
C5941 VDPWR.n330 VGND 0.00847f
C5942 VDPWR.t815 VGND 0.007175f
C5943 VDPWR.n331 VGND 0.009165f
C5944 VDPWR.n332 VGND 0.003488f
C5945 VDPWR.n333 VGND 0.005888f
C5946 VDPWR.n334 VGND 0.004416f
C5947 VDPWR.t1046 VGND 0.007172f
C5948 VDPWR.n335 VGND 0.00847f
C5949 VDPWR.t1099 VGND 0.007175f
C5950 VDPWR.n336 VGND 0.009165f
C5951 VDPWR.n337 VGND 0.001519f
C5952 VDPWR.n338 VGND 0.005888f
C5953 VDPWR.n339 VGND 0.004416f
C5954 VDPWR.n340 VGND 0.00224f
C5955 VDPWR.t596 VGND 0.064097f
C5956 VDPWR.t435 VGND 0.039378f
C5957 VDPWR.t233 VGND 0.016158f
C5958 VDPWR.t237 VGND 0.022364f
C5959 VDPWR.t814 VGND 0.016158f
C5960 VDPWR.t1045 VGND 0.022364f
C5961 VDPWR.t1098 VGND 0.016158f
C5962 VDPWR.t1096 VGND 0.024184f
C5963 VDPWR.n341 VGND 0.026472f
C5964 VDPWR.n342 VGND 0.012237f
C5965 VDPWR.n343 VGND 0.005471f
C5966 VDPWR.t598 VGND 0.004984f
C5967 VDPWR.n344 VGND 0.008777f
C5968 VDPWR.n345 VGND 0.014953f
C5969 VDPWR.n346 VGND 0.002976f
C5970 VDPWR.n347 VGND 0.027044f
C5971 VDPWR.n348 VGND 0.026223f
C5972 VDPWR.n349 VGND 6.08e-19
C5973 VDPWR.t1011 VGND 0.007136f
C5974 VDPWR.n350 VGND 0.013312f
C5975 VDPWR.t850 VGND 0.007172f
C5976 VDPWR.n351 VGND 0.008357f
C5977 VDPWR.t105 VGND 0.002363f
C5978 VDPWR.t111 VGND 0.006281f
C5979 VDPWR.n352 VGND 0.003563f
C5980 VDPWR.t852 VGND 0.007041f
C5981 VDPWR.n353 VGND 0.007429f
C5982 VDPWR.n354 VGND 0.009555f
C5983 VDPWR.n355 VGND 0.001258f
C5984 VDPWR.n356 VGND 0.005888f
C5985 VDPWR.n357 VGND 0.003488f
C5986 VDPWR.n358 VGND 0.002016f
C5987 VDPWR.n359 VGND 0.00224f
C5988 VDPWR.n360 VGND 0.012275f
C5989 VDPWR.n361 VGND 0.032875f
C5990 VDPWR.t108 VGND 0.006226f
C5991 VDPWR.t176 VGND 0.016226f
C5992 VDPWR.t178 VGND 0.018113f
C5993 VDPWR.t989 VGND 0.012641f
C5994 VDPWR.t1089 VGND 0.023585f
C5995 VDPWR.t70 VGND 0.033207f
C5996 VDPWR.t72 VGND 0.016226f
C5997 VDPWR.t188 VGND 0.012641f
C5998 VDPWR.t285 VGND 0.029245f
C5999 VDPWR.t539 VGND 0.020377f
C6000 VDPWR.t61 VGND 0.027547f
C6001 VDPWR.t764 VGND 0.02849f
C6002 VDPWR.n362 VGND 0.019402f
C6003 VDPWR.n363 VGND 0.005637f
C6004 VDPWR.n364 VGND 0.003862f
C6005 VDPWR.n365 VGND 0.009272f
C6006 VDPWR.n366 VGND 0.002696f
C6007 VDPWR.n367 VGND 0.005888f
C6008 VDPWR.n368 VGND 0.004416f
C6009 VDPWR.n369 VGND 0.002625f
C6010 VDPWR.n370 VGND 0.008924f
C6011 VDPWR.n371 VGND 0.006148f
C6012 VDPWR.n372 VGND 0.004064f
C6013 VDPWR.n373 VGND 0.011493f
C6014 VDPWR.n374 VGND 0.089674f
C6015 VDPWR.n375 VGND 0.05908f
C6016 VDPWR.n376 VGND 0.114583f
C6017 VDPWR.n377 VGND 0.318185f
C6018 VDPWR.n378 VGND 0.114492f
C6019 VDPWR.n379 VGND 0.056224f
C6020 VDPWR.n380 VGND 0.076648f
C6021 VDPWR.n381 VGND 0.056138f
C6022 VDPWR.n382 VGND 0.465708f
C6023 VDPWR.t772 VGND 0.619228f
C6024 VDPWR.n385 VGND 0.465708f
C6025 VDPWR.n386 VGND 0.055408f
C6026 VDPWR.n387 VGND 0.036337f
C6027 VDPWR.n388 VGND 0.073206f
C6028 VDPWR.n389 VGND 0.038046f
C6029 VDPWR.n390 VGND 0.114492f
C6030 VDPWR.n391 VGND 0.056224f
C6031 VDPWR.n392 VGND 0.076648f
C6032 VDPWR.n393 VGND 0.056138f
C6033 VDPWR.n394 VGND 0.465708f
C6034 VDPWR.t119 VGND 0.619228f
C6035 VDPWR.n397 VGND 0.465708f
C6036 VDPWR.n398 VGND 0.055408f
C6037 VDPWR.n399 VGND 0.036337f
C6038 VDPWR.n400 VGND 0.073206f
C6039 VDPWR.n401 VGND 0.071425f
C6040 VDPWR.n402 VGND 0.171041f
C6041 VDPWR.n403 VGND 0.073588f
C6042 VDPWR.n404 VGND 0.035269f
C6043 VDPWR.n405 VGND 0.114487f
C6044 VDPWR.n406 VGND 0.055474f
C6045 VDPWR.n407 VGND 0.055474f
C6046 VDPWR.n408 VGND 0.055293f
C6047 VDPWR.n409 VGND 0.076656f
C6048 VDPWR.n410 VGND 0.247132f
C6049 VDPWR.t345 VGND 0.356671f
C6050 VDPWR.n411 VGND 0.344366f
C6051 VDPWR.t1037 VGND 0.356671f
C6052 VDPWR.n412 VGND 0.247132f
C6053 VDPWR.n413 VGND 2.15e-19
C6054 VDPWR.n414 VGND 0.025894f
C6055 VDPWR.n415 VGND 0.035269f
C6056 VDPWR.n416 VGND 0.076656f
C6057 VDPWR.n417 VGND 0.247132f
C6058 VDPWR.n418 VGND 2.38e-19
C6059 VDPWR.n419 VGND 0.247132f
C6060 VDPWR.t958 VGND 0.356671f
C6061 VDPWR.t959 VGND 0.356671f
C6062 VDPWR.n420 VGND 0.055293f
C6063 VDPWR.n421 VGND 0.055474f
C6064 VDPWR.n422 VGND 0.344366f
C6065 VDPWR.n423 VGND 0.055474f
C6066 VDPWR.n424 VGND 0.114487f
C6067 VDPWR.n425 VGND 0.060635f
C6068 VDPWR.n426 VGND 0.018181f
C6069 VDPWR.n427 VGND 0.029454f
C6070 VDPWR.n428 VGND 0.073168f
C6071 VDPWR.n429 VGND 0.084539f
C6072 VDPWR.n430 VGND 0.035235f
C6073 VDPWR.n431 VGND 0.114487f
C6074 VDPWR.n432 VGND 0.00445f
C6075 VDPWR.n433 VGND 0.055474f
C6076 VDPWR.n434 VGND 0.055474f
C6077 VDPWR.n435 VGND 0.055293f
C6078 VDPWR.n436 VGND 0.076656f
C6079 VDPWR.n437 VGND 0.247132f
C6080 VDPWR.t120 VGND 0.356671f
C6081 VDPWR.n438 VGND 0.344366f
C6082 VDPWR.t123 VGND 0.356671f
C6083 VDPWR.n439 VGND 0.247132f
C6084 VDPWR.n440 VGND 0.002025f
C6085 VDPWR.n441 VGND 0.060694f
C6086 VDPWR.n442 VGND 0.018181f
C6087 VDPWR.n443 VGND 0.029169f
C6088 VDPWR.n444 VGND 0.067579f
C6089 VDPWR.n445 VGND 0.082325f
C6090 VDPWR.n446 VGND 0.035121f
C6091 VDPWR.n447 VGND 0.114487f
C6092 VDPWR.n448 VGND 0.004458f
C6093 VDPWR.n449 VGND 0.055474f
C6094 VDPWR.n450 VGND 0.055474f
C6095 VDPWR.n451 VGND 0.055293f
C6096 VDPWR.n452 VGND 0.076656f
C6097 VDPWR.n453 VGND 0.247132f
C6098 VDPWR.t68 VGND 0.356671f
C6099 VDPWR.n454 VGND 0.344366f
C6100 VDPWR.t69 VGND 0.356671f
C6101 VDPWR.n455 VGND 0.247132f
C6102 VDPWR.n456 VGND 0.002138f
C6103 VDPWR.n457 VGND 0.060694f
C6104 VDPWR.n458 VGND 0.018181f
C6105 VDPWR.n459 VGND 0.029169f
C6106 VDPWR.n460 VGND 0.065201f
C6107 VDPWR.n461 VGND 0.075229f
C6108 VDPWR.n462 VGND 0.006257f
C6109 VDPWR.n463 VGND 0.060659f
C6110 VDPWR.n464 VGND 0.018181f
C6111 VDPWR.n465 VGND 0.029431f
C6112 VDPWR.n466 VGND 0.064503f
C6113 VDPWR.n467 VGND 0.08621f
C6114 VDPWR.n468 VGND 0.035269f
C6115 VDPWR.n469 VGND 0.114487f
C6116 VDPWR.n470 VGND 0.055474f
C6117 VDPWR.n471 VGND 0.055474f
C6118 VDPWR.n472 VGND 0.055293f
C6119 VDPWR.n473 VGND 0.076656f
C6120 VDPWR.n474 VGND 0.247132f
C6121 VDPWR.t956 VGND 0.356671f
C6122 VDPWR.n475 VGND 0.344366f
C6123 VDPWR.t957 VGND 0.356671f
C6124 VDPWR.n476 VGND 0.247132f
C6125 VDPWR.n477 VGND 2.38e-19
C6126 VDPWR.n478 VGND 0.006274f
C6127 VDPWR.n479 VGND 0.060635f
C6128 VDPWR.n480 VGND 0.018181f
C6129 VDPWR.n481 VGND 0.029454f
C6130 VDPWR.n482 VGND 0.043811f
C6131 VDPWR.n483 VGND 0.106582f
C6132 VDPWR.n484 VGND 0.035235f
C6133 VDPWR.n485 VGND 0.114487f
C6134 VDPWR.n486 VGND 0.00445f
C6135 VDPWR.n487 VGND 0.055474f
C6136 VDPWR.n488 VGND 0.055474f
C6137 VDPWR.n489 VGND 0.055293f
C6138 VDPWR.n490 VGND 0.076656f
C6139 VDPWR.n491 VGND 0.247132f
C6140 VDPWR.t122 VGND 0.356671f
C6141 VDPWR.n492 VGND 0.344366f
C6142 VDPWR.t121 VGND 0.356671f
C6143 VDPWR.n493 VGND 0.247132f
C6144 VDPWR.n494 VGND 0.002025f
C6145 VDPWR.n495 VGND 0.060694f
C6146 VDPWR.n496 VGND 0.018181f
C6147 VDPWR.n497 VGND 0.029169f
C6148 VDPWR.n498 VGND 0.067579f
C6149 VDPWR.n499 VGND 0.082325f
C6150 VDPWR.n500 VGND 0.035121f
C6151 VDPWR.n501 VGND 0.114487f
C6152 VDPWR.n502 VGND 0.004458f
C6153 VDPWR.n503 VGND 0.055474f
C6154 VDPWR.n504 VGND 0.055474f
C6155 VDPWR.n505 VGND 0.055293f
C6156 VDPWR.n506 VGND 0.076656f
C6157 VDPWR.n507 VGND 0.247132f
C6158 VDPWR.t67 VGND 0.356671f
C6159 VDPWR.n508 VGND 0.344366f
C6160 VDPWR.t13 VGND 0.356671f
C6161 VDPWR.n509 VGND 0.247132f
C6162 VDPWR.n510 VGND 0.002138f
C6163 VDPWR.n511 VGND 0.060694f
C6164 VDPWR.n512 VGND 0.018181f
C6165 VDPWR.n513 VGND 0.029169f
C6166 VDPWR.n514 VGND 0.064853f
C6167 VDPWR.n515 VGND 0.086126f
C6168 VDPWR.n516 VGND 0.035269f
C6169 VDPWR.n517 VGND 0.114487f
C6170 VDPWR.n518 VGND 0.055474f
C6171 VDPWR.n519 VGND 0.055474f
C6172 VDPWR.n520 VGND 0.055293f
C6173 VDPWR.n521 VGND 0.076656f
C6174 VDPWR.n522 VGND 0.247132f
C6175 VDPWR.t1036 VGND 0.356671f
C6176 VDPWR.n523 VGND 0.344366f
C6177 VDPWR.t1035 VGND 0.356671f
C6178 VDPWR.n524 VGND 0.247132f
C6179 VDPWR.n525 VGND 2.15e-19
C6180 VDPWR.n526 VGND 0.006257f
C6181 VDPWR.n527 VGND 0.060659f
C6182 VDPWR.n528 VGND 0.018181f
C6183 VDPWR.n529 VGND 0.029432f
C6184 VDPWR.n530 VGND 0.108553f
C6185 VDPWR.n531 VGND 0.406145f
C6186 VDPWR.n532 VGND 1.02472f
C6187 VDPWR.t951 VGND 0.0028f
C6188 VDPWR.t1202 VGND 0.00165f
C6189 VDPWR.t942 VGND 0.0028f
C6190 VDPWR.t1193 VGND 0.00165f
C6191 VDPWR.n533 VGND 0.004698f
C6192 VDPWR.n534 VGND 0.006946f
C6193 VDPWR.n535 VGND 0.006899f
C6194 VDPWR.n536 VGND 0.002816f
C6195 VDPWR.n537 VGND 0.366828f
C6196 VDPWR.n538 VGND 0.003488f
C6197 VDPWR.t187 VGND 0.007172f
C6198 VDPWR.n539 VGND 0.007983f
C6199 VDPWR.t789 VGND 7.56e-19
C6200 VDPWR.t19 VGND 0.001148f
C6201 VDPWR.n540 VGND 0.001983f
C6202 VDPWR.t185 VGND 0.007175f
C6203 VDPWR.t1165 VGND 0.00704f
C6204 VDPWR.n541 VGND 0.006705f
C6205 VDPWR.n542 VGND 0.003488f
C6206 VDPWR.n543 VGND 0.003158f
C6207 VDPWR.t911 VGND 0.001036f
C6208 VDPWR.n544 VGND 0.00294f
C6209 VDPWR.t965 VGND 0.004259f
C6210 VDPWR.n545 VGND 0.00392f
C6211 VDPWR.n546 VGND 0.003499f
C6212 VDPWR.t1163 VGND 0.007175f
C6213 VDPWR.n547 VGND 5.76e-19
C6214 VDPWR.t146 VGND 0.003015f
C6215 VDPWR.t682 VGND 0.004984f
C6216 VDPWR.n548 VGND 0.004913f
C6217 VDPWR.n549 VGND 0.005888f
C6218 VDPWR.t1207 VGND 0.020799f
C6219 VDPWR.n550 VGND 0.018812f
C6220 VDPWR.t288 VGND 5.64e-19
C6221 VDPWR.t329 VGND 0.001513f
C6222 VDPWR.n551 VGND 0.006904f
C6223 VDPWR.n552 VGND 0.003647f
C6224 VDPWR.t683 VGND 0.004984f
C6225 VDPWR.n553 VGND 0.01361f
C6226 VDPWR.n554 VGND 0.010753f
C6227 VDPWR.n555 VGND 0.013967f
C6228 VDPWR.n556 VGND 0.008065f
C6229 VDPWR.n557 VGND 0.005888f
C6230 VDPWR.n558 VGND 0.004416f
C6231 VDPWR.n559 VGND 0.005354f
C6232 VDPWR.n560 VGND 0.006068f
C6233 VDPWR.n561 VGND 0.013691f
C6234 VDPWR.t28 VGND 0.014151f
C6235 VDPWR.n562 VGND 7.37e-19
C6236 VDPWR.n563 VGND 0.004416f
C6237 VDPWR.n564 VGND 0.00136f
C6238 VDPWR.t856 VGND 7.56e-19
C6239 VDPWR.t31 VGND 0.001148f
C6240 VDPWR.n565 VGND 0.001983f
C6241 VDPWR.n566 VGND 0.005856f
C6242 VDPWR.n567 VGND 0.003488f
C6243 VDPWR.t1261 VGND 0.020799f
C6244 VDPWR.n568 VGND 0.005184f
C6245 VDPWR.n569 VGND 0.003488f
C6246 VDPWR.t5 VGND 5.64e-19
C6247 VDPWR.t1034 VGND 0.001513f
C6248 VDPWR.n570 VGND 0.006904f
C6249 VDPWR.t1214 VGND 0.020799f
C6250 VDPWR.t1024 VGND 0.003047f
C6251 VDPWR.n571 VGND 0.009651f
C6252 VDPWR.n572 VGND 0.005344f
C6253 VDPWR.n573 VGND 0.002933f
C6254 VDPWR.t668 VGND 0.004984f
C6255 VDPWR.n574 VGND 0.004913f
C6256 VDPWR.n575 VGND 0.018812f
C6257 VDPWR.n576 VGND 0.008065f
C6258 VDPWR.n577 VGND 0.013967f
C6259 VDPWR.t1023 VGND 0.02849f
C6260 VDPWR.t1033 VGND 0.027547f
C6261 VDPWR.t667 VGND 0.020377f
C6262 VDPWR.t4 VGND 0.029245f
C6263 VDPWR.t971 VGND 0.02849f
C6264 VDPWR.t924 VGND 0.032453f
C6265 VDPWR.t30 VGND 0.023585f
C6266 VDPWR.t855 VGND 0.012641f
C6267 VDPWR.t979 VGND 0.005849f
C6268 VDPWR.t981 VGND 0.020566f
C6269 VDPWR.n578 VGND 0.026837f
C6270 VDPWR.t982 VGND 0.007137f
C6271 VDPWR.n579 VGND 0.002016f
C6272 VDPWR.n580 VGND 0.0024f
C6273 VDPWR.n581 VGND 0.018611f
C6274 VDPWR.n582 VGND 0.005471f
C6275 VDPWR.t669 VGND 0.004984f
C6276 VDPWR.n583 VGND 0.008777f
C6277 VDPWR.n584 VGND 0.010753f
C6278 VDPWR.n585 VGND 0.003648f
C6279 VDPWR.n586 VGND 0.02906f
C6280 VDPWR.n587 VGND 0.039529f
C6281 VDPWR.t700 VGND 0.004984f
C6282 VDPWR.n588 VGND 0.009746f
C6283 VDPWR.n589 VGND 0.018812f
C6284 VDPWR.n590 VGND 0.011593f
C6285 VDPWR.t944 VGND 0.007172f
C6286 VDPWR.n591 VGND 0.00838f
C6287 VDPWR.n592 VGND 0.003488f
C6288 VDPWR.n593 VGND 0.001519f
C6289 VDPWR.n594 VGND 0.001519f
C6290 VDPWR.n595 VGND 0.1025f
C6291 VDPWR.t517 VGND 0.004984f
C6292 VDPWR.n596 VGND 0.004913f
C6293 VDPWR.n597 VGND 0.005888f
C6294 VDPWR.t1205 VGND 0.020799f
C6295 VDPWR.n598 VGND 0.018812f
C6296 VDPWR.n599 VGND 0.003647f
C6297 VDPWR.t518 VGND 0.004984f
C6298 VDPWR.n600 VGND 0.01361f
C6299 VDPWR.n601 VGND 0.014953f
C6300 VDPWR.n602 VGND 0.011593f
C6301 VDPWR.n603 VGND 0.005888f
C6302 VDPWR.n604 VGND 0.004416f
C6303 VDPWR.n605 VGND 0.005604f
C6304 VDPWR.t58 VGND 0.007175f
C6305 VDPWR.n606 VGND 0.009278f
C6306 VDPWR.n607 VGND 0.003488f
C6307 VDPWR.n608 VGND 0.005888f
C6308 VDPWR.n609 VGND 0.004416f
C6309 VDPWR.t854 VGND 0.007172f
C6310 VDPWR.n610 VGND 0.00847f
C6311 VDPWR.t115 VGND 0.007175f
C6312 VDPWR.n611 VGND 0.009165f
C6313 VDPWR.n612 VGND 0.003488f
C6314 VDPWR.n613 VGND 0.005888f
C6315 VDPWR.n614 VGND 0.004416f
C6316 VDPWR.t117 VGND 0.007172f
C6317 VDPWR.n615 VGND 0.00847f
C6318 VDPWR.t953 VGND 0.007175f
C6319 VDPWR.n616 VGND 0.009165f
C6320 VDPWR.n617 VGND 0.001519f
C6321 VDPWR.n618 VGND 0.005888f
C6322 VDPWR.n619 VGND 0.004416f
C6323 VDPWR.n620 VGND 0.00224f
C6324 VDPWR.t699 VGND 0.064097f
C6325 VDPWR.t516 VGND 0.039378f
C6326 VDPWR.t57 VGND 0.016158f
C6327 VDPWR.t853 VGND 0.022364f
C6328 VDPWR.t114 VGND 0.016158f
C6329 VDPWR.t116 VGND 0.022364f
C6330 VDPWR.t952 VGND 0.016158f
C6331 VDPWR.t943 VGND 0.024184f
C6332 VDPWR.n621 VGND 0.026472f
C6333 VDPWR.n622 VGND 0.012237f
C6334 VDPWR.n623 VGND 0.005471f
C6335 VDPWR.t701 VGND 0.004984f
C6336 VDPWR.n624 VGND 0.008777f
C6337 VDPWR.n625 VGND 0.014953f
C6338 VDPWR.n626 VGND 0.002976f
C6339 VDPWR.n627 VGND 0.027044f
C6340 VDPWR.n628 VGND 0.026223f
C6341 VDPWR.n629 VGND 6.08e-19
C6342 VDPWR.t980 VGND 0.007136f
C6343 VDPWR.n630 VGND 0.013312f
C6344 VDPWR.t970 VGND 0.007172f
C6345 VDPWR.n631 VGND 0.008357f
C6346 VDPWR.t925 VGND 0.002363f
C6347 VDPWR.t29 VGND 0.006281f
C6348 VDPWR.n632 VGND 0.003563f
C6349 VDPWR.t972 VGND 0.007041f
C6350 VDPWR.n633 VGND 0.007429f
C6351 VDPWR.n634 VGND 0.009555f
C6352 VDPWR.n635 VGND 0.001258f
C6353 VDPWR.n636 VGND 0.005888f
C6354 VDPWR.n637 VGND 0.003488f
C6355 VDPWR.n638 VGND 0.002016f
C6356 VDPWR.n639 VGND 0.00224f
C6357 VDPWR.n640 VGND 0.012275f
C6358 VDPWR.n641 VGND 0.032875f
C6359 VDPWR.t788 VGND 0.006226f
C6360 VDPWR.t186 VGND 0.016226f
C6361 VDPWR.t184 VGND 0.018113f
C6362 VDPWR.t18 VGND 0.012641f
C6363 VDPWR.t910 VGND 0.023585f
C6364 VDPWR.t1164 VGND 0.033207f
C6365 VDPWR.t1162 VGND 0.016226f
C6366 VDPWR.t964 VGND 0.012641f
C6367 VDPWR.t287 VGND 0.029245f
C6368 VDPWR.t681 VGND 0.020377f
C6369 VDPWR.t328 VGND 0.027547f
C6370 VDPWR.t145 VGND 0.02849f
C6371 VDPWR.n642 VGND 0.019402f
C6372 VDPWR.n643 VGND 0.005637f
C6373 VDPWR.n644 VGND 0.003862f
C6374 VDPWR.n645 VGND 0.009272f
C6375 VDPWR.n646 VGND 0.002696f
C6376 VDPWR.n647 VGND 0.005888f
C6377 VDPWR.n648 VGND 0.004416f
C6378 VDPWR.n649 VGND 0.002625f
C6379 VDPWR.n650 VGND 0.008924f
C6380 VDPWR.n651 VGND 0.006148f
C6381 VDPWR.n652 VGND 0.004064f
C6382 VDPWR.n653 VGND 0.011493f
C6383 VDPWR.n654 VGND 0.0731f
C6384 VDPWR.n655 VGND 0.037381f
C6385 VDPWR.n656 VGND 0.117598f
C6386 VDPWR.n657 VGND 0.025894f
C6387 VDPWR.n658 VGND 0.035269f
C6388 VDPWR.n659 VGND 0.076656f
C6389 VDPWR.n660 VGND 0.247132f
C6390 VDPWR.n661 VGND 2.38e-19
C6391 VDPWR.n662 VGND 0.247132f
C6392 VDPWR.t763 VGND 0.356671f
C6393 VDPWR.t762 VGND 0.356671f
C6394 VDPWR.n663 VGND 0.055293f
C6395 VDPWR.n664 VGND 0.055474f
C6396 VDPWR.n665 VGND 0.344366f
C6397 VDPWR.n666 VGND 0.055474f
C6398 VDPWR.n667 VGND 0.114487f
C6399 VDPWR.n668 VGND 0.060635f
C6400 VDPWR.n669 VGND 0.018181f
C6401 VDPWR.n670 VGND 0.029454f
C6402 VDPWR.n671 VGND 0.073168f
C6403 VDPWR.n672 VGND 0.084539f
C6404 VDPWR.n673 VGND 0.035235f
C6405 VDPWR.n674 VGND 0.114487f
C6406 VDPWR.n675 VGND 0.00445f
C6407 VDPWR.n676 VGND 0.055474f
C6408 VDPWR.n677 VGND 0.055474f
C6409 VDPWR.n678 VGND 0.055293f
C6410 VDPWR.n679 VGND 0.076656f
C6411 VDPWR.n680 VGND 0.247132f
C6412 VDPWR.t281 VGND 0.356671f
C6413 VDPWR.n681 VGND 0.344366f
C6414 VDPWR.t282 VGND 0.356671f
C6415 VDPWR.n682 VGND 0.247132f
C6416 VDPWR.n683 VGND 0.002025f
C6417 VDPWR.n684 VGND 0.060694f
C6418 VDPWR.n685 VGND 0.018181f
C6419 VDPWR.n686 VGND 0.029169f
C6420 VDPWR.n687 VGND 0.067579f
C6421 VDPWR.n688 VGND 0.082325f
C6422 VDPWR.n689 VGND 0.035121f
C6423 VDPWR.n690 VGND 0.114487f
C6424 VDPWR.n691 VGND 0.004458f
C6425 VDPWR.n692 VGND 0.055474f
C6426 VDPWR.n693 VGND 0.055474f
C6427 VDPWR.n694 VGND 0.055293f
C6428 VDPWR.n695 VGND 0.076656f
C6429 VDPWR.n696 VGND 0.247132f
C6430 VDPWR.t760 VGND 0.356671f
C6431 VDPWR.n697 VGND 0.344366f
C6432 VDPWR.t761 VGND 0.356671f
C6433 VDPWR.n698 VGND 0.247132f
C6434 VDPWR.n699 VGND 0.002138f
C6435 VDPWR.n700 VGND 0.060694f
C6436 VDPWR.n701 VGND 0.018181f
C6437 VDPWR.n702 VGND 0.029169f
C6438 VDPWR.n703 VGND 0.064853f
C6439 VDPWR.n704 VGND 0.086053f
C6440 VDPWR.n705 VGND 0.035269f
C6441 VDPWR.n706 VGND 0.114487f
C6442 VDPWR.n707 VGND 0.055474f
C6443 VDPWR.n708 VGND 0.055474f
C6444 VDPWR.n709 VGND 0.055293f
C6445 VDPWR.n710 VGND 0.076656f
C6446 VDPWR.n711 VGND 0.247132f
C6447 VDPWR.t315 VGND 0.356671f
C6448 VDPWR.n712 VGND 0.344366f
C6449 VDPWR.t314 VGND 0.356671f
C6450 VDPWR.n713 VGND 0.247132f
C6451 VDPWR.n714 VGND 2.15e-19
C6452 VDPWR.n715 VGND 0.006257f
C6453 VDPWR.n716 VGND 0.060659f
C6454 VDPWR.n717 VGND 0.018181f
C6455 VDPWR.n718 VGND 0.029432f
C6456 VDPWR.n719 VGND 0.059483f
C6457 VDPWR.n720 VGND 0.358402f
C6458 VDPWR.n721 VGND 5.33642f
C6459 VDPWR.t373 VGND 0.120007f
C6460 VDPWR.t340 VGND 0.074568f
C6461 VDPWR.t822 VGND 0.019801f
C6462 VDPWR.t219 VGND 0.019801f
C6463 VDPWR.n722 VGND 0.047461f
C6464 VDPWR.n723 VGND 0.423604f
C6465 VDPWR.t344 VGND 0.07455f
C6466 VDPWR.t824 VGND 0.019801f
C6467 VDPWR.t820 VGND 0.019801f
C6468 VDPWR.n724 VGND 0.047461f
C6469 VDPWR.n725 VGND 0.413821f
C6470 VDPWR.t253 VGND 0.019801f
C6471 VDPWR.t342 VGND 0.019801f
C6472 VDPWR.n726 VGND 0.047461f
C6473 VDPWR.n727 VGND 0.158951f
C6474 VDPWR.n728 VGND 0.064745f
C6475 VDPWR.n729 VGND 0.023069f
C6476 VDPWR.n730 VGND 0.03559f
C6477 VDPWR.n731 VGND 0.03559f
C6478 VDPWR.n732 VGND 0.03559f
C6479 VDPWR.n733 VGND 0.034528f
C6480 VDPWR.n734 VGND 0.218283f
C6481 VDPWR.t339 VGND 0.209454f
C6482 VDPWR.t821 VGND 0.143241f
C6483 VDPWR.t218 VGND 0.143241f
C6484 VDPWR.t252 VGND 0.107431f
C6485 VDPWR.n735 VGND 0.071621f
C6486 VDPWR.t341 VGND 0.107431f
C6487 VDPWR.t823 VGND 0.143241f
C6488 VDPWR.t819 VGND 0.143241f
C6489 VDPWR.t343 VGND 0.209454f
C6490 VDPWR.n736 VGND 0.218283f
C6491 VDPWR.n737 VGND 0.034517f
C6492 VDPWR.n738 VGND 0.023068f
C6493 VDPWR.n739 VGND 0.302545f
C6494 VDPWR.n740 VGND 0.014605f
C6495 VDPWR.n741 VGND 0.02803f
C6496 VDPWR.n742 VGND 0.02803f
C6497 VDPWR.t372 VGND 0.269964f
C6498 VDPWR.n743 VGND 0.027307f
C6499 VDPWR.n745 VGND 0.207311f
C6500 VDPWR.n746 VGND 0.02803f
C6501 VDPWR.n748 VGND 0.207311f
C6502 VDPWR.n749 VGND 0.027294f
C6503 VDPWR.n750 VGND 0.014601f
C6504 VDPWR.n751 VGND 0.170811f
C6505 VDPWR.n752 VGND 0.317852f
C6506 VDPWR.n753 VGND 0.465132f
C6507 VDPWR.n754 VGND 0.951569f
C6508 VDPWR.n755 VGND 1.09773f
C6509 VDPWR.n756 VGND 4.26152f
C6510 VDPWR.n757 VGND 3.16295f
C6511 VDPWR.n758 VGND 1.27886f
C6512 VDPWR.n759 VGND 0.16157f
C6513 VDPWR.n760 VGND 0.035269f
C6514 VDPWR.n761 VGND 0.114487f
C6515 VDPWR.n762 VGND 0.055474f
C6516 VDPWR.n763 VGND 0.055474f
C6517 VDPWR.n764 VGND 0.055293f
C6518 VDPWR.n765 VGND 0.076656f
C6519 VDPWR.n766 VGND 0.247132f
C6520 VDPWR.t1012 VGND 0.356671f
C6521 VDPWR.n767 VGND 0.344366f
C6522 VDPWR.t118 VGND 0.356671f
C6523 VDPWR.n768 VGND 0.247132f
C6524 VDPWR.n769 VGND 2.15e-19
C6525 VDPWR.n770 VGND 0.348256f
C6526 VDPWR.n771 VGND 0.012843f
C6527 VDPWR.n772 VGND 0.003054f
C6528 VDPWR.n773 VGND 0.001579f
C6529 VDPWR.n774 VGND 0.001579f
C6530 VDPWR.n775 VGND 0.116061f
C6531 VDPWR.n776 VGND 0.281618f
C6532 VDPWR.n777 VGND 0.096641f
C6533 VDPWR.n778 VGND 0.219213f
C6534 VDPWR.n779 VGND 0.281574f
C6535 VDPWR.n780 VGND 0.060111f
C6536 VDPWR.n781 VGND 0.096641f
C6537 VDPWR.n782 VGND 0.107527f
C6538 VDPWR.n783 VGND 0.001579f
C6539 VDPWR.n784 VGND 0.003054f
C6540 VDPWR.n785 VGND 0.003054f
C6541 VDPWR.n786 VGND 0.001973f
C6542 VDPWR.n787 VGND 0.002048f
C6543 VDPWR.n788 VGND 5.48e-19
C6544 VDPWR.t871 VGND 0.003019f
C6545 VDPWR.n789 VGND 0.006163f
C6546 VDPWR.n790 VGND 0.00224f
C6547 VDPWR.t531 VGND 0.052075f
C6548 VDPWR.t78 VGND 0.028868f
C6549 VDPWR.t938 VGND 0.022453f
C6550 VDPWR.t542 VGND 0.029245f
C6551 VDPWR.t962 VGND 0.03434f
C6552 VDPWR.t757 VGND 0.022453f
C6553 VDPWR.t507 VGND 0.029245f
C6554 VDPWR.t471 VGND 0.031509f
C6555 VDPWR.t248 VGND 0.033585f
C6556 VDPWR.t1146 VGND 0.02283f
C6557 VDPWR.t38 VGND 0.041132f
C6558 VDPWR.t265 VGND 0.016604f
C6559 VDPWR.t874 VGND 0.010566f
C6560 VDPWR.t966 VGND 0.017358f
C6561 VDPWR.t128 VGND 0.055283f
C6562 VDPWR.t998 VGND 0.060189f
C6563 VDPWR.t627 VGND 0.020377f
C6564 VDPWR.t916 VGND 0.027547f
C6565 VDPWR.t868 VGND 0.02849f
C6566 VDPWR.n791 VGND 0.038158f
C6567 VDPWR.t628 VGND 0.004984f
C6568 VDPWR.n792 VGND 0.008777f
C6569 VDPWR.t869 VGND 0.003019f
C6570 VDPWR.t1198 VGND 0.036876f
C6571 VDPWR.n793 VGND 0.011929f
C6572 VDPWR.n794 VGND 0.004416f
C6573 VDPWR.t999 VGND 5.64e-19
C6574 VDPWR.t917 VGND 0.001513f
C6575 VDPWR.n795 VGND 0.006904f
C6576 VDPWR.n796 VGND 0.013967f
C6577 VDPWR.t129 VGND 0.007511f
C6578 VDPWR.n797 VGND 0.016861f
C6579 VDPWR.t629 VGND 0.004984f
C6580 VDPWR.n798 VGND 0.004829f
C6581 VDPWR.t875 VGND 0.001527f
C6582 VDPWR.t39 VGND 0.001527f
C6583 VDPWR.n799 VGND 0.003322f
C6584 VDPWR.n800 VGND 0.007816f
C6585 VDPWR.n801 VGND 0.002048f
C6586 VDPWR.n802 VGND 0.001973f
C6587 VDPWR.n803 VGND 0.001579f
C6588 VDPWR.n804 VGND 0.003054f
C6589 VDPWR.n805 VGND 0.001973f
C6590 VDPWR.n806 VGND 0.002949f
C6591 VDPWR.t266 VGND 0.007332f
C6592 VDPWR.n807 VGND 0.005407f
C6593 VDPWR.n808 VGND 0.001734f
C6594 VDPWR.n809 VGND 0.001472f
C6595 VDPWR.n810 VGND 0.001472f
C6596 VDPWR.n811 VGND 8.32e-19
C6597 VDPWR.n812 VGND 0.001599f
C6598 VDPWR.t1147 VGND 0.001372f
C6599 VDPWR.t249 VGND 0.002267f
C6600 VDPWR.n813 VGND 0.006267f
C6601 VDPWR.n814 VGND 0.008122f
C6602 VDPWR.t1259 VGND 0.029301f
C6603 VDPWR.n815 VGND 0.015457f
C6604 VDPWR.n816 VGND 0.003488f
C6605 VDPWR.t508 VGND 0.005024f
C6606 VDPWR.t1265 VGND 0.010664f
C6607 VDPWR.n818 VGND 0.027341f
C6608 VDPWR.t509 VGND 0.005024f
C6609 VDPWR.n819 VGND 0.013522f
C6610 VDPWR.t543 VGND 0.005019f
C6611 VDPWR.n820 VGND 0.002332f
C6612 VDPWR.t758 VGND 0.001527f
C6613 VDPWR.t963 VGND 0.001527f
C6614 VDPWR.n821 VGND 0.003322f
C6615 VDPWR.n822 VGND 0.011761f
C6616 VDPWR.t1245 VGND 0.03788f
C6617 VDPWR.n823 VGND 0.06464f
C6618 VDPWR.n824 VGND 0.019984f
C6619 VDPWR.t939 VGND 0.001527f
C6620 VDPWR.t79 VGND 0.001527f
C6621 VDPWR.n825 VGND 0.003322f
C6622 VDPWR.n826 VGND 0.021375f
C6623 VDPWR.n827 VGND 7.36e-19
C6624 VDPWR.n828 VGND 0.001973f
C6625 VDPWR.n829 VGND 0.002944f
C6626 VDPWR.t544 VGND 0.004984f
C6627 VDPWR.n830 VGND 0.008777f
C6628 VDPWR.n831 VGND 0.005471f
C6629 VDPWR.t532 VGND 0.005024f
C6630 VDPWR.t1248 VGND 0.010664f
C6631 VDPWR.n833 VGND 0.027341f
C6632 VDPWR.t533 VGND 0.005024f
C6633 VDPWR.n834 VGND 0.014893f
C6634 VDPWR.n835 VGND 0.002048f
C6635 VDPWR.t656 VGND 0.005024f
C6636 VDPWR.t1185 VGND 0.010664f
C6637 VDPWR.n837 VGND 0.027341f
C6638 VDPWR.t657 VGND 0.005024f
C6639 VDPWR.n838 VGND 0.014893f
C6640 VDPWR.n839 VGND 0.001973f
C6641 VDPWR.n840 VGND 0.002112f
C6642 VDPWR.n841 VGND 0.002885f
C6643 VDPWR.n842 VGND 0.001376f
C6644 VDPWR.n843 VGND 0.012553f
C6645 VDPWR.n844 VGND 0.002048f
C6646 VDPWR.n845 VGND 0.001472f
C6647 VDPWR.n846 VGND 0.001973f
C6648 VDPWR.n847 VGND 0.003054f
C6649 VDPWR.n848 VGND 0.002949f
C6650 VDPWR.n849 VGND 0.005152f
C6651 VDPWR.n850 VGND 0.002016f
C6652 VDPWR.n851 VGND 0.015457f
C6653 VDPWR.n852 VGND 0.012685f
C6654 VDPWR.n853 VGND 0.00224f
C6655 VDPWR.n854 VGND 0.006234f
C6656 VDPWR.n855 VGND 0.002016f
C6657 VDPWR.n856 VGND 0.00475f
C6658 VDPWR.t473 VGND 0.005064f
C6659 VDPWR.n857 VGND 0.007505f
C6660 VDPWR.n858 VGND 0.018913f
C6661 VDPWR.n859 VGND 0.020217f
C6662 VDPWR.n860 VGND 0.005888f
C6663 VDPWR.n861 VGND 0.004416f
C6664 VDPWR.n862 VGND 0.0024f
C6665 VDPWR.n863 VGND 0.039775f
C6666 VDPWR.t472 VGND 0.004984f
C6667 VDPWR.n864 VGND 0.008777f
C6668 VDPWR.n865 VGND 0.002829f
C6669 VDPWR.n866 VGND 0.002048f
C6670 VDPWR.n867 VGND 0.001472f
C6671 VDPWR.n868 VGND 0.001973f
C6672 VDPWR.n869 VGND 0.001579f
C6673 VDPWR.n870 VGND 0.128008f
C6674 VDPWR.n871 VGND 0.281618f
C6675 VDPWR.n872 VGND 0.128862f
C6676 VDPWR.n873 VGND 0.003404f
C6677 VDPWR.n874 VGND 0.00352f
C6678 VDPWR.n875 VGND 0.002757f
C6679 VDPWR.n876 VGND 0.001579f
C6680 VDPWR.n877 VGND 0.002944f
C6681 VDPWR.t1270 VGND 0.020799f
C6682 VDPWR.n878 VGND 0.015788f
C6683 VDPWR.t915 VGND 0.003019f
C6684 VDPWR.n879 VGND 0.012345f
C6685 VDPWR.n880 VGND 0.002048f
C6686 VDPWR.n881 VGND 0.001973f
C6687 VDPWR.n882 VGND 0.00352f
C6688 VDPWR.n883 VGND 0.001579f
C6689 VDPWR.t485 VGND 0.004984f
C6690 VDPWR.n884 VGND 0.004325f
C6691 VDPWR.n885 VGND 0.005471f
C6692 VDPWR.t426 VGND 0.052075f
C6693 VDPWR.t876 VGND 0.028868f
C6694 VDPWR.t967 VGND 0.019245f
C6695 VDPWR.t553 VGND 0.017547f
C6696 VDPWR.t392 VGND 0.024906f
C6697 VDPWR.t974 VGND 0.039811f
C6698 VDPWR.t9 VGND 0.009057f
C6699 VDPWR.t1015 VGND 0.016038f
C6700 VDPWR.t294 VGND 0.015849f
C6701 VDPWR.t334 VGND 0.017924f
C6702 VDPWR.t973 VGND 0.035472f
C6703 VDPWR.t250 VGND 0.019434f
C6704 VDPWR.t890 VGND 0.016038f
C6705 VDPWR.t338 VGND 0.024906f
C6706 VDPWR.t271 VGND 0.017924f
C6707 VDPWR.t333 VGND 0.017924f
C6708 VDPWR.t976 VGND 0.019434f
C6709 VDPWR.t864 VGND 0.015849f
C6710 VDPWR.t293 VGND 0.024906f
C6711 VDPWR.t862 VGND 0.021509f
C6712 VDPWR.t212 VGND 0.017924f
C6713 VDPWR.t336 VGND 0.030566f
C6714 VDPWR.t337 VGND 0.024906f
C6715 VDPWR.t36 VGND 0.021509f
C6716 VDPWR.t204 VGND 0.015849f
C6717 VDPWR.t214 VGND 0.039623f
C6718 VDPWR.t269 VGND 0.038868f
C6719 VDPWR.t991 VGND 0.015849f
C6720 VDPWR.t202 VGND 0.035472f
C6721 VDPWR.t1150 VGND 0.025094f
C6722 VDPWR.t1027 VGND 0.020566f
C6723 VDPWR.t730 VGND 0.015849f
C6724 VDPWR.t326 VGND 0.024151f
C6725 VDPWR.t771 VGND 0.023208f
C6726 VDPWR.n886 VGND 0.020611f
C6727 VDPWR.t327 VGND 0.0018f
C6728 VDPWR.t1028 VGND 0.0018f
C6729 VDPWR.n887 VGND 0.003918f
C6730 VDPWR.n888 VGND 0.004957f
C6731 VDPWR.t731 VGND 0.005024f
C6732 VDPWR.t1180 VGND 0.010664f
C6733 VDPWR.n890 VGND 0.027341f
C6734 VDPWR.t732 VGND 0.005024f
C6735 VDPWR.n891 VGND 0.014893f
C6736 VDPWR.t1151 VGND 0.00632f
C6737 VDPWR.n892 VGND 0.001133f
C6738 VDPWR.t203 VGND 0.0018f
C6739 VDPWR.t270 VGND 0.0018f
C6740 VDPWR.n893 VGND 0.004032f
C6741 VDPWR.n894 VGND 0.00519f
C6742 VDPWR.n895 VGND 0.004416f
C6743 VDPWR.t205 VGND 0.002834f
C6744 VDPWR.t215 VGND 0.0018f
C6745 VDPWR.t37 VGND 0.0018f
C6746 VDPWR.n896 VGND 0.004032f
C6747 VDPWR.n897 VGND 0.00519f
C6748 VDPWR.n898 VGND 0.004672f
C6749 VDPWR.t213 VGND 0.002834f
C6750 VDPWR.t863 VGND 0.00135f
C6751 VDPWR.t865 VGND 0.002785f
C6752 VDPWR.n899 VGND 0.00567f
C6753 VDPWR.n900 VGND 0.004406f
C6754 VDPWR.n901 VGND 0.002949f
C6755 VDPWR.n902 VGND 0.002112f
C6756 VDPWR.n903 VGND 0.003083f
C6757 VDPWR.n904 VGND 0.001973f
C6758 VDPWR.n905 VGND 0.001579f
C6759 VDPWR.n906 VGND 0.001973f
C6760 VDPWR.n907 VGND 0.002048f
C6761 VDPWR.n908 VGND 0.005888f
C6762 VDPWR.n909 VGND 0.002944f
C6763 VDPWR.n910 VGND 0.002048f
C6764 VDPWR.n911 VGND 0.001598f
C6765 VDPWR.n912 VGND 0.002085f
C6766 VDPWR.t272 VGND 0.00135f
C6767 VDPWR.t891 VGND 0.002785f
C6768 VDPWR.n913 VGND 0.00567f
C6769 VDPWR.n914 VGND 0.005888f
C6770 VDPWR.t251 VGND 0.002776f
C6771 VDPWR.t335 VGND 0.001152f
C6772 VDPWR.t1016 VGND 0.001152f
C6773 VDPWR.n915 VGND 0.002399f
C6774 VDPWR.n916 VGND 0.006924f
C6775 VDPWR.t10 VGND 0.002776f
C6776 VDPWR.t554 VGND 0.004984f
C6777 VDPWR.n917 VGND 0.008777f
C6778 VDPWR.n918 VGND 0.003488f
C6779 VDPWR.t1250 VGND 0.029301f
C6780 VDPWR.t975 VGND 0.001152f
C6781 VDPWR.t393 VGND 0.001152f
C6782 VDPWR.n919 VGND 0.002373f
C6783 VDPWR.n920 VGND 0.014953f
C6784 VDPWR.n921 VGND 7.36e-19
C6785 VDPWR.n922 VGND 0.001973f
C6786 VDPWR.n923 VGND 0.116061f
C6787 VDPWR.n924 VGND 0.003404f
C6788 VDPWR.n925 VGND 0.003083f
C6789 VDPWR.n926 VGND 0.00352f
C6790 VDPWR.n927 VGND 0.001973f
C6791 VDPWR.n928 VGND 0.002048f
C6792 VDPWR.n929 VGND 0.007329f
C6793 VDPWR.t676 VGND 0.005024f
C6794 VDPWR.t1190 VGND 0.010664f
C6795 VDPWR.n931 VGND 0.027341f
C6796 VDPWR.t677 VGND 0.005024f
C6797 VDPWR.n932 VGND 0.014893f
C6798 VDPWR.n933 VGND 0.005888f
C6799 VDPWR.t1247 VGND 0.029301f
C6800 VDPWR.n934 VGND 0.044937f
C6801 VDPWR.n935 VGND 0.005445f
C6802 VDPWR.t154 VGND 0.001152f
C6803 VDPWR.t391 VGND 0.001152f
C6804 VDPWR.n936 VGND 0.002373f
C6805 VDPWR.n937 VGND 0.008042f
C6806 VDPWR.n938 VGND 0.0048f
C6807 VDPWR.t978 VGND 0.002755f
C6808 VDPWR.t716 VGND 0.005483f
C6809 VDPWR.n939 VGND 0.00426f
C6810 VDPWR.n940 VGND 0.002944f
C6811 VDPWR.n941 VGND 0.001973f
C6812 VDPWR.n942 VGND 0.00352f
C6813 VDPWR.n943 VGND 0.116061f
C6814 VDPWR.n944 VGND 0.00352f
C6815 VDPWR.n945 VGND 0.002949f
C6816 VDPWR.n946 VGND 0.001579f
C6817 VDPWR.n947 VGND 0.002048f
C6818 VDPWR.n948 VGND 0.005687f
C6819 VDPWR.n949 VGND 0.005888f
C6820 VDPWR.t1178 VGND 0.072626f
C6821 VDPWR.n950 VGND 0.033923f
C6822 VDPWR.n951 VGND 0.005888f
C6823 VDPWR.t813 VGND 0.00281f
C6824 VDPWR.t811 VGND 0.0018f
C6825 VDPWR.t158 VGND 0.0018f
C6826 VDPWR.n952 VGND 0.004032f
C6827 VDPWR.n953 VGND 0.007616f
C6828 VDPWR.n954 VGND 0.01243f
C6829 VDPWR.n955 VGND 0.002048f
C6830 VDPWR.n956 VGND 0.001973f
C6831 VDPWR.n957 VGND 0.00352f
C6832 VDPWR.n958 VGND 0.001579f
C6833 VDPWR.n959 VGND 0.002048f
C6834 VDPWR.n960 VGND 0.002944f
C6835 VDPWR.t1236 VGND 0.020799f
C6836 VDPWR.n961 VGND 0.007141f
C6837 VDPWR.t796 VGND 0.007646f
C6838 VDPWR.n962 VGND 0.011292f
C6839 VDPWR.n963 VGND 0.005888f
C6840 VDPWR.t54 VGND 0.0018f
C6841 VDPWR.t378 VGND 0.0018f
C6842 VDPWR.n964 VGND 0.004032f
C6843 VDPWR.t380 VGND 0.002834f
C6844 VDPWR.n965 VGND 0.006409f
C6845 VDPWR.n966 VGND 0.005344f
C6846 VDPWR.n967 VGND 0.001099f
C6847 VDPWR.n968 VGND 0.002949f
C6848 VDPWR.n969 VGND 0.002763f
C6849 VDPWR.n970 VGND 0.00288f
C6850 VDPWR.n971 VGND 0.001579f
C6851 VDPWR.n972 VGND 0.00352f
C6852 VDPWR.n973 VGND 0.116061f
C6853 VDPWR.n974 VGND 0.128008f
C6854 VDPWR.n975 VGND 0.00352f
C6855 VDPWR.n976 VGND 0.002949f
C6856 VDPWR.n977 VGND 0.001973f
C6857 VDPWR.n978 VGND 0.001579f
C6858 VDPWR.t1149 VGND 0.001148f
C6859 VDPWR.t367 VGND -7.28e-19
C6860 VDPWR.n979 VGND 0.007328f
C6861 VDPWR.n980 VGND 0.005643f
C6862 VDPWR.t1135 VGND 0.002776f
C6863 VDPWR.n981 VGND 0.001349f
C6864 VDPWR.n982 VGND 0.001151f
C6865 VDPWR.t1105 VGND 0.001867f
C6866 VDPWR.t1107 VGND 0.001867f
C6867 VDPWR.n983 VGND 0.003854f
C6868 VDPWR.n984 VGND 0.001131f
C6869 VDPWR.n985 VGND 0.002048f
C6870 VDPWR.n986 VGND 0.001973f
C6871 VDPWR.n987 VGND 0.00352f
C6872 VDPWR.n988 VGND 0.116061f
C6873 VDPWR.n989 VGND 0.128008f
C6874 VDPWR.n990 VGND 0.00352f
C6875 VDPWR.n991 VGND 0.002949f
C6876 VDPWR.n992 VGND 0.001579f
C6877 VDPWR.n993 VGND 0.002048f
C6878 VDPWR.n994 VGND 0.002944f
C6879 VDPWR.t1043 VGND 0.001036f
C6880 VDPWR.t226 VGND 0.001036f
C6881 VDPWR.n995 VGND 0.002169f
C6882 VDPWR.t1129 VGND 0.001867f
C6883 VDPWR.t1103 VGND 0.001867f
C6884 VDPWR.n996 VGND 0.003854f
C6885 VDPWR.t1121 VGND 0.0018f
C6886 VDPWR.t1125 VGND 0.001867f
C6887 VDPWR.n997 VGND 0.003787f
C6888 VDPWR.n998 VGND 0.005527f
C6889 VDPWR.n999 VGND 0.004432f
C6890 VDPWR.t1131 VGND 0.001867f
C6891 VDPWR.t1123 VGND 0.001867f
C6892 VDPWR.n1000 VGND 0.003881f
C6893 VDPWR.n1001 VGND 0.006736f
C6894 VDPWR.n1002 VGND 0.005888f
C6895 VDPWR.t1119 VGND 0.00659f
C6896 VDPWR.n1003 VGND 0.008378f
C6897 VDPWR.n1004 VGND 0.005344f
C6898 VDPWR.t901 VGND 0.001527f
C6899 VDPWR.t955 VGND 0.001527f
C6900 VDPWR.n1005 VGND 0.003322f
C6901 VDPWR.n1006 VGND 0.019777f
C6902 VDPWR.n1007 VGND 0.001973f
C6903 VDPWR.n1008 VGND 0.00352f
C6904 VDPWR.n1009 VGND 0.140809f
C6905 VDPWR.n1010 VGND 0.167264f
C6906 VDPWR.n1011 VGND 0.281618f
C6907 VDPWR.n1012 VGND 0.116061f
C6908 VDPWR.n1013 VGND 0.003404f
C6909 VDPWR.n1014 VGND 0.00352f
C6910 VDPWR.n1015 VGND 0.002757f
C6911 VDPWR.n1016 VGND 0.001579f
C6912 VDPWR.n1017 VGND 0.002944f
C6913 VDPWR.t1273 VGND 0.020799f
C6914 VDPWR.n1018 VGND 0.021306f
C6915 VDPWR.t729 VGND 0.004984f
C6916 VDPWR.n1019 VGND 0.011445f
C6917 VDPWR.n1020 VGND 0.002048f
C6918 VDPWR.n1021 VGND 0.001973f
C6919 VDPWR.n1022 VGND 0.00352f
C6920 VDPWR.n1023 VGND 0.001579f
C6921 VDPWR.t583 VGND 0.052075f
C6922 VDPWR.t696 VGND 0.085094f
C6923 VDPWR.t1081 VGND 0.069434f
C6924 VDPWR.t589 VGND 0.016226f
C6925 VDPWR.t1077 VGND 0.018868f
C6926 VDPWR.t1055 VGND 0.032453f
C6927 VDPWR.t1083 VGND 0.032453f
C6928 VDPWR.t1059 VGND 0.032453f
C6929 VDPWR.t1057 VGND 0.032453f
C6930 VDPWR.t1085 VGND 0.032453f
C6931 VDPWR.t1079 VGND 0.025849f
C6932 VDPWR.t1063 VGND 0.022642f
C6933 VDPWR.t1073 VGND 0.032453f
C6934 VDPWR.t1069 VGND 0.032453f
C6935 VDPWR.t1065 VGND 0.032453f
C6936 VDPWR.t1075 VGND 0.032453f
C6937 VDPWR.t1071 VGND 0.027358f
C6938 VDPWR.t630 VGND 0.016226f
C6939 VDPWR.t1067 VGND 0.021321f
C6940 VDPWR.t1061 VGND 0.032453f
C6941 VDPWR.t1154 VGND 0.032453f
C6942 VDPWR.t779 VGND 0.032453f
C6943 VDPWR.t1152 VGND 0.032453f
C6944 VDPWR.t1156 VGND 0.022264f
C6945 VDPWR.n1024 VGND 0.037412f
C6946 VDPWR.n1025 VGND 0.008952f
C6947 VDPWR.n1026 VGND 0.002791f
C6948 VDPWR.n1027 VGND 0.005888f
C6949 VDPWR.t1157 VGND 0.006898f
C6950 VDPWR.n1028 VGND 0.006782f
C6951 VDPWR.t631 VGND 0.005483f
C6952 VDPWR.n1029 VGND 0.004139f
C6953 VDPWR.t1153 VGND 0.001867f
C6954 VDPWR.t780 VGND 0.001867f
C6955 VDPWR.n1030 VGND 0.004011f
C6956 VDPWR.t1216 VGND 0.073477f
C6957 VDPWR.n1031 VGND 0.030131f
C6958 VDPWR.n1032 VGND 0.005888f
C6959 VDPWR.t1155 VGND 0.001867f
C6960 VDPWR.t1062 VGND 0.001867f
C6961 VDPWR.n1033 VGND 0.004002f
C6962 VDPWR.n1034 VGND 0.008485f
C6963 VDPWR.t1068 VGND 0.001867f
C6964 VDPWR.t1072 VGND 0.001867f
C6965 VDPWR.n1035 VGND 0.003854f
C6966 VDPWR.n1036 VGND 0.005775f
C6967 VDPWR.n1037 VGND 0.002949f
C6968 VDPWR.t1076 VGND 0.001867f
C6969 VDPWR.t1066 VGND 0.001867f
C6970 VDPWR.n1038 VGND 0.003854f
C6971 VDPWR.n1039 VGND 0.008648f
C6972 VDPWR.t1070 VGND 0.001867f
C6973 VDPWR.t1074 VGND 0.001867f
C6974 VDPWR.n1040 VGND 0.003854f
C6975 VDPWR.n1041 VGND 0.008648f
C6976 VDPWR.n1042 VGND 0.002112f
C6977 VDPWR.n1043 VGND 0.003083f
C6978 VDPWR.n1044 VGND 0.001973f
C6979 VDPWR.n1045 VGND 0.00352f
C6980 VDPWR.n1046 VGND 0.116061f
C6981 VDPWR.n1047 VGND 0.001579f
C6982 VDPWR.n1048 VGND 0.001973f
C6983 VDPWR.n1049 VGND 0.005888f
C6984 VDPWR.t1064 VGND 0.001867f
C6985 VDPWR.t1080 VGND 0.0018f
C6986 VDPWR.n1050 VGND 0.003797f
C6987 VDPWR.t632 VGND 0.005483f
C6988 VDPWR.n1051 VGND 0.004291f
C6989 VDPWR.n1052 VGND 0.005694f
C6990 VDPWR.n1053 VGND 0.002048f
C6991 VDPWR.n1054 VGND 0.002944f
C6992 VDPWR.n1055 VGND 0.001504f
C6993 VDPWR.n1056 VGND 0.001321f
C6994 VDPWR.n1057 VGND 0.006783f
C6995 VDPWR.t1086 VGND 0.001867f
C6996 VDPWR.t1058 VGND 0.001867f
C6997 VDPWR.n1058 VGND 0.003854f
C6998 VDPWR.n1059 VGND 0.003782f
C6999 VDPWR.n1060 VGND 0.005888f
C7000 VDPWR.t1230 VGND 0.072626f
C7001 VDPWR.t1060 VGND 0.001867f
C7002 VDPWR.t1084 VGND 0.001867f
C7003 VDPWR.n1061 VGND 0.003854f
C7004 VDPWR.n1062 VGND 0.00661f
C7005 VDPWR.n1063 VGND 0.033913f
C7006 VDPWR.t1056 VGND 0.001867f
C7007 VDPWR.t1078 VGND 0.001867f
C7008 VDPWR.n1064 VGND 0.003854f
C7009 VDPWR.t1082 VGND 0.006558f
C7010 VDPWR.n1065 VGND 0.009583f
C7011 VDPWR.t697 VGND 0.004984f
C7012 VDPWR.n1066 VGND 0.006247f
C7013 VDPWR.n1067 VGND 0.005696f
C7014 VDPWR.t1284 VGND 0.020799f
C7015 VDPWR.n1068 VGND 0.021306f
C7016 VDPWR.t698 VGND 0.004984f
C7017 VDPWR.t584 VGND 0.005024f
C7018 VDPWR.t1234 VGND 0.010664f
C7019 VDPWR.n1070 VGND 0.027341f
C7020 VDPWR.t585 VGND 0.005024f
C7021 VDPWR.n1071 VGND 0.014893f
C7022 VDPWR.t692 VGND 0.005024f
C7023 VDPWR.t1167 VGND 0.010664f
C7024 VDPWR.n1073 VGND 0.027341f
C7025 VDPWR.t693 VGND 0.005024f
C7026 VDPWR.n1074 VGND 0.014893f
C7027 VDPWR.n1075 VGND 0.012551f
C7028 VDPWR.n1076 VGND 0.002949f
C7029 VDPWR.n1077 VGND 0.002048f
C7030 VDPWR.n1078 VGND 0.003083f
C7031 VDPWR.n1079 VGND 0.001973f
C7032 VDPWR.n1080 VGND 0.003404f
C7033 VDPWR.n1081 VGND 0.001579f
C7034 VDPWR.n1082 VGND 0.001973f
C7035 VDPWR.n1083 VGND 0.002944f
C7036 VDPWR.n1084 VGND 0.002048f
C7037 VDPWR.n1085 VGND 0.002112f
C7038 VDPWR.n1086 VGND 0.001376f
C7039 VDPWR.n1087 VGND 0.002885f
C7040 VDPWR.n1088 VGND 0.003083f
C7041 VDPWR.n1089 VGND 0.140809f
C7042 VDPWR.n1090 VGND 0.532156f
C7043 VDPWR.n1091 VGND 0.140809f
C7044 VDPWR.n1092 VGND 0.003404f
C7045 VDPWR.n1093 VGND 0.00352f
C7046 VDPWR.n1094 VGND 0.002949f
C7047 VDPWR.n1095 VGND 0.001579f
C7048 VDPWR.n1096 VGND 0.002048f
C7049 VDPWR.n1097 VGND 0.00288f
C7050 VDPWR.t425 VGND 0.001867f
C7051 VDPWR.t397 VGND 0.001867f
C7052 VDPWR.n1098 VGND 0.003854f
C7053 VDPWR.t1283 VGND 0.072626f
C7054 VDPWR.t411 VGND 0.001867f
C7055 VDPWR.t421 VGND 0.001867f
C7056 VDPWR.n1099 VGND 0.003854f
C7057 VDPWR.n1100 VGND 0.008648f
C7058 VDPWR.n1101 VGND 0.005888f
C7059 VDPWR.t257 VGND 0.001867f
C7060 VDPWR.t417 VGND 0.001867f
C7061 VDPWR.n1102 VGND 0.004002f
C7062 VDPWR.n1103 VGND 0.005793f
C7063 VDPWR.t255 VGND 0.006898f
C7064 VDPWR.n1104 VGND 0.006887f
C7065 VDPWR.n1105 VGND 0.005836f
C7066 VDPWR.t1240 VGND 0.020636f
C7067 VDPWR.n1106 VGND 0.010252f
C7068 VDPWR.n1107 VGND 0.003941f
C7069 VDPWR.t563 VGND 0.004984f
C7070 VDPWR.n1108 VGND 0.002657f
C7071 VDPWR.t525 VGND 0.066226f
C7072 VDPWR.t678 VGND 0.055472f
C7073 VDPWR.t556 VGND 0.092264f
C7074 VDPWR.t492 VGND 0.063962f
C7075 VDPWR.t640 VGND 0.109622f
C7076 VDPWR.t704 VGND 0.098679f
C7077 VDPWR.t727 VGND 0.063962f
C7078 VDPWR.t736 VGND 0.040566f
C7079 VDPWR.t418 VGND 0.048868f
C7080 VDPWR.t414 VGND 0.032453f
C7081 VDPWR.t404 VGND 0.032453f
C7082 VDPWR.t408 VGND 0.032453f
C7083 VDPWR.t406 VGND 0.022453f
C7084 VDPWR.t412 VGND 0.026226f
C7085 VDPWR.t402 VGND 0.032453f
C7086 VDPWR.t398 VGND 0.032264f
C7087 VDPWR.t394 VGND 0.032264f
C7088 VDPWR.t422 VGND 0.032453f
C7089 VDPWR.t400 VGND 0.023962f
C7090 VDPWR.t432 VGND 0.016226f
C7091 VDPWR.t396 VGND 0.024717f
C7092 VDPWR.t424 VGND 0.032453f
C7093 VDPWR.t420 VGND 0.032453f
C7094 VDPWR.t410 VGND 0.032453f
C7095 VDPWR.t416 VGND 0.032453f
C7096 VDPWR.t256 VGND 0.032453f
C7097 VDPWR.t258 VGND 0.02f
C7098 VDPWR.t1019 VGND 0.028679f
C7099 VDPWR.t254 VGND 0.016792f
C7100 VDPWR.t562 VGND 0.006038f
C7101 VDPWR.n1109 VGND 0.037412f
C7102 VDPWR.n1110 VGND 0.017118f
C7103 VDPWR.n1111 VGND 0.002949f
C7104 VDPWR.n1112 VGND 0.012758f
C7105 VDPWR.n1113 VGND 0.002048f
C7106 VDPWR.n1114 VGND 0.001579f
C7107 VDPWR.n1115 VGND 0.00352f
C7108 VDPWR.n1116 VGND 0.116061f
C7109 VDPWR.n1117 VGND 0.003404f
C7110 VDPWR.n1118 VGND 0.00352f
C7111 VDPWR.n1119 VGND 0.002949f
C7112 VDPWR.n1120 VGND 0.001579f
C7113 VDPWR.n1121 VGND 0.002048f
C7114 VDPWR.n1122 VGND 0.002048f
C7115 VDPWR.n1123 VGND 0.003083f
C7116 VDPWR.n1124 VGND 0.002949f
C7117 VDPWR.n1125 VGND 0.012758f
C7118 VDPWR.n1126 VGND 0.015948f
C7119 VDPWR.t547 VGND 0.005499f
C7120 VDPWR.n1127 VGND 0.016304f
C7121 VDPWR.n1128 VGND 0.009681f
C7122 VDPWR.n1129 VGND 0.005888f
C7123 VDPWR.n1130 VGND 0.010659f
C7124 VDPWR.n1131 VGND 0.015934f
C7125 VDPWR.t1271 VGND 0.072626f
C7126 VDPWR.n1132 VGND 0.03993f
C7127 VDPWR.t449 VGND 0.004984f
C7128 VDPWR.n1133 VGND 0.005908f
C7129 VDPWR.t665 VGND 0.005483f
C7130 VDPWR.n1134 VGND 0.006928f
C7131 VDPWR.n1135 VGND 0.002048f
C7132 VDPWR.n1136 VGND 0.001973f
C7133 VDPWR.n1137 VGND 0.001579f
C7134 VDPWR.n1138 VGND 0.001579f
C7135 VDPWR.n1139 VGND 0.001973f
C7136 VDPWR.n1140 VGND 0.002048f
C7137 VDPWR.n1141 VGND 0.005888f
C7138 VDPWR.t1172 VGND 0.072626f
C7139 VDPWR.n1142 VGND 0.012342f
C7140 VDPWR.n1143 VGND 0.002944f
C7141 VDPWR.n1144 VGND 0.002112f
C7142 VDPWR.n1145 VGND 0.001973f
C7143 VDPWR.n1146 VGND 0.00288f
C7144 VDPWR.n1147 VGND 0.002048f
C7145 VDPWR.n1148 VGND 0.012758f
C7146 VDPWR.n1149 VGND 0.009777f
C7147 VDPWR.n1150 VGND 0.036592f
C7148 VDPWR.n1151 VGND 0.005756f
C7149 VDPWR.n1152 VGND 0.005888f
C7150 VDPWR.t644 VGND 0.005483f
C7151 VDPWR.n1153 VGND 0.006928f
C7152 VDPWR.t1184 VGND 0.072626f
C7153 VDPWR.n1154 VGND 0.036175f
C7154 VDPWR.t666 VGND 0.005483f
C7155 VDPWR.n1155 VGND 0.003531f
C7156 VDPWR.t659 VGND 0.005483f
C7157 VDPWR.n1156 VGND 0.006928f
C7158 VDPWR.n1157 VGND 0.005888f
C7159 VDPWR.t1174 VGND 0.072626f
C7160 VDPWR.n1158 VGND 0.036592f
C7161 VDPWR.n1159 VGND 0.00224f
C7162 VDPWR.n1160 VGND 0.001973f
C7163 VDPWR.n1161 VGND 0.00352f
C7164 VDPWR.n1162 VGND 0.116061f
C7165 VDPWR.n1163 VGND 0.00352f
C7166 VDPWR.n1164 VGND 0.001973f
C7167 VDPWR.n1165 VGND 0.002048f
C7168 VDPWR.t441 VGND 0.066226f
C7169 VDPWR.t616 VGND 0.072641f
C7170 VDPWR.t477 VGND 0.109622f
C7171 VDPWR.t577 VGND 0.063962f
C7172 VDPWR.t559 VGND 0.109622f
C7173 VDPWR.t545 VGND 0.098679f
C7174 VDPWR.n1166 VGND 0.072506f
C7175 VDPWR.t447 VGND 0.086792f
C7176 VDPWR.t749 VGND 0.109622f
C7177 VDPWR.t664 VGND 0.098679f
C7178 VDPWR.t643 VGND 0.109622f
C7179 VDPWR.t658 VGND 0.098679f
C7180 VDPWR.t513 VGND 0.052075f
C7181 VDPWR.t47 VGND 0.046226f
C7182 VDPWR.t932 VGND 0.033019f
C7183 VDPWR.t759 VGND 0.017358f
C7184 VDPWR.t605 VGND 0.006604f
C7185 VDPWR.t994 VGND 0.047358f
C7186 VDPWR.t992 VGND 0.038302f
C7187 VDPWR.t996 VGND 0.012264f
C7188 VDPWR.t934 VGND 0.021509f
C7189 VDPWR.t132 VGND 0.015849f
C7190 VDPWR.t1017 VGND 0.015849f
C7191 VDPWR.t135 VGND 0.017547f
C7192 VDPWR.t44 VGND 0.017924f
C7193 VDPWR.t65 VGND 0.017924f
C7194 VDPWR.t94 VGND 0.024906f
C7195 VDPWR.t1002 VGND 0.023208f
C7196 VDPWR.t1004 VGND 0.013019f
C7197 VDPWR.t134 VGND 0.017924f
C7198 VDPWR.t346 VGND 0.017924f
C7199 VDPWR.t133 VGND 0.015849f
C7200 VDPWR.t348 VGND 0.016038f
C7201 VDPWR.t918 VGND 0.023396f
C7202 VDPWR.t6 VGND 0.01283f
C7203 VDPWR.t136 VGND 0.013585f
C7204 VDPWR.t102 VGND 0.015849f
C7205 VDPWR.t1013 VGND 0.008868f
C7206 VDPWR.t739 VGND 0.072641f
C7207 VDPWR.n1167 VGND 0.060619f
C7208 VDPWR.n1168 VGND 0.009361f
C7209 VDPWR.n1169 VGND 0.002048f
C7210 VDPWR.n1170 VGND 0.001579f
C7211 VDPWR.n1171 VGND 0.001579f
C7212 VDPWR.n1172 VGND 0.001973f
C7213 VDPWR.n1173 VGND 0.002944f
C7214 VDPWR.n1174 VGND 0.002944f
C7215 VDPWR.n1175 VGND 0.002048f
C7216 VDPWR.n1176 VGND 0.012342f
C7217 VDPWR.t645 VGND 0.005483f
C7218 VDPWR.n1177 VGND 0.006928f
C7219 VDPWR.n1178 VGND 0.006017f
C7220 VDPWR.t740 VGND 0.004984f
C7221 VDPWR.n1179 VGND 0.006247f
C7222 VDPWR.n1180 VGND 0.005888f
C7223 VDPWR.t1275 VGND 0.020799f
C7224 VDPWR.n1181 VGND 0.021306f
C7225 VDPWR.t741 VGND 0.004984f
C7226 VDPWR.t103 VGND 0.007187f
C7227 VDPWR.n1182 VGND 0.012163f
C7228 VDPWR.n1183 VGND 0.003456f
C7229 VDPWR.t919 VGND 0.002754f
C7230 VDPWR.t349 VGND 0.006295f
C7231 VDPWR.n1184 VGND 0.005479f
C7232 VDPWR.n1185 VGND 0.004672f
C7233 VDPWR.n1186 VGND 0.001598f
C7234 VDPWR.n1187 VGND 0.002949f
C7235 VDPWR.n1188 VGND 0.003083f
C7236 VDPWR.n1189 VGND 0.001973f
C7237 VDPWR.n1190 VGND 0.00352f
C7238 VDPWR.n1191 VGND 0.140809f
C7239 VDPWR.n1192 VGND 0.281618f
C7240 VDPWR.n1193 VGND 0.116061f
C7241 VDPWR.n1194 VGND 0.003404f
C7242 VDPWR.n1195 VGND 0.003083f
C7243 VDPWR.n1196 VGND 0.00352f
C7244 VDPWR.n1197 VGND 0.001973f
C7245 VDPWR.n1198 VGND 0.002048f
C7246 VDPWR.t747 VGND 0.004984f
C7247 VDPWR.t1166 VGND 0.020982f
C7248 VDPWR.n1200 VGND 0.036453f
C7249 VDPWR.t748 VGND 0.004984f
C7250 VDPWR.n1201 VGND 0.020917f
C7251 VDPWR.t614 VGND 0.004984f
C7252 VDPWR.t1237 VGND 0.020982f
C7253 VDPWR.n1203 VGND 0.036453f
C7254 VDPWR.t615 VGND 0.004984f
C7255 VDPWR.n1204 VGND 0.020917f
C7256 VDPWR.n1205 VGND 0.018023f
C7257 VDPWR.t742 VGND 0.005024f
C7258 VDPWR.t1220 VGND 0.010664f
C7259 VDPWR.n1207 VGND 0.027341f
C7260 VDPWR.t743 VGND 0.005024f
C7261 VDPWR.n1208 VGND 0.014893f
C7262 VDPWR.n1209 VGND 0.001133f
C7263 VDPWR.n1210 VGND 0.005888f
C7264 VDPWR.t43 VGND 0.00632f
C7265 VDPWR.n1211 VGND 0.002085f
C7266 VDPWR.n1212 VGND 0.002405f
C7267 VDPWR.t455 VGND 0.005483f
C7268 VDPWR.n1213 VGND 0.002283f
C7269 VDPWR.n1214 VGND 0.002048f
C7270 VDPWR.n1215 VGND 0.001579f
C7271 VDPWR.n1216 VGND 0.001579f
C7272 VDPWR.n1217 VGND 0.002949f
C7273 VDPWR.n1218 VGND 0.007422f
C7274 VDPWR.n1219 VGND 0.005888f
C7275 VDPWR.t175 VGND 0.002754f
C7276 VDPWR.t826 VGND 0.001152f
C7277 VDPWR.t164 VGND 0.001152f
C7278 VDPWR.n1220 VGND 0.002373f
C7279 VDPWR.n1221 VGND 0.006065f
C7280 VDPWR.t454 VGND 0.0055f
C7281 VDPWR.t746 VGND 0.005055f
C7282 VDPWR.n1222 VGND 0.035589f
C7283 VDPWR.t602 VGND 0.052075f
C7284 VDPWR.t613 VGND 0.069811f
C7285 VDPWR.t46 VGND 0.014151f
C7286 VDPWR.t0 VGND 0.015849f
C7287 VDPWR.t940 VGND 0.015849f
C7288 VDPWR.t906 VGND 0.015849f
C7289 VDPWR.t936 VGND 0.031321f
C7290 VDPWR.t42 VGND 0.024151f
C7291 VDPWR.t2 VGND 0.029811f
C7292 VDPWR.t25 VGND 0.02717f
C7293 VDPWR.t857 VGND 0.015849f
C7294 VDPWR.t166 VGND 0.024717f
C7295 VDPWR.t26 VGND 0.028302f
C7296 VDPWR.t168 VGND 0.04434f
C7297 VDPWR.t165 VGND 0.037358f
C7298 VDPWR.t24 VGND 0.033962f
C7299 VDPWR.t174 VGND 0.033019f
C7300 VDPWR.t453 VGND 0.035472f
C7301 VDPWR.t163 VGND 0.03434f
C7302 VDPWR.t825 VGND 0.021698f
C7303 VDPWR.t744 VGND 0.052075f
C7304 VDPWR.n1223 VGND 0.037789f
C7305 VDPWR.n1224 VGND 0.006017f
C7306 VDPWR.n1225 VGND 0.002048f
C7307 VDPWR.n1226 VGND 0.001973f
C7308 VDPWR.n1227 VGND 0.00352f
C7309 VDPWR.n1228 VGND 0.116061f
C7310 VDPWR.n1229 VGND 0.00352f
C7311 VDPWR.n1230 VGND 0.002757f
C7312 VDPWR.n1231 VGND 0.001579f
C7313 VDPWR.n1232 VGND 0.001579f
C7314 VDPWR.n1233 VGND 0.001973f
C7315 VDPWR.n1234 VGND 0.002944f
C7316 VDPWR.n1235 VGND 0.012758f
C7317 VDPWR.n1236 VGND 0.005888f
C7318 VDPWR.t1177 VGND 0.072626f
C7319 VDPWR.t1223 VGND 0.072626f
C7320 VDPWR.n1237 VGND 0.036592f
C7321 VDPWR.n1238 VGND 0.005344f
C7322 VDPWR.t612 VGND 0.005501f
C7323 VDPWR.n1239 VGND 0.011251f
C7324 VDPWR.n1240 VGND 0.005888f
C7325 VDPWR.n1241 VGND 0.012758f
C7326 VDPWR.n1242 VGND 0.002048f
C7327 VDPWR.n1243 VGND 0.001973f
C7328 VDPWR.n1244 VGND 0.00352f
C7329 VDPWR.n1245 VGND 0.116061f
C7330 VDPWR.n1246 VGND 0.116061f
C7331 VDPWR.n1247 VGND 0.00352f
C7332 VDPWR.n1248 VGND 0.002949f
C7333 VDPWR.n1249 VGND 0.001579f
C7334 VDPWR.n1250 VGND 0.002048f
C7335 VDPWR.n1251 VGND 0.002112f
C7336 VDPWR.n1252 VGND 0.001579f
C7337 VDPWR.n1253 VGND 0.001973f
C7338 VDPWR.n1254 VGND 0.00288f
C7339 VDPWR.t1235 VGND 0.072626f
C7340 VDPWR.n1255 VGND 0.009361f
C7341 VDPWR.n1256 VGND 0.004416f
C7342 VDPWR.t726 VGND 0.005059f
C7343 VDPWR.n1257 VGND 0.01476f
C7344 VDPWR.n1258 VGND 0.015674f
C7345 VDPWR.t1189 VGND 0.021124f
C7346 VDPWR.n1259 VGND 0.020912f
C7347 VDPWR.t725 VGND 0.004984f
C7348 VDPWR.n1260 VGND 0.005999f
C7349 VDPWR.n1261 VGND 0.006f
C7350 VDPWR.t536 VGND 0.066226f
C7351 VDPWR.t519 VGND 0.072641f
C7352 VDPWR.t717 VGND 0.109622f
C7353 VDPWR.t580 VGND 0.063962f
C7354 VDPWR.t468 VGND 0.109622f
C7355 VDPWR.t550 VGND 0.098679f
C7356 VDPWR.t574 VGND 0.098679f
C7357 VDPWR.t650 VGND 0.109622f
C7358 VDPWR.t610 VGND 0.098679f
C7359 VDPWR.t752 VGND 0.109622f
C7360 VDPWR.t724 VGND 0.034717f
C7361 VDPWR.n1262 VGND 0.037412f
C7362 VDPWR.n1263 VGND 0.006017f
C7363 VDPWR.n1264 VGND 0.002048f
C7364 VDPWR.n1265 VGND 0.001973f
C7365 VDPWR.n1266 VGND 0.00352f
C7366 VDPWR.n1267 VGND 0.116061f
C7367 VDPWR.n1268 VGND 0.00352f
C7368 VDPWR.n1269 VGND 0.002949f
C7369 VDPWR.n1270 VGND 0.001579f
C7370 VDPWR.n1271 VGND 0.002048f
C7371 VDPWR.n1272 VGND 0.002944f
C7372 VDPWR.t1260 VGND 0.072626f
C7373 VDPWR.n1273 VGND 0.012758f
C7374 VDPWR.n1274 VGND 0.005344f
C7375 VDPWR.t1286 VGND 0.074001f
C7376 VDPWR.t582 VGND 0.005483f
C7377 VDPWR.n1275 VGND 0.006928f
C7378 VDPWR.n1276 VGND 0.005888f
C7379 VDPWR.n1277 VGND 0.008742f
C7380 VDPWR.n1278 VGND 0.005888f
C7381 VDPWR.t1246 VGND 0.072626f
C7382 VDPWR.n1279 VGND 0.040608f
C7383 VDPWR.n1280 VGND 0.00288f
C7384 VDPWR.n1281 VGND 0.001973f
C7385 VDPWR.n1282 VGND 0.00352f
C7386 VDPWR.n1283 VGND 0.155317f
C7387 VDPWR.n1284 VGND 0.167264f
C7388 VDPWR.n1285 VGND 0.003404f
C7389 VDPWR.n1286 VGND 0.00352f
C7390 VDPWR.n1287 VGND 0.001477f
C7391 VDPWR.n1288 VGND 0.001579f
C7392 VDPWR.n1289 VGND 0.002048f
C7393 VDPWR.n1290 VGND 0.003083f
C7394 VDPWR.t1088 VGND 0.001527f
C7395 VDPWR.t41 VGND 0.001527f
C7396 VDPWR.n1291 VGND 0.003322f
C7397 VDPWR.t686 VGND 0.004984f
C7398 VDPWR.n1292 VGND 0.011445f
C7399 VDPWR.n1293 VGND 0.005888f
C7400 VDPWR.n1294 VGND 0.015256f
C7401 VDPWR.n1295 VGND 0.005888f
C7402 VDPWR.t1171 VGND 0.036876f
C7403 VDPWR.t654 VGND 0.005483f
C7404 VDPWR.n1296 VGND 0.003947f
C7405 VDPWR.n1297 VGND 0.022156f
C7406 VDPWR.n1298 VGND 0.002048f
C7407 VDPWR.n1299 VGND 0.001973f
C7408 VDPWR.n1300 VGND 0.00352f
C7409 VDPWR.n1301 VGND 0.00352f
C7410 VDPWR.n1302 VGND 0.002757f
C7411 VDPWR.n1303 VGND 0.001579f
C7412 VDPWR.n1304 VGND 0.001579f
C7413 VDPWR.n1305 VGND 0.001973f
C7414 VDPWR.n1306 VGND 0.002944f
C7415 VDPWR.n1307 VGND 0.012758f
C7416 VDPWR.n1308 VGND 0.005888f
C7417 VDPWR.t1191 VGND 0.072626f
C7418 VDPWR.t1168 VGND 0.072626f
C7419 VDPWR.n1309 VGND 0.066804f
C7420 VDPWR.n1310 VGND 0.005888f
C7421 VDPWR.t466 VGND 0.005483f
C7422 VDPWR.t622 VGND 0.005483f
C7423 VDPWR.n1311 VGND 0.007477f
C7424 VDPWR.t567 VGND 0.005483f
C7425 VDPWR.t710 VGND 0.005483f
C7426 VDPWR.n1312 VGND 0.007477f
C7427 VDPWR.n1313 VGND 0.003904f
C7428 VDPWR.n1314 VGND 0.012758f
C7429 VDPWR.n1315 VGND 0.002112f
C7430 VDPWR.n1316 VGND 0.001973f
C7431 VDPWR.n1317 VGND 0.00352f
C7432 VDPWR.n1318 VGND 0.00352f
C7433 VDPWR.n1319 VGND 0.002949f
C7434 VDPWR.n1320 VGND 0.001579f
C7435 VDPWR.n1321 VGND 0.009361f
C7436 VDPWR.n1322 VGND 0.005888f
C7437 VDPWR.t566 VGND 0.005483f
C7438 VDPWR.t709 VGND 0.005483f
C7439 VDPWR.n1323 VGND 0.007477f
C7440 VDPWR.t487 VGND 0.005024f
C7441 VDPWR.t1244 VGND 0.010664f
C7442 VDPWR.n1325 VGND 0.027341f
C7443 VDPWR.t488 VGND 0.005024f
C7444 VDPWR.n1326 VGND 0.014893f
C7445 VDPWR.t675 VGND 0.005499f
C7446 VDPWR.n1327 VGND 0.016304f
C7447 VDPWR.t621 VGND 0.005483f
C7448 VDPWR.n1328 VGND 0.006928f
C7449 VDPWR.n1329 VGND 0.002048f
C7450 VDPWR.n1330 VGND 0.001973f
C7451 VDPWR.n1331 VGND 0.00352f
C7452 VDPWR.n1332 VGND 0.00352f
C7453 VDPWR.n1333 VGND 0.002949f
C7454 VDPWR.n1334 VGND 0.001579f
C7455 VDPWR.n1335 VGND 0.002048f
C7456 VDPWR.n1336 VGND 0.002944f
C7457 VDPWR.t1213 VGND 0.072626f
C7458 VDPWR.n1337 VGND 0.012758f
C7459 VDPWR.n1338 VGND 0.005344f
C7460 VDPWR.t1192 VGND 0.074001f
C7461 VDPWR.t524 VGND 0.005483f
C7462 VDPWR.n1339 VGND 0.006928f
C7463 VDPWR.n1340 VGND 0.005888f
C7464 VDPWR.n1341 VGND 0.008742f
C7465 VDPWR.n1342 VGND 0.005888f
C7466 VDPWR.t1272 VGND 0.072626f
C7467 VDPWR.n1343 VGND 0.040608f
C7468 VDPWR.n1344 VGND 0.00288f
C7469 VDPWR.n1345 VGND 0.001973f
C7470 VDPWR.n1346 VGND 0.00352f
C7471 VDPWR.n1347 VGND 0.001579f
C7472 VDPWR.n1348 VGND 0.002048f
C7473 VDPWR.t1239 VGND 0.036234f
C7474 VDPWR.n1349 VGND 0.027337f
C7475 VDPWR.t523 VGND 0.005483f
C7476 VDPWR.t505 VGND 0.004984f
C7477 VDPWR.n1350 VGND 0.011995f
C7478 VDPWR.t457 VGND 0.005024f
C7479 VDPWR.t1258 VGND 0.010664f
C7480 VDPWR.n1352 VGND 0.027341f
C7481 VDPWR.t458 VGND 0.005024f
C7482 VDPWR.n1353 VGND 0.014893f
C7483 VDPWR.t646 VGND 0.005024f
C7484 VDPWR.t1225 VGND 0.010664f
C7485 VDPWR.n1355 VGND 0.027341f
C7486 VDPWR.t647 VGND 0.005024f
C7487 VDPWR.n1356 VGND 0.014893f
C7488 VDPWR.n1357 VGND 0.01227f
C7489 VDPWR.t430 VGND 0.005024f
C7490 VDPWR.t1262 VGND 0.010664f
C7491 VDPWR.n1359 VGND 0.027341f
C7492 VDPWR.t431 VGND 0.005024f
C7493 VDPWR.n1360 VGND 0.014893f
C7494 VDPWR.n1361 VGND 0.003844f
C7495 VDPWR.n1362 VGND 0.004957f
C7496 VDPWR.t633 VGND 0.005024f
C7497 VDPWR.t1233 VGND 0.010664f
C7498 VDPWR.n1364 VGND 0.027341f
C7499 VDPWR.t634 VGND 0.005024f
C7500 VDPWR.n1365 VGND 0.014893f
C7501 VDPWR.n1366 VGND 0.013462f
C7502 VDPWR.n1367 VGND 0.00331f
C7503 VDPWR.n1368 VGND 0.003842f
C7504 VDPWR.n1369 VGND 0.004416f
C7505 VDPWR.n1370 VGND 0.002368f
C7506 VDPWR.n1371 VGND 0.001973f
C7507 VDPWR.n1372 VGND 0.003404f
C7508 VDPWR.n1373 VGND 0.003083f
C7509 VDPWR.n1374 VGND 0.002629f
C7510 VDPWR.n1375 VGND 0.00352f
C7511 VDPWR.n1376 VGND 0.015256f
C7512 VDPWR.n1377 VGND 0.025685f
C7513 VDPWR.n1378 VGND 0.015256f
C7514 VDPWR.n1379 VGND 0.015934f
C7515 VDPWR.n1380 VGND 0.002048f
C7516 VDPWR.n1381 VGND 0.002944f
C7517 VDPWR.n1382 VGND 0.001973f
C7518 VDPWR.n1383 VGND 0.001579f
C7519 VDPWR.n1384 VGND 0.00352f
C7520 VDPWR.n1385 VGND 0.003404f
C7521 VDPWR.n1386 VGND 0.003083f
C7522 VDPWR.n1387 VGND 0.002117f
C7523 VDPWR.n1388 VGND 0.003008f
C7524 VDPWR.n1389 VGND 0.015256f
C7525 VDPWR.n1390 VGND 0.020793f
C7526 VDPWR.t506 VGND 0.004984f
C7527 VDPWR.n1391 VGND 0.011445f
C7528 VDPWR.n1392 VGND 0.020115f
C7529 VDPWR.n1393 VGND 0.005888f
C7530 VDPWR.n1394 VGND 0.003488f
C7531 VDPWR.n1395 VGND 0.004416f
C7532 VDPWR.n1396 VGND 0.005612f
C7533 VDPWR.t620 VGND 0.005483f
C7534 VDPWR.n1397 VGND 0.006928f
C7535 VDPWR.n1398 VGND 0.012342f
C7536 VDPWR.n1399 VGND 0.012342f
C7537 VDPWR.n1400 VGND 0.005888f
C7538 VDPWR.n1401 VGND 0.003488f
C7539 VDPWR.n1402 VGND 0.003209f
C7540 VDPWR.n1403 VGND 0.034322f
C7541 VDPWR.n1404 VGND 0.002865f
C7542 VDPWR.t674 VGND 0.005483f
C7543 VDPWR.n1405 VGND 0.006928f
C7544 VDPWR.n1406 VGND 0.012342f
C7545 VDPWR.n1407 VGND 0.005888f
C7546 VDPWR.n1408 VGND 0.005888f
C7547 VDPWR.n1409 VGND 0.004544f
C7548 VDPWR.n1410 VGND 0.009777f
C7549 VDPWR.n1411 VGND 0.036592f
C7550 VDPWR.n1412 VGND 0.009361f
C7551 VDPWR.n1413 VGND 0.012342f
C7552 VDPWR.n1414 VGND 0.012758f
C7553 VDPWR.n1415 VGND 0.002048f
C7554 VDPWR.n1416 VGND 0.001579f
C7555 VDPWR.n1417 VGND 0.001973f
C7556 VDPWR.n1418 VGND 0.00224f
C7557 VDPWR.n1419 VGND 0.002752f
C7558 VDPWR.n1420 VGND 0.001973f
C7559 VDPWR.n1421 VGND 0.003083f
C7560 VDPWR.n1422 VGND 0.003404f
C7561 VDPWR.n1423 VGND 0.155317f
C7562 VDPWR.n1424 VGND 0.003404f
C7563 VDPWR.n1425 VGND 0.003083f
C7564 VDPWR.n1426 VGND 0.002949f
C7565 VDPWR.n1427 VGND 0.002528f
C7566 VDPWR.n1428 VGND 0.006017f
C7567 VDPWR.t456 VGND 0.066226f
C7568 VDPWR.t429 VGND 0.072641f
C7569 VDPWR.t504 VGND 0.109622f
C7570 VDPWR.t522 VGND 0.063962f
C7571 VDPWR.t619 VGND 0.109622f
C7572 VDPWR.t673 VGND 0.098679f
C7573 VDPWR.t450 VGND 0.052075f
C7574 VDPWR.t459 VGND 0.208301f
C7575 VDPWR.t40 VGND 0.028868f
C7576 VDPWR.t1087 VGND 0.022453f
C7577 VDPWR.t653 VGND 0.063962f
C7578 VDPWR.t684 VGND 0.092075f
C7579 VDPWR.n1429 VGND 0.040844f
C7580 VDPWR.t465 VGND 0.208301f
C7581 VDPWR.t565 VGND 0.208301f
C7582 VDPWR.t486 VGND 0.055283f
C7583 VDPWR.n1430 VGND 0.05194f
C7584 VDPWR.n1431 VGND 0.015948f
C7585 VDPWR.n1432 VGND 0.003168f
C7586 VDPWR.n1433 VGND 0.004953f
C7587 VDPWR.n1434 VGND 0.010348f
C7588 VDPWR.n1435 VGND 0.004425f
C7589 VDPWR.n1436 VGND 0.004416f
C7590 VDPWR.n1437 VGND 0.005888f
C7591 VDPWR.n1438 VGND 0.012342f
C7592 VDPWR.n1439 VGND 0.012758f
C7593 VDPWR.t1281 VGND 0.072626f
C7594 VDPWR.t1252 VGND 0.072626f
C7595 VDPWR.n1440 VGND 0.066804f
C7596 VDPWR.n1441 VGND 0.009777f
C7597 VDPWR.n1442 VGND 0.005888f
C7598 VDPWR.n1443 VGND 0.005888f
C7599 VDPWR.n1444 VGND 0.005568f
C7600 VDPWR.n1445 VGND 0.012758f
C7601 VDPWR.n1446 VGND 0.012758f
C7602 VDPWR.n1447 VGND 0.002048f
C7603 VDPWR.n1448 VGND 0.001579f
C7604 VDPWR.n1449 VGND 0.001973f
C7605 VDPWR.n1450 VGND 0.00288f
C7606 VDPWR.n1451 VGND 0.002048f
C7607 VDPWR.n1452 VGND 0.002944f
C7608 VDPWR.n1453 VGND 0.001973f
C7609 VDPWR.n1454 VGND 0.003083f
C7610 VDPWR.n1455 VGND 0.003404f
C7611 VDPWR.n1456 VGND 0.155317f
C7612 VDPWR.n1457 VGND 0.003404f
C7613 VDPWR.n1458 VGND 0.003083f
C7614 VDPWR.n1459 VGND 0.002949f
C7615 VDPWR.n1460 VGND 0.002048f
C7616 VDPWR.n1461 VGND 0.012758f
C7617 VDPWR.n1462 VGND 0.012758f
C7618 VDPWR.n1463 VGND 0.012342f
C7619 VDPWR.n1464 VGND 0.005888f
C7620 VDPWR.n1465 VGND 0.004818f
C7621 VDPWR.n1466 VGND 0.004712f
C7622 VDPWR.n1467 VGND 0.005344f
C7623 VDPWR.n1468 VGND 0.005888f
C7624 VDPWR.n1469 VGND 0.012342f
C7625 VDPWR.n1470 VGND 0.012758f
C7626 VDPWR.n1471 VGND 0.009777f
C7627 VDPWR.n1472 VGND 0.005888f
C7628 VDPWR.n1473 VGND 0.005888f
C7629 VDPWR.n1474 VGND 0.009361f
C7630 VDPWR.n1475 VGND 0.012758f
C7631 VDPWR.n1476 VGND 0.012758f
C7632 VDPWR.n1477 VGND 0.005888f
C7633 VDPWR.n1478 VGND 0.005888f
C7634 VDPWR.n1479 VGND 0.003648f
C7635 VDPWR.n1480 VGND 0.012758f
C7636 VDPWR.t467 VGND 0.005483f
C7637 VDPWR.n1481 VGND 0.00453f
C7638 VDPWR.t623 VGND 0.005483f
C7639 VDPWR.n1482 VGND 0.007477f
C7640 VDPWR.n1483 VGND 0.002944f
C7641 VDPWR.n1484 VGND 0.002048f
C7642 VDPWR.n1485 VGND 0.012342f
C7643 VDPWR.n1486 VGND 0.012758f
C7644 VDPWR.n1487 VGND 0.002048f
C7645 VDPWR.n1488 VGND 0.00224f
C7646 VDPWR.n1489 VGND 0.001973f
C7647 VDPWR.n1490 VGND 0.003083f
C7648 VDPWR.n1491 VGND 0.003404f
C7649 VDPWR.n1492 VGND 0.155317f
C7650 VDPWR.n1493 VGND 0.003404f
C7651 VDPWR.n1494 VGND 0.003083f
C7652 VDPWR.n1495 VGND 5.48e-19
C7653 VDPWR.n1496 VGND 0.003168f
C7654 VDPWR.n1497 VGND 0.00224f
C7655 VDPWR.n1498 VGND 0.001642f
C7656 VDPWR.n1499 VGND 0.003023f
C7657 VDPWR.n1500 VGND 0.002272f
C7658 VDPWR.n1501 VGND 0.004416f
C7659 VDPWR.n1502 VGND 0.008674f
C7660 VDPWR.t685 VGND 0.004984f
C7661 VDPWR.n1503 VGND 0.011445f
C7662 VDPWR.n1504 VGND 0.015143f
C7663 VDPWR.n1505 VGND 0.052403f
C7664 VDPWR.t1222 VGND 0.072626f
C7665 VDPWR.n1506 VGND 0.040608f
C7666 VDPWR.n1507 VGND 0.010509f
C7667 VDPWR.n1508 VGND 0.005888f
C7668 VDPWR.n1509 VGND 0.005888f
C7669 VDPWR.n1510 VGND 0.005888f
C7670 VDPWR.n1511 VGND 0.020793f
C7671 VDPWR.n1512 VGND 0.020793f
C7672 VDPWR.n1513 VGND 0.020115f
C7673 VDPWR.n1514 VGND 0.005888f
C7674 VDPWR.n1515 VGND 0.003488f
C7675 VDPWR.n1516 VGND 0.008952f
C7676 VDPWR.n1517 VGND 0.00176f
C7677 VDPWR.n1518 VGND 0.007073f
C7678 VDPWR.n1519 VGND 0.013601f
C7679 VDPWR.t655 VGND 0.005483f
C7680 VDPWR.n1520 VGND 0.00426f
C7681 VDPWR.t460 VGND 0.005483f
C7682 VDPWR.t608 VGND 0.005483f
C7683 VDPWR.n1521 VGND 0.007477f
C7684 VDPWR.n1522 VGND 9.32e-19
C7685 VDPWR.n1523 VGND 0.005888f
C7686 VDPWR.t1195 VGND 0.072626f
C7687 VDPWR.t1170 VGND 0.072626f
C7688 VDPWR.n1524 VGND 0.066804f
C7689 VDPWR.n1525 VGND 0.005888f
C7690 VDPWR.n1526 VGND 0.012758f
C7691 VDPWR.n1527 VGND 0.005888f
C7692 VDPWR.t461 VGND 0.005483f
C7693 VDPWR.t609 VGND 0.005483f
C7694 VDPWR.n1528 VGND 0.007477f
C7695 VDPWR.n1529 VGND 7.36e-19
C7696 VDPWR.n1530 VGND 0.001973f
C7697 VDPWR.n1531 VGND 0.155317f
C7698 VDPWR.n1532 VGND 0.00352f
C7699 VDPWR.n1533 VGND 0.001579f
C7700 VDPWR.n1534 VGND 0.0024f
C7701 VDPWR.n1535 VGND 0.002048f
C7702 VDPWR.n1536 VGND 0.002112f
C7703 VDPWR.n1537 VGND 0.00453f
C7704 VDPWR.t451 VGND 0.005024f
C7705 VDPWR.t1257 VGND 0.010664f
C7706 VDPWR.n1539 VGND 0.027341f
C7707 VDPWR.t452 VGND 0.005024f
C7708 VDPWR.n1540 VGND 0.014893f
C7709 VDPWR.t648 VGND 0.005024f
C7710 VDPWR.t1226 VGND 0.010664f
C7711 VDPWR.n1542 VGND 0.027341f
C7712 VDPWR.t649 VGND 0.005024f
C7713 VDPWR.n1543 VGND 0.014893f
C7714 VDPWR.n1544 VGND 0.001973f
C7715 VDPWR.n1545 VGND 0.003404f
C7716 VDPWR.n1546 VGND 0.003083f
C7717 VDPWR.n1547 VGND 0.002885f
C7718 VDPWR.n1548 VGND 0.001376f
C7719 VDPWR.n1549 VGND 0.012555f
C7720 VDPWR.n1550 VGND 0.002048f
C7721 VDPWR.n1551 VGND 0.002944f
C7722 VDPWR.n1552 VGND 0.001973f
C7723 VDPWR.n1553 VGND 0.001579f
C7724 VDPWR.n1554 VGND 0.00352f
C7725 VDPWR.n1555 VGND 0.003404f
C7726 VDPWR.n1556 VGND 0.003083f
C7727 VDPWR.n1557 VGND 0.002949f
C7728 VDPWR.n1558 VGND 0.005696f
C7729 VDPWR.n1559 VGND 0.012342f
C7730 VDPWR.n1560 VGND 0.012758f
C7731 VDPWR.n1561 VGND 0.012758f
C7732 VDPWR.n1562 VGND 0.005888f
C7733 VDPWR.n1563 VGND 0.005888f
C7734 VDPWR.n1564 VGND 0.005888f
C7735 VDPWR.n1565 VGND 0.012758f
C7736 VDPWR.n1566 VGND 0.012758f
C7737 VDPWR.n1567 VGND 0.009361f
C7738 VDPWR.n1568 VGND 0.005888f
C7739 VDPWR.n1569 VGND 0.005888f
C7740 VDPWR.n1570 VGND 0.009777f
C7741 VDPWR.n1571 VGND 0.012758f
C7742 VDPWR.n1572 VGND 0.012342f
C7743 VDPWR.n1573 VGND 0.005888f
C7744 VDPWR.n1574 VGND 0.004416f
C7745 VDPWR.n1575 VGND 0.004739f
C7746 VDPWR.n1576 VGND 0.002934f
C7747 VDPWR.n1577 VGND 0.001504f
C7748 VDPWR.n1578 VGND 0.002944f
C7749 VDPWR.n1579 VGND 0.001973f
C7750 VDPWR.n1580 VGND 0.00352f
C7751 VDPWR.n1581 VGND 0.001579f
C7752 VDPWR.n1582 VGND 0.001973f
C7753 VDPWR.n1583 VGND 0.002112f
C7754 VDPWR.n1584 VGND 0.002336f
C7755 VDPWR.n1585 VGND 0.001973f
C7756 VDPWR.n1586 VGND 0.003083f
C7757 VDPWR.n1587 VGND 0.003404f
C7758 VDPWR.n1588 VGND 0.155317f
C7759 VDPWR.n1589 VGND 0.116061f
C7760 VDPWR.n1590 VGND 0.281618f
C7761 VDPWR.n1591 VGND 0.281618f
C7762 VDPWR.n1592 VGND 0.281618f
C7763 VDPWR.n1593 VGND 0.532156f
C7764 VDPWR.n1594 VGND 0.194931f
C7765 VDPWR.n1595 VGND 0.003404f
C7766 VDPWR.n1596 VGND 0.194931f
C7767 VDPWR.n1597 VGND 0.00352f
C7768 VDPWR.n1598 VGND 0.002629f
C7769 VDPWR.n1599 VGND 0.001579f
C7770 VDPWR.n1600 VGND 0.002944f
C7771 VDPWR.n1601 VGND 0.015256f
C7772 VDPWR.t578 VGND 0.005483f
C7773 VDPWR.t478 VGND 0.004984f
C7774 VDPWR.n1602 VGND 0.011995f
C7775 VDPWR.n1603 VGND 0.003842f
C7776 VDPWR.t617 VGND 0.005024f
C7777 VDPWR.t1186 VGND 0.010664f
C7778 VDPWR.n1605 VGND 0.027341f
C7779 VDPWR.t618 VGND 0.005024f
C7780 VDPWR.n1606 VGND 0.014893f
C7781 VDPWR.n1607 VGND 0.00352f
C7782 VDPWR.n1608 VGND 0.004416f
C7783 VDPWR.n1609 VGND 0.004957f
C7784 VDPWR.t694 VGND 0.005024f
C7785 VDPWR.t1169 VGND 0.010664f
C7786 VDPWR.n1611 VGND 0.027341f
C7787 VDPWR.t695 VGND 0.005024f
C7788 VDPWR.n1612 VGND 0.014893f
C7789 VDPWR.t442 VGND 0.005024f
C7790 VDPWR.t1251 VGND 0.010664f
C7791 VDPWR.n1614 VGND 0.027341f
C7792 VDPWR.t443 VGND 0.005024f
C7793 VDPWR.n1615 VGND 0.014893f
C7794 VDPWR.n1616 VGND 0.003844f
C7795 VDPWR.t534 VGND 0.005024f
C7796 VDPWR.t1229 VGND 0.010664f
C7797 VDPWR.n1618 VGND 0.027341f
C7798 VDPWR.t535 VGND 0.005024f
C7799 VDPWR.n1619 VGND 0.014893f
C7800 VDPWR.n1620 VGND 0.01227f
C7801 VDPWR.n1621 VGND 0.013462f
C7802 VDPWR.n1622 VGND 0.00331f
C7803 VDPWR.t1241 VGND 0.036234f
C7804 VDPWR.n1623 VGND 0.027337f
C7805 VDPWR.n1624 VGND 0.025685f
C7806 VDPWR.t1210 VGND 0.072626f
C7807 VDPWR.n1625 VGND 0.040608f
C7808 VDPWR.n1626 VGND 0.005888f
C7809 VDPWR.t479 VGND 0.004984f
C7810 VDPWR.n1627 VGND 0.011445f
C7811 VDPWR.t560 VGND 0.005483f
C7812 VDPWR.n1628 VGND 0.006928f
C7813 VDPWR.n1629 VGND 0.005888f
C7814 VDPWR.t1208 VGND 0.074001f
C7815 VDPWR.n1630 VGND 0.034322f
C7816 VDPWR.n1631 VGND 0.005888f
C7817 VDPWR.t1224 VGND 0.072626f
C7818 VDPWR.n1632 VGND 0.009361f
C7819 VDPWR.n1633 VGND 0.036592f
C7820 VDPWR.n1634 VGND 0.009777f
C7821 VDPWR.n1635 VGND 0.004544f
C7822 VDPWR.n1636 VGND 0.005888f
C7823 VDPWR.n1637 VGND 0.012758f
C7824 VDPWR.n1638 VGND 0.012342f
C7825 VDPWR.t546 VGND 0.005483f
C7826 VDPWR.n1639 VGND 0.006928f
C7827 VDPWR.n1640 VGND 0.002865f
C7828 VDPWR.n1641 VGND 0.005344f
C7829 VDPWR.n1642 VGND 0.003488f
C7830 VDPWR.n1643 VGND 0.003209f
C7831 VDPWR.t579 VGND 0.005483f
C7832 VDPWR.n1644 VGND 0.006928f
C7833 VDPWR.n1645 VGND 0.012342f
C7834 VDPWR.n1646 VGND 0.012342f
C7835 VDPWR.n1647 VGND 0.005888f
C7836 VDPWR.n1648 VGND 0.004416f
C7837 VDPWR.n1649 VGND 0.005612f
C7838 VDPWR.n1650 VGND 0.008742f
C7839 VDPWR.n1651 VGND 0.003488f
C7840 VDPWR.n1652 VGND 0.005888f
C7841 VDPWR.n1653 VGND 0.020115f
C7842 VDPWR.n1654 VGND 0.020793f
C7843 VDPWR.n1655 VGND 0.015256f
C7844 VDPWR.n1656 VGND 0.003008f
C7845 VDPWR.n1657 VGND 0.002117f
C7846 VDPWR.n1658 VGND 0.001973f
C7847 VDPWR.n1659 VGND 0.00352f
C7848 VDPWR.n1660 VGND 0.001579f
C7849 VDPWR.n1661 VGND 0.003083f
C7850 VDPWR.n1662 VGND 0.001973f
C7851 VDPWR.n1663 VGND 0.00288f
C7852 VDPWR.n1664 VGND 0.002048f
C7853 VDPWR.n1665 VGND 0.015934f
C7854 VDPWR.n1666 VGND 0.015256f
C7855 VDPWR.n1667 VGND 0.002048f
C7856 VDPWR.n1668 VGND 0.002368f
C7857 VDPWR.n1669 VGND 0.001973f
C7858 VDPWR.n1670 VGND 0.003083f
C7859 VDPWR.n1671 VGND 0.003404f
C7860 VDPWR.n1672 VGND 0.140809f
C7861 VDPWR.n1673 VGND 0.281618f
C7862 VDPWR.n1674 VGND 0.532156f
C7863 VDPWR.n1675 VGND 0.194931f
C7864 VDPWR.n1676 VGND 0.00352f
C7865 VDPWR.n1677 VGND 0.002629f
C7866 VDPWR.n1678 VGND 0.001579f
C7867 VDPWR.n1679 VGND 0.001579f
C7868 VDPWR.n1680 VGND 0.001973f
C7869 VDPWR.n1681 VGND 0.002944f
C7870 VDPWR.t1199 VGND 0.036234f
C7871 VDPWR.n1682 VGND 0.027337f
C7872 VDPWR.t581 VGND 0.005483f
C7873 VDPWR.t718 VGND 0.004984f
C7874 VDPWR.n1683 VGND 0.011995f
C7875 VDPWR.t690 VGND 0.005024f
C7876 VDPWR.t1221 VGND 0.010664f
C7877 VDPWR.n1685 VGND 0.027341f
C7878 VDPWR.t691 VGND 0.005024f
C7879 VDPWR.n1686 VGND 0.014893f
C7880 VDPWR.t537 VGND 0.005024f
C7881 VDPWR.t1266 VGND 0.010664f
C7882 VDPWR.n1688 VGND 0.027341f
C7883 VDPWR.t538 VGND 0.005024f
C7884 VDPWR.n1689 VGND 0.014893f
C7885 VDPWR.n1690 VGND 0.01227f
C7886 VDPWR.t520 VGND 0.005024f
C7887 VDPWR.t1227 VGND 0.010664f
C7888 VDPWR.n1692 VGND 0.027341f
C7889 VDPWR.t521 VGND 0.005024f
C7890 VDPWR.n1693 VGND 0.014893f
C7891 VDPWR.n1694 VGND 0.003844f
C7892 VDPWR.n1695 VGND 0.004957f
C7893 VDPWR.t702 VGND 0.005024f
C7894 VDPWR.t1197 VGND 0.010664f
C7895 VDPWR.n1697 VGND 0.027341f
C7896 VDPWR.t703 VGND 0.005024f
C7897 VDPWR.n1698 VGND 0.014893f
C7898 VDPWR.n1699 VGND 0.013462f
C7899 VDPWR.n1700 VGND 0.00331f
C7900 VDPWR.n1701 VGND 0.003842f
C7901 VDPWR.n1702 VGND 0.004416f
C7902 VDPWR.n1703 VGND 0.00352f
C7903 VDPWR.n1704 VGND 0.015256f
C7904 VDPWR.n1705 VGND 0.025685f
C7905 VDPWR.n1706 VGND 0.002048f
C7906 VDPWR.n1707 VGND 0.015934f
C7907 VDPWR.n1708 VGND 0.015256f
C7908 VDPWR.n1709 VGND 0.002048f
C7909 VDPWR.n1710 VGND 0.002368f
C7910 VDPWR.n1711 VGND 0.001973f
C7911 VDPWR.n1712 VGND 0.003083f
C7912 VDPWR.n1713 VGND 0.003404f
C7913 VDPWR.n1714 VGND 0.140809f
C7914 VDPWR.n1715 VGND 0.003404f
C7915 VDPWR.n1716 VGND 0.003083f
C7916 VDPWR.n1717 VGND 0.002117f
C7917 VDPWR.n1718 VGND 0.003008f
C7918 VDPWR.n1719 VGND 0.015256f
C7919 VDPWR.n1720 VGND 0.020793f
C7920 VDPWR.t719 VGND 0.004984f
C7921 VDPWR.n1721 VGND 0.011445f
C7922 VDPWR.n1722 VGND 0.020115f
C7923 VDPWR.n1723 VGND 0.005888f
C7924 VDPWR.n1724 VGND 0.003488f
C7925 VDPWR.n1725 VGND 0.004416f
C7926 VDPWR.n1726 VGND 0.005612f
C7927 VDPWR.t469 VGND 0.005483f
C7928 VDPWR.n1727 VGND 0.006928f
C7929 VDPWR.n1728 VGND 0.012342f
C7930 VDPWR.n1729 VGND 0.012342f
C7931 VDPWR.n1730 VGND 0.005888f
C7932 VDPWR.n1731 VGND 0.003488f
C7933 VDPWR.n1732 VGND 0.003209f
C7934 VDPWR.n1733 VGND 0.034322f
C7935 VDPWR.n1734 VGND 0.002865f
C7936 VDPWR.t551 VGND 0.005483f
C7937 VDPWR.n1735 VGND 0.006928f
C7938 VDPWR.n1736 VGND 0.012342f
C7939 VDPWR.n1737 VGND 0.005888f
C7940 VDPWR.n1738 VGND 0.005888f
C7941 VDPWR.n1739 VGND 0.004544f
C7942 VDPWR.n1740 VGND 0.009777f
C7943 VDPWR.n1741 VGND 0.036592f
C7944 VDPWR.n1742 VGND 0.009361f
C7945 VDPWR.t470 VGND 0.005483f
C7946 VDPWR.n1743 VGND 0.006928f
C7947 VDPWR.n1744 VGND 0.012342f
C7948 VDPWR.n1745 VGND 0.012758f
C7949 VDPWR.n1746 VGND 0.002048f
C7950 VDPWR.n1747 VGND 0.001579f
C7951 VDPWR.n1748 VGND 0.001973f
C7952 VDPWR.n1749 VGND 0.00224f
C7953 VDPWR.n1750 VGND 0.002752f
C7954 VDPWR.n1751 VGND 0.001973f
C7955 VDPWR.n1752 VGND 0.003083f
C7956 VDPWR.n1753 VGND 0.003404f
C7957 VDPWR.n1754 VGND 0.140809f
C7958 VDPWR.n1755 VGND 0.003404f
C7959 VDPWR.n1756 VGND 0.003083f
C7960 VDPWR.n1757 VGND 0.002949f
C7961 VDPWR.n1758 VGND 0.002528f
C7962 VDPWR.n1759 VGND 0.003168f
C7963 VDPWR.n1760 VGND 0.017118f
C7964 VDPWR.t552 VGND 0.0055f
C7965 VDPWR.n1761 VGND 0.011274f
C7966 VDPWR.n1762 VGND 0.006252f
C7967 VDPWR.n1763 VGND 0.00224f
C7968 VDPWR.n1764 VGND 0.003146f
C7969 VDPWR.n1765 VGND 0.00425f
C7970 VDPWR.n1766 VGND 0.007049f
C7971 VDPWR.t753 VGND 0.0055f
C7972 VDPWR.n1767 VGND 0.011154f
C7973 VDPWR.n1768 VGND 0.004646f
C7974 VDPWR.t611 VGND 0.005483f
C7975 VDPWR.n1769 VGND 0.006928f
C7976 VDPWR.t1175 VGND 0.072626f
C7977 VDPWR.n1770 VGND 0.036592f
C7978 VDPWR.n1771 VGND 0.009361f
C7979 VDPWR.n1772 VGND 0.005888f
C7980 VDPWR.n1773 VGND 0.005888f
C7981 VDPWR.n1774 VGND 0.005568f
C7982 VDPWR.n1775 VGND 0.009777f
C7983 VDPWR.n1776 VGND 0.036592f
C7984 VDPWR.n1777 VGND 0.009361f
C7985 VDPWR.n1778 VGND 0.012758f
C7986 VDPWR.n1779 VGND 0.002048f
C7987 VDPWR.n1780 VGND 0.002944f
C7988 VDPWR.n1781 VGND 0.001973f
C7989 VDPWR.n1782 VGND 0.003083f
C7990 VDPWR.n1783 VGND 0.003404f
C7991 VDPWR.n1784 VGND 0.140809f
C7992 VDPWR.n1785 VGND 0.003404f
C7993 VDPWR.n1786 VGND 0.003083f
C7994 VDPWR.n1787 VGND 0.002949f
C7995 VDPWR.n1788 VGND 0.003904f
C7996 VDPWR.n1789 VGND 0.012758f
C7997 VDPWR.n1790 VGND 0.012342f
C7998 VDPWR.t754 VGND 0.005483f
C7999 VDPWR.n1791 VGND 0.006928f
C8000 VDPWR.n1792 VGND 0.004736f
C8001 VDPWR.n1793 VGND 0.003488f
C8002 VDPWR.n1794 VGND 0.00425f
C8003 VDPWR.n1795 VGND 0.004321f
C8004 VDPWR.t651 VGND 0.0055f
C8005 VDPWR.n1796 VGND 0.011154f
C8006 VDPWR.n1797 VGND 0.004646f
C8007 VDPWR.t575 VGND 0.005483f
C8008 VDPWR.n1798 VGND 0.006928f
C8009 VDPWR.n1799 VGND 0.009361f
C8010 VDPWR.n1800 VGND 0.005888f
C8011 VDPWR.n1801 VGND 0.005888f
C8012 VDPWR.n1802 VGND 0.009361f
C8013 VDPWR.n1803 VGND 0.009777f
C8014 VDPWR.n1804 VGND 0.036592f
C8015 VDPWR.n1805 VGND 0.009361f
C8016 VDPWR.n1806 VGND 0.005888f
C8017 VDPWR.n1807 VGND 0.005888f
C8018 VDPWR.n1808 VGND 0.003648f
C8019 VDPWR.n1809 VGND 0.012758f
C8020 VDPWR.t652 VGND 0.005483f
C8021 VDPWR.n1810 VGND 0.006928f
C8022 VDPWR.n1811 VGND 0.002944f
C8023 VDPWR.n1812 VGND 0.002048f
C8024 VDPWR.n1813 VGND 0.012342f
C8025 VDPWR.n1814 VGND 0.012758f
C8026 VDPWR.n1815 VGND 0.002048f
C8027 VDPWR.n1816 VGND 0.00224f
C8028 VDPWR.n1817 VGND 0.001973f
C8029 VDPWR.n1818 VGND 0.003083f
C8030 VDPWR.n1819 VGND 0.003404f
C8031 VDPWR.n1820 VGND 0.140809f
C8032 VDPWR.n1821 VGND 0.003404f
C8033 VDPWR.n1822 VGND 0.003083f
C8034 VDPWR.n1823 VGND 5.48e-19
C8035 VDPWR.n1824 VGND 0.003168f
C8036 VDPWR.n1825 VGND 0.015948f
C8037 VDPWR.t576 VGND 0.005504f
C8038 VDPWR.n1826 VGND 0.00626f
C8039 VDPWR.n1827 VGND 0.008018f
C8040 VDPWR.t1181 VGND 0.021195f
C8041 VDPWR.n1828 VGND 0.007844f
C8042 VDPWR.t745 VGND 0.004984f
C8043 VDPWR.n1829 VGND 0.003662f
C8044 VDPWR.n1830 VGND 0.002301f
C8045 VDPWR.n1831 VGND 0.002016f
C8046 VDPWR.n1832 VGND 0.006108f
C8047 VDPWR.n1833 VGND 0.012813f
C8048 VDPWR.n1834 VGND 0.016328f
C8049 VDPWR.t1219 VGND 0.072626f
C8050 VDPWR.n1835 VGND 0.033842f
C8051 VDPWR.n1836 VGND 0.004517f
C8052 VDPWR.n1837 VGND 0.002016f
C8053 VDPWR.n1838 VGND 0.005344f
C8054 VDPWR.n1839 VGND 0.003792f
C8055 VDPWR.n1840 VGND 0.007139f
C8056 VDPWR.n1841 VGND 0.007119f
C8057 VDPWR.n1842 VGND 0.003993f
C8058 VDPWR.n1843 VGND 0.005888f
C8059 VDPWR.n1844 VGND 0.005888f
C8060 VDPWR.n1845 VGND 0.004672f
C8061 VDPWR.n1846 VGND 0.007422f
C8062 VDPWR.t169 VGND 0.002785f
C8063 VDPWR.t27 VGND 0.00135f
C8064 VDPWR.n1847 VGND 0.00567f
C8065 VDPWR.n1848 VGND 0.006831f
C8066 VDPWR.n1849 VGND 0.005687f
C8067 VDPWR.n1850 VGND 0.007422f
C8068 VDPWR.n1851 VGND 0.002048f
C8069 VDPWR.n1852 VGND 0.001973f
C8070 VDPWR.n1853 VGND 0.002112f
C8071 VDPWR.n1854 VGND 0.00288f
C8072 VDPWR.n1855 VGND 0.001973f
C8073 VDPWR.n1856 VGND 0.003083f
C8074 VDPWR.n1857 VGND 0.003404f
C8075 VDPWR.n1858 VGND 0.00352f
C8076 VDPWR.n1859 VGND 0.00352f
C8077 VDPWR.n1860 VGND 0.003404f
C8078 VDPWR.n1861 VGND 0.003083f
C8079 VDPWR.n1862 VGND 0.001973f
C8080 VDPWR.n1863 VGND 0.002944f
C8081 VDPWR.n1864 VGND 0.001504f
C8082 VDPWR.n1865 VGND 0.003079f
C8083 VDPWR.n1866 VGND 0.001972f
C8084 VDPWR.n1867 VGND 0.0048f
C8085 VDPWR.n1868 VGND 0.005888f
C8086 VDPWR.n1869 VGND 0.005888f
C8087 VDPWR.n1870 VGND 0.001247f
C8088 VDPWR.n1871 VGND 0.00338f
C8089 VDPWR.t3 VGND 0.002834f
C8090 VDPWR.n1872 VGND 0.00693f
C8091 VDPWR.t937 VGND 0.0018f
C8092 VDPWR.t941 VGND 0.0018f
C8093 VDPWR.n1873 VGND 0.003905f
C8094 VDPWR.t907 VGND 0.0018f
C8095 VDPWR.t1 VGND 0.0018f
C8096 VDPWR.n1874 VGND 0.004032f
C8097 VDPWR.n1875 VGND 0.005167f
C8098 VDPWR.n1876 VGND 0.004501f
C8099 VDPWR.n1877 VGND 9.41e-19
C8100 VDPWR.n1878 VGND 0.005888f
C8101 VDPWR.n1879 VGND 0.005888f
C8102 VDPWR.n1880 VGND 0.003488f
C8103 VDPWR.n1881 VGND 0.002085f
C8104 VDPWR.n1882 VGND 0.001757f
C8105 VDPWR.n1883 VGND 0.00224f
C8106 VDPWR.n1884 VGND 0.007808f
C8107 VDPWR.n1885 VGND 7.36e-19
C8108 VDPWR.n1886 VGND 0.006896f
C8109 VDPWR.n1887 VGND 0.003083f
C8110 VDPWR.n1888 VGND 0.001579f
C8111 VDPWR.n1889 VGND 0.001973f
C8112 VDPWR.n1890 VGND 0.001472f
C8113 VDPWR.n1891 VGND 0.002944f
C8114 VDPWR.n1892 VGND 0.002048f
C8115 VDPWR.t603 VGND 0.005024f
C8116 VDPWR.t1242 VGND 0.010664f
C8117 VDPWR.n1894 VGND 0.027341f
C8118 VDPWR.t604 VGND 0.005024f
C8119 VDPWR.n1895 VGND 0.014893f
C8120 VDPWR.n1896 VGND 0.012262f
C8121 VDPWR.n1897 VGND 0.001376f
C8122 VDPWR.n1898 VGND 0.002885f
C8123 VDPWR.n1899 VGND 0.002112f
C8124 VDPWR.n1900 VGND 0.001973f
C8125 VDPWR.n1901 VGND 0.001579f
C8126 VDPWR.n1902 VGND 0.00352f
C8127 VDPWR.n1903 VGND 0.003404f
C8128 VDPWR.n1904 VGND 0.140809f
C8129 VDPWR.n1905 VGND 0.116061f
C8130 VDPWR.n1906 VGND 0.167264f
C8131 VDPWR.n1907 VGND 0.281618f
C8132 VDPWR.n1908 VGND 0.116061f
C8133 VDPWR.n1909 VGND 0.001579f
C8134 VDPWR.n1910 VGND 0.001973f
C8135 VDPWR.n1911 VGND 0.001472f
C8136 VDPWR.n1912 VGND 0.002048f
C8137 VDPWR.n1913 VGND 0.002944f
C8138 VDPWR.n1914 VGND 0.002048f
C8139 VDPWR.n1915 VGND 0.004863f
C8140 VDPWR.t45 VGND 0.00112f
C8141 VDPWR.t95 VGND -0.001177f
C8142 VDPWR.n1916 VGND 0.007456f
C8143 VDPWR.t1003 VGND 0.002785f
C8144 VDPWR.t66 VGND 0.00135f
C8145 VDPWR.n1917 VGND 0.00567f
C8146 VDPWR.n1918 VGND 0.004338f
C8147 VDPWR.n1919 VGND 0.00438f
C8148 VDPWR.n1920 VGND 0.001111f
C8149 VDPWR.t993 VGND 0.0018f
C8150 VDPWR.t995 VGND 0.0018f
C8151 VDPWR.n1921 VGND 0.004044f
C8152 VDPWR.n1922 VGND 0.017119f
C8153 VDPWR.t997 VGND 0.002834f
C8154 VDPWR.n1923 VGND 0.005888f
C8155 VDPWR.n1924 VGND 0.01283f
C8156 VDPWR.t1196 VGND 0.037391f
C8157 VDPWR.t606 VGND 0.004984f
C8158 VDPWR.n1925 VGND 0.06261f
C8159 VDPWR.n1926 VGND 0.016449f
C8160 VDPWR.t933 VGND 0.001867f
C8161 VDPWR.t48 VGND 0.002067f
C8162 VDPWR.n1927 VGND 0.003981f
C8163 VDPWR.t607 VGND 0.004984f
C8164 VDPWR.n1928 VGND 0.008777f
C8165 VDPWR.n1929 VGND 7.36e-19
C8166 VDPWR.n1930 VGND 0.001973f
C8167 VDPWR.n1931 VGND 0.00352f
C8168 VDPWR.n1932 VGND 0.001579f
C8169 VDPWR.n1933 VGND 0.001472f
C8170 VDPWR.n1934 VGND 0.002048f
C8171 VDPWR.n1935 VGND 0.002112f
C8172 VDPWR.n1936 VGND 0.005471f
C8173 VDPWR.t514 VGND 0.005024f
C8174 VDPWR.t1232 VGND 0.010664f
C8175 VDPWR.n1938 VGND 0.027341f
C8176 VDPWR.t515 VGND 0.005024f
C8177 VDPWR.n1939 VGND 0.014893f
C8178 VDPWR.t592 VGND 0.005024f
C8179 VDPWR.t1203 VGND 0.010664f
C8180 VDPWR.n1941 VGND 0.027341f
C8181 VDPWR.t593 VGND 0.005024f
C8182 VDPWR.n1942 VGND 0.014893f
C8183 VDPWR.n1943 VGND 0.001973f
C8184 VDPWR.n1944 VGND 0.003404f
C8185 VDPWR.n1945 VGND 0.003083f
C8186 VDPWR.n1946 VGND 0.002885f
C8187 VDPWR.n1947 VGND 0.001376f
C8188 VDPWR.n1948 VGND 0.012553f
C8189 VDPWR.n1949 VGND 0.002048f
C8190 VDPWR.n1950 VGND 0.002944f
C8191 VDPWR.n1951 VGND 0.001973f
C8192 VDPWR.n1952 VGND 0.001579f
C8193 VDPWR.n1953 VGND 0.00352f
C8194 VDPWR.n1954 VGND 0.003404f
C8195 VDPWR.n1955 VGND 0.003083f
C8196 VDPWR.n1956 VGND 0.001477f
C8197 VDPWR.n1957 VGND 0.004416f
C8198 VDPWR.n1958 VGND 0.014953f
C8199 VDPWR.n1959 VGND 0.007897f
C8200 VDPWR.n1960 VGND 0.009969f
C8201 VDPWR.n1961 VGND 0.012517f
C8202 VDPWR.n1962 VGND 0.005344f
C8203 VDPWR.n1963 VGND 0.002016f
C8204 VDPWR.n1964 VGND 0.006234f
C8205 VDPWR.n1965 VGND 0.00224f
C8206 VDPWR.n1966 VGND 0.006477f
C8207 VDPWR.t1018 VGND 7.56e-19
C8208 VDPWR.t935 VGND 7.56e-19
C8209 VDPWR.n1967 VGND 0.00175f
C8210 VDPWR.n1968 VGND 0.016544f
C8211 VDPWR.n1969 VGND 0.002085f
C8212 VDPWR.n1970 VGND 0.006766f
C8213 VDPWR.n1971 VGND 0.002949f
C8214 VDPWR.n1972 VGND 0.003083f
C8215 VDPWR.n1973 VGND 0.003404f
C8216 VDPWR.n1974 VGND 0.140809f
C8217 VDPWR.n1975 VGND 0.003404f
C8218 VDPWR.n1976 VGND 0.00352f
C8219 VDPWR.n1977 VGND 0.001579f
C8220 VDPWR.n1978 VGND 0.001973f
C8221 VDPWR.n1979 VGND 9.28e-19
C8222 VDPWR.n1980 VGND 0.001711f
C8223 VDPWR.t347 VGND 0.002467f
C8224 VDPWR.t1005 VGND 0.001867f
C8225 VDPWR.n1981 VGND 0.00469f
C8226 VDPWR.n1982 VGND 0.009342f
C8227 VDPWR.n1983 VGND 0.001643f
C8228 VDPWR.n1984 VGND 0.005888f
C8229 VDPWR.n1985 VGND 0.004416f
C8230 VDPWR.n1986 VGND 1.47e-19
C8231 VDPWR.n1987 VGND 0.004452f
C8232 VDPWR.n1988 VGND 0.001655f
C8233 VDPWR.t1014 VGND 0.001152f
C8234 VDPWR.t137 VGND 0.001152f
C8235 VDPWR.n1989 VGND 0.002399f
C8236 VDPWR.n1990 VGND 0.006697f
C8237 VDPWR.n1991 VGND 0.005344f
C8238 VDPWR.n1992 VGND 0.002016f
C8239 VDPWR.n1993 VGND 0.003488f
C8240 VDPWR.n1994 VGND 0.007364f
C8241 VDPWR.t660 VGND 0.005483f
C8242 VDPWR.n1995 VGND 0.011995f
C8243 VDPWR.n1996 VGND 0.020115f
C8244 VDPWR.n1997 VGND 0.015595f
C8245 VDPWR.n1998 VGND 0.005888f
C8246 VDPWR.n1999 VGND 0.004416f
C8247 VDPWR.n2000 VGND 0.008952f
C8248 VDPWR.n2001 VGND 0.016769f
C8249 VDPWR.n2002 VGND 0.003168f
C8250 VDPWR.n2003 VGND 5.48e-19
C8251 VDPWR.n2004 VGND 0.003083f
C8252 VDPWR.n2005 VGND 0.003404f
C8253 VDPWR.n2006 VGND 0.140809f
C8254 VDPWR.n2007 VGND 0.003404f
C8255 VDPWR.n2008 VGND 0.003083f
C8256 VDPWR.n2009 VGND 0.002757f
C8257 VDPWR.n2010 VGND 0.003648f
C8258 VDPWR.n2011 VGND 0.009777f
C8259 VDPWR.n2012 VGND 0.012758f
C8260 VDPWR.n2013 VGND 0.012342f
C8261 VDPWR.n2014 VGND 0.005888f
C8262 VDPWR.n2015 VGND 0.005344f
C8263 VDPWR.n2016 VGND 0.005756f
C8264 VDPWR.n2017 VGND 0.005803f
C8265 VDPWR.n2018 VGND 0.003488f
C8266 VDPWR.n2019 VGND 0.005888f
C8267 VDPWR.n2020 VGND 0.009777f
C8268 VDPWR.n2021 VGND 0.012758f
C8269 VDPWR.n2022 VGND 0.012342f
C8270 VDPWR.n2023 VGND 0.005888f
C8271 VDPWR.n2024 VGND 0.005344f
C8272 VDPWR.n2025 VGND 0.003488f
C8273 VDPWR.n2026 VGND 0.005803f
C8274 VDPWR.t751 VGND 0.005483f
C8275 VDPWR.n2027 VGND 0.006928f
C8276 VDPWR.n2028 VGND 0.012342f
C8277 VDPWR.n2029 VGND 0.009361f
C8278 VDPWR.n2030 VGND 0.003904f
C8279 VDPWR.n2031 VGND 0.002949f
C8280 VDPWR.n2032 VGND 0.003083f
C8281 VDPWR.n2033 VGND 0.003404f
C8282 VDPWR.n2034 VGND 0.00352f
C8283 VDPWR.n2035 VGND 0.00352f
C8284 VDPWR.n2036 VGND 0.003404f
C8285 VDPWR.n2037 VGND 0.003083f
C8286 VDPWR.n2038 VGND 0.002949f
C8287 VDPWR.n2039 VGND 0.004096f
C8288 VDPWR.n2040 VGND 0.005612f
C8289 VDPWR.n2041 VGND 0.008742f
C8290 VDPWR.n2042 VGND 0.003488f
C8291 VDPWR.n2043 VGND 0.005888f
C8292 VDPWR.n2044 VGND 0.005888f
C8293 VDPWR.n2045 VGND 0.020793f
C8294 VDPWR.n2046 VGND 0.020115f
C8295 VDPWR.t750 VGND 0.005483f
C8296 VDPWR.n2047 VGND 0.010606f
C8297 VDPWR.n2048 VGND 0.013537f
C8298 VDPWR.t448 VGND 0.004984f
C8299 VDPWR.n2049 VGND 0.029901f
C8300 VDPWR.t1249 VGND 0.017526f
C8301 VDPWR.n2050 VGND 0.03397f
C8302 VDPWR.n2051 VGND 0.007752f
C8303 VDPWR.n2052 VGND 0.001735f
C8304 VDPWR.n2053 VGND 0.009861f
C8305 VDPWR.n2054 VGND 0.005344f
C8306 VDPWR.n2055 VGND 0.004953f
C8307 VDPWR.n2056 VGND 0.003168f
C8308 VDPWR.n2057 VGND 0.002528f
C8309 VDPWR.n2058 VGND 0.006017f
C8310 VDPWR.t561 VGND 0.005483f
C8311 VDPWR.n2059 VGND 0.006928f
C8312 VDPWR.n2060 VGND 0.012342f
C8313 VDPWR.n2061 VGND 0.002048f
C8314 VDPWR.n2062 VGND 0.002944f
C8315 VDPWR.n2063 VGND 0.001973f
C8316 VDPWR.n2064 VGND 0.00352f
C8317 VDPWR.n2065 VGND 0.001579f
C8318 VDPWR.n2066 VGND 0.001973f
C8319 VDPWR.n2067 VGND 0.00224f
C8320 VDPWR.n2068 VGND 0.002752f
C8321 VDPWR.n2069 VGND 0.001973f
C8322 VDPWR.n2070 VGND 0.003083f
C8323 VDPWR.n2071 VGND 0.003404f
C8324 VDPWR.n2072 VGND 0.140809f
C8325 VDPWR.n2073 VGND 0.116061f
C8326 VDPWR.n2074 VGND 0.00352f
C8327 VDPWR.n2075 VGND 0.002949f
C8328 VDPWR.n2076 VGND 0.001579f
C8329 VDPWR.t1279 VGND 0.072626f
C8330 VDPWR.n2077 VGND 0.036592f
C8331 VDPWR.n2078 VGND 0.005888f
C8332 VDPWR.t1209 VGND 0.072626f
C8333 VDPWR.n2079 VGND 0.036175f
C8334 VDPWR.t494 VGND 0.005483f
C8335 VDPWR.n2080 VGND 0.006928f
C8336 VDPWR.n2081 VGND 0.004416f
C8337 VDPWR.t558 VGND 0.004984f
C8338 VDPWR.n2082 VGND 0.011445f
C8339 VDPWR.n2083 VGND 0.005888f
C8340 VDPWR.n2084 VGND 0.015256f
C8341 VDPWR.n2085 VGND 0.00288f
C8342 VDPWR.n2086 VGND 0.001973f
C8343 VDPWR.n2087 VGND 0.00352f
C8344 VDPWR.n2088 VGND 0.001579f
C8345 VDPWR.n2089 VGND 0.002368f
C8346 VDPWR.t1243 VGND 0.036876f
C8347 VDPWR.t557 VGND 0.004984f
C8348 VDPWR.n2090 VGND 0.011445f
C8349 VDPWR.t680 VGND 0.005101f
C8350 VDPWR.n2091 VGND 0.002138f
C8351 VDPWR.n2092 VGND 0.011656f
C8352 VDPWR.t1188 VGND 0.010699f
C8353 VDPWR.n2093 VGND 0.020574f
C8354 VDPWR.t679 VGND 0.005024f
C8355 VDPWR.n2094 VGND 0.007271f
C8356 VDPWR.n2095 VGND 0.007169f
C8357 VDPWR.t526 VGND 0.005024f
C8358 VDPWR.t1254 VGND 0.010664f
C8359 VDPWR.n2097 VGND 0.027341f
C8360 VDPWR.t527 VGND 0.005024f
C8361 VDPWR.n2098 VGND 0.014893f
C8362 VDPWR.t635 VGND 0.005024f
C8363 VDPWR.t1183 VGND 0.010664f
C8364 VDPWR.n2100 VGND 0.027341f
C8365 VDPWR.t636 VGND 0.005024f
C8366 VDPWR.n2101 VGND 0.014893f
C8367 VDPWR.n2102 VGND 0.01227f
C8368 VDPWR.n2103 VGND 0.003844f
C8369 VDPWR.n2104 VGND 0.003523f
C8370 VDPWR.n2105 VGND 0.002016f
C8371 VDPWR.n2106 VGND 0.002762f
C8372 VDPWR.t493 VGND 0.005503f
C8373 VDPWR.n2107 VGND 0.006102f
C8374 VDPWR.n2108 VGND 0.007518f
C8375 VDPWR.n2109 VGND 0.004416f
C8376 VDPWR.n2110 VGND 0.001973f
C8377 VDPWR.n2111 VGND 0.003404f
C8378 VDPWR.n2112 VGND 0.003083f
C8379 VDPWR.n2113 VGND 0.002629f
C8380 VDPWR.n2114 VGND 0.00352f
C8381 VDPWR.n2115 VGND 0.015143f
C8382 VDPWR.n2116 VGND 0.052403f
C8383 VDPWR.t1238 VGND 0.072626f
C8384 VDPWR.n2117 VGND 0.040608f
C8385 VDPWR.n2118 VGND 0.010509f
C8386 VDPWR.n2119 VGND 0.002048f
C8387 VDPWR.n2120 VGND 0.002048f
C8388 VDPWR.n2121 VGND 0.002944f
C8389 VDPWR.n2122 VGND 0.001973f
C8390 VDPWR.n2123 VGND 0.001579f
C8391 VDPWR.n2124 VGND 0.00352f
C8392 VDPWR.n2125 VGND 0.003404f
C8393 VDPWR.n2126 VGND 0.003083f
C8394 VDPWR.n2127 VGND 0.002117f
C8395 VDPWR.n2128 VGND 0.003008f
C8396 VDPWR.n2129 VGND 0.020793f
C8397 VDPWR.n2130 VGND 0.020793f
C8398 VDPWR.n2131 VGND 0.020115f
C8399 VDPWR.n2132 VGND 0.005888f
C8400 VDPWR.n2133 VGND 0.003488f
C8401 VDPWR.n2134 VGND 0.008742f
C8402 VDPWR.n2135 VGND 0.005612f
C8403 VDPWR.t641 VGND 0.005483f
C8404 VDPWR.n2136 VGND 0.006928f
C8405 VDPWR.n2137 VGND 0.011926f
C8406 VDPWR.n2138 VGND 0.005888f
C8407 VDPWR.n2139 VGND 0.003488f
C8408 VDPWR.n2140 VGND 0.005803f
C8409 VDPWR.t705 VGND 0.005483f
C8410 VDPWR.n2141 VGND 0.003947f
C8411 VDPWR.n2142 VGND 0.005756f
C8412 VDPWR.n2143 VGND 0.005344f
C8413 VDPWR.n2144 VGND 0.005888f
C8414 VDPWR.n2145 VGND 0.009361f
C8415 VDPWR.n2146 VGND 0.012758f
C8416 VDPWR.n2147 VGND 0.009777f
C8417 VDPWR.n2148 VGND 0.005888f
C8418 VDPWR.n2149 VGND 0.004544f
C8419 VDPWR.n2150 VGND 0.009361f
C8420 VDPWR.n2151 VGND 0.012758f
C8421 VDPWR.n2152 VGND 0.002048f
C8422 VDPWR.n2153 VGND 0.001973f
C8423 VDPWR.n2154 VGND 0.00224f
C8424 VDPWR.n2155 VGND 0.002752f
C8425 VDPWR.n2156 VGND 0.001973f
C8426 VDPWR.n2157 VGND 0.003083f
C8427 VDPWR.n2158 VGND 0.003404f
C8428 VDPWR.n2159 VGND 0.140809f
C8429 VDPWR.n2160 VGND 0.003404f
C8430 VDPWR.n2161 VGND 0.003083f
C8431 VDPWR.n2162 VGND 0.001973f
C8432 VDPWR.n2163 VGND 0.002944f
C8433 VDPWR.n2164 VGND 0.002048f
C8434 VDPWR.n2165 VGND 0.012342f
C8435 VDPWR.t642 VGND 0.005483f
C8436 VDPWR.n2166 VGND 0.006928f
C8437 VDPWR.n2167 VGND 0.006017f
C8438 VDPWR.n2168 VGND 0.002528f
C8439 VDPWR.n2169 VGND 0.003168f
C8440 VDPWR.n2170 VGND 0.00224f
C8441 VDPWR.n2171 VGND 0.006252f
C8442 VDPWR.t706 VGND 0.005503f
C8443 VDPWR.n2172 VGND 0.006241f
C8444 VDPWR.n2173 VGND 0.00232f
C8445 VDPWR.n2174 VGND 0.002016f
C8446 VDPWR.n2175 VGND 0.002944f
C8447 VDPWR.n2176 VGND 0.00168f
C8448 VDPWR.n2177 VGND 0.014269f
C8449 VDPWR.t1020 VGND 0.001867f
C8450 VDPWR.t259 VGND 0.001867f
C8451 VDPWR.n2178 VGND 0.004011f
C8452 VDPWR.t564 VGND 0.004984f
C8453 VDPWR.n2179 VGND 0.014116f
C8454 VDPWR.n2180 VGND 0.014701f
C8455 VDPWR.n2181 VGND 0.005344f
C8456 VDPWR.n2182 VGND 0.003488f
C8457 VDPWR.n2183 VGND 0.004416f
C8458 VDPWR.n2184 VGND 0.002878f
C8459 VDPWR.t433 VGND 0.005483f
C8460 VDPWR.n2185 VGND 0.003532f
C8461 VDPWR.n2186 VGND 0.008738f
C8462 VDPWR.n2187 VGND 0.004474f
C8463 VDPWR.n2188 VGND 0.006263f
C8464 VDPWR.n2189 VGND 0.005888f
C8465 VDPWR.n2190 VGND 0.005568f
C8466 VDPWR.n2191 VGND 0.003213f
C8467 VDPWR.n2192 VGND 0.033954f
C8468 VDPWR.n2193 VGND 0.003782f
C8469 VDPWR.n2194 VGND 0.008648f
C8470 VDPWR.t401 VGND 0.001867f
C8471 VDPWR.t423 VGND 0.001867f
C8472 VDPWR.n2195 VGND 0.003854f
C8473 VDPWR.n2196 VGND 0.008648f
C8474 VDPWR.n2197 VGND 0.002112f
C8475 VDPWR.n2198 VGND 0.005888f
C8476 VDPWR.t395 VGND 0.001867f
C8477 VDPWR.t399 VGND 0.0018f
C8478 VDPWR.n2199 VGND 0.003787f
C8479 VDPWR.n2200 VGND 0.00427f
C8480 VDPWR.t403 VGND 0.001867f
C8481 VDPWR.t413 VGND 0.001867f
C8482 VDPWR.n2201 VGND 0.003854f
C8483 VDPWR.n2202 VGND 0.008115f
C8484 VDPWR.t434 VGND 0.005483f
C8485 VDPWR.n2203 VGND 0.003762f
C8486 VDPWR.t407 VGND 0.001867f
C8487 VDPWR.t409 VGND 0.001867f
C8488 VDPWR.n2204 VGND 0.003854f
C8489 VDPWR.n2205 VGND 0.004861f
C8490 VDPWR.n2206 VGND 0.005888f
C8491 VDPWR.t737 VGND 0.005483f
C8492 VDPWR.n2207 VGND 0.00425f
C8493 VDPWR.t405 VGND 0.001867f
C8494 VDPWR.t415 VGND 0.001867f
C8495 VDPWR.n2208 VGND 0.003854f
C8496 VDPWR.t1173 VGND 0.072626f
C8497 VDPWR.n2209 VGND 0.033277f
C8498 VDPWR.t419 VGND 0.006558f
C8499 VDPWR.n2210 VGND 0.007607f
C8500 VDPWR.t728 VGND 0.004984f
C8501 VDPWR.n2211 VGND 0.006247f
C8502 VDPWR.n2212 VGND 0.008952f
C8503 VDPWR.n2213 VGND 0.002176f
C8504 VDPWR.n2214 VGND 0.00224f
C8505 VDPWR.n2215 VGND 0.007073f
C8506 VDPWR.n2216 VGND 0.004356f
C8507 VDPWR.n2217 VGND 0.004416f
C8508 VDPWR.n2218 VGND 0.005888f
C8509 VDPWR.n2219 VGND 0.005683f
C8510 VDPWR.n2220 VGND 0.004131f
C8511 VDPWR.n2221 VGND 0.008552f
C8512 VDPWR.n2222 VGND 0.006832f
C8513 VDPWR.n2223 VGND 0.005888f
C8514 VDPWR.n2224 VGND 0.005344f
C8515 VDPWR.n2225 VGND 0.002741f
C8516 VDPWR.n2226 VGND 0.002996f
C8517 VDPWR.n2227 VGND 0.003488f
C8518 VDPWR.n2228 VGND 0.005888f
C8519 VDPWR.n2229 VGND 0.005888f
C8520 VDPWR.n2230 VGND 0.006466f
C8521 VDPWR.n2231 VGND 0.008359f
C8522 VDPWR.n2232 VGND 0.004758f
C8523 VDPWR.n2233 VGND 0.005938f
C8524 VDPWR.n2234 VGND 0.003904f
C8525 VDPWR.n2235 VGND 0.001973f
C8526 VDPWR.n2236 VGND 0.00352f
C8527 VDPWR.n2237 VGND 0.001579f
C8528 VDPWR.n2238 VGND 0.001973f
C8529 VDPWR.n2239 VGND 0.003083f
C8530 VDPWR.n2240 VGND 0.002949f
C8531 VDPWR.n2241 VGND 0.002048f
C8532 VDPWR.n2242 VGND 0.005287f
C8533 VDPWR.n2243 VGND 0.00545f
C8534 VDPWR.n2244 VGND 0.002048f
C8535 VDPWR.n2245 VGND 0.002944f
C8536 VDPWR.n2246 VGND 0.001973f
C8537 VDPWR.n2247 VGND 0.003083f
C8538 VDPWR.n2248 VGND 0.003404f
C8539 VDPWR.n2249 VGND 0.140809f
C8540 VDPWR.n2250 VGND 0.116061f
C8541 VDPWR.n2251 VGND 0.281618f
C8542 VDPWR.n2252 VGND 0.281618f
C8543 VDPWR.n2253 VGND 0.281618f
C8544 VDPWR.n2254 VGND 0.167264f
C8545 VDPWR.n2255 VGND 0.116061f
C8546 VDPWR.n2256 VGND 0.140809f
C8547 VDPWR.n2257 VGND 0.003404f
C8548 VDPWR.n2258 VGND 0.00352f
C8549 VDPWR.n2259 VGND 0.00352f
C8550 VDPWR.n2260 VGND 0.001579f
C8551 VDPWR.n2261 VGND 0.001973f
C8552 VDPWR.n2262 VGND 0.001472f
C8553 VDPWR.n2263 VGND 7.36e-19
C8554 VDPWR.n2264 VGND 0.007329f
C8555 VDPWR.t591 VGND 0.005483f
C8556 VDPWR.n2265 VGND 0.011995f
C8557 VDPWR.n2266 VGND 0.020115f
C8558 VDPWR.n2267 VGND 0.015595f
C8559 VDPWR.n2268 VGND 0.005888f
C8560 VDPWR.n2269 VGND 0.004416f
C8561 VDPWR.n2270 VGND 0.008952f
C8562 VDPWR.n2271 VGND 0.004007f
C8563 VDPWR.n2272 VGND 0.004416f
C8564 VDPWR.n2273 VGND 0.005888f
C8565 VDPWR.n2274 VGND 0.006773f
C8566 VDPWR.n2275 VGND 0.004131f
C8567 VDPWR.n2276 VGND 0.008552f
C8568 VDPWR.n2277 VGND 0.005084f
C8569 VDPWR.n2278 VGND 0.005888f
C8570 VDPWR.n2279 VGND 0.005888f
C8571 VDPWR.n2280 VGND 0.005888f
C8572 VDPWR.n2281 VGND 0.006954f
C8573 VDPWR.n2282 VGND 0.008359f
C8574 VDPWR.n2283 VGND 0.004026f
C8575 VDPWR.t590 VGND 0.005483f
C8576 VDPWR.n2284 VGND 0.004291f
C8577 VDPWR.n2285 VGND 0.002441f
C8578 VDPWR.n2286 VGND 0.0048f
C8579 VDPWR.n2287 VGND 0.002405f
C8580 VDPWR.n2288 VGND 0.003083f
C8581 VDPWR.n2289 VGND 0.003404f
C8582 VDPWR.n2290 VGND 0.140809f
C8583 VDPWR.n2291 VGND 0.003404f
C8584 VDPWR.n2292 VGND 0.00352f
C8585 VDPWR.n2293 VGND 0.001579f
C8586 VDPWR.n2294 VGND 0.001973f
C8587 VDPWR.n2295 VGND 0.00288f
C8588 VDPWR.n2296 VGND 0.002048f
C8589 VDPWR.n2297 VGND 0.005287f
C8590 VDPWR.n2298 VGND 0.00545f
C8591 VDPWR.n2299 VGND 0.004672f
C8592 VDPWR.n2300 VGND 0.005888f
C8593 VDPWR.n2301 VGND 0.005888f
C8594 VDPWR.n2302 VGND 0.004962f
C8595 VDPWR.n2303 VGND 0.008648f
C8596 VDPWR.n2304 VGND 0.006263f
C8597 VDPWR.n2305 VGND 0.004474f
C8598 VDPWR.n2306 VGND 0.005888f
C8599 VDPWR.n2307 VGND 0.005888f
C8600 VDPWR.n2308 VGND 0.006418f
C8601 VDPWR.n2309 VGND 0.003953f
C8602 VDPWR.n2310 VGND 0.009049f
C8603 VDPWR.n2311 VGND 0.006938f
C8604 VDPWR.n2312 VGND 0.005344f
C8605 VDPWR.n2313 VGND 0.002016f
C8606 VDPWR.n2314 VGND 0.002016f
C8607 VDPWR.n2315 VGND 0.002963f
C8608 VDPWR.t738 VGND 0.005483f
C8609 VDPWR.n2316 VGND 0.00426f
C8610 VDPWR.n2317 VGND 0.016735f
C8611 VDPWR.n2318 VGND 0.00224f
C8612 VDPWR.n2319 VGND 5.48e-19
C8613 VDPWR.n2320 VGND 0.003083f
C8614 VDPWR.n2321 VGND 0.001973f
C8615 VDPWR.n2322 VGND 0.002944f
C8616 VDPWR.n2323 VGND 0.002048f
C8617 VDPWR.n2324 VGND 0.020115f
C8618 VDPWR.n2325 VGND 0.015595f
C8619 VDPWR.n2326 VGND 0.002048f
C8620 VDPWR.n2327 VGND 0.00224f
C8621 VDPWR.n2328 VGND 0.001973f
C8622 VDPWR.n2329 VGND 0.003083f
C8623 VDPWR.n2330 VGND 0.003404f
C8624 VDPWR.n2331 VGND 0.140809f
C8625 VDPWR.n2332 VGND 0.116061f
C8626 VDPWR.n2333 VGND 0.281618f
C8627 VDPWR.n2334 VGND 0.281618f
C8628 VDPWR.n2335 VGND 0.532156f
C8629 VDPWR.n2336 VGND 0.194931f
C8630 VDPWR.n2338 VGND 0.003432f
C8631 VDPWR.n2339 VGND 0.107527f
C8632 VDPWR.n2340 VGND 0.097681f
C8633 VDPWR.n2341 VGND 0.001579f
C8634 VDPWR.n2342 VGND 0.003054f
C8635 VDPWR.n2343 VGND 0.427843f
C8636 VDPWR.n2344 VGND 0.003054f
C8637 VDPWR.n2345 VGND 0.001973f
C8638 VDPWR.n2346 VGND 0.002949f
C8639 VDPWR.t802 VGND 0.001527f
C8640 VDPWR.t8 VGND 0.001527f
C8641 VDPWR.n2347 VGND 0.003322f
C8642 VDPWR.t1052 VGND 0.003924f
C8643 VDPWR.t374 VGND 0.002867f
C8644 VDPWR.n2348 VGND 0.010151f
C8645 VDPWR.n2349 VGND 0.005906f
C8646 VDPWR.n2350 VGND 0.005344f
C8647 VDPWR.t834 VGND 0.002741f
C8648 VDPWR.t1194 VGND 0.029301f
C8649 VDPWR.n2351 VGND 0.039775f
C8650 VDPWR.t353 VGND 0.0022f
C8651 VDPWR.t913 VGND 0.0022f
C8652 VDPWR.n2352 VGND 0.004485f
C8653 VDPWR.n2353 VGND 0.006511f
C8654 VDPWR.n2354 VGND 0.004416f
C8655 VDPWR.t296 VGND 0.001527f
C8656 VDPWR.t301 VGND 0.001527f
C8657 VDPWR.n2355 VGND 0.003394f
C8658 VDPWR.t21 VGND 0.002267f
C8659 VDPWR.t1050 VGND 0.002333f
C8660 VDPWR.n2356 VGND 0.005483f
C8661 VDPWR.t440 VGND 0.004984f
C8662 VDPWR.n2357 VGND 0.008777f
C8663 VDPWR.n2358 VGND 0.003008f
C8664 VDPWR.t1269 VGND 0.020799f
C8665 VDPWR.t389 VGND 0.00632f
C8666 VDPWR.n2359 VGND 0.005918f
C8667 VDPWR.n2360 VGND 0.001472f
C8668 VDPWR.n2361 VGND 0.002117f
C8669 VDPWR.n2362 VGND 0.001579f
C8670 VDPWR.n2363 VGND 0.001973f
C8671 VDPWR.n2364 VGND 0.001579f
C8672 VDPWR.n2365 VGND 0.002629f
C8673 VDPWR.t809 VGND 0.0018f
C8674 VDPWR.t806 VGND 0.0018f
C8675 VDPWR.n2366 VGND 0.003944f
C8676 VDPWR.n2367 VGND 0.00352f
C8677 VDPWR.t97 VGND 0.001527f
C8678 VDPWR.t808 VGND 0.001527f
C8679 VDPWR.n2368 VGND 0.003394f
C8680 VDPWR.n2369 VGND 0.001711f
C8681 VDPWR.t836 VGND 0.001527f
C8682 VDPWR.t141 VGND 0.001527f
C8683 VDPWR.n2370 VGND 0.003394f
C8684 VDPWR.t475 VGND 0.005024f
C8685 VDPWR.t1274 VGND 0.010664f
C8686 VDPWR.n2372 VGND 0.027341f
C8687 VDPWR.t476 VGND 0.005024f
C8688 VDPWR.n2373 VGND 0.014893f
C8689 VDPWR.t594 VGND 0.005024f
C8690 VDPWR.t1211 VGND 0.010664f
C8691 VDPWR.n2375 VGND 0.027341f
C8692 VDPWR.t595 VGND 0.005024f
C8693 VDPWR.n2376 VGND 0.014893f
C8694 VDPWR.n2377 VGND 0.012599f
C8695 VDPWR.n2378 VGND 0.003844f
C8696 VDPWR.n2379 VGND 0.002016f
C8697 VDPWR.n2380 VGND 0.001383f
C8698 VDPWR.n2381 VGND 0.009183f
C8699 VDPWR.n2382 VGND 0.0032f
C8700 VDPWR.n2383 VGND 0.002016f
C8701 VDPWR.n2384 VGND 0.004416f
C8702 VDPWR.n2385 VGND 0.001711f
C8703 VDPWR.n2386 VGND 0.012693f
C8704 VDPWR.n2387 VGND 8.61e-19
C8705 VDPWR.n2388 VGND 0.001792f
C8706 VDPWR.n2389 VGND 0.002368f
C8707 VDPWR.n2390 VGND 0.001973f
C8708 VDPWR.n2391 VGND 0.003054f
C8709 VDPWR.n2392 VGND 0.24535f
C8710 VDPWR.n2393 VGND 0.003054f
C8711 VDPWR.n2394 VGND 0.001973f
C8712 VDPWR.n2395 VGND 0.00288f
C8713 VDPWR.n2396 VGND 0.002048f
C8714 VDPWR.n2397 VGND 0.002847f
C8715 VDPWR.t439 VGND 0.004984f
C8716 VDPWR.n2398 VGND 0.004913f
C8717 VDPWR.n2399 VGND 0.018812f
C8718 VDPWR.n2400 VGND 0.011593f
C8719 VDPWR.n2401 VGND 0.014953f
C8720 VDPWR.n2402 VGND 0.004416f
C8721 VDPWR.n2403 VGND 0.002016f
C8722 VDPWR.n2404 VGND 0.005635f
C8723 VDPWR.n2405 VGND 0.008623f
C8724 VDPWR.n2406 VGND 0.008617f
C8725 VDPWR.n2407 VGND 0.005888f
C8726 VDPWR.n2408 VGND 0.004416f
C8727 VDPWR.n2409 VGND 0.00224f
C8728 VDPWR.n2410 VGND 0.001408f
C8729 VDPWR.t638 VGND 0.004984f
C8730 VDPWR.n2411 VGND 0.008777f
C8731 VDPWR.n2412 VGND 0.005906f
C8732 VDPWR.n2413 VGND 0.004416f
C8733 VDPWR.n2414 VGND 0.004416f
C8734 VDPWR.n2415 VGND 0.002016f
C8735 VDPWR.n2416 VGND 0.008233f
C8736 VDPWR.n2417 VGND 0.011294f
C8737 VDPWR.n2418 VGND 0.014953f
C8738 VDPWR.t1041 VGND 0.001036f
C8739 VDPWR.t357 VGND 0.001036f
C8740 VDPWR.n2419 VGND 0.002169f
C8741 VDPWR.t639 VGND 0.004984f
C8742 VDPWR.n2420 VGND 0.007433f
C8743 VDPWR.n2421 VGND 0.013464f
C8744 VDPWR.n2422 VGND 0.009073f
C8745 VDPWR.n2423 VGND 0.004544f
C8746 VDPWR.n2424 VGND 0.002949f
C8747 VDPWR.n2425 VGND 0.001888f
C8748 VDPWR.n2426 VGND 0.001973f
C8749 VDPWR.n2427 VGND 9.28e-19
C8750 VDPWR.n2428 VGND 0.001472f
C8751 VDPWR.n2429 VGND 7.36e-19
C8752 VDPWR.n2430 VGND 0.001782f
C8753 VDPWR.n2431 VGND 0.007807f
C8754 VDPWR.t474 VGND 0.052075f
C8755 VDPWR.t835 VGND 0.017547f
C8756 VDPWR.t140 VGND 0.01717f
C8757 VDPWR.t387 VGND 0.023208f
C8758 VDPWR.t96 VGND 0.031698f
C8759 VDPWR.t805 VGND 0.016604f
C8760 VDPWR.t807 VGND 0.013019f
C8761 VDPWR.t388 VGND 0.038302f
C8762 VDPWR.t167 VGND 0.037358f
C8763 VDPWR.t438 VGND 0.031132f
C8764 VDPWR.t20 VGND 0.01717f
C8765 VDPWR.t295 VGND 0.007358f
C8766 VDPWR.t1049 VGND 0.016604f
C8767 VDPWR.t300 VGND 0.017736f
C8768 VDPWR.t352 VGND 0.020755f
C8769 VDPWR.t912 VGND 0.026604f
C8770 VDPWR.t837 VGND 0.052453f
C8771 VDPWR.t637 VGND 0.005849f
C8772 VDPWR.t833 VGND 0.019245f
C8773 VDPWR.t1040 VGND 0.038491f
C8774 VDPWR.t356 VGND 0.027358f
C8775 VDPWR.t1051 VGND 0.017358f
C8776 VDPWR.t801 VGND 0.022453f
C8777 VDPWR.t7 VGND 0.043019f
C8778 VDPWR.t51 VGND 0.019057f
C8779 VDPWR.t870 VGND 0.016604f
C8780 VDPWR.t124 VGND 0.01566f
C8781 VDPWR.t126 VGND 0.017358f
C8782 VDPWR.t846 VGND 0.029245f
C8783 VDPWR.t733 VGND 0.031509f
C8784 VDPWR.t63 VGND 0.045849f
C8785 VDPWR.t159 VGND 0.022453f
C8786 VDPWR.t510 VGND 0.017358f
C8787 VDPWR.t670 VGND 0.103962f
C8788 VDPWR.t922 VGND 0.045849f
C8789 VDPWR.t223 VGND 0.017358f
C8790 VDPWR.t229 VGND 0.005849f
C8791 VDPWR.t297 VGND 0.025094f
C8792 VDPWR.t799 VGND 0.035849f
C8793 VDPWR.t227 VGND 0.021509f
C8794 VDPWR.t480 VGND 0.018868f
C8795 VDPWR.t324 VGND 0.02283f
C8796 VDPWR.n2432 VGND 0.053108f
C8797 VDPWR.n2433 VGND 0.022154f
C8798 VDPWR.t1255 VGND 0.029301f
C8799 VDPWR.t325 VGND 0.002741f
C8800 VDPWR.n2434 VGND 0.011294f
C8801 VDPWR.n2435 VGND 0.005888f
C8802 VDPWR.t228 VGND 0.001036f
C8803 VDPWR.t800 VGND 0.001036f
C8804 VDPWR.n2436 VGND 0.002169f
C8805 VDPWR.t482 VGND 0.004984f
C8806 VDPWR.n2437 VGND 0.008777f
C8807 VDPWR.t298 VGND 0.003924f
C8808 VDPWR.t230 VGND 0.002867f
C8809 VDPWR.n2438 VGND 0.010226f
C8810 VDPWR.n2439 VGND 0.002016f
C8811 VDPWR.n2440 VGND 0.003872f
C8812 VDPWR.t224 VGND 0.001527f
C8813 VDPWR.t923 VGND 0.001527f
C8814 VDPWR.n2441 VGND 0.003394f
C8815 VDPWR.n2442 VGND 0.002505f
C8816 VDPWR.n2443 VGND 0.001088f
C8817 VDPWR.n2444 VGND 0.001973f
C8818 VDPWR.n2445 VGND 0.001579f
C8819 VDPWR.n2446 VGND 0.003054f
C8820 VDPWR.n2447 VGND 0.001472f
C8821 VDPWR.n2448 VGND 0.002048f
C8822 VDPWR.n2449 VGND 0.002949f
C8823 VDPWR.t671 VGND 0.004984f
C8824 VDPWR.t511 VGND 0.005483f
C8825 VDPWR.n2450 VGND 0.011995f
C8826 VDPWR.n2451 VGND 0.003842f
C8827 VDPWR.n2452 VGND 0.003295f
C8828 VDPWR.t1182 VGND 0.029107f
C8829 VDPWR.n2453 VGND 0.015278f
C8830 VDPWR.n2454 VGND 0.015934f
C8831 VDPWR.n2455 VGND 0.003488f
C8832 VDPWR.t1264 VGND 0.072626f
C8833 VDPWR.n2456 VGND 0.040608f
C8834 VDPWR.n2457 VGND 0.004416f
C8835 VDPWR.t160 VGND 0.001527f
C8836 VDPWR.t64 VGND 0.001527f
C8837 VDPWR.n2458 VGND 0.003322f
C8838 VDPWR.t512 VGND 0.005501f
C8839 VDPWR.n2459 VGND 0.011323f
C8840 VDPWR.n2460 VGND 0.00425f
C8841 VDPWR.t127 VGND 0.001513f
C8842 VDPWR.t847 VGND 5.64e-19
C8843 VDPWR.n2461 VGND 0.006953f
C8844 VDPWR.t125 VGND 0.001527f
C8845 VDPWR.t52 VGND 0.001527f
C8846 VDPWR.n2462 VGND 0.003322f
C8847 VDPWR.n2463 VGND 0.008065f
C8848 VDPWR.n2464 VGND 9.32e-19
C8849 VDPWR.n2465 VGND 0.001973f
C8850 VDPWR.n2466 VGND 0.001472f
C8851 VDPWR.n2467 VGND 0.0024f
C8852 VDPWR.n2468 VGND 7.36e-19
C8853 VDPWR.n2469 VGND 0.001235f
C8854 VDPWR.n2470 VGND 0.015495f
C8855 VDPWR.t735 VGND 0.005058f
C8856 VDPWR.n2471 VGND 0.005913f
C8857 VDPWR.n2472 VGND 0.023007f
C8858 VDPWR.t1280 VGND 0.021124f
C8859 VDPWR.n2473 VGND 0.020912f
C8860 VDPWR.t734 VGND 0.004984f
C8861 VDPWR.n2474 VGND 0.005999f
C8862 VDPWR.n2475 VGND 0.00595f
C8863 VDPWR.n2476 VGND 0.003146f
C8864 VDPWR.n2477 VGND 0.00224f
C8865 VDPWR.n2478 VGND 0.006252f
C8866 VDPWR.n2479 VGND 0.007422f
C8867 VDPWR.n2480 VGND 0.013157f
C8868 VDPWR.n2481 VGND 0.005888f
C8869 VDPWR.n2482 VGND 0.004416f
C8870 VDPWR.n2483 VGND 0.004047f
C8871 VDPWR.n2484 VGND 0.008952f
C8872 VDPWR.t672 VGND 0.004984f
C8873 VDPWR.n2485 VGND 0.011445f
C8874 VDPWR.n2486 VGND 0.014578f
C8875 VDPWR.n2487 VGND 0.005888f
C8876 VDPWR.n2488 VGND 0.005888f
C8877 VDPWR.n2489 VGND 0.003904f
C8878 VDPWR.n2490 VGND 0.02068f
C8879 VDPWR.n2491 VGND 0.020136f
C8880 VDPWR.n2492 VGND 0.009831f
C8881 VDPWR.n2493 VGND 0.002048f
C8882 VDPWR.n2494 VGND 0.001973f
C8883 VDPWR.n2495 VGND 0.002112f
C8884 VDPWR.n2496 VGND 0.00288f
C8885 VDPWR.n2497 VGND 0.001973f
C8886 VDPWR.n2498 VGND 0.001579f
C8887 VDPWR.n2499 VGND 0.116061f
C8888 VDPWR.n2500 VGND 0.097057f
C8889 VDPWR.n2501 VGND 0.139727f
C8890 VDPWR.n2502 VGND 0.293684f
C8891 VDPWR.n2503 VGND 0.061977f
C8892 VDPWR.n2504 VGND 0.532156f
C8893 VDPWR.n2505 VGND 0.281618f
C8894 VDPWR.n2506 VGND 0.063151f
C8895 VDPWR.n2507 VGND 0.140809f
C8896 VDPWR.n2508 VGND 0.078917f
C8897 VDPWR.n2509 VGND 0.003054f
C8898 VDPWR.n2510 VGND 0.001477f
C8899 VDPWR.n2511 VGND 0.002944f
C8900 VDPWR.n2512 VGND 0.001711f
C8901 VDPWR.n2513 VGND 0.008968f
C8902 VDPWR.n2514 VGND 0.009333f
C8903 VDPWR.n2515 VGND 0.005043f
C8904 VDPWR.n2516 VGND 0.003488f
C8905 VDPWR.n2517 VGND 0.005888f
C8906 VDPWR.n2518 VGND 0.013609f
C8907 VDPWR.n2519 VGND 0.013968f
C8908 VDPWR.n2520 VGND 0.009073f
C8909 VDPWR.n2521 VGND 0.014953f
C8910 VDPWR.n2522 VGND 0.005344f
C8911 VDPWR.n2523 VGND 0.002016f
C8912 VDPWR.n2524 VGND 0.03255f
C8913 VDPWR.t481 VGND 0.004984f
C8914 VDPWR.n2525 VGND 0.008777f
C8915 VDPWR.n2526 VGND 0.005471f
C8916 VDPWR.n2527 VGND 0.00224f
C8917 VDPWR.n2528 VGND 0.00224f
C8918 VDPWR.n2529 VGND 0.003456f
C8919 VDPWR.n2530 VGND 0.001757f
C8920 VDPWR.n2531 VGND 0.007623f
C8921 VDPWR.n2532 VGND 0.002048f
C8922 VDPWR.n2533 VGND 0.0024f
C8923 VDPWR.n2534 VGND 0.001973f
C8924 VDPWR.n2535 VGND 0.001579f
C8925 VDPWR.n2536 VGND 0.081339f
C8926 VDPWR.n2537 VGND 0.107527f
C8927 VDPWR.n2538 VGND 0.116061f
C8928 VDPWR.n2539 VGND 0.532156f
C8929 VDPWR.n2540 VGND 0.194931f
C8930 VDPWR.n2541 VGND 0.00352f
C8931 VDPWR.n2542 VGND 0.001973f
C8932 VDPWR.n2543 VGND 0.00288f
C8933 VDPWR.n2544 VGND 0.005888f
C8934 VDPWR.t832 VGND 0.0018f
C8935 VDPWR.t321 VGND 0.0018f
C8936 VDPWR.n2545 VGND 0.004032f
C8937 VDPWR.t1144 VGND 0.0018f
C8938 VDPWR.t330 VGND 0.0018f
C8939 VDPWR.n2546 VGND 0.004032f
C8940 VDPWR.n2547 VGND 0.009337f
C8941 VDPWR.n2548 VGND 0.002048f
C8942 VDPWR.n2549 VGND 0.003054f
C8943 VDPWR.t707 VGND 0.005024f
C8944 VDPWR.t1179 VGND 0.010664f
C8945 VDPWR.n2551 VGND 0.027341f
C8946 VDPWR.t708 VGND 0.005024f
C8947 VDPWR.n2552 VGND 0.014893f
C8948 VDPWR.t490 VGND 0.005024f
C8949 VDPWR.t1278 VGND 0.010664f
C8950 VDPWR.n2554 VGND 0.027341f
C8951 VDPWR.t491 VGND 0.005024f
C8952 VDPWR.n2555 VGND 0.014893f
C8953 VDPWR.n2556 VGND 0.01227f
C8954 VDPWR.t720 VGND 0.004984f
C8955 VDPWR.t1176 VGND 0.020982f
C8956 VDPWR.n2558 VGND 0.036453f
C8957 VDPWR.t721 VGND 0.004984f
C8958 VDPWR.n2559 VGND 0.020917f
C8959 VDPWR.n2560 VGND 0.003844f
C8960 VDPWR.n2561 VGND 0.006902f
C8961 VDPWR.t499 VGND 0.004984f
C8962 VDPWR.t1276 VGND 0.020982f
C8963 VDPWR.n2563 VGND 0.036453f
C8964 VDPWR.t500 VGND 0.004984f
C8965 VDPWR.n2564 VGND 0.020917f
C8966 VDPWR.n2565 VGND 0.018023f
C8967 VDPWR.n2566 VGND 0.001133f
C8968 VDPWR.n2567 VGND 0.001757f
C8969 VDPWR.n2568 VGND 0.002048f
C8970 VDPWR.n2569 VGND 0.002629f
C8971 VDPWR.n2570 VGND 0.002368f
C8972 VDPWR.n2571 VGND 0.001973f
C8973 VDPWR.n2572 VGND 0.00352f
C8974 VDPWR.n2573 VGND 0.001579f
C8975 VDPWR.n2574 VGND 0.001579f
C8976 VDPWR.n2575 VGND 0.001973f
C8977 VDPWR.n2576 VGND 0.002944f
C8978 VDPWR.n2577 VGND 0.002048f
C8979 VDPWR.n2578 VGND 0.00187f
C8980 VDPWR.t830 VGND 0.002834f
C8981 VDPWR.t1145 VGND 0.002834f
C8982 VDPWR.n2579 VGND 0.002085f
C8983 VDPWR.n2580 VGND 0.005888f
C8984 VDPWR.t818 VGND 0.00135f
C8985 VDPWR.t794 VGND 0.002785f
C8986 VDPWR.n2581 VGND 0.00567f
C8987 VDPWR.t199 VGND 0.00135f
C8988 VDPWR.t201 VGND 0.002785f
C8989 VDPWR.n2582 VGND 0.00567f
C8990 VDPWR.n2583 VGND 0.002085f
C8991 VDPWR.n2584 VGND 0.005888f
C8992 VDPWR.t12 VGND 0.002776f
C8993 VDPWR.t264 VGND 0.002776f
C8994 VDPWR.t770 VGND 0.001152f
C8995 VDPWR.t787 VGND 0.001152f
C8996 VDPWR.n2585 VGND 0.002399f
C8997 VDPWR.t148 VGND 0.001152f
C8998 VDPWR.t784 VGND 0.001152f
C8999 VDPWR.n2586 VGND 0.002399f
C9000 VDPWR.n2587 VGND 0.011445f
C9001 VDPWR.n2588 VGND 0.001888f
C9002 VDPWR.n2589 VGND 0.001973f
C9003 VDPWR.n2590 VGND 0.001579f
C9004 VDPWR.n2591 VGND 0.001579f
C9005 VDPWR.n2592 VGND 0.001973f
C9006 VDPWR.n2593 VGND 0.002048f
C9007 VDPWR.n2594 VGND 0.00136f
C9008 VDPWR.t496 VGND 0.005024f
C9009 VDPWR.t1267 VGND 0.010664f
C9010 VDPWR.n2596 VGND 0.027341f
C9011 VDPWR.t497 VGND 0.005024f
C9012 VDPWR.n2597 VGND 0.014893f
C9013 VDPWR.n2598 VGND 9.28e-19
C9014 VDPWR.n2599 VGND 0.001973f
C9015 VDPWR.n2600 VGND 0.001472f
C9016 VDPWR.n2601 VGND 0.002944f
C9017 VDPWR.n2602 VGND 0.002048f
C9018 VDPWR.t319 VGND 0.0018f
C9019 VDPWR.t769 VGND 0.0018f
C9020 VDPWR.n2603 VGND 0.004047f
C9021 VDPWR.n2604 VGND 0.00224f
C9022 VDPWR.t317 VGND 0.00281f
C9023 VDPWR.n2605 VGND 0.001133f
C9024 VDPWR.n2606 VGND 0.005888f
C9025 VDPWR.t384 VGND 0.0018f
C9026 VDPWR.t1140 VGND 0.0018f
C9027 VDPWR.n2607 VGND 0.004032f
C9028 VDPWR.n2608 VGND 0.00519f
C9029 VDPWR.t382 VGND 0.00281f
C9030 VDPWR.t284 VGND 0.00135f
C9031 VDPWR.t376 VGND 0.002785f
C9032 VDPWR.n2609 VGND 0.00567f
C9033 VDPWR.n2610 VGND 0.002085f
C9034 VDPWR.n2611 VGND 0.005888f
C9035 VDPWR.t139 VGND 0.00135f
C9036 VDPWR.t1001 VGND 0.002785f
C9037 VDPWR.n2612 VGND 0.00567f
C9038 VDPWR.n2613 VGND 0.001349f
C9039 VDPWR.n2614 VGND 0.002048f
C9040 VDPWR.n2615 VGND 0.001973f
C9041 VDPWR.n2616 VGND 0.001579f
C9042 VDPWR.n2617 VGND 0.001579f
C9043 VDPWR.n2618 VGND 0.001973f
C9044 VDPWR.t82 VGND 0.001152f
C9045 VDPWR.t786 VGND 0.001152f
C9046 VDPWR.n2619 VGND 0.002399f
C9047 VDPWR.n2620 VGND 0.006924f
C9048 VDPWR.t35 VGND 0.002765f
C9049 VDPWR.n2621 VGND 0.001723f
C9050 VDPWR.n2622 VGND 0.007854f
C9051 VDPWR.t359 VGND 0.002333f
C9052 VDPWR.t193 VGND 0.002267f
C9053 VDPWR.n2623 VGND 0.005406f
C9054 VDPWR.n2624 VGND 0.004863f
C9055 VDPWR.t351 VGND 7.56e-19
C9056 VDPWR.t101 VGND 7.56e-19
C9057 VDPWR.n2625 VGND 0.00175f
C9058 VDPWR.t355 VGND 0.001513f
C9059 VDPWR.t1133 VGND 5.64e-19
C9060 VDPWR.n2626 VGND 0.006904f
C9061 VDPWR.n2627 VGND 0.009598f
C9062 VDPWR.t484 VGND 0.004984f
C9063 VDPWR.n2628 VGND 0.004577f
C9064 VDPWR.n2629 VGND 0.005906f
C9065 VDPWR.n2630 VGND 0.002176f
C9066 VDPWR.n2631 VGND 0.001984f
C9067 VDPWR.n2632 VGND 0.001612f
C9068 VDPWR.n2633 VGND 0.023712f
C9069 VDPWR.t1026 VGND 0.0022f
C9070 VDPWR.t99 VGND 0.0022f
C9071 VDPWR.n2634 VGND 0.004485f
C9072 VDPWR.n2635 VGND 0.006669f
C9073 VDPWR.t756 VGND 0.00112f
C9074 VDPWR.t33 VGND -0.001177f
C9075 VDPWR.n2636 VGND 0.007481f
C9076 VDPWR.n2637 VGND 0.005999f
C9077 VDPWR.n2638 VGND 0.005888f
C9078 VDPWR.n2639 VGND 0.004416f
C9079 VDPWR.n2640 VGND 0.002944f
C9080 VDPWR.n2641 VGND 0.001723f
C9081 VDPWR.t798 VGND 0.00112f
C9082 VDPWR.t791 VGND -0.001177f
C9083 VDPWR.n2642 VGND 0.007481f
C9084 VDPWR.n2643 VGND 0.006135f
C9085 VDPWR.n2644 VGND 0.003488f
C9086 VDPWR.n2645 VGND 0.005888f
C9087 VDPWR.n2646 VGND 0.005344f
C9088 VDPWR.t1030 VGND 7.56e-19
C9089 VDPWR.t222 VGND 7.56e-19
C9090 VDPWR.n2647 VGND 0.00175f
C9091 VDPWR.t144 VGND 0.001152f
C9092 VDPWR.t323 VGND 0.001152f
C9093 VDPWR.n2648 VGND 0.002399f
C9094 VDPWR.n2649 VGND 0.007139f
C9095 VDPWR.n2650 VGND 0.002944f
C9096 VDPWR.n2651 VGND 0.002048f
C9097 VDPWR.n2652 VGND 0.001973f
C9098 VDPWR.n2653 VGND 0.00288f
C9099 VDPWR.n2654 VGND 0.002112f
C9100 VDPWR.n2655 VGND 6.08e-19
C9101 VDPWR.n2656 VGND 0.00136f
C9102 VDPWR.n2657 VGND 0.020179f
C9103 VDPWR.n2658 VGND 0.001504f
C9104 VDPWR.n2659 VGND 0.001477f
C9105 VDPWR.n2660 VGND 0.003083f
C9106 VDPWR.n2661 VGND 0.003404f
C9107 VDPWR.n2662 VGND 0.00352f
C9108 VDPWR.n2663 VGND 0.00352f
C9109 VDPWR.n2664 VGND 0.003404f
C9110 VDPWR.n2665 VGND 0.003083f
C9111 VDPWR.n2666 VGND 0.002949f
C9112 VDPWR.n2667 VGND 0.005568f
C9113 VDPWR.t1161 VGND 0.002776f
C9114 VDPWR.n2668 VGND 0.005585f
C9115 VDPWR.n2669 VGND 0.00419f
C9116 VDPWR.n2670 VGND 0.00153f
C9117 VDPWR.n2671 VGND 0.002085f
C9118 VDPWR.n2672 VGND 0.005888f
C9119 VDPWR.n2673 VGND 0.005888f
C9120 VDPWR.n2674 VGND 0.005888f
C9121 VDPWR.n2675 VGND 0.001598f
C9122 VDPWR.n2676 VGND 0.004168f
C9123 VDPWR.n2677 VGND 0.004846f
C9124 VDPWR.n2678 VGND 0.001281f
C9125 VDPWR.n2679 VGND 0.001995f
C9126 VDPWR.n2680 VGND 0.005888f
C9127 VDPWR.n2681 VGND 0.005888f
C9128 VDPWR.n2682 VGND 0.004416f
C9129 VDPWR.n2683 VGND 0.001847f
C9130 VDPWR.n2684 VGND 0.005401f
C9131 VDPWR.t489 VGND 0.074905f
C9132 VDPWR.t498 VGND 0.09f
C9133 VDPWR.t831 VGND 0.040943f
C9134 VDPWR.t320 VGND 0.055472f
C9135 VDPWR.t829 VGND 0.061132f
C9136 VDPWR.t152 VGND 0.037358f
C9137 VDPWR.t150 VGND 0.033774f
C9138 VDPWR.t198 VGND 0.04283f
C9139 VDPWR.t200 VGND 0.04434f
C9140 VDPWR.t149 VGND 0.037358f
C9141 VDPWR.t151 VGND 0.033962f
C9142 VDPWR.t11 VGND 0.051509f
C9143 VDPWR.t147 VGND 0.051321f
C9144 VDPWR.t783 VGND 0.024906f
C9145 VDPWR.t318 VGND 0.031509f
C9146 VDPWR.t495 VGND 0.015849f
C9147 VDPWR.t768 VGND 0.020566f
C9148 VDPWR.t914 VGND 0.029245f
C9149 VDPWR.t483 VGND 0.015849f
C9150 VDPWR.t354 VGND 0.026038f
C9151 VDPWR.t1132 VGND 0.034717f
C9152 VDPWR.t192 VGND 0.01717f
C9153 VDPWR.t100 VGND 0.013774f
C9154 VDPWR.t358 VGND 0.015849f
C9155 VDPWR.t350 VGND 0.017736f
C9156 VDPWR.t98 VGND 0.017547f
C9157 VDPWR.t755 VGND 0.018113f
C9158 VDPWR.t1025 VGND 0.017924f
C9159 VDPWR.t32 VGND 0.018113f
C9160 VDPWR.t220 VGND 0.035472f
C9161 VDPWR.t790 VGND 0.036415f
C9162 VDPWR.t785 VGND 0.009623f
C9163 VDPWR.t797 VGND 0.015849f
C9164 VDPWR.t81 VGND 0.017547f
C9165 VDPWR.t221 VGND 0.018113f
C9166 VDPWR.t1029 VGND 0.021698f
C9167 VDPWR.t34 VGND 0.017358f
C9168 VDPWR.t816 VGND 0.009057f
C9169 VDPWR.t322 VGND 0.017924f
C9170 VDPWR.t80 VGND 0.035283f
C9171 VDPWR.t1000 VGND 0.035472f
C9172 VDPWR.t1160 VGND 0.024906f
C9173 VDPWR.t138 VGND 0.016038f
C9174 VDPWR.t766 VGND 0.017924f
C9175 VDPWR.t83 VGND 0.017924f
C9176 VDPWR.t143 VGND 0.015849f
C9177 VDPWR.t817 VGND 0.019434f
C9178 VDPWR.t375 VGND 0.021509f
C9179 VDPWR.t381 VGND 0.024906f
C9180 VDPWR.t283 VGND 0.032075f
C9181 VDPWR.t142 VGND 0.025472f
C9182 VDPWR.t1139 VGND 0.015849f
C9183 VDPWR.t767 VGND 0.015849f
C9184 VDPWR.t383 VGND 0.021509f
C9185 VDPWR.t316 VGND 0.028302f
C9186 VDPWR.n2685 VGND 0.031563f
C9187 VDPWR.n2686 VGND 0.010857f
C9188 VDPWR.n2687 VGND 0.014434f
C9189 VDPWR.n2688 VGND 0.002528f
C9190 VDPWR.n2689 VGND 0.002949f
C9191 VDPWR.n2690 VGND 0.003083f
C9192 VDPWR.n2691 VGND 0.003404f
C9193 VDPWR.n2692 VGND 0.00352f
C9194 VDPWR.n2693 VGND 0.00352f
C9195 VDPWR.n2694 VGND 0.003404f
C9196 VDPWR.n2695 VGND 0.003083f
C9197 VDPWR.n2696 VGND 0.002949f
C9198 VDPWR.n2697 VGND 0.004544f
C9199 VDPWR.n2698 VGND 0.005888f
C9200 VDPWR.n2699 VGND 0.001349f
C9201 VDPWR.n2700 VGND 0.009459f
C9202 VDPWR.n2701 VGND 0.00187f
C9203 VDPWR.n2702 VGND 0.005888f
C9204 VDPWR.n2703 VGND 0.005888f
C9205 VDPWR.n2704 VGND 0.005888f
C9206 VDPWR.n2705 VGND 0.002085f
C9207 VDPWR.n2706 VGND 0.001598f
C9208 VDPWR.n2707 VGND 0.007769f
C9209 VDPWR.n2708 VGND 0.00153f
C9210 VDPWR.n2709 VGND 0.005888f
C9211 VDPWR.n2710 VGND 0.005888f
C9212 VDPWR.n2711 VGND 0.005888f
C9213 VDPWR.n2712 VGND 0.002085f
C9214 VDPWR.n2713 VGND 0.001496f
C9215 VDPWR.n2714 VGND 0.011469f
C9216 VDPWR.n2715 VGND 0.003008f
C9217 VDPWR.n2716 VGND 0.002117f
C9218 VDPWR.n2717 VGND 0.003054f
C9219 VDPWR.n2718 VGND 0.003432f
C9220 VDPWR.n2719 VGND 0.128008f
C9221 VDPWR.n2720 VGND 0.00352f
C9222 VDPWR.n2721 VGND 0.007212f
C9223 VDPWR.n2722 VGND 0.001579f
C9224 VDPWR.n2723 VGND 0.001579f
C9225 VDPWR.n2724 VGND 0.001973f
C9226 VDPWR.n2725 VGND 0.002944f
C9227 VDPWR.n2726 VGND 0.016028f
C9228 VDPWR.t1204 VGND 0.037597f
C9229 VDPWR.n2727 VGND 0.067773f
C9230 VDPWR.t572 VGND 0.004984f
C9231 VDPWR.n2728 VGND 0.016028f
C9232 VDPWR.t625 VGND 0.005024f
C9233 VDPWR.t1218 VGND 0.010664f
C9234 VDPWR.n2730 VGND 0.027341f
C9235 VDPWR.t626 VGND 0.005024f
C9236 VDPWR.n2731 VGND 0.014893f
C9237 VDPWR.t722 VGND 0.005024f
C9238 VDPWR.t1277 VGND 0.010664f
C9239 VDPWR.n2733 VGND 0.027341f
C9240 VDPWR.t723 VGND 0.005024f
C9241 VDPWR.n2734 VGND 0.014893f
C9242 VDPWR.n2735 VGND 0.012599f
C9243 VDPWR.n2736 VGND 0.003844f
C9244 VDPWR.n2737 VGND 0.00224f
C9245 VDPWR.n2738 VGND 0.001428f
C9246 VDPWR.n2739 VGND 0.017613f
C9247 VDPWR.t588 VGND 0.004984f
C9248 VDPWR.n2740 VGND 0.030163f
C9249 VDPWR.t1231 VGND 0.028799f
C9250 VDPWR.n2741 VGND 0.019432f
C9251 VDPWR.n2742 VGND 0.00833f
C9252 VDPWR.t587 VGND 0.004984f
C9253 VDPWR.n2743 VGND 0.003892f
C9254 VDPWR.n2744 VGND 0.004088f
C9255 VDPWR.n2745 VGND 0.002272f
C9256 VDPWR.n2746 VGND 0.005f
C9257 VDPWR.n2747 VGND 9.28e-19
C9258 VDPWR.n2748 VGND 0.00176f
C9259 VDPWR.n2749 VGND 0.021585f
C9260 VDPWR.n2750 VGND 0.002048f
C9261 VDPWR.n2751 VGND 0.002368f
C9262 VDPWR.n2752 VGND 0.001973f
C9263 VDPWR.n2753 VGND 0.003083f
C9264 VDPWR.n2754 VGND 0.003404f
C9265 VDPWR.n2755 VGND 0.128862f
C9266 VDPWR.n2756 VGND 0.003404f
C9267 VDPWR.n2757 VGND 0.003083f
C9268 VDPWR.n2758 VGND 0.001477f
C9269 VDPWR.n2759 VGND 6.08e-19
C9270 VDPWR.n2760 VGND 0.013021f
C9271 VDPWR.n2761 VGND 0.021375f
C9272 VDPWR.t573 VGND 0.004984f
C9273 VDPWR.n2762 VGND 0.008777f
C9274 VDPWR.n2763 VGND 0.005754f
C9275 VDPWR.n2764 VGND 0.003488f
C9276 VDPWR.n2765 VGND 0.004416f
C9277 VDPWR.n2766 VGND 0.005888f
C9278 VDPWR.n2767 VGND 0.00245f
C9279 VDPWR.n2768 VGND 0.003286f
C9280 VDPWR.t268 VGND 0.004259f
C9281 VDPWR.n2769 VGND 0.00392f
C9282 VDPWR.t969 VGND 0.001036f
C9283 VDPWR.n2770 VGND 0.002948f
C9284 VDPWR.n2771 VGND 0.005781f
C9285 VDPWR.t1113 VGND 0.001867f
C9286 VDPWR.t1115 VGND 0.001867f
C9287 VDPWR.n2772 VGND 0.003889f
C9288 VDPWR.n2773 VGND 0.006022f
C9289 VDPWR.n2774 VGND 0.001365f
C9290 VDPWR.n2775 VGND 0.005888f
C9291 VDPWR.t867 VGND 0.001148f
C9292 VDPWR.t386 VGND 7.56e-19
C9293 VDPWR.n2776 VGND 0.001983f
C9294 VDPWR.n2777 VGND 0.004651f
C9295 VDPWR.n2778 VGND 0.005888f
C9296 VDPWR.n2779 VGND 0.003488f
C9297 VDPWR.n2780 VGND 0.001306f
C9298 VDPWR.t1127 VGND 0.001867f
C9299 VDPWR.t1117 VGND 0.001867f
C9300 VDPWR.n2781 VGND 0.003889f
C9301 VDPWR.n2782 VGND 0.007282f
C9302 VDPWR.t263 VGND 0.002867f
C9303 VDPWR.t361 VGND 0.003924f
C9304 VDPWR.n2783 VGND 0.010151f
C9305 VDPWR.n2784 VGND 0.007557f
C9306 VDPWR.n2785 VGND 0.001096f
C9307 VDPWR.n2786 VGND 0.005888f
C9308 VDPWR.n2787 VGND 0.004544f
C9309 VDPWR.n2788 VGND 0.001353f
C9310 VDPWR.n2789 VGND 0.001703f
C9311 VDPWR.n2790 VGND 0.005793f
C9312 VDPWR.n2791 VGND 0.006683f
C9313 VDPWR.t1101 VGND 0.001867f
C9314 VDPWR.t1111 VGND 0.001867f
C9315 VDPWR.n2792 VGND 0.003854f
C9316 VDPWR.t162 VGND 0.002741f
C9317 VDPWR.n2793 VGND 0.004148f
C9318 VDPWR.n2794 VGND 0.005921f
C9319 VDPWR.n2795 VGND 0.001563f
C9320 VDPWR.n2796 VGND 0.001259f
C9321 VDPWR.n2797 VGND 0.002048f
C9322 VDPWR.n2798 VGND 0.001579f
C9323 VDPWR.n2799 VGND 0.001973f
C9324 VDPWR.n2800 VGND 0.00224f
C9325 VDPWR.n2801 VGND 0.002752f
C9326 VDPWR.n2802 VGND 0.001973f
C9327 VDPWR.n2803 VGND 0.003083f
C9328 VDPWR.n2804 VGND 0.003404f
C9329 VDPWR.n2805 VGND 0.128862f
C9330 VDPWR.n2806 VGND 0.003404f
C9331 VDPWR.n2807 VGND 0.003083f
C9332 VDPWR.n2808 VGND 0.002949f
C9333 VDPWR.n2809 VGND 0.002528f
C9334 VDPWR.n2810 VGND 0.00224f
C9335 VDPWR.t624 VGND 0.051698f
C9336 VDPWR.t586 VGND 0.074717f
C9337 VDPWR.t571 VGND 0.046604f
C9338 VDPWR.t900 VGND 0.022453f
C9339 VDPWR.t954 VGND 0.028868f
C9340 VDPWR.t267 VGND 0.026604f
C9341 VDPWR.t1118 VGND 0.019623f
C9342 VDPWR.t1112 VGND 0.030189f
C9343 VDPWR.t968 VGND 0.016226f
C9344 VDPWR.t1114 VGND 0.016604f
C9345 VDPWR.t866 VGND 0.016226f
C9346 VDPWR.t1130 VGND 0.018113f
C9347 VDPWR.t1122 VGND 0.016604f
C9348 VDPWR.t385 VGND 0.012641f
C9349 VDPWR.t1126 VGND 0.019811f
C9350 VDPWR.t1116 VGND 0.019623f
C9351 VDPWR.t262 VGND 0.016226f
C9352 VDPWR.t1120 VGND 0.028868f
C9353 VDPWR.t1124 VGND 0.01849f
C9354 VDPWR.t360 VGND 0.016226f
C9355 VDPWR.t1128 VGND 0.016226f
C9356 VDPWR.t1042 VGND 0.016226f
C9357 VDPWR.t1102 VGND 0.019623f
C9358 VDPWR.t225 VGND 0.016226f
C9359 VDPWR.t1100 VGND 0.018868f
C9360 VDPWR.t161 VGND 0.016226f
C9361 VDPWR.t1110 VGND 0.012264f
C9362 VDPWR.t1104 VGND 0.014151f
C9363 VDPWR.t444 VGND 0.052075f
C9364 VDPWR.t462 VGND 0.098679f
C9365 VDPWR.t687 VGND 0.057736f
C9366 VDPWR.t1044 VGND 0.02566f
C9367 VDPWR.t872 VGND 0.039811f
C9368 VDPWR.t390 VGND 0.024906f
C9369 VDPWR.t153 VGND 0.039811f
C9370 VDPWR.t977 VGND 0.027547f
C9371 VDPWR.t804 VGND 0.033962f
C9372 VDPWR.t155 VGND 0.037358f
C9373 VDPWR.t1053 VGND 0.04434f
C9374 VDPWR.t920 VGND 0.033774f
C9375 VDPWR.t714 VGND 0.017924f
C9376 VDPWR.t156 VGND 0.024906f
C9377 VDPWR.t803 VGND 0.037358f
C9378 VDPWR.t812 VGND 0.061132f
C9379 VDPWR.t157 VGND 0.055472f
C9380 VDPWR.t810 VGND 0.023396f
C9381 VDPWR.n2811 VGND 0.038158f
C9382 VDPWR.t1141 VGND 0.029245f
C9383 VDPWR.t501 VGND 0.01849f
C9384 VDPWR.t22 VGND 0.018113f
C9385 VDPWR.t194 VGND 0.039057f
C9386 VDPWR.t14 VGND 0.036981f
C9387 VDPWR.t795 VGND 0.037358f
C9388 VDPWR.t377 VGND 0.013585f
C9389 VDPWR.t1143 VGND 0.015849f
C9390 VDPWR.t53 VGND 0.018113f
C9391 VDPWR.t308 VGND 0.039623f
C9392 VDPWR.t379 VGND 0.042641f
C9393 VDPWR.t362 VGND 0.021509f
C9394 VDPWR.t828 VGND 0.021321f
C9395 VDPWR.t1006 VGND 0.013019f
C9396 VDPWR.t986 VGND 0.020755f
C9397 VDPWR.t190 VGND 0.026792f
C9398 VDPWR.t364 VGND 0.022453f
C9399 VDPWR.t299 VGND 0.016038f
C9400 VDPWR.t231 VGND 0.017736f
C9401 VDPWR.t92 VGND 0.019434f
C9402 VDPWR.t983 VGND 0.022075f
C9403 VDPWR.t827 VGND 0.028868f
C9404 VDPWR.t1047 VGND 0.016038f
C9405 VDPWR.t1134 VGND 0.020755f
C9406 VDPWR.t1148 VGND 0.033962f
C9407 VDPWR.t366 VGND 0.019811f
C9408 VDPWR.t984 VGND 0.00566f
C9409 VDPWR.t1158 VGND 0.017547f
C9410 VDPWR.t773 VGND 0.025472f
C9411 VDPWR.t775 VGND 0.01717f
C9412 VDPWR.t331 VGND 0.016226f
C9413 VDPWR.t781 VGND 0.016604f
C9414 VDPWR.t16 VGND 0.00717f
C9415 VDPWR.t777 VGND 0.01717f
C9416 VDPWR.t1108 VGND 0.02434f
C9417 VDPWR.t1106 VGND 0.03f
C9418 VDPWR.n2812 VGND 0.019299f
C9419 VDPWR.n2813 VGND 0.011327f
C9420 VDPWR.n2814 VGND 0.00598f
C9421 VDPWR.t1109 VGND 0.001867f
C9422 VDPWR.t778 VGND 0.001867f
C9423 VDPWR.n2815 VGND 0.004076f
C9424 VDPWR.n2816 VGND 0.006757f
C9425 VDPWR.n2817 VGND 0.001703f
C9426 VDPWR.n2818 VGND 0.004416f
C9427 VDPWR.n2819 VGND 0.003744f
C9428 VDPWR.n2820 VGND 0.002016f
C9429 VDPWR.n2821 VGND 0.001213f
C9430 VDPWR.t17 VGND 0.001527f
C9431 VDPWR.t332 VGND 0.001527f
C9432 VDPWR.n2822 VGND 0.003394f
C9433 VDPWR.t782 VGND 0.001867f
C9434 VDPWR.t776 VGND 0.001867f
C9435 VDPWR.n2823 VGND 0.004071f
C9436 VDPWR.n2824 VGND 0.014462f
C9437 VDPWR.n2825 VGND 0.005344f
C9438 VDPWR.n2826 VGND 0.004416f
C9439 VDPWR.n2827 VGND 0.002016f
C9440 VDPWR.t774 VGND 0.006972f
C9441 VDPWR.n2828 VGND 0.008825f
C9442 VDPWR.t1159 VGND 0.001152f
C9443 VDPWR.t985 VGND 0.001152f
C9444 VDPWR.n2829 VGND 0.002399f
C9445 VDPWR.n2830 VGND 0.006436f
C9446 VDPWR.n2831 VGND 0.002048f
C9447 VDPWR.n2832 VGND 0.005312f
C9448 VDPWR.n2833 VGND 0.005568f
C9449 VDPWR.n2834 VGND 0.005721f
C9450 VDPWR.t1048 VGND 0.002195f
C9451 VDPWR.t93 VGND 0.002658f
C9452 VDPWR.n2835 VGND 0.006308f
C9453 VDPWR.n2836 VGND 0.003819f
C9454 VDPWR.n2837 VGND 0.001702f
C9455 VDPWR.n2838 VGND 0.002048f
C9456 VDPWR.n2839 VGND 0.002048f
C9457 VDPWR.n2840 VGND 0.002944f
C9458 VDPWR.n2841 VGND 0.001973f
C9459 VDPWR.n2842 VGND 0.003083f
C9460 VDPWR.n2843 VGND 0.003404f
C9461 VDPWR.n2844 VGND 0.128862f
C9462 VDPWR.n2845 VGND 0.003404f
C9463 VDPWR.n2846 VGND 0.003083f
C9464 VDPWR.n2847 VGND 0.001973f
C9465 VDPWR.n2848 VGND 0.002112f
C9466 VDPWR.n2849 VGND 0.002048f
C9467 VDPWR.n2850 VGND 0.002024f
C9468 VDPWR.t232 VGND 0.002785f
C9469 VDPWR.t191 VGND 0.00135f
C9470 VDPWR.n2851 VGND 0.00567f
C9471 VDPWR.t365 VGND 0.002864f
C9472 VDPWR.n2852 VGND 0.008079f
C9473 VDPWR.n2853 VGND 0.004349f
C9474 VDPWR.n2854 VGND 0.001598f
C9475 VDPWR.n2855 VGND 0.003904f
C9476 VDPWR.n2856 VGND 0.004416f
C9477 VDPWR.n2857 VGND 0.002016f
C9478 VDPWR.n2858 VGND 0.00187f
C9479 VDPWR.t363 VGND 0.001372f
C9480 VDPWR.t1007 VGND 0.002267f
C9481 VDPWR.n2859 VGND 0.006283f
C9482 VDPWR.n2860 VGND 0.007702f
C9483 VDPWR.n2861 VGND 7.82e-19
C9484 VDPWR.n2862 VGND 0.005888f
C9485 VDPWR.n2863 VGND 0.005888f
C9486 VDPWR.n2864 VGND 0.005888f
C9487 VDPWR.t309 VGND 0.007351f
C9488 VDPWR.n2865 VGND 0.006963f
C9489 VDPWR.n2866 VGND 0.005167f
C9490 VDPWR.n2867 VGND 0.001133f
C9491 VDPWR.n2868 VGND 0.001179f
C9492 VDPWR.n2869 VGND 0.004416f
C9493 VDPWR.n2870 VGND 0.002944f
C9494 VDPWR.n2871 VGND 0.001089f
C9495 VDPWR.t15 VGND 0.004259f
C9496 VDPWR.t195 VGND 0.001036f
C9497 VDPWR.n2872 VGND 0.002948f
C9498 VDPWR.n2873 VGND 0.00392f
C9499 VDPWR.n2874 VGND 0.002688f
C9500 VDPWR.n2875 VGND 0.003005f
C9501 VDPWR.n2876 VGND 0.00224f
C9502 VDPWR.n2877 VGND 0.00224f
C9503 VDPWR.n2878 VGND 0.001973f
C9504 VDPWR.n2879 VGND 0.003404f
C9505 VDPWR.n2880 VGND 0.003083f
C9506 VDPWR.n2881 VGND 0.002757f
C9507 VDPWR.n2882 VGND 0.002176f
C9508 VDPWR.n2883 VGND 0.003702f
C9509 VDPWR.t502 VGND 0.004984f
C9510 VDPWR.n2884 VGND 0.004913f
C9511 VDPWR.n2885 VGND 0.018812f
C9512 VDPWR.n2886 VGND 0.011593f
C9513 VDPWR.t23 VGND 0.001148f
C9514 VDPWR.t1142 VGND 7.56e-19
C9515 VDPWR.n2887 VGND 0.00196f
C9516 VDPWR.n2888 VGND 0.005471f
C9517 VDPWR.t503 VGND 0.004984f
C9518 VDPWR.n2889 VGND 0.008609f
C9519 VDPWR.n2890 VGND 0.011129f
C9520 VDPWR.n2891 VGND 0.007897f
C9521 VDPWR.n2892 VGND 0.002048f
C9522 VDPWR.n2893 VGND 0.002944f
C9523 VDPWR.n2894 VGND 0.001973f
C9524 VDPWR.n2895 VGND 0.001579f
C9525 VDPWR.n2896 VGND 0.00352f
C9526 VDPWR.n2897 VGND 0.003404f
C9527 VDPWR.n2898 VGND 0.003083f
C9528 VDPWR.n2899 VGND 5.48e-19
C9529 VDPWR.n2900 VGND 0.00224f
C9530 VDPWR.n2901 VGND 0.002272f
C9531 VDPWR.n2902 VGND 0.001642f
C9532 VDPWR.t715 VGND 0.005483f
C9533 VDPWR.n2903 VGND 8.72e-19
C9534 VDPWR.n2904 VGND 0.003023f
C9535 VDPWR.n2905 VGND 0.004416f
C9536 VDPWR.n2906 VGND 0.005888f
C9537 VDPWR.n2907 VGND 0.007099f
C9538 VDPWR.n2908 VGND 0.004558f
C9539 VDPWR.n2909 VGND 0.008069f
C9540 VDPWR.n2910 VGND 0.00484f
C9541 VDPWR.n2911 VGND 0.005888f
C9542 VDPWR.n2912 VGND 0.005888f
C9543 VDPWR.n2913 VGND 0.005445f
C9544 VDPWR.n2914 VGND 0.007422f
C9545 VDPWR.t921 VGND 0.00135f
C9546 VDPWR.t1054 VGND 0.002785f
C9547 VDPWR.n2915 VGND 0.00567f
C9548 VDPWR.n2916 VGND 0.007073f
C9549 VDPWR.n2917 VGND 0.005445f
C9550 VDPWR.n2918 VGND 0.005888f
C9551 VDPWR.n2919 VGND 0.005888f
C9552 VDPWR.n2920 VGND 0.004672f
C9553 VDPWR.n2921 VGND 0.007422f
C9554 VDPWR.n2922 VGND 0.007422f
C9555 VDPWR.n2923 VGND 0.00718f
C9556 VDPWR.n2924 VGND 0.002048f
C9557 VDPWR.n2925 VGND 0.001579f
C9558 VDPWR.n2926 VGND 0.001973f
C9559 VDPWR.n2927 VGND 0.002112f
C9560 VDPWR.n2928 VGND 0.00288f
C9561 VDPWR.n2929 VGND 0.001973f
C9562 VDPWR.n2930 VGND 0.003083f
C9563 VDPWR.n2931 VGND 0.003404f
C9564 VDPWR.n2932 VGND 0.128862f
C9565 VDPWR.n2933 VGND 0.003404f
C9566 VDPWR.n2934 VGND 0.003083f
C9567 VDPWR.n2935 VGND 0.002405f
C9568 VDPWR.n2936 VGND 0.001504f
C9569 VDPWR.n2937 VGND 9.22e-19
C9570 VDPWR.n2938 VGND 0.005576f
C9571 VDPWR.n2939 VGND 0.002784f
C9572 VDPWR.t688 VGND 0.005483f
C9573 VDPWR.n2940 VGND 0.00426f
C9574 VDPWR.n2941 VGND 0.00355f
C9575 VDPWR.n2942 VGND 0.005888f
C9576 VDPWR.n2943 VGND 0.003488f
C9577 VDPWR.n2944 VGND 0.007341f
C9578 VDPWR.t873 VGND 0.007047f
C9579 VDPWR.t1187 VGND 0.072626f
C9580 VDPWR.n2945 VGND 0.033681f
C9581 VDPWR.n2946 VGND 0.011895f
C9582 VDPWR.n2947 VGND 0.003953f
C9583 VDPWR.n2948 VGND 0.004416f
C9584 VDPWR.n2949 VGND 0.005888f
C9585 VDPWR.n2950 VGND 0.003456f
C9586 VDPWR.n2951 VGND 0.007073f
C9587 VDPWR.t463 VGND 0.004984f
C9588 VDPWR.n2952 VGND 0.011445f
C9589 VDPWR.n2953 VGND 0.008952f
C9590 VDPWR.n2954 VGND 0.004416f
C9591 VDPWR.n2955 VGND 0.005888f
C9592 VDPWR.n2956 VGND 0.005888f
C9593 VDPWR.n2957 VGND 0.020793f
C9594 VDPWR.n2958 VGND 0.020793f
C9595 VDPWR.t464 VGND 0.004984f
C9596 VDPWR.t689 VGND 0.005483f
C9597 VDPWR.n2959 VGND 0.011995f
C9598 VDPWR.n2960 VGND 0.020115f
C9599 VDPWR.n2961 VGND 0.005696f
C9600 VDPWR.n2962 VGND 7.36e-19
C9601 VDPWR.n2963 VGND 0.002949f
C9602 VDPWR.n2964 VGND 0.003083f
C9603 VDPWR.n2965 VGND 0.001579f
C9604 VDPWR.n2966 VGND 0.001973f
C9605 VDPWR.n2967 VGND 0.001472f
C9606 VDPWR.n2968 VGND 0.002944f
C9607 VDPWR.n2969 VGND 0.002048f
C9608 VDPWR.t445 VGND 0.005024f
C9609 VDPWR.t1253 VGND 0.010664f
C9610 VDPWR.n2971 VGND 0.027341f
C9611 VDPWR.t446 VGND 0.005024f
C9612 VDPWR.n2972 VGND 0.014893f
C9613 VDPWR.n2973 VGND 0.012551f
C9614 VDPWR.n2974 VGND 0.001376f
C9615 VDPWR.n2975 VGND 0.002885f
C9616 VDPWR.n2976 VGND 0.002112f
C9617 VDPWR.n2977 VGND 0.001973f
C9618 VDPWR.n2978 VGND 0.001579f
C9619 VDPWR.n2979 VGND 0.00352f
C9620 VDPWR.n2980 VGND 0.003404f
C9621 VDPWR.n2981 VGND 0.128862f
C9622 VDPWR.n2982 VGND 0.128008f
C9623 VDPWR.n2983 VGND 0.001579f
C9624 VDPWR.n2984 VGND 0.001579f
C9625 VDPWR.n2985 VGND 0.001973f
C9626 VDPWR.n2986 VGND 0.002112f
C9627 VDPWR.t877 VGND 0.007047f
C9628 VDPWR.t555 VGND 0.004984f
C9629 VDPWR.n2987 VGND 0.018696f
C9630 VDPWR.n2988 VGND 0.005471f
C9631 VDPWR.t427 VGND 0.005024f
C9632 VDPWR.t1285 VGND 0.010664f
C9633 VDPWR.n2990 VGND 0.027341f
C9634 VDPWR.t428 VGND 0.005024f
C9635 VDPWR.n2991 VGND 0.014893f
C9636 VDPWR.n2992 VGND 0.001472f
C9637 VDPWR.n2993 VGND 0.002048f
C9638 VDPWR.n2994 VGND 0.001973f
C9639 VDPWR.n2995 VGND 0.002944f
C9640 VDPWR.n2996 VGND 0.002048f
C9641 VDPWR.t548 VGND 0.005024f
C9642 VDPWR.t1256 VGND 0.010664f
C9643 VDPWR.n2998 VGND 0.027341f
C9644 VDPWR.t549 VGND 0.005024f
C9645 VDPWR.n2999 VGND 0.014893f
C9646 VDPWR.n3000 VGND 0.012553f
C9647 VDPWR.n3001 VGND 0.001376f
C9648 VDPWR.n3002 VGND 0.002885f
C9649 VDPWR.n3003 VGND 0.003083f
C9650 VDPWR.n3004 VGND 0.003404f
C9651 VDPWR.n3005 VGND 0.00352f
C9652 VDPWR.n3006 VGND 0.00352f
C9653 VDPWR.n3007 VGND 0.003404f
C9654 VDPWR.n3008 VGND 0.003083f
C9655 VDPWR.n3009 VGND 0.002949f
C9656 VDPWR.n3010 VGND 0.00512f
C9657 VDPWR.n3011 VGND 0.002048f
C9658 VDPWR.n3012 VGND 0.015457f
C9659 VDPWR.n3013 VGND 0.015289f
C9660 VDPWR.n3014 VGND 0.01206f
C9661 VDPWR.n3015 VGND 0.032215f
C9662 VDPWR.n3016 VGND 0.005888f
C9663 VDPWR.n3017 VGND 0.004416f
C9664 VDPWR.n3018 VGND 0.005376f
C9665 VDPWR.n3019 VGND 0.005676f
C9666 VDPWR.n3020 VGND 0.003488f
C9667 VDPWR.n3021 VGND 0.005888f
C9668 VDPWR.n3022 VGND 0.005888f
C9669 VDPWR.n3023 VGND 0.001349f
C9670 VDPWR.n3024 VGND 0.006073f
C9671 VDPWR.n3025 VGND 0.001383f
C9672 VDPWR.n3026 VGND 0.004406f
C9673 VDPWR.n3027 VGND 0.00153f
C9674 VDPWR.n3028 VGND 0.0048f
C9675 VDPWR.n3029 VGND 0.002949f
C9676 VDPWR.n3030 VGND 0.003083f
C9677 VDPWR.n3031 VGND 0.003404f
C9678 VDPWR.n3032 VGND 0.00352f
C9679 VDPWR.n3033 VGND 0.003404f
C9680 VDPWR.n3034 VGND 0.00352f
C9681 VDPWR.n3035 VGND 0.001579f
C9682 VDPWR.n3036 VGND 0.001973f
C9683 VDPWR.n3037 VGND 0.00288f
C9684 VDPWR.n3038 VGND 0.002048f
C9685 VDPWR.n3039 VGND 9.41e-19
C9686 VDPWR.n3040 VGND 0.007134f
C9687 VDPWR.n3041 VGND 0.00187f
C9688 VDPWR.n3042 VGND 0.005888f
C9689 VDPWR.n3043 VGND 0.005888f
C9690 VDPWR.n3044 VGND 5.44e-19
C9691 VDPWR.n3045 VGND 0.007134f
C9692 VDPWR.n3046 VGND 0.00187f
C9693 VDPWR.n3047 VGND 0.004416f
C9694 VDPWR.n3048 VGND 0.005888f
C9695 VDPWR.n3049 VGND 0.004416f
C9696 VDPWR.n3050 VGND 0.001247f
C9697 VDPWR.n3051 VGND 0.00364f
C9698 VDPWR.n3052 VGND 0.013305f
C9699 VDPWR.n3053 VGND 0.012101f
C9700 VDPWR.n3054 VGND 0.002016f
C9701 VDPWR.n3055 VGND 5.48e-19
C9702 VDPWR.n3056 VGND 0.003083f
C9703 VDPWR.n3057 VGND 0.001973f
C9704 VDPWR.n3058 VGND 0.002944f
C9705 VDPWR.n3059 VGND 0.002048f
C9706 VDPWR.n3060 VGND 0.012181f
C9707 VDPWR.n3061 VGND 0.011593f
C9708 VDPWR.n3062 VGND 0.002048f
C9709 VDPWR.n3063 VGND 0.00224f
C9710 VDPWR.n3064 VGND 0.001973f
C9711 VDPWR.n3065 VGND 0.003083f
C9712 VDPWR.n3066 VGND 0.003404f
C9713 VDPWR.n3067 VGND 0.128008f
C9714 VDPWR.n3068 VGND 0.116061f
C9715 VDPWR.n3069 VGND 0.281618f
C9716 VDPWR.n3070 VGND 0.167264f
C9717 VDPWR.n3071 VGND 0.281618f
C9718 VDPWR.n3072 VGND 0.116061f
C9719 VDPWR.n3073 VGND 0.107527f
C9720 VDPWR.n3074 VGND 0.078829f
C9721 VDPWR.n3075 VGND 0.003054f
C9722 VDPWR.n3076 VGND 0.002949f
C9723 VDPWR.n3077 VGND 0.004128f
C9724 VDPWR.n3078 VGND 0.002016f
C9725 VDPWR.n3079 VGND 0.001941f
C9726 VDPWR.n3080 VGND 0.005906f
C9727 VDPWR.n3081 VGND 0.003488f
C9728 VDPWR.n3082 VGND 0.004416f
C9729 VDPWR.n3083 VGND 0.011677f
C9730 VDPWR.n3084 VGND 0.015457f
C9731 VDPWR.n3085 VGND 0.011257f
C9732 VDPWR.n3086 VGND 0.005888f
C9733 VDPWR.n3087 VGND 0.005888f
C9734 VDPWR.n3088 VGND 0.005344f
C9735 VDPWR.n3089 VGND 0.011425f
C9736 VDPWR.n3090 VGND 0.046459f
C9737 VDPWR.n3091 VGND 0.009153f
C9738 VDPWR.n3092 VGND 0.010501f
C9739 VDPWR.n3093 VGND 0.002016f
C9740 VDPWR.n3094 VGND 0.002272f
C9741 VDPWR.n3095 VGND 0.005471f
C9742 VDPWR.n3096 VGND 0.01243f
C9743 VDPWR.n3097 VGND 0.001156f
C9744 VDPWR.n3098 VGND 0.002048f
C9745 VDPWR.n3099 VGND 0.002944f
C9746 VDPWR.n3100 VGND 0.001973f
C9747 VDPWR.n3101 VGND 0.001579f
C9748 VDPWR.n3102 VGND 0.078408f
C9749 VDPWR.n3103 VGND 0.272304f
C9750 VDPWR.n3104 VGND 0.13926f
C9751 VDPWR.n3105 VGND 0.13926f
C9752 VDPWR.n3106 VGND 0.209943f
C9753 VDPWR.n3107 VGND 0.292729f
C9754 VDPWR.n3108 VGND 0.060111f
C9755 VDPWR.n3109 VGND 0.281618f
C9756 VDPWR.n3110 VGND 0.167264f
C9757 VDPWR.n3111 VGND 0.060111f
C9758 VDPWR.n3112 VGND 0.096641f
C9759 VDPWR.n3113 VGND 0.107527f
C9760 VDPWR.n3114 VGND 0.02543f
C9761 VDPWR.n3115 VGND 0.067982f
C9762 VDPWR.n3116 VGND 1.57447f
C9763 VDPWR.n3117 VGND 3.32341f
C9764 VDPWR.n3118 VGND 0.390779f
C9765 VDPWR.n3119 VGND 0.035269f
C9766 VDPWR.n3120 VGND 0.114487f
C9767 VDPWR.n3121 VGND 0.055474f
C9768 VDPWR.n3122 VGND 0.055474f
C9769 VDPWR.n3123 VGND 0.055293f
C9770 VDPWR.n3124 VGND 0.076656f
C9771 VDPWR.n3125 VGND 0.247132f
C9772 VDPWR.t1094 VGND 0.356671f
C9773 VDPWR.n3126 VGND 0.344366f
C9774 VDPWR.t1095 VGND 0.356671f
C9775 VDPWR.n3127 VGND 0.247132f
C9776 VDPWR.n3128 VGND 2.38e-19
C9777 VDPWR.n3129 VGND 0.006274f
C9778 VDPWR.n3130 VGND 0.060635f
C9779 VDPWR.n3131 VGND 0.018181f
C9780 VDPWR.n3132 VGND 0.030678f
C9781 VDPWR.n3133 VGND 0.156059f
C9782 VDPWR.n3134 VGND 0.169072f
C9783 VDPWR.n3135 VGND 0.035235f
C9784 VDPWR.n3136 VGND 0.114487f
C9785 VDPWR.n3137 VGND 0.00445f
C9786 VDPWR.n3138 VGND 0.055474f
C9787 VDPWR.n3139 VGND 0.055474f
C9788 VDPWR.n3140 VGND 0.055293f
C9789 VDPWR.n3141 VGND 0.076656f
C9790 VDPWR.n3142 VGND 0.247132f
C9791 VDPWR.t49 VGND 0.356671f
C9792 VDPWR.n3143 VGND 0.344366f
C9793 VDPWR.t50 VGND 0.356671f
C9794 VDPWR.n3144 VGND 0.247132f
C9795 VDPWR.n3145 VGND 0.002025f
C9796 VDPWR.n3146 VGND 0.060694f
C9797 VDPWR.n3147 VGND 0.018181f
C9798 VDPWR.n3148 VGND 0.029169f
C9799 VDPWR.n3149 VGND 0.160902f
C9800 VDPWR.n3150 VGND 0.183546f
C9801 VDPWR.n3151 VGND 0.035121f
C9802 VDPWR.n3152 VGND 0.114487f
C9803 VDPWR.n3153 VGND 0.004458f
C9804 VDPWR.n3154 VGND 0.055474f
C9805 VDPWR.n3155 VGND 0.055474f
C9806 VDPWR.n3156 VGND 0.055293f
C9807 VDPWR.n3157 VGND 0.076656f
C9808 VDPWR.n3158 VGND 0.247132f
C9809 VDPWR.t239 VGND 0.356671f
C9810 VDPWR.n3159 VGND 0.344366f
C9811 VDPWR.t1093 VGND 0.356671f
C9812 VDPWR.n3160 VGND 0.247132f
C9813 VDPWR.n3161 VGND 0.002138f
C9814 VDPWR.n3162 VGND 0.060694f
C9815 VDPWR.n3163 VGND 0.018181f
C9816 VDPWR.n3164 VGND 0.029169f
C9817 VDPWR.n3165 VGND 0.162708f
C9818 VDPWR.n3166 VGND 0.166655f
C9819 VDPWR.n3167 VGND 0.006257f
C9820 VDPWR.n3168 VGND 0.060659f
C9821 VDPWR.n3169 VGND 0.018181f
C9822 VDPWR.n3170 VGND 0.029432f
C9823 VDPWR.n3171 VGND 0.060236f
C9824 VDPWR.n3172 VGND 0.674934f
C9825 VDPWR.t945 VGND 0.0028f
C9826 VDPWR.t1212 VGND 0.00165f
C9827 VDPWR.t948 VGND 0.0028f
C9828 VDPWR.t1206 VGND 0.00165f
C9829 VDPWR.n3173 VGND 0.004698f
C9830 VDPWR.n3174 VGND 0.006946f
C9831 VDPWR.n3175 VGND 0.006899f
C9832 VDPWR.n3176 VGND 0.030149f
C9833 VDPWR.n3177 VGND 0.092595f
C9834 VDPWR.n3178 VGND 0.037419f
C9835 ringtest_0.x4.net2.t7 VGND 0.015381f
C9836 ringtest_0.x4.net2.t8 VGND 0.026101f
C9837 ringtest_0.x4.net2.n0 VGND 0.037026f
C9838 ringtest_0.x4.net2.t4 VGND 0.015381f
C9839 ringtest_0.x4.net2.t3 VGND 0.026101f
C9840 ringtest_0.x4.net2.n1 VGND 0.033335f
C9841 ringtest_0.x4.net2.n2 VGND 0.017289f
C9842 ringtest_0.x4.net2.n3 VGND 0.0837f
C9843 ringtest_0.x4.net2.t5 VGND 0.026101f
C9844 ringtest_0.x4.net2.t2 VGND 0.016278f
C9845 ringtest_0.x4.net2.n4 VGND 0.052479f
C9846 ringtest_0.x4.net2.n5 VGND 0.259642f
C9847 ringtest_0.x4.net2.t9 VGND 0.013842f
C9848 ringtest_0.x4.net2.t11 VGND 0.011454f
C9849 ringtest_0.x4.net2.n6 VGND 0.060494f
C9850 ringtest_0.x4.net2.n7 VGND 0.03533f
C9851 ringtest_0.x4.net2.n8 VGND 0.650991f
C9852 ringtest_0.x4.net2.t6 VGND 0.017756f
C9853 ringtest_0.x4.net2.t10 VGND 0.028277f
C9854 ringtest_0.x4.net2.n9 VGND 0.038818f
C9855 ringtest_0.x4.net2.n10 VGND 0.03575f
C9856 ringtest_0.x4.net2.n11 VGND 0.11929f
C9857 ringtest_0.x4.net2.n12 VGND 0.278364f
C9858 ringtest_0.x4.net2.n13 VGND 0.037886f
C9859 ringtest_0.x4.net2.t1 VGND 0.08709f
C9860 ringtest_0.x4.net2.n14 VGND 0.10636f
C9861 ringtest_0.x4.net2.t0 VGND 0.032833f
.ends

