* NGSPICE file created from ringtest_parax.ext - technology: sky130A

.subckt ringtest_parax enable_ring select0 mux_out enable_counter select1 VSS VDD
X0 a_17405_n2032# x3.x1.nSEL1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X1 VDD VSS.t967 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X2 VSS.t5 x4.clknet_1_0__leaf_clk.t32 a_23339_n9259# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 a_21119_n968.t0 ring_out.t10 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=2.026362 ps=18.53074 w=9 l=0.15
**devattr s=104400,3716 d=104400,3716
X4 a_28197_n9259# a_28031_n9259# VSS.t177 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X5 x3.x2.GP4.t3 x3.x2.GN4 VSS.t241 VSS.t240 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X6 a_29021_n8337# a_28031_n8709# a_28895_n8715# VSS.t901 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X7 VSS.t672 VDD VSS.t671 VSS.t670 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X8 VDD x4.clknet_1_0__leaf_clk.t33 a_23339_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X9 VDD VSS.t968 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X10 VDD VSS.t969 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X11 a_26295_n7249# a_26159_n7409# a_25875_n7395# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.078615 pd=0.771795 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4380,215
X12 VSS.t669 VDD VSS.t668 VSS.t373 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X13 a_28197_n9259# a_28031_n9259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X14 VSS.t667 VDD VSS.t666 VSS.t639 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X15 x4._13_ x4._11_.t4 VSS.t336 VSS.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X16 a_24053_n8337# a_23063_n8709# a_23927_n8715# VSS.t160 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X17 VDD x1.sky130_fd_sc_hd__inv_2_12.A x1.sky130_fd_sc_hd__inv_2_13.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X18 VDD x4.net4 a_23421_n7921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X19 VSS.t949 a_26798_n8741# a_26756_n8337# VSS.t948 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X20 drv_out.t19 a_21119_n968.t2 VSS.t136 VSS.t135 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X21 VDD VSS.t970 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X22 drv_out.t1 x3.x2.GN2 mux_out.t11 VSS.t749 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X23 a_23633_n4541# a_23295_n4755# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4452,274 d=3528,168
X24 a_26159_n7409# x4.clknet_1_1__leaf_clk.t32 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X25 VSS.t116 a_25709_n7109# x4.clknet_0_clk.t31 VSS.t115 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X26 VDD VSS.t971 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X27 VDD a_23851_n9829# x4._03_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=7430,283
X28 VSS.t665 VDD VSS.t664 VSS.t663 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X29 a_24287_n8893# a_23505_n9259# a_24203_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X30 VSS.t662 VDD VSS.t661 VSS.t660 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X31 VDD VSS.t972 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X32 VSS.t659 VDD VSS.t658 VSS.t657 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X33 VDD a_25709_n7109# x4.clknet_0_clk.t15 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X34 a_28197_n8709# a_28031_n8709# VSS.t900 VSS.t899 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X35 x4.counter[9] a_29319_n10347# VSS.t962 VSS.t961 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X36 VDD x1.sky130_fd_sc_hd__inv_2_13.A x1.sky130_fd_sc_hd__inv_2_14.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X37 a_27755_n7261# x4._11_.t5 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X38 VSS.t725 a_27423_n8893# a_27591_n8991# VSS.t724 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X39 VSS.t173 a_24095_n8741# a_24053_n8337# VSS.t172 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X40 VSS.t656 VDD VSS.t655 VSS.t654 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X41 a_28638_n9147# a_28470_n8893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.168863 ps=1.544228 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X42 VDD VSS.t973 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X43 x4._17_ a_27755_n7261# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X44 VDD a_29063_n8991# a_28979_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X45 x4.net4 a_24095_n8741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X46 VSS.t193 x1.sky130_fd_sc_hd__inv_2_16.A x1.sky130_fd_sc_hd__inv_2_17.A VSS.t26 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X47 VDD VSS.t974 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X48 VDD x4.net2.t2 a_23615_n5995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X49 VDD a_24203_n8893# a_24371_n8991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X50 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t15 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X51 a_18409_n2290# select1.t0 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X52 x4.net11 a_29063_n8991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X53 a_23697_n5995# x4.net2.t3 a_23615_n5995# VSS.t916 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X54 VSS.t653 VDD VSS.t652 VSS.t651 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X55 x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_8.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X56 x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_8.Y VSS.t920 VSS.t750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X57 x4.net6.t1 a_24647_n7903# VSS.t154 VSS.t153 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X58 VSS.t918 x4.net2.t4 a_23255_n4363# VSS.t917 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X59 x4._06_ a_25834_n7921# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=7430,283 d=10400,504
X60 a_22837_n10182# x4.net2.t5 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X61 VSS.t650 VDD VSS.t649 VSS.t648 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X62 VDD a_28895_n8715# a_29063_n8741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X63 VSS.t647 VDD VSS.t646 VSS.t645 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X64 a_23295_n5219# a_23391_n5219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X65 a_25875_n7395# a_26159_n7409# a_26094_n7261# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2736,148
X66 VDD VSS.t975 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X67 VSS.t114 a_25709_n7109# x4.clknet_0_clk.t30 VSS.t113 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X68 VSS.t941 select0.t0 a_18585_n1958# VSS.t940 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X69 VDD a_18033_n1958# a_17857_n2290# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X70 VDD VSS.t976 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X71 drv_out.t18 a_21119_n968.t3 VSS.t138 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X72 VDD VSS.t977 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X73 x4.clknet_0_clk.t14 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X74 x4.clknet_0_clk.t13 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X75 VSS.t73 a_26159_n7409# a_26166_n7505# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X76 a_28999_n7408# x4._25_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X77 VSS.t768 select1.t1 x3.x1.nSEL1 VSS.t767 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X78 VSS.t209 a_23941_n3056# x4.net1 VSS.t208 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X79 VSS.t343 a_24371_n8991# a_24329_n9259# VSS.t342 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X80 a_26094_n7261# a_25779_n7395# VSS.t805 VSS.t804 sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X81 a_28725_n10182# x4.net9 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X82 x4._01_ x4._12_ VSS.t211 VSS.t210 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X83 VSS.t58 a_26147_n9107# x4._20_ VSS.t57 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=5266,228
X84 VDD a_25709_n7109# x4.clknet_0_clk.t12 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X85 VSS.t706 a_23225_n7109# x4.clknet_1_0__leaf_clk.t31 VSS.t705 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X86 VDD VSS.t978 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X87 a_28470_n8893# a_28197_n9259# a_28385_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X88 a_27423_n8893# a_26559_n9259# a_27166_n9147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X89 VSS.t644 VDD VSS.t643 VSS.t642 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X90 VDD x4.clknet_0_clk.t32 a_23225_n7109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X91 a_27093_n8893# a_26559_n9259# a_26998_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X92 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t15 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X93 a_23769_n5995# x4.net3.t2 a_23697_n5995# VSS.t878 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X94 a_24605_n8171# a_23615_n8171# a_24479_n7805# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X95 VDD a_26147_n9107# x4._20_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5689,267
X96 VSS.t641 VDD VSS.t640 VSS.t639 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X97 a_24525_n5745# x4._12_ x4._01_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X98 x4.net8 a_27223_n8741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X99 counter7.t3 x3.x2.GN4 mux_out.t2 VSS.t239 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X100 VSS.t638 VDD VSS.t637 VSS.t636 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X101 VSS.t187 a_26366_n7350# a_26295_n7249# VSS.t186 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.126592 ps=1.2736 w=0.64 l=0.15
**devattr s=3956,199 d=4838,217
X102 x4.clknet_1_1__leaf_clk.t14 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X103 VDD a_27166_n9147# a_27093_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X104 a_27139_n8715# a_26357_n8709# a_27055_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X105 VDD VSS.t979 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X106 a_26885_n10182# x4.net7 VSS.t818 VSS.t817 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X107 VSS.t635 VDD VSS.t634 VSS.t633 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X108 VDD VSS.t980 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X109 x4.clknet_0_clk.t29 a_25709_n7109# VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X110 x4.clknet_0_clk.t28 a_25709_n7109# VSS.t110 VSS.t109 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X111 VSS.t295 a_24479_n7805# a_24647_n7903# VSS.t294 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X112 a_26309_n9259# x4.net8 VSS.t859 VSS.t858 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0 ps=0 w=0.42 l=0.15
**devattr s=5266,228 d=1764,126
X113 VSS.t150 x4._18_ a_25449_n7261# VSS.t149 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X114 VSS.t122 a_18409_n2290# x3.x2.GN3 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X115 x4._25_ a_28579_n7627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X116 x4.net4 a_24095_n8741# VSS.t171 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X117 x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_2.A VSS.t922 VSS.t196 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X118 a_26913_n9259# x4._07_ VSS.t801 VSS.t800 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X119 VDD VSS.t981 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X120 a_23391_n5219# a_23675_n5233# a_23610_n5085# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2736,148
X121 VSS.t108 a_25709_n7109# x4.clknet_0_clk.t27 VSS.t107 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X122 VDD VSS.t982 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.97
**devattr d=9048,452
X123 x4.clknet_0_clk.t11 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X124 a_29645_n10182# x4.net10 VSS.t300 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X125 VDD x4._20_ a_25639_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X126 x1.sky130_fd_sc_hd__inv_2_14.A x1.sky130_fd_sc_hd__inv_2_13.A VSS.t261 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X127 VSS.t909 x4.clknet_0_clk.t33 a_23225_n7109# VSS.t908 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X128 a_25779_n7395# a_25875_n7395# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X129 a_23904_n9259# a_23505_n9259# a_23778_n8893# VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X130 a_25823_n8395# x4._11_.t6 a_25729_n8395# VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
**devattr s=4160,194 d=4290,196
X131 VSS.t293 a_27194_n8171# x4.clknet_1_1__leaf_clk.t31 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X132 x3.x1.nSEL1 select1.t2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X133 a_26457_n7849# x4._21_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X134 x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_3.A VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X135 VDD x4._11_.t7 a_24525_n5745# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X136 VDD VSS.t983 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X137 x4._06_ a_25834_n7921# VSS.t755 VSS.t754 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X138 a_28895_n8715# a_28197_n8709# a_28638_n8741# VSS.t894 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X139 VDD x1.sky130_fd_sc_hd__inv_2_17.A x1.sky130_fd_sc_hd__inv_2_17.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X140 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t14 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X141 a_29133_n9803# a_29103_n9829# x4._09_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.3 ps=2.6 w=1 l=0.15
**devattr s=12000,520 d=10400,504
X142 x4.clknet_1_1__leaf_clk.t30 a_27194_n8171# VSS.t291 VSS.t290 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X143 VDD x4.clknet_0_clk.t34 a_23225_n7109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X144 VSS.t632 VDD VSS.t631 VSS.t630 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X145 VSS.t629 VDD VSS.t628 VSS.t627 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X146 VSS.t799 a_28638_n9147# a_28596_n9259# VSS.t798 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X147 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t13 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X148 VDD VSS.t984 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X149 VDD x1.sky130_fd_sc_hd__inv_2_14.A x1.sky130_fd_sc_hd__inv_2_15.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X150 a_25875_n7395# a_26166_n7505# a_26117_n7627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=2268,138
X151 VSS.t626 VDD VSS.t625 VSS.t406 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X152 a_27805_n10182# x4.net8 VSS.t857 VSS.t856 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X153 x4.clknet_1_1__leaf_clk.t12 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X154 VSS.t624 VDD VSS.t623 VSS.t564 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X155 VDD VSS.t985 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X156 VSS.t347 a_28999_n7408# x4._08_ VSS.t346 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X157 VSS.t674 a_17857_n2290# x3.x2.GN2 VSS.t673 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X158 VDD VSS.t986 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X159 VSS.t308 x4._10_ a_24075_n5995# VSS.t307 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=2730,149
X160 a_26159_n7409# x4.clknet_1_1__leaf_clk.t33 VSS.t874 VSS.t873 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X161 a_27423_n8893# a_26725_n9259# a_27166_n9147# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X162 x4.clknet_0_clk.t26 a_25709_n7109# VSS.t106 VSS.t105 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
X163 a_26798_n8741# a_26630_n8715# VSS.t249 VSS.t248 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X164 VDD x3.x2.GN2 x3.x2.GP2.t1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X165 a_25709_n7109# drv_out.t20 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X166 VDD a_23941_n3056# x4.net1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X167 VDD x4._10_ a_24075_n5995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6500,265
X168 VSS.t622 VDD VSS.t621 VSS.t550 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X169 a_23502_n8715# a_23063_n8709# a_23417_n8715# VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X170 VDD x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_5.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X171 VSS.t785 a_28638_n8741# a_28596_n8337# VSS.t784 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X172 VSS.t704 a_23225_n7109# x4.clknet_1_0__leaf_clk.t30 VSS.t703 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X173 VSS.t911 x4.clknet_0_clk.t35 a_23225_n7109# VSS.t910 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X174 VSS.t289 a_27194_n8171# x4.clknet_1_1__leaf_clk.t29 VSS.t288 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X175 VSS.t789 x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_6.A VSS.t788 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X176 VSS.t753 x1.sky130_fd_sc_hd__inv_2_17.Y x1.sky130_fd_sc_hd__inv_2_8.Y VSS.t752 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X177 x4.clknet_1_0__leaf_clk.t13 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X178 a_28647_n9483# x4._11_.t8 a_28457_n9803# VSS.t895 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X179 a_24220_n9483# x4.net5 VSS.t835 VSS.t834 sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6890,366
X180 a_28895_n8715# a_28031_n8709# a_28638_n8741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X181 VDD VSS.t987 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X182 a_26998_n8893# a_26559_n9259# a_26913_n9259# VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X183 a_28565_n8715# a_28031_n8709# a_28470_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X184 VDD a_23927_n8715# a_24095_n8741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X185 VSS.t620 VDD VSS.t619 VSS.t618 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X186 VDD VSS.t988 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X187 x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_5.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X188 x4._19_ a_25359_n7627# VSS.t233 VSS.t232 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X189 VDD VSS.t989 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X190 x4.clknet_1_1__leaf_clk.t28 a_27194_n8171# VSS.t287 VSS.t286 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X191 VSS.t225 a_21119_n968.t4 drv_out.t17 VSS.t224 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X192 VSS.t617 VDD VSS.t616 VSS.t615 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X193 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t12 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X194 VDD x4.clknet_0_clk.t36 a_27194_n8171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X195 a_23505_n9259# a_23339_n9259# VSS.t120 VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X196 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t11 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X197 VSS.t614 VDD VSS.t613 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X198 VDD a_25229_n10182# counter3.t2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X199 a_25359_n7627# a_25179_n7627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X200 VDD VSS.t990 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X201 VDD a_28638_n8741# a_28565_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X202 VSS.t33 x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_7.A VSS.t32 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X203 x1.sky130_fd_sc_hd__nand2_2_0.B x1.sky130_fd_sc_hd__inv_2_9.A VSS.t223 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X204 VDD x3.x2.GN4 x3.x2.GP4.t1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X205 VDD VSS.t991 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X206 a_23505_n9259# a_23339_n9259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X207 a_25709_n7109# drv_out.t21 VSS.t880 VSS.t879 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X208 a_24125_n10182# x4.net4 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X209 VSS.t803 a_25779_n7395# x4.net7 VSS.t802 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X210 x1.sky130_fd_sc_hd__inv_2_11.A ring_out.t11 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X211 VSS.t46 a_27251_n7408# x4._05_ VSS.t45 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X212 VSS.t766 x4.net4 x4._13_ VSS.t765 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X213 VSS.t612 VDD VSS.t611 VSS.t610 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X214 VDD x4._11_.t9 a_25729_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6400,264 d=6600,266
X215 VDD x4._24_ a_28579_n7627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X216 VSS.t609 VDD VSS.t608 VSS.t607 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X217 VSS.t606 VDD VSS.t605 VSS.t604 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X218 x4.clknet_0_clk.t10 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X219 a_25709_n7109# drv_out.t22 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X220 VSS.t213 a_27055_n8715# a_27223_n8741# VSS.t212 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X221 x4.clknet_1_0__leaf_clk.t29 a_23225_n7109# VSS.t702 VSS.t701 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X222 VDD x4.net5 a_25211_n9465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X223 VDD VSS.t992 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X224 VSS.t939 x4._21_ a_25900_n8197# VSS.t938 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4010,197
X225 a_26630_n8715# a_26191_n8709# a_26545_n8715# VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X226 VSS.t603 VDD VSS.t602 VSS.t601 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X227 VDD VSS.t993 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X228 a_23610_n4907# a_23295_n4755# VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X229 VSS.t700 a_23225_n7109# x4.clknet_1_0__leaf_clk.t28 VSS.t699 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X230 VSS.t600 VDD VSS.t599 VSS.t598 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X231 VSS.t285 a_27194_n8171# x4.clknet_1_1__leaf_clk.t27 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X232 VSS.t144 x4.clknet_0_clk.t37 a_27194_n8171# VSS.t143 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X233 x4.clknet_1_0__leaf_clk.t11 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X234 a_24054_n7805# a_23615_n8171# a_23969_n8171# VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X235 a_24479_n7805# a_23781_n8171# a_24222_n8059# VSS.t737 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X236 VDD VSS.t994 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X237 a_21119_n968.t1 ring_out.t12 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=34800,1316 d=34800,1316
X238 VSS.t84 x4._14_ a_24220_n9483# VSS.t83 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=4290,196 d=3510,184
X239 VDD a_19061_n2032# x3.x2.GN4 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X240 x4._12_ x4.net3.t3 a_22879_n5451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X241 VSS.t774 a_28895_n8893# a_29063_n8991# VSS.t773 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X242 VDD a_24371_n8991# a_24287_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X243 x1.sky130_fd_sc_hd__inv_2_15.A x1.sky130_fd_sc_hd__inv_2_14.A VSS.t964 VSS.t786 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X244 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t10 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X245 VDD x4._15_ a_27807_n9829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=3108,158
X246 VSS.t597 VDD VSS.t596 VSS.t595 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X247 VDD x4.clknet_0_clk.t38 a_27194_n8171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X248 x4.net5 a_24371_n8991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X249 VSS.t954 x4._22_ a_28743_n9483# VSS.t953 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.104 ps=0.97 w=0.65 l=0.15
**devattr s=4160,194 d=4485,199
X250 VDD x1.sky130_fd_sc_hd__inv_2_9.A x1.sky130_fd_sc_hd__nand2_2_0.B VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X251 VDD x4.net1 a_23615_n5995# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X252 x1.sky130_fd_sc_hd__inv_2_12.A x1.sky130_fd_sc_hd__inv_2_11.A VSS.t320 VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X253 VDD select1.t3 a_19061_n2032# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X254 x3.x2.GP4.t0 x3.x2.GN4 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X255 VSS.t594 VDD VSS.t593 VSS.t592 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X256 x4.clknet_0_clk.t25 a_25709_n7109# VSS.t104 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X257 a_25709_n7109# drv_out.t23 VSS.t882 VSS.t881 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X258 VDD x4._16_.t2 a_26593_n7906# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.129 ps=1.18 w=0.42 l=0.15
**devattr s=5160,236 d=5830,267
X259 VSS.t591 VDD VSS.t590 VSS.t518 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X260 a_23505_n4043# x4.net2.t6 VSS.t843 VSS.t842 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X261 VSS.t1 a_23295_n4755# x4.net2.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X262 a_22837_n10182# x4.net2.t7 VSS.t845 VSS.t844 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X263 a_23927_n8715# a_23229_n8709# a_23670_n8741# VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X264 VDD x1.sky130_fd_sc_hd__inv_2_15.A x1.sky130_fd_sc_hd__inv_2_16.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X265 x4.net10 a_29063_n8741# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X266 VDD x4._11_.t10 a_28551_n9803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6600,266 d=6600,266
X267 x4.clknet_0_clk.t9 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X268 VSS.t870 a_27807_n9829# x4._23_ VSS.t869 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=7851,266
X269 VSS.t589 VDD VSS.t588 VSS.t587 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X270 x4.clknet_1_0__leaf_clk.t27 a_23225_n7109# VSS.t698 VSS.t697 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X271 a_25211_n9465# x4.net4 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X272 a_23205_n10182# x4.net3.t4 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X273 VDD a_24095_n8741# a_24011_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X274 mux_out.t15 x3.x2.GP4.t4 counter7.t5 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X275 a_27549_n9259# a_26559_n9259# a_27423_n8893# VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X276 VDD x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X277 counter3.t5 x3.x2.GN3 mux_out.t9 VSS.t735 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X278 VSS.t586 VDD VSS.t585 VSS.t584 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X279 VSS.t696 a_23225_n7109# x4.clknet_1_0__leaf_clk.t26 VSS.t695 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X280 VSS.t897 x4._11_.t11 x4._01_ VSS.t896 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X281 a_27124_n9259# a_26725_n9259# a_26998_n8893# VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X282 VSS.t884 x4.clknet_0_clk.t39 a_27194_n8171# VSS.t883 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X283 a_23882_n5174# a_23675_n5233# a_24058_n5451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=2730,149
X284 VDD VSS.t995 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X285 x4.clknet_1_0__leaf_clk.t9 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X286 VDD a_27805_n10182# x4.counter[6] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X287 x4.clknet_1_0__leaf_clk.t8 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X288 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t10 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X289 ring_out.t9 x3.x2.GN1 mux_out.t7 VSS.t358 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X290 a_27507_n8893# a_26725_n9259# a_27423_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X291 x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X292 VSS.t583 VDD VSS.t582 VSS.t558 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X293 VDD x4._21_ a_25900_n8197# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=7430,283
X294 a_28743_n9483# x4._15_ a_28647_n9483# VSS.t868 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4160,194
X295 a_25965_n10182# x4.net6.t2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X296 VSS.t227 a_21119_n968.t5 drv_out.t16 VSS.t226 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X297 VDD VSS.t996 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X298 VDD VSS.t997 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X299 VDD VSS.t998 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X300 VDD x4.net1 a_22879_n5451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=10600,506 d=5900,259
X301 VDD x4._15_ a_27755_n7261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X302 a_27925_n7261# x4.net7 a_27837_n7261# VSS.t816 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X303 x4.clknet_0_clk.t24 a_25709_n7109# VSS.t102 VSS.t101 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X304 VSS.t312 a_25600_n8741# x4._18_ VSS.t311 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=4485,199
X305 VSS.t581 VDD VSS.t580 VSS.t579 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X306 a_24031_n4907# a_23811_n4907# VSS.t333 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.074954 pd=0.823846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4838,217 d=2784,153
X307 VDD x4._05_ a_26713_n7249# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=4368,272
X308 a_24054_n7805# a_23781_n8171# a_23969_n8171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X309 a_18585_n1958# select0.t1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X310 a_23675_n4933# x4.clknet_1_0__leaf_clk.t34 VSS.t247 VSS.t246 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X311 VDD a_25965_n10182# x4.counter[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X312 a_23994_n9687# x4._16_.t3 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=7430,283 d=4704,280
X313 VSS.t578 VDD VSS.t577 VSS.t576 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X314 VSS.t349 a_23255_n4363# x4._00_ VSS.t348 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X315 a_23502_n8715# a_23229_n8709# a_23417_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X316 a_17405_n2032# x3.x1.nSEL0 a_17579_n1926# VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X317 a_23882_n4933# a_23675_n4933# a_24058_n4541# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=2730,149
X318 VDD VSS.t999 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X319 x4._12_ x4.net2.t8 a_22962_n5131# VSS.t846 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
**devattr s=3835,189 d=3640,186
X320 a_24316_n9803# x4._14_ a_23851_n9829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=4200,242
X321 a_17857_n2290# select0.t2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X322 x4.clknet_1_0__leaf_clk.t25 a_23225_n7109# VSS.t694 VSS.t693 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X323 x4._02_ x4._13_ VSS.t330 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X324 VSS.t575 VDD VSS.t574 VSS.t573 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X325 x4.clknet_1_0__leaf_clk.t24 a_23225_n7109# VSS.t692 VSS.t691 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X326 VDD a_27223_n8741# a_27139_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X327 VSS.t283 a_27194_n8171# x4.clknet_1_1__leaf_clk.t26 VSS.t282 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X328 a_23781_n8171# a_23615_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X329 VDD a_28725_n10182# counter7.t0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X330 a_26816_n8171# x4._22_ a_26593_n7906# VSS.t952 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2646,147
X331 VDD a_21119_n968.t6 drv_out.t11 VDD sky130_fd_pr__pfet_01v8 ad=2.026362 pd=18.53074 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X332 VDD VSS.t1000 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X333 VDD x4._22_ a_28551_n9803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6400,264 d=6900,269
X334 a_28638_n8741# a_28470_n8715# VSS.t251 VSS.t250 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X335 VDD select1.t4 x3.x1.nSEL1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X336 VDD VSS.t1001 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X337 a_26542_n7627# a_26295_n7249# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=7155,252 d=3066,157
X338 VSS.t759 select1.t5 a_18033_n1958# VSS.t758 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X339 a_24595_n9571# x4.net4 a_24769_n9465# VSS.t764 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X340 a_29021_n9259# a_28031_n9259# a_28895_n8893# VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X341 VSS.t199 a_23946_n9147# a_23904_n9259# VSS.t198 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X342 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_17.Y VSS.t751 VSS.t750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X343 VDD a_21119_n968.t7 drv_out.t10 VDD sky130_fd_pr__pfet_01v8 ad=2.026362 pd=18.53074 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X344 a_26366_n7350# a_26159_n7409# a_26542_n7627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=2730,149
X345 a_19207_65# x1.sky130_fd_sc_hd__nand2_2_0.B VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X346 a_23295_n5219# a_23391_n5219# VSS.t781 VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X347 VDD x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__inv_2_9.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X348 VDD enable_ring.t0 ring_out.t0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X349 x1.sky130_fd_sc_hd__inv_2_16.A x1.sky130_fd_sc_hd__inv_2_15.A VSS.t306 VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X350 VDD a_27807_n9829# x4._23_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=12498,336
X351 VSS.t572 VDD VSS.t571 VSS.t570 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X352 VDD a_26885_n10182# x4.counter[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X353 VDD VSS.t1002 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X354 drv_out.t9 a_21119_n968.t8 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=2.026362 ps=18.53074 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X355 VDD a_21119_n968.t9 drv_out.t8 VDD sky130_fd_pr__pfet_01v8 ad=2.026362 pd=18.53074 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=111600,3724
X356 VSS.t860 a_23882_n4933# a_23811_n4907# VSS.t794 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.126592 ps=1.2736 w=0.64 l=0.15
**devattr s=3956,199 d=4838,217
X357 VSS.t569 VDD VSS.t568 VSS.t567 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X358 VDD VSS.t1003 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X359 VDD x4.net5 a_24316_n9803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=11200,512
X360 x1.sky130_fd_sc_hd__inv_2_13.A x1.sky130_fd_sc_hd__inv_2_12.A VSS.t316 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X361 x1.sky130_fd_sc_hd__nand2_2_0.B x1.sky130_fd_sc_hd__inv_2_9.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X362 VSS.t921 x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_3.A VSS.t194 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X363 VSS.t220 a_23675_n4933# a_23682_n4633# VSS.t39 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X364 VSS.t566 VDD VSS.t565 VSS.t564 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X365 a_26798_n8741# a_26630_n8715# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.168863 ps=1.544228 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X366 VSS.t357 x3.x2.GN1 x3.x2.GP1.t3 VSS.t356 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X367 a_26630_n8715# a_26357_n8709# a_26545_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X368 a_19207_65# enable_ring.t1 ring_out.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X369 drv_out.t7 a_21119_n968.t10 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=2.026362 ps=18.53074 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X370 VDD x1.sky130_fd_sc_hd__inv_2_16.A x1.sky130_fd_sc_hd__inv_2_17.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X371 a_17579_n1926# x3.x1.nSEL1 VSS.t928 VSS.t927 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X372 VDD a_25709_n7109# x4.clknet_0_clk.t8 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X373 a_28551_n9803# x4._15_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=6600,266 d=6400,264
X374 VDD a_29645_n10182# x4.counter[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X375 VSS.t563 VDD VSS.t562 VSS.t561 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X376 a_23946_n9147# a_23778_n8893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.168863 ps=1.544228 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X377 x1.sky130_fd_sc_hd__inv_2_17.A x1.sky130_fd_sc_hd__inv_2_16.A VSS.t192 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X378 VDD a_24647_n7903# a_24563_n7805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X379 a_29321_n9483# x4._23_ x4._09_ VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=3510,184
X380 VSS.t560 VDD VSS.t559 VSS.t558 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X381 VDD x4.clknet_1_0__leaf_clk.t35 a_23615_n8171# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X382 a_23628_n8337# a_23229_n8709# a_23502_n8715# VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X383 VDD x4.net2.t9 a_23337_n4363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X384 a_28979_n8715# a_28197_n8709# a_28895_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X385 VSS.t903 a_28895_n8715# a_29063_n8741# VSS.t902 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X386 VDD VSS.t1004 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X387 VDD VSS.t1005 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X388 VDD a_25600_n8741# x4._18_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6900,269
X389 VDD VSS.t1006 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X390 a_28470_n8715# a_28031_n8709# a_28385_n8715# VSS.t898 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X391 mux_out.t5 x3.x2.GP3 counter3.t1 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X392 a_28031_n7261# x4._11_.t12 a_27925_n7261# VSS.t740 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X393 a_24769_n9465# x4._11_.t13 VSS.t742 VSS.t741 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X394 a_19061_n2032# select0.t3 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X395 mux_out.t4 x3.x2.GP3 counter3.t0 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X396 a_26979_n9829# x4.net6.t3 a_27377_n9437# VSS.t824 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=4368,272
X397 VDD VSS.t1007 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X398 VSS.t326 a_25229_n10182# counter3.t3 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X399 a_24813_n8395# x4._16_.t4 x4._04_ VSS.t877 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=3510,184
X400 a_23811_n5073# a_23675_n5233# a_23391_n5219# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.078615 pd=0.771795 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4380,215
X401 VSS.t64 x4._01_ a_24229_n5073# VSS.t63 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.087554 ps=0.893846 w=0.42 l=0.15
**devattr s=3252,166 d=4368,272
X402 a_24125_n10182# x4.net4 VSS.t763 VSS.t762 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X403 a_25779_n7395# a_25875_n7395# VSS.t183 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X404 VSS.t557 VDD VSS.t556 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X405 VDD VSS.t1008 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.97
**devattr d=9048,452
X406 VSS.t100 a_25709_n7109# x4.clknet_0_clk.t23 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X407 VSS.t867 x4._15_ a_28031_n7261# VSS.t866 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X408 a_18409_n2290# a_18585_n1958# a_18537_n1898# VSS.t823 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X409 VDD a_26366_n7350# a_26295_n7249# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.168863 pd=1.544228 as=0.140385 ps=1.378205 w=0.75 l=0.15
**devattr s=4380,215 d=7155,252
X410 a_25229_n10182# x4.net5 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X411 VSS.t134 x4._05_ a_26713_n7249# VSS.t133 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.087554 ps=0.893846 w=0.42 l=0.15
**devattr s=3252,166 d=4368,272
X412 x4.net8 a_27223_n8741# VSS.t945 VSS.t944 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X413 x3.x2.GP1.t2 x3.x2.GN1 VSS.t355 VSS.t354 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X414 VSS.t554 VDD VSS.t553 VSS.t536 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X415 x1.sky130_fd_sc_hd__inv_2_9.A x1.sky130_fd_sc_hd__inv_2_7.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X416 x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_6.A VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X417 VDD a_25709_n7109# x4.clknet_0_clk.t7 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X418 a_27807_n9829# x4.net10 a_28205_n9437# VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=4368,272
X419 a_27175_n9437# x4.net9 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0 ps=0 w=0.42 l=0.15
**devattr s=7851,266 d=2772,150
X420 VDD VSS.t1009 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X421 a_25729_n8395# x4._15_ VSS.t865 VSS.t864 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0 ps=0 w=0.65 l=0.15
**devattr s=4485,199 d=4160,194
X422 VDD VSS.t1010 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X423 VDD VSS.t1011 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X424 a_23811_n4907# a_23675_n4933# a_23391_n4933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.078615 pd=0.771795 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4380,215
X425 x4.clknet_0_clk.t6 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X426 a_26756_n8337# a_26357_n8709# a_26630_n8715# VSS.t205 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X427 VSS.t552 VDD VSS.t551 VSS.t550 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X428 VSS.t181 a_24203_n8893# a_24371_n8991# VSS.t180 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X429 x4._00_ a_23255_n4363# a_23505_n4363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X430 VSS.t549 VDD VSS.t548 VSS.t547 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X431 VSS.t546 VDD VSS.t545 VSS.t460 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X432 x4._16_.t1 a_25211_n9231# VSS.t219 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X433 VDD x4._17_ a_25179_n7627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X434 a_24180_n8171# a_23781_n8171# a_24054_n7805# VSS.t736 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X435 x4.net11 a_29063_n8991# VSS.t245 VSS.t244 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X436 a_28385_n9259# x4._09_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X437 x4.clknet_1_1__leaf_clk.t9 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X438 VDD x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_7.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X439 x1.sky130_fd_sc_hd__inv_2_14.A x1.sky130_fd_sc_hd__inv_2_13.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X440 VSS.t544 VDD VSS.t543 VSS.t542 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X441 a_23255_n4363# x4.net1 VSS.t258 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X442 a_23391_n5219# a_23682_n5329# a_23633_n5451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=2268,138
X443 x4._16_.t0 a_25211_n9231# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X444 a_23670_n8741# a_23502_n8715# VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X445 VDD VSS.t1012 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X446 x4._24_ a_28457_n9803# VSS.t837 VSS.t836 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0 ps=0 w=0.65 l=0.15
**devattr s=4485,199 d=6890,366
X447 VSS.t541 VDD VSS.t540 VSS.t539 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X448 VDD VSS.t1013 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X449 x4._00_ x4.net1 a_23505_n4043# VSS.t256 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X450 a_25449_n7261# a_25179_n7627# a_25359_n7627# VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X451 VSS.t538 VDD VSS.t537 VSS.t536 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X452 VDD a_23295_n5219# x4.net3.t0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X453 a_29133_n9803# x4._23_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X454 a_26725_n9259# a_26559_n9259# VSS.t66 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X455 ring_out.t4 enable_ring.t2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X456 VSS.t98 a_25709_n7109# x4.clknet_0_clk.t22 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X457 a_27251_n7408# x4._19_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X458 a_28579_n7627# a_28399_n7627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X459 VDD VSS.t1014 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X460 a_26725_n9259# a_26559_n9259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X461 VSS.t535 VDD VSS.t534 VSS.t533 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X462 VDD VSS.t1015 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X463 VSS.t532 VDD VSS.t531 VSS.t530 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X464 x4.clknet_0_clk.t21 a_25709_n7109# VSS.t96 VSS.t95 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X465 a_26366_n7350# a_26166_n7505# a_26515_n7261# VSS.t822 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.064246 ps=0.706154 w=0.36 l=0.15
**devattr s=2784,153 d=2484,141
X466 VDD VSS.t1016 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X467 a_23205_n10182# x4.net3.t5 VSS.t777 VSS.t776 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X468 VDD VSS.t1017 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X469 VDD a_25709_n7109# x4.clknet_0_clk.t5 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X470 a_28895_n8893# a_28197_n9259# a_28638_n9147# VSS.t930 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X471 VSS.t9 ring_out.t13 x1.sky130_fd_sc_hd__inv_2_11.A VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X472 a_24625_n8715# x4._16_.t5 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X473 a_23417_n8715# x4._02_ VSS.t217 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X474 x4.clknet_1_1__leaf_clk.t25 a_27194_n8171# VSS.t281 VSS.t280 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X475 VSS.t772 a_27805_n10182# x4.counter[6] VSS.t771 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X476 x1.sky130_fd_sc_hd__inv_2_17.Y x1.sky130_fd_sc_hd__inv_2_17.A VSS.t197 VSS.t196 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X477 VDD VSS.t1018 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X478 a_23391_n4933# a_23682_n4633# a_23633_n4541# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=2268,138
X479 VSS.t363 VDD x3.nselect2 VSS.t362 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X480 VDD VSS.t1019 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X481 a_25600_n8741# x4.net6.t4 a_25823_n8395# VSS.t825 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X482 VDD a_18409_n2290# x3.x2.GN3 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X483 a_23225_n7109# x4.clknet_0_clk.t40 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X484 a_25965_n10182# x4.net6.t5 VSS.t827 VSS.t826 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X485 VSS.t70 a_27166_n9147# a_27124_n9259# VSS.t69 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X486 VDD a_29063_n8741# a_28979_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X487 VSS.t529 VDD VSS.t528 VSS.t527 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X488 VSS.t932 a_21119_n968.t11 drv_out.t15 VSS.t931 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X489 VDD VSS.t1020 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X490 VSS.t526 VDD VSS.t525 VSS.t524 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X491 VSS.t523 VDD VSS.t522 VSS.t521 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X492 VSS.t152 a_24647_n7903# a_24605_n8171# VSS.t151 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X493 VDD x1.sky130_fd_sc_hd__inv_2_17.Y x1.sky130_fd_sc_hd__inv_2_8.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X494 VDD a_27591_n8991# a_27507_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X495 VDD a_22837_n10182# x4.counter[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X496 VSS.t797 a_25965_n10182# x4.counter[4] VSS.t796 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X497 VSS.t351 a_23927_n8715# a_24095_n8741# VSS.t350 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X498 a_25729_n8715# x4._15_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=6900,269 d=6400,264
X499 counter7.t2 x3.x2.GN4 mux_out.t3 VSS.t238 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X500 x4.net9 a_27591_n8991# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X501 VSS.t94 a_25709_n7109# x4.clknet_0_clk.t20 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X502 x4._19_ a_25359_n7627# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X503 a_23882_n4933# a_23682_n4633# a_24031_n4907# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.064246 ps=0.706154 w=0.36 l=0.15
**devattr s=2784,153 d=2484,141
X504 VDD VSS.t1021 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X505 VSS.t520 VDD VSS.t519 VSS.t518 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X506 VDD drv_out.t24 a_25709_n7109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X507 VSS.t517 VDD VSS.t516 VSS.t515 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X508 x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__inv_2_7.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X509 VSS.t82 x4._14_ x4._02_ VSS.t81 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X510 VDD VSS.t1022 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X511 VSS.t514 VDD VSS.t513 VSS.t512 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X512 a_23295_n4755# a_23391_n4933# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X513 a_24058_n5451# a_23811_n5073# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=7155,252 d=3066,157
X514 VDD x4.clknet_1_1__leaf_clk.t34 a_26191_n8709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X515 VSS.t23 a_28725_n10182# counter7.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X516 VSS.t721 select0.t4 x3.x1.nSEL0 VSS.t720 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X517 a_23225_n7109# x4.clknet_0_clk.t41 VSS.t886 VSS.t885 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X518 a_23969_n8171# x4._04_ VSS.t807 VSS.t806 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X519 a_28638_n8741# a_28470_n8715# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.168863 ps=1.544228 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X520 a_26545_n8715# x4._06_ VSS.t757 VSS.t756 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X521 VDD a_17857_n2290# x3.x2.GN2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X522 mux_out.t12 x3.x2.GP2.t4 drv_out.t2 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X523 a_27271_n9437# x4.net8 a_27175_n9437# VSS.t855 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3192,160
X524 a_28470_n8715# a_28197_n8709# a_28385_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X525 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t7 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X526 VSS.t511 VDD VSS.t510 VSS.t509 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X527 a_23778_n8893# a_23505_n9259# a_23693_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X528 VDD x1.sky130_fd_sc_hd__nand2_2_0.B ring_out.t3 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X529 VDD a_26593_n7906# a_26529_n7849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0672 ps=0.74 w=0.42 l=0.15
**devattr s=2688,148 d=8370,269
X530 x4._24_ a_28457_n9803# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=6900,269 d=10600,506
X531 x4._21_ a_25639_n9259# VSS.t148 VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X532 VSS.t508 VDD VSS.t507 VSS.t506 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X533 x3.nselect2 VDD VSS.t505 VSS.t504 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X534 VSS.t734 x3.x2.GN3 x3.x2.GP3 VSS.t733 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X535 x4.clknet_1_0__leaf_clk.t6 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X536 x4._04_ a_24595_n8741# VSS.t215 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0 ps=0 w=0.65 l=0.15
**devattr s=8320,388 d=10010,284
X537 a_24595_n8741# x4.net6.t6 VSS.t142 VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X538 a_25179_n7627# x4._17_ VSS.t915 VSS.t914 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X539 x4._21_ a_25639_n9259# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X540 VSS.t820 a_26885_n10182# x4.counter[5] VSS.t819 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X541 a_27166_n9147# a_26998_n8893# VSS.t185 VSS.t184 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X542 mux_out.t0 x3.x2.GP1.t4 ring_out.t6 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X543 VSS.t888 drv_out.t25 a_25709_n7109# VSS.t887 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X544 VSS.t503 VDD VSS.t502 VSS.t477 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X545 a_24058_n4541# a_23811_n4907# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=7155,252 d=3066,157
X546 a_24203_n8893# a_23505_n9259# a_23946_n9147# VSS.t178 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X547 VSS.t713 a_17405_n2032# x3.x2.GN1 VSS.t712 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X548 x4._11_.t3 a_24075_n5995# VSS.t191 VSS.t190 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2730,149 d=2268,138
X549 a_22885_n8715# x4._13_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X550 VSS.t76 x1.sky130_fd_sc_hd__nand2_2_0.B a_19207_65# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X551 x1.sky130_fd_sc_hd__inv_2_15.A x1.sky130_fd_sc_hd__inv_2_14.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X552 VDD a_25709_n7109# x4.clknet_0_clk.t4 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X553 a_28003_n9437# x4._22_ VSS.t951 VSS.t950 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0 ps=0 w=0.42 l=0.15
**devattr s=7851,266 d=2772,150
X554 a_26529_n7849# a_26593_n7906# a_26375_n8171# VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X555 VDD drv_out.t26 a_25709_n7109# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X556 VDD VSS.t1023 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X557 VDD VSS.t1024 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X558 VSS.t690 a_23225_n7109# x4.clknet_1_0__leaf_clk.t23 VSS.t689 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X559 a_28999_n7408# x4._25_ VSS.t852 VSS.t851 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X560 a_25729_n8715# x4.net6.t7 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=6600,266 d=6600,266
X561 VSS.t302 a_29645_n10182# x4.counter[8] VSS.t301 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X562 x1.sky130_fd_sc_hd__inv_2_12.A x1.sky130_fd_sc_hd__inv_2_11.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X563 VSS.t128 x4.net11 a_29321_n9483# VSS.t127 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X564 x4._11_.t1 a_24075_n5995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=6500,265 d=5400,254
X565 x4.clknet_1_0__leaf_clk.t22 a_23225_n7109# VSS.t688 VSS.t687 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X566 drv_out.t6 a_21119_n968.t12 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=2.026362 ps=18.53074 w=9 l=0.15
**devattr s=111600,3724 d=59400,1866
X567 a_18033_n1958# select1.t6 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X568 x3.x1.nSEL0 select0.t5 VSS.t723 VSS.t722 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X569 a_23505_n4363# x4.net2.t10 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X570 x4.net10 a_29063_n8741# VSS.t56 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X571 VSS.t715 x4._16_.t6 a_26816_n8171# VSS.t714 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2646,147 d=3945,196
X572 VDD VSS.t1025 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X573 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t5 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X574 VDD x4.net6.t8 a_26979_n9829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=4368,272
X575 VSS.t318 x1.sky130_fd_sc_hd__inv_2_11.A x1.sky130_fd_sc_hd__inv_2_12.A VSS.t317 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X576 VSS.t924 a_24595_n9571# x4._14_ VSS.t923 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X577 VSS.t501 VDD VSS.t500 VSS.t499 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X578 VDD x4._01_ a_24229_n5073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=4368,272
X579 a_26117_n7627# a_25779_n7395# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4452,274 d=3528,168
X580 a_26593_n7906# x4._22_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=8370,269 d=5160,236
X581 ring_out.t5 enable_ring.t3 a_19207_65# VSS.t203 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X582 drv_out.t5 a_21119_n968.t13 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=2.026362 ps=18.53074 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X583 VDD VSS.t1026 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X584 VSS.t815 x4.net7 a_25600_n8741# VSS.t814 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=8320,388
X585 VSS.t872 x4.net6.t9 a_24813_n8395# VSS.t871 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X586 a_28596_n8337# a_28197_n8709# a_28470_n8715# VSS.t893 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X587 VSS.t498 VDD VSS.t497 VSS.t463 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X588 VSS.t496 VDD VSS.t495 VSS.t494 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X589 x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_3.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X590 VDD VSS.t1027 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X591 VSS.t876 x4.clknet_1_1__leaf_clk.t35 a_26559_n9259# VSS.t875 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X592 VSS.t493 VDD VSS.t492 VSS.t491 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X593 VSS.t854 x4.net8 a_25667_n8171# VSS.t853 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=6890,366 d=3510,184
X594 x4._02_ x4._14_ a_22885_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X595 VDD a_21119_n968.t14 drv_out.t4 VDD sky130_fd_pr__pfet_01v8 ad=2.026362 pd=18.53074 as=0 ps=0 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X596 VDD VSS.t1028 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X597 VSS.t92 a_25709_n7109# x4.clknet_0_clk.t19 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X598 VSS.t890 drv_out.t27 a_25709_n7109# VSS.t889 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X599 VDD a_23205_n10182# x4.counter[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X600 a_23675_n4933# x4.clknet_1_0__leaf_clk.t36 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X601 VSS.t490 VDD VSS.t489 VSS.t422 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X602 VDD x4.clknet_1_1__leaf_clk.t36 a_26559_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X603 VDD VSS.t1029 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X604 mux_out.t14 x3.x2.GP4.t5 counter7.t4 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X605 a_25229_n10182# x4.net5 VSS.t833 VSS.t832 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X606 VDD VSS.t1030 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X607 VDD x4.net10 a_27807_n9829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=4368,272
X608 a_26979_n9829# x4.net9 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=12498,336 d=2352,140
X609 a_23781_n8171# a_23615_n8171# VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X610 VDD x3.x2.GN1 x3.x2.GP1.t1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X611 VSS.t686 a_23225_n7109# x4.clknet_1_0__leaf_clk.t21 VSS.t685 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X612 x4.net6.t0 a_24647_n7903# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X613 VDD x4._00_ a_24229_n4907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=4368,272
X614 a_24222_n8059# a_24054_n7805# VSS.t140 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X615 VDD VSS.t1031 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X616 VDD x4.net11 a_29319_n10347# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X617 a_24981_n8715# x4.net6.t10 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X618 VDD x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X619 a_19061_n2032# select1.t7 a_19235_n1926# VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X620 VSS.t488 VDD VSS.t487 VSS.t486 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X621 VSS.t485 VDD VSS.t484 VSS.t483 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X622 VSS.t717 x4._16_.t7 a_24595_n8741# VSS.t716 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X623 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t4 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X624 VDD a_23225_n7109# x4.clknet_1_0__leaf_clk.t3 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X625 a_24229_n4907# a_23675_n4933# a_23882_n4933# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.075046 pd=0.766154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=3252,166
X626 x4.net5 a_24371_n8991# VSS.t341 VSS.t340 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X627 a_23693_n9259# x4._03_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X628 VDD VSS.t1032 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X629 VSS.t27 x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_4.A VSS.t26 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X630 a_22879_n5451# x4.net2.t11 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5900,259 d=5600,256
X631 a_27166_n9147# a_26998_n8893# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.168863 ps=1.544228 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X632 VSS.t482 VDD VSS.t481 VSS.t480 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
**devattr d=5720,324
X633 VSS.t831 x4.net5 a_25297_n9465# VSS.t830 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X634 VDD VSS.t1033 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X635 a_27377_n9437# x4.net7 a_27271_n9437# VSS.t813 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2436,142
X636 VSS.t479 VDD VSS.t478 VSS.t477 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X637 ring_out.t2 x1.sky130_fd_sc_hd__nand2_2_0.B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X638 x4._07_ a_26529_n7849# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5830,267 d=10400,504
X639 VDD a_24125_n10182# x4.counter[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X640 VSS.t476 VDD VSS.t475 VSS.t474 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X641 VDD a_27423_n8893# a_27591_n8991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X642 a_23670_n8741# a_23502_n8715# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.168863 ps=1.544228 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X643 VDD VSS.t1034 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X644 VSS.t770 x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_5.A VSS.t303 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X645 VSS.t473 VDD VSS.t472 VSS.t446 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X646 VDD x4.net11 a_29133_n9803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X647 VSS.t471 VDD VSS.t470 VSS.t469 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X648 VDD a_23675_n4933# a_23682_n4633# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X649 a_28385_n9259# x4._09_ VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X650 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_17.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X651 VDD a_28999_n7408# x4._08_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X652 VDD VSS.t1035 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X653 VDD a_24595_n9571# x4._14_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X654 VSS.t468 VDD VSS.t467 VSS.t466 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X655 a_23417_n8715# x4._02_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X656 VDD VSS.t1036 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X657 VDD VSS.t1037 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X658 VSS.t684 a_23225_n7109# x4.clknet_1_0__leaf_clk.t20 VSS.t683 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X659 VSS.t682 a_23225_n7109# x4.clknet_1_0__leaf_clk.t19 VSS.t681 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X660 VSS.t48 x4.clknet_1_0__leaf_clk.t37 a_23615_n8171# VSS.t47 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X661 a_24329_n9259# a_23339_n9259# a_24203_n8893# VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X662 VSS.t839 x4.clknet_1_1__leaf_clk.t37 a_26191_n8709# VSS.t838 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X663 x1.sky130_fd_sc_hd__inv_2_16.A x1.sky130_fd_sc_hd__inv_2_15.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X664 x3.x2.GP1.t0 x3.x2.GN1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X665 VDD a_24479_n7805# a_24647_n7903# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X666 a_28205_n9437# x4._11_.t14 a_28099_n9437# VSS.t743 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2436,142
X667 VDD x4._11_.t15 a_25639_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X668 a_23229_n8709# a_23063_n8709# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X669 a_26979_n9829# x4.net7 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=3108,158 d=2940,154
X670 a_25600_n8741# x4.net7 a_25729_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6600,266 d=12800,528
X671 VDD x4.net6.t11 a_24625_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X672 a_17857_n2290# a_18033_n1958# a_17985_n1898# VSS.t793 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X673 VDD VSS.t1038 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X674 a_26713_n7249# a_26159_n7409# a_26366_n7350# VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.075046 pd=0.766154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=3252,166
X675 a_25721_n9259# x4._11_.t16 a_25639_n9259# VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X676 VDD VSS.t1039 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X677 x1.sky130_fd_sc_hd__inv_2_13.A x1.sky130_fd_sc_hd__inv_2_12.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X678 x3.x2.GP3 x3.x2.GN3 VSS.t732 VSS.t731 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X679 VSS.t729 a_27591_n8991# a_27549_n9259# VSS.t728 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X680 a_26725_n8715# a_26191_n8709# a_26630_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X681 VDD x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_2.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X682 VSS.t465 VDD VSS.t464 VSS.t463 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X683 x4._07_ a_26529_n7849# VSS.t761 VSS.t760 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3945,196 d=6760,364
X684 counter3.t4 x3.x2.GN3 mux_out.t8 VSS.t730 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X685 VDD x4.clknet_1_1__leaf_clk.t38 a_28031_n8709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X686 VSS.t314 x1.sky130_fd_sc_hd__inv_2_12.A x1.sky130_fd_sc_hd__inv_2_13.A VSS.t313 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X687 VDD x4.net7 a_27755_n7261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X688 a_28385_n8715# x4._08_ VSS.t345 VSS.t344 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X689 a_25297_n9465# x4.net4 a_25211_n9465# VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X690 VDD a_26798_n8741# a_26725_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X691 VDD VSS.t1040 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X692 x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__inv_2_7.A VSS.t339 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X693 VSS.t462 VDD VSS.t461 VSS.t460 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X694 x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_2.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X695 x1.sky130_fd_sc_hd__inv_2_17.A x1.sky130_fd_sc_hd__inv_2_16.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X696 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t8 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X697 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t7 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X698 VDD x4._23_ a_28399_n7627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X699 a_27807_n9829# x4._11_.t17 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=3108,158 d=2940,154
X700 VDD a_23882_n4933# a_23811_n4907# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.168863 pd=1.544228 as=0.140385 ps=1.378205 w=0.75 l=0.15
**devattr s=4380,215 d=7155,252
X701 VSS.t207 a_22837_n10182# x4.counter[0] VSS.t206 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X702 a_26375_n8171# x4.net9 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X703 a_23994_n9687# x4._16_.t8 VSS.t719 VSS.t718 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=4010,197 d=4368,272
X704 a_24595_n8741# x4._16_.t9 a_24981_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X705 VDD VSS.t1041 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X706 VDD a_27251_n7408# x4._05_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.17787 pd=1.626587 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X707 drv_out.t14 a_21119_n968.t15 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X708 a_23941_n3056# enable_counter VSS.t780 VSS.t779 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X709 x1.sky130_fd_sc_hd__inv_2_9.A x1.sky130_fd_sc_hd__inv_2_7.Y VSS.t324 VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X710 x3.x2.GP2.t3 x3.x2.GN2 VSS.t748 VSS.t747 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X711 VDD a_23882_n5174# a_23811_n5073# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.168863 pd=1.544228 as=0.140385 ps=1.378205 w=0.75 l=0.15
**devattr s=4380,215 d=7155,252
X712 VSS.t459 VDD VSS.t458 VSS.t457 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X713 VDD VSS.t1042 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X714 VSS.t322 x4._24_ a_28669_n7261# VSS.t321 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X715 VSS.t456 VDD VSS.t455 VSS.t454 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X716 a_25793_n9259# x4._15_ a_25721_n9259# VSS.t863 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X717 a_26545_n8715# x4._06_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X718 VSS.t260 x1.sky130_fd_sc_hd__inv_2_13.A x1.sky130_fd_sc_hd__inv_2_14.A VSS.t32 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X719 x4.clknet_0_clk.t3 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X720 VSS.t164 x4._23_ a_29103_n9829# VSS.t163 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X721 a_27181_n8337# a_26191_n8709# a_27055_n8715# VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X722 VSS.t453 VDD VSS.t452 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X723 VDD VSS.t1043 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X724 x4._17_ a_27755_n7261# VSS.t966 VSS.t965 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X725 a_28669_n7261# a_28399_n7627# a_28579_n7627# VSS.t775 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X726 VDD a_24222_n8059# a_24149_n7805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X727 a_25762_n7921# x4.net8 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=11200,512 d=4200,242
X728 a_26357_n8709# a_26191_n8709# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X729 VDD VSS.t1044 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X730 VDD VSS.t1045 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X731 a_28470_n8893# a_28031_n9259# a_28385_n9259# VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X732 VDD VSS.t1046 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X733 VDD a_23670_n8741# a_23597_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X734 a_26147_n9107# x4.net8 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=5689,267 d=2646,147
X735 VDD VSS.t1047 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X736 VSS.t783 a_23295_n5219# x4.net3.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X737 VSS.t451 VDD VSS.t450 VSS.t449 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X738 VDD VDD x3.nselect2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X739 VDD VSS.t1048 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X740 VSS.t279 a_27194_n8171# x4.clknet_1_1__leaf_clk.t24 VSS.t278 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X741 VSS.t277 a_27194_n8171# x4.clknet_1_1__leaf_clk.t23 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X742 a_28895_n8893# a_28031_n9259# a_28638_n9147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X743 x4.clknet_1_1__leaf_clk.t6 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X744 VSS.t448 VDD VSS.t447 VSS.t446 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X745 a_28565_n8893# a_28031_n9259# a_28470_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X746 VSS.t445 VDD VSS.t444 VSS.t443 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X747 VDD VSS.t1049 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X748 a_23811_n4907# a_23682_n4633# a_23391_n4933# VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.071208 pd=0.7164 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=3956,199
X749 a_26713_n7249# a_26166_n7505# a_26366_n7350# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=2310,139
X750 a_23882_n5174# a_23682_n5329# a_24031_n5085# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.064246 ps=0.706154 w=0.36 l=0.15
**devattr s=2784,153 d=2484,141
X751 VSS.t943 a_27223_n8741# a_27181_n8337# VSS.t942 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X752 VSS.t442 VDD VSS.t441 VSS.t440 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X753 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t5 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X754 a_27807_n9829# x4._22_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=12498,336 d=2352,140
X755 a_18537_n1898# select1.t8 VSS.t202 VSS.t201 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X756 VDD a_28638_n9147# a_28565_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X757 VDD x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_7.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X758 x4.clknet_0_clk.t18 a_25709_n7109# VSS.t90 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X759 VSS.t60 x4._20_ a_25793_n9259# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X760 VSS.t937 x4._21_ a_26375_n8171# VSS.t936 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X761 VSS.t439 VDD VSS.t438 VSS.t437 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X762 VSS.t436 VDD VSS.t435 VSS.t434 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X763 VSS.t433 VDD VSS.t432 VSS.t431 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X764 VSS.t189 a_24075_n5995# x4._11_.t2 VSS.t188 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X765 a_25834_n7921# x4._17_ a_25762_n7921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=6600,266
X766 VDD VSS.t1050 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X767 a_19235_n1926# select0.t6 VSS.t958 VSS.t957 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X768 VDD VSS.t1051 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X769 drv_out.t13 a_21119_n968.t16 VSS.t905 VSS.t904 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=37200,1324 d=19800,666
X770 a_23675_n5233# x4.clknet_1_0__leaf_clk.t38 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X771 x4.clknet_0_clk.t2 a_25709_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X772 a_23969_n8171# x4._04_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X773 a_23337_n4363# x4.net1 a_23255_n4363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X774 VDD a_24075_n5995# x4._11_.t0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X775 a_29103_n9829# x4.net11 VSS.t126 VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X776 VSS.t430 VDD VSS.t429 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X777 VDD x4.net1 a_23505_n4363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X778 x4.clknet_1_1__leaf_clk.t22 a_27194_n8171# VSS.t275 VSS.t274 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X779 VDD select0.t7 x3.x1.nSEL0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X780 VDD VSS.t1052 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X781 a_27755_n7261# x4.net6.t12 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X782 x4.clknet_1_0__leaf_clk.t2 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X783 VDD VSS.t1053 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X784 VSS.t273 a_27194_n8171# x4.clknet_1_1__leaf_clk.t21 VSS.t272 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X785 x3.nselect2 VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X786 VDD x3.x2.GN3 x3.x2.GP3 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X787 VSS.t707 x4._00_ a_24229_n4907# VSS.t63 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.087554 ps=0.893846 w=0.42 l=0.15
**devattr s=3252,166 d=4368,272
X788 x4._25_ a_28579_n7627# VSS.t231 VSS.t230 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X789 x4.clknet_1_1__leaf_clk.t4 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X790 x4.clknet_1_1__leaf_clk.t3 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X791 VSS.t907 a_21119_n968.t17 drv_out.t12 VSS.t906 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
**devattr s=19800,666 d=37200,1324
X792 VDD VSS.t1054 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X793 VDD ring_out.t14 x1.sky130_fd_sc_hd__inv_2_11.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X794 a_17985_n1898# select0.t8 VSS.t960 VSS.t959 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X795 a_24222_n8059# a_24054_n7805# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.168863 ps=1.544228 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X796 a_25667_n8171# x4._17_ VSS.t913 VSS.t912 sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=4290,196
X797 a_26998_n8893# a_26725_n9259# a_26913_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X798 mux_out.t1 x3.x2.GP1.t5 ring_out.t7 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X799 VSS.t709 x4.clknet_1_1__leaf_clk.t39 a_28031_n9259# VSS.t708 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X800 VDD a_18585_n1958# a_18409_n2290# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X801 VDD a_27194_n8171# x4.clknet_1_1__leaf_clk.t2 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X802 a_29103_n9829# x4._23_ a_29489_n9803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X803 VSS.t829 a_23205_n10182# x4.counter[1] VSS.t828 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X804 VDD VSS.t1055 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X805 VSS.t427 VDD VSS.t426 VSS.t425 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X806 x1.sky130_fd_sc_hd__inv_2_17.Y x1.sky130_fd_sc_hd__inv_2_17.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X807 a_23941_n3056# enable_counter VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X808 VDD x4.clknet_1_1__leaf_clk.t40 a_28031_n9259# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X809 x4.clknet_0_clk.t17 a_25709_n7109# VSS.t88 VSS.t87 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X810 a_28099_n9437# x4._15_ a_28003_n9437# VSS.t862 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3192,160
X811 a_28399_n7627# x4._23_ VSS.t162 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X812 VDD x4.clknet_1_0__leaf_clk.t39 a_23063_n8709# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X813 VSS.t424 VDD VSS.t423 VSS.t422 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X814 VSS.t421 VDD VSS.t420 VSS.t419 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X815 VSS.t195 x1.sky130_fd_sc_hd__inv_2_17.A x1.sky130_fd_sc_hd__inv_2_17.Y VSS.t194 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X816 a_24625_n8715# a_24595_n8741# x4._04_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.3 ps=2.6 w=1 l=0.15
**devattr s=12000,520 d=10400,504
X817 a_23229_n8709# a_23063_n8709# VSS.t158 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X818 VSS.t861 x4._15_ a_25297_n9231# VSS.t830 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X819 VSS.t124 x4.net11 a_29319_n10347# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X820 VSS.t963 x1.sky130_fd_sc_hd__inv_2_14.A x1.sky130_fd_sc_hd__inv_2_15.A VSS.t788 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X821 VDD a_23675_n5233# a_23682_n5329# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X822 x4.clknet_1_0__leaf_clk.t18 a_23225_n7109# VSS.t680 VSS.t679 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
X823 a_24203_n8893# a_23339_n9259# a_23946_n9147# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X824 a_28457_n9803# x4.net10 VSS.t297 VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0 ps=0 w=0.65 l=0.15
**devattr s=8320,388 d=4290,196
X825 x4.clknet_1_1__leaf_clk.t20 a_27194_n8171# VSS.t271 VSS.t270 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X826 VSS.t418 VDD VSS.t417 VSS.t416 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X827 a_26529_n7849# x4.net9 a_26457_n7849# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2688,148
X828 VDD VSS.t1056 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.97
**devattr d=9048,452
X829 x4.clknet_1_1__leaf_clk.t19 a_27194_n8171# VSS.t269 VSS.t268 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X830 x3.x1.nSEL0 select0.t9 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X831 VSS.t711 x4.clknet_1_1__leaf_clk.t41 a_28031_n8709# VSS.t710 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X832 VDD VSS.t1057 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X833 a_23610_n5085# a_23295_n5219# VSS.t782 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.071077 pd=0.802308 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X834 VSS.t415 VDD VSS.t414 VSS.t391 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X835 x4.counter[9] a_29319_n10347# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X836 VSS.t267 a_27194_n8171# x4.clknet_1_1__leaf_clk.t18 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X837 x4.clknet_1_0__leaf_clk.t1 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X838 VSS.t413 VDD VSS.t412 VSS.t411 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X839 VDD VSS.t1058 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X840 a_27194_n8171# x4.clknet_0_clk.t42 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X841 VSS.t947 a_24125_n10182# x4.counter[2] VSS.t946 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X842 x4.clknet_1_1__leaf_clk.t1 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X843 VDD VSS.t1059 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.97
**devattr d=9048,452
X844 VDD a_28895_n8893# a_29063_n8991# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X845 drv_out.t0 x3.x2.GN2 mux_out.t10 VSS.t746 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X846 a_23693_n9259# x4._03_ VSS.t850 VSS.t849 sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X847 VDD x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_6.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X848 VSS.t795 a_23882_n5174# a_23811_n5073# VSS.t794 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.126592 ps=1.2736 w=0.64 l=0.15
**devattr s=3956,199 d=4838,217
X849 a_29489_n9803# x4.net11 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X850 a_27055_n8715# a_26357_n8709# a_26798_n8741# VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X851 x4._09_ a_29103_n9829# VSS.t130 VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0 ps=0 w=0.65 l=0.15
**devattr s=8320,388 d=10010,284
X852 x4._15_ a_25211_n9465# VSS.t156 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X853 a_28638_n9147# a_28470_n8893# VSS.t892 VSS.t891 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X854 mux_out.t13 x3.x2.GP2.t5 drv_out.t3 VDD sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X855 VDD a_25709_n7109# x4.clknet_0_clk.t1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X856 VDD a_25900_n8197# a_25834_n7921# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=12000,520
X857 a_26357_n8709# a_26191_n8709# VSS.t167 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X858 VSS.t332 a_19061_n2032# x3.x2.GN4 VSS.t331 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X859 a_23295_n4755# a_23391_n4933# VSS.t132 VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X860 a_24229_n5073# a_23675_n5233# a_23882_n5174# VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.075046 pd=0.766154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=3252,166
X861 VDD VSS.t1060 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X862 a_25639_n9259# x4._15_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X863 x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_6.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X864 a_25297_n9231# x4._11_.t18 a_25211_n9231# VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X865 ring_out.t8 x3.x2.GN1 mux_out.t6 VSS.t353 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X866 x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_4.A VSS.t769 VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X867 VDD VSS.t1061 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X868 VSS.t919 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_2.A VSS.t752 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X869 x3.x1.nSEL1 select1.t9 VSS.t926 VSS.t925 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X870 a_23225_n7109# x4.clknet_0_clk.t43 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X871 x4.clknet_1_0__leaf_clk.t17 a_23225_n7109# VSS.t678 VSS.t677 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X872 a_24220_n9483# a_23994_n9687# a_23851_n9829# VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X873 VSS.t410 VDD VSS.t409 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X874 VSS.t255 x4.net1 a_23769_n5995# VSS.t254 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X875 a_28725_n10182# x4.net9 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X876 VSS.t243 a_29063_n8991# a_29021_n9259# VSS.t242 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X877 a_28385_n8715# x4._08_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X878 a_27194_n8171# x4.clknet_0_clk.t44 VSS.t841 VSS.t840 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X879 x4.clknet_1_1__leaf_clk.t17 a_27194_n8171# VSS.t265 VSS.t264 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
X880 x1.sky130_fd_sc_hd__inv_2_11.A ring_out.t15 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X881 a_23391_n4933# a_23675_n4933# a_23610_n4907# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.060923 ps=0.687692 w=0.36 l=0.15
**devattr s=2640,149 d=2736,148
X882 a_28197_n8709# a_28031_n8709# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.144097 ps=1.317742 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X883 VSS.t408 VDD VSS.t407 VSS.t406 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X884 a_27837_n7261# x4.net6.t13 a_27755_n7261# VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X885 VDD VSS.t1062 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X886 x4.clknet_1_0__leaf_clk.t0 a_23225_n7109# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X887 VDD VSS.t1063 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.97
**devattr d=9048,452
X888 x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_5.A VSS.t787 VSS.t786 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X889 VSS.t405 VDD VSS.t404 VSS.t403 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X890 VSS.t402 VDD VSS.t401 VSS.t400 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X891 a_27194_n8171# x4.clknet_0_clk.t45 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X892 VSS.t739 a_24222_n8059# a_24180_n8171# VSS.t738 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X893 x4.net9 a_27591_n8991# VSS.t727 VSS.t726 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X894 a_26913_n9259# x4._07_ VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X895 VDD a_27055_n8715# a_27223_n8741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X896 VSS.t328 a_26979_n9829# x4._22_ VSS.t327 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=7851,266
X897 VSS.t848 a_23851_n9829# x4._03_ VSS.t847 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4010,197
X898 a_26381_n9259# x4.net7 a_26309_n9259# VSS.t812 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X899 VSS.t86 a_25709_n7109# x4.clknet_0_clk.t16 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X900 a_25834_n7921# a_25900_n8197# a_25667_n8171# VSS.t778 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=4290,196 d=6760,364
X901 VDD x1.sky130_fd_sc_hd__inv_2_11.A x1.sky130_fd_sc_hd__inv_2_12.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X902 VDD VSS.t1064 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X903 a_26885_n10182# x4.net7 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X904 a_27055_n8715# a_26191_n8709# a_26798_n8741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X905 VSS.t399 VDD VSS.t398 VSS.t397 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X906 a_24563_n7805# a_23781_n8171# a_24479_n7805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X907 x4._10_ a_23615_n5995# VSS.t310 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X908 a_28551_n9803# x4.net10 a_28457_n9803# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.32 ps=2.64 w=1 l=0.15
**devattr s=12800,528 d=6600,266
X909 VSS.t396 VDD VSS.t395 VSS.t394 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X910 VSS.t745 x3.x2.GN2 x3.x2.GP2.t2 VSS.t744 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X911 VDD a_23295_n4755# x4.net2.t0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X912 a_24031_n5085# a_23811_n5073# VSS.t25 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.074954 pd=0.823846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4838,217 d=2784,153
X913 VSS.t54 a_29063_n8741# a_29021_n8337# VSS.t53 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X914 VDD VSS.t1065 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X915 a_23675_n5233# x4.clknet_1_0__leaf_clk.t40 VSS.t933 VSS.t246 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X916 a_23225_n7109# x4.clknet_0_clk.t46 VSS.t809 VSS.t808 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X917 VDD x4.net4 a_24595_n9571# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X918 VDD x4._15_ a_25211_n9231# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X919 a_24011_n8715# a_23229_n8709# a_23927_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X920 VDD VSS.t1066 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X921 VSS.t35 x4.net3.t6 x4._12_ VSS.t34 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X922 a_23778_n8893# a_23339_n9259# a_23693_n9259# VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X923 x4._10_ a_23615_n5995# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X924 VDD VSS.t1067 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X925 a_29645_n10182# x4.net10 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X926 VSS.t393 VDD VSS.t392 VSS.t391 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X927 VDD a_25779_n7395# x4.net7 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X928 a_26295_n7249# a_26166_n7505# a_25875_n7395# VSS.t821 sky130_fd_pr__nfet_01v8 ad=0.071208 pd=0.7164 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=3956,199
X929 VDD a_26159_n7409# a_26166_n7505# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.144097 pd=1.317742 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X930 VDD a_17405_n2032# x3.x2.GN1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X931 x3.x2.GP3 x3.x2.GN3 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X932 x4.clknet_1_0__leaf_clk.t16 a_23225_n7109# VSS.t676 VSS.t675 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X933 a_26515_n7261# a_26295_n7249# VSS.t792 VSS.t791 sky130_fd_pr__nfet_01v8 ad=0.074954 pd=0.823846 as=0 ps=0 w=0.42 l=0.15
**devattr s=4838,217 d=2784,153
X934 VSS.t390 VDD VSS.t389 VSS.t388 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X935 a_28596_n9259# a_28197_n9259# a_28470_n8893# VSS.t929 sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X936 a_26147_n9107# x4.net6.t14 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X937 a_27194_n8171# x4.clknet_0_clk.t47 VSS.t811 VSS.t810 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X938 x4.clknet_1_1__leaf_clk.t0 a_27194_n8171# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X939 VDD VSS.t1068 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X940 VDD VSS.t1069 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X941 VDD VSS.t1070 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.97
**devattr d=9048,452
X942 a_23873_n8893# a_23339_n9259# a_23778_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X943 a_24229_n5073# a_23682_n5329# a_23882_n5174# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=2310,139
X944 a_28979_n8893# a_28197_n9259# a_28895_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X945 a_26147_n9107# x4.net6.t15 a_26381_n9259# VSS.t790 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=4368,272
X946 VSS.t338 x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_7.Y VSS.t313 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X947 VSS.t304 x1.sky130_fd_sc_hd__inv_2_15.A x1.sky130_fd_sc_hd__inv_2_16.A VSS.t303 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X948 VDD x3.x1.nSEL0 a_17405_n2032# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X949 VDD VSS.t1071 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=4.73
**devattr d=9048,452
X950 x4._15_ a_25211_n9465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X951 VSS.t237 x3.x2.GN4 x3.x2.GP4.t2 VSS.t236 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X952 VDD x4._18_ a_25359_n7627# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X953 a_23946_n9147# a_23778_n8893# VSS.t229 VSS.t228 sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0 ps=0 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X954 VDD a_23946_n9147# a_23873_n8893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X955 VDD VSS.t1072 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=2.89
**devattr d=9048,452
X956 a_27805_n10182# x4.net8 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.17787 ps=1.626587 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X957 a_27251_n7408# x4._19_ VSS.t235 VSS.t234 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X958 VSS.t387 VDD VSS.t386 VSS.t385 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X959 VSS.t323 x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__inv_2_9.A VSS.t317 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X960 VSS.t384 VDD VSS.t383 VSS.t382 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X961 VSS.t381 VDD VSS.t380 VSS.t379 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
**devattr d=5720,324
X962 VSS.t378 VDD VSS.t377 VSS.t376 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X963 VSS.t935 x4.clknet_1_0__leaf_clk.t41 a_23063_n8709# VSS.t934 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X964 a_24479_n7805# a_23615_n8171# a_24222_n8059# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X965 VDD x4.net8 a_26979_n9829# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=3108,158
X966 a_23851_n9829# a_23994_n9687# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=12000,520 d=6600,266
X967 VSS.t956 a_23670_n8741# a_23628_n8337# VSS.t955 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X968 a_24149_n7805# a_23615_n8171# a_24054_n7805# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X969 VSS.t375 VDD VSS.t374 VSS.t373 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X970 x3.x2.GP2.t0 x3.x2.GN2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.225151 ps=2.058971 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X971 VSS.t372 VDD VSS.t371 VSS.t370 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
**devattr d=5720,324
X972 VSS.t40 a_23675_n5233# a_23682_n5329# VSS.t39 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X973 VSS.t369 VDD VSS.t368 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X974 a_24595_n9571# x4._11_.t19 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X975 a_25211_n9231# x4._11_.t20 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X976 a_23927_n8715# a_23063_n8709# a_23670_n8741# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X977 VDD VSS.t1073 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.05
**devattr d=9048,452
X978 a_23597_n8715# a_23063_n8709# a_23502_n8715# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X979 VSS.t366 VDD VSS.t365 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X980 a_24229_n4907# a_23682_n4633# a_23882_n4933# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=2310,139
X981 a_23421_n7921# x4._11_.t21 x4._13_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X982 x4.clknet_1_1__leaf_clk.t16 a_27194_n8171# VSS.t263 VSS.t262 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X983 VSS.t222 x1.sky130_fd_sc_hd__inv_2_9.A x1.sky130_fd_sc_hd__nand2_2_0.B VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X984 a_22962_n5131# x4.net1 VSS.t253 VSS.t252 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0 ps=0 w=0.65 l=0.15
**devattr s=6890,366 d=3835,189
X985 a_23633_n5451# a_23295_n5219# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=4452,274 d=3528,168
X986 VDD a_25709_n7109# x4.clknet_0_clk.t0 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0 ps=0 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X987 VSS.t361 VDD VSS.t360 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X988 VDD VSS.t1074 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=0.59
**devattr d=9048,452
X989 a_23811_n5073# a_23682_n5329# a_23391_n5219# VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.071208 pd=0.7164 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=3956,199
X990 VDD a_26979_n9829# x4._22_ VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225151 pd=2.058971 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=12498,336
X991 VDD VSS.t1075 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195882 pd=1.791305 as=0.195882 ps=1.791305 w=0.87 l=1.97
**devattr d=9048,452
X992 VDD x4.net7 a_26147_n9107# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.094564 pd=0.864768 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=2268,138
X993 a_23615_n5995# x4.net3.t7 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0.094564 ps=0.864768 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
R0 VSS.n2759 VSS.n2754 3.3176e+06
R1 VSS.n2759 VSS.n2758 2.3386e+06
R2 VSS.n2758 VSS.n2757 2.1446e+06
R3 VSS.n2758 VSS.t240 1.17707e+06
R4 VSS.n2767 VSS.n2754 396385
R5 VSS.n2754 VSS.n2753 391216
R6 VSS.n2865 VSS.n5 53736.2
R7 VSS.n2856 VSS.n64 38301.6
R8 VSS.n2691 VSS.n3 35421.6
R9 VSS.n2858 VSS.n2856 29605.7
R10 VSS.n2683 VSS 23608
R11 VSS.n2683 VSS.n3 15966.1
R12 VSS.t906 VSS.n2683 13977.5
R13 VSS.n2756 VSS.n2728 11744.7
R14 VSS.n2781 VSS.n2728 11744.7
R15 VSS.n2756 VSS.n2729 11744.7
R16 VSS.n2781 VSS.n2729 11744.7
R17 VSS.n2752 VSS.n2740 11744.7
R18 VSS.n2746 VSS.n2740 11744.7
R19 VSS.n2752 VSS.n2741 11744.7
R20 VSS.n2746 VSS.n2741 11744.7
R21 VSS.n2768 VSS.n2738 11744.7
R22 VSS.n2764 VSS.n2738 11744.7
R23 VSS.n2768 VSS.n2739 11744.7
R24 VSS.n2764 VSS.n2739 11744.7
R25 VSS.n2790 VSS.n2722 11744.7
R26 VSS.n2790 VSS.n2723 11744.7
R27 VSS.n2785 VSS.n2722 11744.7
R28 VSS.n2785 VSS.n2723 11744.7
R29 VSS.n2761 VSS.n2760 10248.5
R30 VSS.n2859 VSS.n2858 9243.96
R31 VSS.n2868 VSS.n2867 8555.7
R32 VSS.n1929 VSS 8554.54
R33 VSS.n2867 VSS.n3 8490.24
R34 VSS.n2499 VSS 8079.51
R35 VSS.n2499 VSS.n267 7881.01
R36 VSS.n1333 VSS.n267 7881.01
R37 VSS.n1334 VSS.n1333 7881.01
R38 VSS.n1334 VSS.n1030 7881.01
R39 VSS.n1929 VSS.n1030 7881.01
R40 VSS.n2767 VSS.t239 7088.89
R41 VSS.t238 VSS.n2765 7088.89
R42 VSS.n2753 VSS.t735 6925.66
R43 VSS.n2745 VSS.t730 6925.66
R44 VSS.n2757 VSS.t746 6925.66
R45 VSS.n2782 VSS.t749 6925.66
R46 VSS.t239 VSS.n2766 6733.33
R47 VSS.n2766 VSS.t238 6733.33
R48 VSS.n2744 VSS.t735 6578.29
R49 VSS.t730 VSS.n2744 6578.29
R50 VSS.t746 VSS.n2755 6578.29
R51 VSS.n2755 VSS.t749 6578.29
R52 VSS.n2684 VSS.n119 5434.88
R53 VSS.n2689 VSS.n119 5434.88
R54 VSS.n2689 VSS.n120 5434.88
R55 VSS.n2684 VSS.n120 5434.88
R56 VSS.n2784 VSS.n2783 5125.3
R57 VSS VSS.t446 4888.89
R58 VSS.n2761 VSS.n2727 4823.17
R59 VSS.n2783 VSS.n2727 4705.56
R60 VSS.n2765 VSS.n2761 4474.07
R61 VSS.t446 VSS 4408.43
R62 VSS.n2783 VSS.n2782 4363.82
R63 VSS.n2745 VSS.n2727 4320.4
R64 VSS.n2867 VSS.n2866 4049.09
R65 VSS.t443 VSS.t648 3877.39
R66 VSS.t651 VSS.t561 3877.39
R67 VSS.n118 VSS.n116 3464.88
R68 VSS.n2694 VSS.n116 3464.88
R69 VSS.n2693 VSS.n118 3464.88
R70 VSS.n2694 VSS.n2693 3464.88
R71 VSS.t595 VSS 3346.36
R72 VSS VSS.t530 3346.36
R73 VSS VSS.t499 3346.36
R74 VSS VSS.t400 3346.36
R75 VSS.t379 VSS 3346.36
R76 VSS VSS.t428 3346.36
R77 VSS VSS.t642 3346.36
R78 VSS.t440 VSS.t425 3101.92
R79 VSS.t657 VSS.t584 3101.92
R80 VSS.t533 VSS.t512 3101.92
R81 VSS VSS.t547 2857.47
R82 VSS.t587 VSS 2857.47
R83 VSS.t416 VSS 2857.47
R84 VSS.t660 VSS 2857.47
R85 VSS.t437 VSS 2857.47
R86 VSS.t573 VSS 2857.47
R87 VSS.t693 VSS.t567 2495.02
R88 VSS VSS.n523 2469.73
R89 VSS VSS.t550 2452.87
R90 VSS VSS.t536 2452.87
R91 VSS.t367 VSS.t558 2326.44
R92 VSS.t422 VSS.t555 2326.44
R93 VSS.t463 VSS.t639 2326.44
R94 VSS VSS.n267 2183.14
R95 VSS.n1333 VSS 2183.14
R96 VSS VSS.n1334 2183.14
R97 VSS VSS.n1030 2183.14
R98 VSS VSS.n1929 2183.14
R99 VSS VSS.n2499 2183.14
R100 VSS VSS.t515 2081.99
R101 VSS.t483 VSS 2081.99
R102 VSS.n594 VSS.t370 1938.7
R103 VSS.t515 VSS 1812.26
R104 VSS.t425 VSS 1795.4
R105 VSS VSS.t657 1795.4
R106 VSS VSS.t466 1795.4
R107 VSS.t512 VSS 1795.4
R108 VSS VSS.t419 1786.97
R109 VSS.t518 VSS 1786.97
R110 VSS VSS.t579 1786.97
R111 VSS VSS.t406 1702.68
R112 VSS.n1336 VSS 1677.39
R113 VSS.t2 VSS.t131 1593.1
R114 VSS.t53 VSS.t902 1593.1
R115 VSS.t180 VSS.t342 1593.1
R116 VSS.t39 VSS.t63 1584.67
R117 VSS.t230 VSS.t346 1584.67
R118 VSS.t454 VSS.t147 1567.82
R119 VSS.t615 VSS.t595 1550.96
R120 VSS.t530 VSS.t457 1550.96
R121 VSS.t499 VSS.t587 1550.96
R122 VSS.t400 VSS.t416 1550.96
R123 VSS.t419 VSS.t660 1550.96
R124 VSS.t397 VSS.t379 1550.96
R125 VSS.t428 VSS.t437 1550.96
R126 VSS.t642 VSS.t573 1550.96
R127 VSS.t348 VSS.t256 1550.96
R128 VSS VSS.t576 1502.01
R129 VSS.t129 VSS.t773 1416.09
R130 VSS VSS.t564 1407.66
R131 VSS VSS.t460 1407.66
R132 VSS VSS.t359 1407.66
R133 VSS VSS.t155 1407.66
R134 VSS VSS.t373 1407.66
R135 VSS VSS.t477 1407.66
R136 VSS VSS.t391 1399.23
R137 VSS.t866 VSS.t965 1399.23
R138 VSS.t0 VSS 1390.8
R139 VSS VSS.t615 1306.51
R140 VSS VSS.t440 1306.51
R141 VSS.t370 VSS 1306.51
R142 VSS.t521 VSS 1306.51
R143 VSS.t457 VSS 1306.51
R144 VSS.t584 VSS 1306.51
R145 VSS.t376 VSS 1306.51
R146 VSS.t527 VSS 1306.51
R147 VSS.t567 VSS 1306.51
R148 VSS VSS.t610 1306.51
R149 VSS VSS.t518 1306.51
R150 VSS VSS.t397 1306.51
R151 VSS VSS.t533 1306.51
R152 VSS.t542 VSS 1306.51
R153 VSS.t579 VSS 1306.51
R154 VSS.n2634 VSS.n2579 1294.86
R155 VSS VSS.t940 1289.66
R156 VSS.t800 VSS 1272.8
R157 VSS.n2682 VSS.n2681 1198.25
R158 VSS.n1928 VSS.n1927 1198.25
R159 VSS.n1335 VSS.n866 1198.25
R160 VSS.n1930 VSS.n984 1198.25
R161 VSS.n1872 VSS.n1073 1198.25
R162 VSS.n2805 VSS.n2792 1198.25
R163 VSS.n65 VSS.n6 1198.25
R164 VSS.n2864 VSS.n2863 1198.25
R165 VSS.n2845 VSS.n70 1198.25
R166 VSS.n2498 VSS.n2497 1198.25
R167 VSS.n595 VSS.n594 1196.22
R168 VSS.n2359 VSS.n523 1196.22
R169 VSS.n1497 VSS.n1486 1194.5
R170 VSS.n1332 VSS.n1331 1194.5
R171 VSS.n2310 VSS.n549 1194.5
R172 VSS.n1337 VSS.n1336 1194.5
R173 VSS.n1559 VSS.n1443 1194.5
R174 VSS.n1932 VSS.n1931 1194.5
R175 VSS.n2565 VSS.n226 1194.5
R176 VSS.n2501 VSS.n2500 1194.5
R177 VSS.n2855 VSS.n2854 1194.5
R178 VSS.t814 VSS.t938 1188.51
R179 VSS.n2830 VSS.n96 1171.32
R180 VSS.n1931 VSS.t724 1146.36
R181 VSS VSS.t348 1137.93
R182 VSS.n64 VSS.n2 1105.32
R183 VSS.t55 VSS 1104.21
R184 VSS VSS.t157 1078.93
R185 VSS.t858 VSS.t57 1078.93
R186 VSS.t147 VSS.t59 1078.93
R187 VSS.n1073 VSS.t388 1076.6
R188 VSS VSS.t896 1070.5
R189 VSS VSS.t309 1036.78
R190 VSS.t965 VSS 1036.78
R191 VSS.t547 VSS 1019.92
R192 VSS.t648 VSS 1019.92
R193 VSS.t561 VSS 1019.92
R194 VSS VSS.t527 1019.92
R195 VSS.t24 VSS.t794 1003.07
R196 VSS.t161 VSS 1003.07
R197 VSS.t228 VSS.t198 1003.07
R198 VSS.n501 VSS.n500 999.607
R199 VSS.n1233 VSS.n1232 999.607
R200 VSS.n2460 VSS.n2398 999.607
R201 VSS.t111 VSS.t232 960.92
R202 VSS.t877 VSS.t151 952.49
R203 VSS.t63 VSS.t41 944.062
R204 VSS.t61 VSS.t174 944.062
R205 VSS.t117 VSS.t849 944.062
R206 VSS.n1332 VSS 927.203
R207 VSS.n2500 VSS 927.203
R208 VSS VSS.t367 918.774
R209 VSS.t391 VSS 918.774
R210 VSS.t555 VSS 918.774
R211 VSS.n549 VSS 918.774
R212 VSS.t564 VSS 918.774
R213 VSS.t460 VSS 918.774
R214 VSS.t359 VSS 918.774
R215 VSS.t630 VSS 918.774
R216 VSS.t373 VSS 918.774
R217 VSS.n2857 VSS 918.774
R218 VSS.n2855 VSS 918.774
R219 VSS.t712 VSS 918.774
R220 VSS VSS.t463 918.774
R221 VSS.n226 VSS 918.774
R222 VSS.t477 VSS 918.774
R223 VSS.t155 VSS.t830 910.346
R224 VSS.n1335 VSS 901.917
R225 VSS.n1930 VSS 901.917
R226 VSS.t36 VSS.t42 893.487
R227 VSS.t52 VSS.t737 893.487
R228 VSS.t388 VSS 881.561
R229 VSS.n2208 VSS.n2207 870.4
R230 VSS.t794 VSS.t36 851.341
R231 VSS.t80 VSS.t14 851.341
R232 VSS.t146 VSS 851.341
R233 VSS.t166 VSS.t936 842.913
R234 VSS.n1928 VSS.t645 837.352
R235 VSS.t41 VSS.t37 834.484
R236 VSS.t37 VSS.t24 834.484
R237 VSS.t169 VSS.t205 834.484
R238 VSS.t311 VSS.t864 834.484
R239 VSS.t738 VSS.t736 834.484
R240 VSS.t79 VSS.t159 834.484
R241 VSS.t43 VSS.t68 834.484
R242 VSS.t321 VSS.t230 826.054
R243 VSS.t218 VSS.t598 826.054
R244 VSS.t259 VSS.t228 826.054
R245 VSS.t201 VSS.t121 826.054
R246 VSS.t959 VSS.t673 826.054
R247 VSS.t740 VSS.t866 809.196
R248 VSS.t327 VSS.t800 809.196
R249 VSS.t42 VSS.t2 800.766
R250 VSS.t190 VSS.t307 800.766
R251 VSS.t901 VSS.t53 800.766
R252 VSS.t175 VSS.t242 800.766
R253 VSS.t592 VSS.t188 792.337
R254 VSS.t816 VSS.t394 792.337
R255 VSS.t758 VSS.t767 792.337
R256 VSS VSS.t633 790.544
R257 VSS.t663 VSS 790.544
R258 VSS VSS.t670 790.544
R259 VSS.t83 VSS.t178 783.909
R260 VSS.t466 VSS.t483 775.48
R261 VSS.n2780 VSS.n2779 763.09
R262 VSS.n2748 VSS.n2747 763.09
R263 VSS.n2763 VSS.n2762 763.09
R264 VSS.n2787 VSS.n2786 763.09
R265 VSS.t598 VSS.t914 758.621
R266 VSS.t718 VSS.t179 758.621
R267 VSS.t846 VSS.t252 750.192
R268 VSS.t346 VSS.t851 741.763
R269 VSS.t221 VSS.t816 741.763
R270 VSS.t278 VSS.t894 741.763
R271 VSS.t743 VSS.t298 741.763
R272 VSS.n2779 VSS.n2778 732.236
R273 VSS.n2750 VSS.n2748 732.236
R274 VSS.n2762 VSS.n2736 732.236
R275 VSS.n2788 VSS.n2787 732.236
R276 VSS.t34 VSS.t846 724.904
R277 VSS.t887 VSS.t879 724.904
R278 VSS.t89 VSS.t99 724.904
R279 VSS.t93 VSS.t105 724.904
R280 VSS.t101 VSS.t113 724.904
R281 VSS.t113 VSS.t95 724.904
R282 VSS.t908 VSS.t885 724.904
R283 VSS.t885 VSS.t910 724.904
R284 VSS.t910 VSS.t808 724.904
R285 VSS.t808 VSS.t689 724.904
R286 VSS.t689 VSS.t701 724.904
R287 VSS.t685 VSS.t697 724.904
R288 VSS.t697 VSS.t681 724.904
R289 VSS.t681 VSS.t691 724.904
R290 VSS.t691 VSS.t705 724.904
R291 VSS.t705 VSS.t679 724.904
R292 VSS.t703 VSS.t687 724.904
R293 VSS.t687 VSS.t699 724.904
R294 VSS.t699 VSS.t677 724.904
R295 VSS.t677 VSS.t695 724.904
R296 VSS.t695 VSS.t675 724.904
R297 VSS.t675 VSS.t683 724.904
R298 VSS.t268 VSS.t288 724.904
R299 VSS.t264 VSS.t284 724.904
R300 VSS.t290 VSS.t276 724.904
R301 VSS.t840 VSS.t143 724.904
R302 VSS.t883 VSS.t840 724.904
R303 VSS.t726 VSS.t950 724.904
R304 VSS.t45 VSS.t889 716.476
R305 VSS.t272 VSS.t494 716.476
R306 VSS.t778 VSS.t814 716.476
R307 VSS.t912 VSS.t825 716.476
R308 VSS.t246 VSS.t39 708.047
R309 VSS.t131 VSS.t0 708.047
R310 VSS.t896 VSS.t210 708.047
R311 VSS.t188 VSS.t190 708.047
R312 VSS.t936 VSS.t16 708.047
R313 VSS.t716 VSS.t141 708.047
R314 VSS.t160 VSS.t806 708.047
R315 VSS.t765 VSS.t335 708.047
R316 VSS.t157 VSS.t934 708.047
R317 VSS.t81 VSS.t329 708.047
R318 VSS.t127 VSS.t125 708.047
R319 VSS.t708 VSS.t176 708.047
R320 VSS.t65 VSS.t875 708.047
R321 VSS.t830 VSS.t146 708.047
R322 VSS.t119 VSS.t4 708.047
R323 VSS.n2858 VSS.n2857 708.047
R324 VSS.t8 VSS.t10 708.047
R325 VSS.t317 VSS.t319 708.047
R326 VSS.t313 VSS.t315 708.047
R327 VSS.t32 VSS.t30 708.047
R328 VSS.t788 VSS.t786 708.047
R329 VSS.t303 VSS.t305 708.047
R330 VSS.t26 VSS.t28 708.047
R331 VSS.t194 VSS.t196 708.047
R332 VSS.t752 VSS.t750 708.047
R333 VSS.n2869 VSS.n2868 708.047
R334 VSS.n2856 VSS.n2855 708.047
R335 VSS.t362 VSS.t504 708.047
R336 VSS.t767 VSS.t925 708.047
R337 VSS.t720 VSS.t722 708.047
R338 VSS.t334 VSS.t927 708.047
R339 VSS.t256 VSS.t842 708.047
R340 VSS.t842 VSS.t917 708.047
R341 VSS.t917 VSS.t257 708.047
R342 VSS.t109 VSS.t791 699.617
R343 VSS.t802 VSS.t111 691.188
R344 VSS.t449 VSS.t55 691.188
R345 VSS.t810 VSS.t942 691.188
R346 VSS.t847 VSS 682.76
R347 VSS.n96 VSS.t524 681.482
R348 VSS.t182 VSS.t107 674.331
R349 VSS.t276 VSS 674.331
R350 VSS.t756 VSS.t352 674.331
R351 VSS.t869 VSS.t726 674.331
R352 VSS.t775 VSS.t321 657.471
R353 VSS.t149 VSS.t218 657.471
R354 VSS.t737 VSS.t170 657.471
R355 VSS.t953 VSS.t930 657.471
R356 VSS VSS.t474 649.043
R357 VSS.t633 VSS 642.317
R358 VSS VSS.t645 642.317
R359 VSS VSS.t663 642.317
R360 VSS.t670 VSS 642.317
R361 VSS.t153 VSS.t871 640.614
R362 VSS.t294 VSS.t877 640.614
R363 VSS.t558 VSS 632.184
R364 VSS.n523 VSS 632.184
R365 VSS.n594 VSS 632.184
R366 VSS VSS.t422 632.184
R367 VSS VSS.n1332 632.184
R368 VSS VSS.n549 632.184
R369 VSS.t406 VSS 632.184
R370 VSS.n1336 VSS 632.184
R371 VSS.t85 VSS.t804 632.184
R372 VSS VSS.n1335 632.184
R373 VSS.t550 VSS 632.184
R374 VSS.t944 VSS.t266 632.184
R375 VSS.n1486 VSS 632.184
R376 VSS.t536 VSS 632.184
R377 VSS VSS.n1930 632.184
R378 VSS.n2869 VSS 632.184
R379 VSS.t639 VSS 632.184
R380 VSS.n2500 VSS 632.184
R381 VSS VSS.n226 632.184
R382 VSS.t284 VSS.t344 623.755
R383 VSS.n2784 VSS.t358 620.971
R384 VSS.t280 VSS.t250 615.327
R385 VSS.t266 VSS.n1443 615.327
R386 VSS.t212 VSS.t270 615.327
R387 VSS.t853 VSS.t337 615.327
R388 VSS.t254 VSS.t878 606.898
R389 VSS.t878 VSS.t916 606.898
R390 VSS.t636 VSS.t693 606.898
R391 VSS.t898 VSS.t274 606.898
R392 VSS.t790 VSS.t812 606.898
R393 VSS.t812 VSS.t858 606.898
R394 VSS.t59 VSS.t863 606.898
R395 VSS.t863 VSS.t145 606.898
R396 VSS.t741 VSS.t340 606.898
R397 VSS.t206 VSS.t385 603.311
R398 VSS.n2857 VSS.n63 599.125
R399 VSS.n2870 VSS.n2869 599.125
R400 VSS.t72 VSS.t89 598.467
R401 VSS.t151 VSS.t214 598.467
R402 VSS.t868 VSS.t891 598.467
R403 VSS.t184 VSS.t855 598.467
R404 VSS.t834 VSS.t118 598.467
R405 VSS.t97 VSS.t822 590.038
R406 VSS VSS.t775 581.61
R407 VSS.t873 VSS.t115 581.61
R408 VSS.t329 VSS 581.61
R409 VSS.t165 VSS.t244 573.181
R410 VSS.n2683 VSS 564.751
R411 VSS VSS.t254 564.751
R412 VSS.n2683 VSS 564.751
R413 VSS.n2683 VSS 564.751
R414 VSS.t172 VSS.t51 564.751
R415 VSS.n2683 VSS 564.751
R416 VSS VSS.t764 564.751
R417 VSS.n2683 VSS 564.751
R418 VSS.t10 VSS 564.751
R419 VSS.t319 VSS 564.751
R420 VSS.t315 VSS 564.751
R421 VSS.t30 VSS 564.751
R422 VSS.t786 VSS 564.751
R423 VSS.t305 VSS 564.751
R424 VSS.t28 VSS 564.751
R425 VSS.t196 VSS 564.751
R426 VSS.t750 VSS 564.751
R427 VSS.t504 VSS 564.751
R428 VSS.t722 VSS 564.751
R429 VSS VSS.t334 564.751
R430 VSS VSS.n64 564.751
R431 VSS.n2683 VSS 564.751
R432 VSS VSS.t654 559.102
R433 VSS.t307 VSS 556.322
R434 VSS.t103 VSS.t74 556.322
R435 VSS.t44 VSS.t813 556.322
R436 VSS.t627 VSS 551.301
R437 VSS.t916 VSS 547.894
R438 VSS VSS.t161 547.894
R439 VSS VSS.t221 547.894
R440 VSS.t914 VSS 547.894
R441 VSS.t714 VSS.t248 547.894
R442 VSS VSS.t311 547.894
R443 VSS.t14 VSS.t49 547.894
R444 VSS.t145 VSS 547.894
R445 VSS.t210 VSS 539.465
R446 VSS.t480 VSS 539.465
R447 VSS VSS.t443 531.034
R448 VSS VSS.t651 531.034
R449 VSS VSS.t539 531.034
R450 VSS.t604 VSS 531.034
R451 VSS.t469 VSS 527.896
R452 VSS.t232 VSS 522.606
R453 VSS.t286 VSS 522.606
R454 VSS.t927 VSS.t607 522.606
R455 VSS.t309 VSS 514.177
R456 VSS.t139 VSS.t350 514.177
R457 VSS VSS.t61 514.177
R458 VSS.t205 VSS.t952 505.748
R459 VSS.t216 VSS 505.748
R460 VSS.t506 VSS.t685 497.318
R461 VSS.t893 VSS.t292 497.318
R462 VSS VSS.t741 497.318
R463 VSS.t364 VSS.t208 495.106
R464 VSS.t350 VSS.t738 488.889
R465 VSS.t301 VSS.t961 488.889
R466 VSS.t87 VSS.t71 480.461
R467 VSS.t282 VSS.t899 480.461
R468 VSS VSS.t166 480.461
R469 VSS.t728 VSS 480.461
R470 VSS.t793 VSS 480.461
R471 VSS.t889 VSS 463.603
R472 VSS.t133 VSS.t87 463.603
R473 VSS.t186 VSS.t91 463.603
R474 VSS.t524 VSS 459.26
R475 VSS.t948 VSS.t714 455.173
R476 VSS.t49 VSS.t955 455.173
R477 VSS VSS.t175 455.173
R478 VSS.t174 VSS.t296 455.173
R479 VSS VSS.t901 446.743
R480 VSS.t894 VSS 446.743
R481 VSS.t204 VSS 446.743
R482 VSS VSS.t163 446.743
R483 VSS.n1931 VSS.t728 446.743
R484 VSS.t67 VSS 446.743
R485 VSS VSS.t618 445.288
R486 VSS VSS.t509 445.288
R487 VSS VSS.t411 445.288
R488 VSS.t938 VSS 438.315
R489 VSS VSS.t703 429.885
R490 VSS.t929 VSS.t895 429.885
R491 VSS.t18 VSS.t43 429.885
R492 VSS.t22 VSS 410.875
R493 VSS VSS.t819 410.875
R494 VSS VSS.t796 410.875
R495 VSS.t946 VSS 410.875
R496 VSS.t828 VSS 410.875
R497 VSS VSS.t710 404.599
R498 VSS.t47 VSS 404.599
R499 VSS.t934 VSS 404.599
R500 VSS.t798 VSS.t868 404.599
R501 VSS.t895 VSS.t798 404.599
R502 VSS.t855 VSS.t69 404.599
R503 VSS.t69 VSS.t18 404.599
R504 VSS.t875 VSS 404.599
R505 VSS.t923 VSS.t180 404.599
R506 VSS.t4 VSS 404.599
R507 VSS.t654 VSS 403.074
R508 VSS VSS.t627 403.074
R509 VSS.t618 VSS 400.837
R510 VSS.t509 VSS 400.837
R511 VSS.t411 VSS 400.837
R512 VSS VSS.t364 400.837
R513 VSS.t91 VSS.t821 387.74
R514 VSS.t784 VSS.t280 387.74
R515 VSS.t607 VSS.t712 387.74
R516 VSS.t296 VSS.t929 379.31
R517 VSS.t950 VSS 379.31
R518 VSS.t849 VSS.t630 370.882
R519 VSS VSS.t733 370.37
R520 VSS VSS.t356 370.37
R521 VSS.t771 VSS.n1928 364.067
R522 VSS.n1073 VSS.t325 364.067
R523 VSS.n2685 VSS.n121 353.13
R524 VSS.n2688 VSS.n121 353.13
R525 VSS.n2051 VSS.n969 352
R526 VSS.t821 VSS.t103 337.166
R527 VSS.t292 VSS.t784 337.166
R528 VSS VSS.t204 337.166
R529 VSS.n70 VSS.t823 337.166
R530 VSS.n2792 VSS.n2791 334.815
R531 VSS.n2688 VSS.n2687 330.486
R532 VSS.t952 VSS.t948 328.736
R533 VSS VSS.t716 328.736
R534 VSS.t163 VSS 328.736
R535 VSS.n2686 VSS.n2685 324.425
R536 VSS VSS.t67 320.307
R537 VSS.n70 VSS.t201 320.307
R538 VSS VSS.t65 311.877
R539 VSS.t382 VSS 305.8
R540 VSS.n2780 VSS.n2730 304.553
R541 VSS.n2747 VSS.n2743 304.553
R542 VSS.n2763 VSS.n2737 304.553
R543 VSS.n2786 VSS.n2726 304.553
R544 VSS VSS.t486 304.269
R545 VSS VSS.t149 303.449
R546 VSS VSS.t168 303.449
R547 VSS.t340 VSS.t923 303.449
R548 VSS.n2868 VSS.t358 303.42
R549 VSS.t813 VSS.t184 295.019
R550 VSS VSS.t119 295.019
R551 VSS.t823 VSS 295.019
R552 VSS.n2693 VSS.n114 292.5
R553 VSS.n2693 VSS.t6 292.5
R554 VSS.n116 VSS.n115 292.5
R555 VSS.t6 VSS.n116 292.5
R556 VSS VSS.t34 286.591
R557 VSS.t679 VSS 286.591
R558 VSS VSS.t862 286.591
R559 VSS.t385 VSS 283.452
R560 VSS.n2866 VSS.n4 281.377
R561 VSS.n722 VSS.t35 281.25
R562 VSS VSS.t8 278.161
R563 VSS VSS.t317 278.161
R564 VSS VSS.t313 278.161
R565 VSS VSS.t32 278.161
R566 VSS VSS.t788 278.161
R567 VSS VSS.t303 278.161
R568 VSS VSS.t26 278.161
R569 VSS VSS.t194 278.161
R570 VSS VSS.t752 278.161
R571 VSS.n472 VSS.t971 276.531
R572 VSS.n1202 VSS.t968 276.531
R573 VSS.n2409 VSS.t1047 276.531
R574 VSS.n1496 VSS.t717 275.293
R575 VSS.n1647 VSS.t164 275.293
R576 VSS.n2594 VSS.t258 275.293
R577 VSS VSS.t908 269.733
R578 VSS.t352 VSS.t169 269.733
R579 VSS.t736 VSS.t172 269.733
R580 VSS.n2361 VSS.t1025 269.488
R581 VSS.n681 VSS.t1051 269.445
R582 VSS.n2776 VSS.n2730 266.349
R583 VSS.n2743 VSS.n2742 266.349
R584 VSS.n2770 VSS.n2737 266.349
R585 VSS.n2726 VSS.n2724 266.349
R586 VSS.n2275 VSS.t1023 265.317
R587 VSS.n2611 VSS.t974 265.317
R588 VSS.n1188 VSS.t1024 265.298
R589 VSS.n265 VSS.t997 265.298
R590 VSS.n476 VSS.t981 262.784
R591 VSS.n477 VSS.t978 262.784
R592 VSS.n727 VSS.t1037 262.784
R593 VSS.n729 VSS.t1032 262.784
R594 VSS.n479 VSS.t1041 262.784
R595 VSS.n499 VSS.t1038 262.784
R596 VSS.n810 VSS.t1034 262.784
R597 VSS.n812 VSS.t1031 262.784
R598 VSS.n1206 VSS.t979 262.784
R599 VSS.n1207 VSS.t977 262.784
R600 VSS.n1209 VSS.t1040 262.784
R601 VSS.n1231 VSS.t1035 262.784
R602 VSS.n1138 VSS.t1006 262.784
R603 VSS.n1386 VSS.t1003 262.784
R604 VSS.n2262 VSS.t1069 262.784
R605 VSS.n2263 VSS.t1064 262.784
R606 VSS.n1400 VSS.t1065 262.784
R607 VSS.n1402 VSS.t1033 262.784
R608 VSS.n948 VSS.t1014 262.784
R609 VSS.n949 VSS.t989 262.784
R610 VSS.n1125 VSS.t990 262.784
R611 VSS.n1128 VSS.t1067 262.784
R612 VSS.n2060 VSS.t1049 262.784
R613 VSS.n2061 VSS.t1017 262.784
R614 VSS.n2399 VSS.t1057 262.784
R615 VSS.n2468 VSS.t1055 262.784
R616 VSS.n2598 VSS.t1005 262.784
R617 VSS.n2599 VSS.t1002 262.784
R618 VSS.n2396 VSS.t1009 262.784
R619 VSS.n2397 VSS.t1007 262.784
R620 VSS.n186 VSS.t1046 262.719
R621 VSS.n361 VSS.t1028 262.719
R622 VSS.n395 VSS.t996 262.719
R623 VSS.n609 VSS.t1062 262.719
R624 VSS.n606 VSS.t1013 262.719
R625 VSS.n598 VSS.t991 262.719
R626 VSS.n519 VSS.t1021 262.719
R627 VSS.n808 VSS.t995 262.719
R628 VSS.n785 VSS.t1043 262.719
R629 VSS.n1267 VSS.t1020 262.719
R630 VSS.n1307 VSS.t1061 262.719
R631 VSS.n1296 VSS.t1048 262.719
R632 VSS.n546 VSS.t988 262.719
R633 VSS.n2315 VSS.t998 262.719
R634 VSS.n2234 VSS.t969 262.719
R635 VSS.n1362 VSS.t1058 262.719
R636 VSS.n1177 VSS.t985 262.719
R637 VSS.n1971 VSS.t987 262.719
R638 VSS.n246 VSS.t1029 262.719
R639 VSS.n2530 VSS.t1015 262.719
R640 VSS.n229 VSS.t1066 262.719
R641 VSS.n2560 VSS.t972 262.719
R642 VSS.n2641 VSS.t1012 262.719
R643 VSS.n2641 VSS.t1018 262.719
R644 VSS.n2424 VSS.t993 262.719
R645 VSS.n272 VSS.t1071 262.719
R646 VSS VSS.t246 261.303
R647 VSS VSS.t234 261.303
R648 VSS.t99 VSS.t133 261.303
R649 VSS.t610 VSS 261.303
R650 VSS.t248 VSS.t760 261.303
R651 VSS.t539 VSS 261.303
R652 VSS.t125 VSS 261.303
R653 VSS.t836 VSS 261.303
R654 VSS.t298 VSS 261.303
R655 VSS VSS.t824 261.303
R656 VSS VSS.t790 261.303
R657 VSS VSS.t758 261.303
R658 VSS.t486 VSS 259.815
R659 VSS VSS.t382 259.815
R660 VSS.n191 VSS.t976 259.082
R661 VSS.n327 VSS.t1074 259.082
R662 VSS.n1706 VSS.t1019 259.082
R663 VSS.n1562 VSS.t975 259.082
R664 VSS.n2003 VSS.t1011 259.082
R665 VSS.n2045 VSS.t1030 259.082
R666 VSS.n1812 VSS.t1053 259.082
R667 VSS.n451 VSS.t980 259.082
R668 VSS.n303 VSS.t1022 259.082
R669 VSS VSS.t592 252.875
R670 VSS.t105 VSS.t186 252.875
R671 VSS.t760 VSS 252.875
R672 VSS.t955 VSS.t47 252.875
R673 VSS VSS.t81 252.875
R674 VSS.n719 VSS.t3 251
R675 VSS.n719 VSS.t782 251
R676 VSS.n1490 VSS.t152 251
R677 VSS.n2108 VSS.t173 251
R678 VSS.n1657 VSS.t243 251
R679 VSS.n2026 VSS.t343 251
R680 VSS.n2868 VSS.n2 249.105
R681 VSS.t733 VSS.t731 248.889
R682 VSS.t744 VSS.t747 248.889
R683 VSS.t356 VSS.t354 248.889
R684 VSS.n2167 VSS.t805 245.82
R685 VSS.n1602 VSS.t54 245.82
R686 VSS.n1461 VSS.t943 245.82
R687 VSS.n1029 VSS.t729 245.82
R688 VSS VSS.t376 244.445
R689 VSS.t491 VSS 244.445
R690 VSS.t71 VSS.t97 244.445
R691 VSS VSS.t480 244.445
R692 VSS.t434 VSS 244.445
R693 VSS VSS.t542 244.445
R694 VSS.n706 VSS.t707 243.028
R695 VSS.n706 VSS.t64 243.028
R696 VSS.n1529 VSS.t757 243.028
R697 VSS.n2103 VSS.t807 243.028
R698 VSS.n1093 VSS.t62 243.028
R699 VSS.n1011 VSS.t801 243.028
R700 VSS.n869 VSS.t112 242.067
R701 VSS.n1418 VSS.t279 242.067
R702 VSS.n893 VSS.t888 240.948
R703 VSS.n1540 VSS.t811 240.948
R704 VSS.n74 VSS.t759 240.575
R705 VSS.n2152 VSS.t134 238.675
R706 VSS.n1576 VSS.t345 238.675
R707 VSS.n940 VSS.t217 238.675
R708 VSS.n2046 VSS.t850 238.675
R709 VSS.n2866 VSS.t38 238.468
R710 VSS.n2258 VSS.t694 238.44
R711 VSS.n2200 VSS.t915 237.327
R712 VSS.n1171 VSS.t162 237.327
R713 VSS.n68 VSS.t941 237.327
R714 VSS.t899 VSS.t264 236.016
R715 VSS VSS.t754 236.016
R716 VSS.t51 VSS.t160 236.016
R717 VSS.n784 VSS.t189 235.607
R718 VSS.n1957 VSS.n1010 234.667
R719 VSS.n1522 VSS.t815 230.977
R720 VSS.n1666 VSS.t297 230.977
R721 VSS.n735 VSS.t253 229.833
R722 VSS.t299 VSS.t301 228.843
R723 VSS.t961 VSS.t123 228.843
R724 VSS.t20 VSS.t22 228.843
R725 VSS.t856 VSS.t771 228.843
R726 VSS.t819 VSS.t817 228.843
R727 VSS.t796 VSS.t826 228.843
R728 VSS.t325 VSS.t832 228.843
R729 VSS.t762 VSS.t946 228.843
R730 VSS.t776 VSS.t828 228.843
R731 VSS.t844 VSS.t206 228.843
R732 VSS.n1474 VSS.n1473 228.294
R733 VSS.n2037 VSS.n2036 228.294
R734 VSS.t701 VSS.t506 227.587
R735 VSS.t274 VSS.t893 227.587
R736 VSS.t710 VSS.t282 227.587
R737 VSS.t838 VSS 227.587
R738 VSS.n527 VSS.t649 227.256
R739 VSS.n2208 VSS.t909 226.708
R740 VSS.n2695 VSS.n115 225.13
R741 VSS.n117 VSS.n115 225.13
R742 VSS.n1613 VSS.t1039 224.196
R743 VSS.n1279 VSS.t1010 224.102
R744 VSS.n251 VSS.t986 224.102
R745 VSS.n550 VSS.t418 223.282
R746 VSS.n2187 VSS.n2186 222.691
R747 VSS.n2792 VSS 222.222
R748 VSS VSS.n96 222.222
R749 VSS.n551 VSS.t1052 221.972
R750 VSS.n1489 VSS.n1487 221.804
R751 VSS.n1483 VSS.t967 220.952
R752 VSS.n1484 VSS.t1044 220.952
R753 VSS.n2306 VSS.t528 219.972
R754 VSS.n721 VSS.n572 218.506
R755 VSS.n721 VSS.n573 218.506
R756 VSS.n1607 VSS.n1413 218.506
R757 VSS.n1554 VSS.n1447 218.506
R758 VSS.n919 VSS.n918 218.506
R759 VSS.n1119 VSS.n1118 218.506
R760 VSS.n977 VSS.n976 218.506
R761 VSS.n1101 VSS.n1100 218.506
R762 VSS.n1734 VSS.t1060 218.308
R763 VSS.n1880 VSS.t1073 218.308
R764 VSS.n725 VSS.t1001 218.308
R765 VSS.n688 VSS.t1054 218.308
R766 VSS.n2269 VSS.t1027 218.308
R767 VSS.n2198 VSS.t1016 218.308
R768 VSS.n1646 VSS.t994 218.308
R769 VSS.n2605 VSS.t970 218.308
R770 VSS.n2716 VSS.t1045 218.308
R771 VSS.n2820 VSS.t1000 218.308
R772 VSS.n2848 VSS.t1026 218.308
R773 VSS.n83 VSS.t973 218.308
R774 VSS.n1466 VSS.n1465 218.13
R775 VSS.n543 VSS.t401 217.977
R776 VSS.n1291 VSS.t500 217.977
R777 VSS.n2537 VSS.t643 217.977
R778 VSS.n2516 VSS.t429 217.977
R779 VSS.n1278 VSS.t586 217.953
R780 VSS.n264 VSS.t535 217.953
R781 VSS.n1299 VSS.t589 217.892
R782 VSS.n2535 VSS.t439 217.892
R783 VSS.n1377 VSS.t516 216.933
R784 VSS.n1280 VSS.t377 216.589
R785 VSS.n252 VSS.t543 216.589
R786 VSS.n552 VSS.t593 216.579
R787 VSS.n1411 VSS.t450 215.992
R788 VSS.n1279 VSS.t378 214.487
R789 VSS.n251 VSS.t544 214.487
R790 VSS.n125 VSS.t383 214.456
R791 VSS.n144 VSS.t384 214.456
R792 VSS.n187 VSS.t366 214.456
R793 VSS.n175 VSS.t365 214.456
R794 VSS.n190 VSS.t578 214.456
R795 VSS.n188 VSS.t577 214.456
R796 VSS.n304 VSS.t433 214.456
R797 VSS.n302 VSS.t432 214.456
R798 VSS.n450 VSS.t572 214.456
R799 VSS.n453 VSS.t571 214.456
R800 VSS.n289 VSS.t487 214.456
R801 VSS.n435 VSS.t488 214.456
R802 VSS.n270 VSS.t620 214.456
R803 VSS.n420 VSS.t619 214.456
R804 VSS.n326 VSS.t603 214.456
R805 VSS.n325 VSS.t602 214.456
R806 VSS.n389 VSS.t511 214.456
R807 VSS.n340 VSS.t510 214.456
R808 VSS.n362 VSS.t413 214.456
R809 VSS.n345 VSS.t412 214.456
R810 VSS.n2437 VSS.t534 214.456
R811 VSS.n2425 VSS.t514 214.456
R812 VSS.n2420 VSS.t399 214.456
R813 VSS.n2451 VSS.t513 214.456
R814 VSS.n2405 VSS.t381 214.456
R815 VSS.n2459 VSS.t398 214.456
R816 VSS.n2459 VSS.t380 214.456
R817 VSS.n2396 VSS.t498 214.456
R818 VSS.n2396 VSS.t497 214.456
R819 VSS.n2397 VSS.t465 214.456
R820 VSS.n2397 VSS.t464 214.456
R821 VSS.n1697 VSS.t471 214.456
R822 VSS.n1705 VSS.t470 214.456
R823 VSS.n1733 VSS.t656 214.456
R824 VSS.n1731 VSS.t655 214.456
R825 VSS.n1757 VSS.t634 214.456
R826 VSS.n1744 VSS.t635 214.456
R827 VSS.n1811 VSS.t387 214.456
R828 VSS.n1809 VSS.t386 214.456
R829 VSS.n1790 VSS.t672 214.456
R830 VSS.n1789 VSS.t671 214.456
R831 VSS.n1848 VSS.t390 214.456
R832 VSS.n1075 VSS.t389 214.456
R833 VSS.n1879 VSS.t629 214.456
R834 VSS.n1068 VSS.t628 214.456
R835 VSS.n1051 VSS.t665 214.456
R836 VSS.n1050 VSS.t664 214.456
R837 VSS.n1035 VSS.t647 214.456
R838 VSS.n1034 VSS.t646 214.456
R839 VSS.n1179 VSS.t396 214.456
R840 VSS.n1170 VSS.t395 214.456
R841 VSS.n1160 VSS.t493 214.456
R842 VSS.n1142 VSS.t492 214.456
R843 VSS.n1144 VSS.t517 214.456
R844 VSS.n517 VSS.t441 214.456
R845 VSS.n521 VSS.t427 214.456
R846 VSS.n516 VSS.t617 214.456
R847 VSS.n513 VSS.t426 214.456
R848 VSS.n506 VSS.t597 214.456
R849 VSS.n475 VSS.t616 214.456
R850 VSS.n475 VSS.t596 214.456
R851 VSS.n479 VSS.t410 214.456
R852 VSS.n479 VSS.t409 214.456
R853 VSS.n499 VSS.t369 214.456
R854 VSS.n499 VSS.t368 214.456
R855 VSS.n476 VSS.t583 214.456
R856 VSS.n476 VSS.t582 214.456
R857 VSS.n477 VSS.t560 214.456
R858 VSS.n477 VSS.t559 214.456
R859 VSS.n596 VSS.t563 214.456
R860 VSS.n668 VSS.t652 214.456
R861 VSS.n689 VSS.t372 214.456
R862 VSS.n682 VSS.t371 214.456
R863 VSS.n689 VSS.t653 214.456
R864 VSS.n726 VSS.t523 214.456
R865 VSS.n737 VSS.t522 214.456
R866 VSS.n727 VSS.t415 214.456
R867 VSS.n727 VSS.t414 214.456
R868 VSS.n729 VSS.t393 214.456
R869 VSS.n729 VSS.t392 214.456
R870 VSS.n644 VSS.t562 214.456
R871 VSS.n655 VSS.t445 214.456
R872 VSS.n607 VSS.t650 214.456
R873 VSS.n633 VSS.t444 214.456
R874 VSS.n614 VSS.t549 214.456
R875 VSS.n2354 VSS.t442 214.456
R876 VSS.n525 VSS.t548 214.456
R877 VSS.n548 VSS.t402 214.456
R878 VSS.n2334 VSS.t417 214.456
R879 VSS.n551 VSS.t529 214.456
R880 VSS.n766 VSS.t594 214.456
R881 VSS.n797 VSS.t420 214.456
R882 VSS.n809 VSS.t662 214.456
R883 VSS.n804 VSS.t661 214.456
R884 VSS.n809 VSS.t421 214.456
R885 VSS.n810 VSS.t566 214.456
R886 VSS.n810 VSS.t565 214.456
R887 VSS.n812 VSS.t624 214.456
R888 VSS.n812 VSS.t623 214.456
R889 VSS.n1301 VSS.t501 214.456
R890 VSS.n1315 VSS.t588 214.456
R891 VSS.n1193 VSS.t585 214.456
R892 VSS.n1274 VSS.t659 214.456
R893 VSS.n1194 VSS.t459 214.456
R894 VSS.n1245 VSS.t658 214.456
R895 VSS.n1238 VSS.t532 214.456
R896 VSS.n1205 VSS.t458 214.456
R897 VSS.n1205 VSS.t531 214.456
R898 VSS.n1206 VSS.t424 214.456
R899 VSS.n1206 VSS.t423 214.456
R900 VSS.n1207 VSS.t490 214.456
R901 VSS.n1207 VSS.t489 214.456
R902 VSS.n1209 VSS.t557 214.456
R903 VSS.n1209 VSS.t556 214.456
R904 VSS.n1231 VSS.t614 214.456
R905 VSS.n1231 VSS.t613 214.456
R906 VSS.n1138 VSS.t626 214.456
R907 VSS.n1138 VSS.t625 214.456
R908 VSS.n1386 VSS.t408 214.456
R909 VSS.n1386 VSS.t407 214.456
R910 VSS.n2199 VSS.t600 214.456
R911 VSS.n868 VSS.t599 214.456
R912 VSS.n849 VSS.t508 214.456
R913 VSS.n2210 VSS.t507 214.456
R914 VSS.n2248 VSS.t637 214.456
R915 VSS.n2268 VSS.t569 214.456
R916 VSS.n2260 VSS.t568 214.456
R917 VSS.n2268 VSS.t638 214.456
R918 VSS.n2262 VSS.t462 214.456
R919 VSS.n2262 VSS.t461 214.456
R920 VSS.n2263 VSS.t546 214.456
R921 VSS.n2263 VSS.t545 214.456
R922 VSS.n944 VSS.t482 214.456
R923 VSS.n942 VSS.t481 214.456
R924 VSS.n1561 VSS.t496 214.456
R925 VSS.n1440 VSS.t495 214.456
R926 VSS.n1598 VSS.t451 214.456
R927 VSS.n1613 VSS.t612 214.456
R928 VSS.n1403 VSS.t611 214.456
R929 VSS.n1400 VSS.t552 214.456
R930 VSS.n1400 VSS.t551 214.456
R931 VSS.n1402 VSS.t622 214.456
R932 VSS.n1402 VSS.t621 214.456
R933 VSS.n1483 VSS.t520 214.456
R934 VSS.n1483 VSS.t519 214.456
R935 VSS.n1484 VSS.t591 214.456
R936 VSS.n1484 VSS.t590 214.456
R937 VSS.n948 VSS.t361 214.456
R938 VSS.n948 VSS.t360 214.456
R939 VSS.n949 VSS.t453 214.456
R940 VSS.n949 VSS.t452 214.456
R941 VSS.n1122 VSS.t541 214.456
R942 VSS.n1123 VSS.t540 214.456
R943 VSS.n1125 VSS.t554 214.456
R944 VSS.n1125 VSS.t553 214.456
R945 VSS.n1128 VSS.t538 214.456
R946 VSS.n1128 VSS.t537 214.456
R947 VSS.n2065 VSS.t485 214.456
R948 VSS.n2055 VSS.t484 214.456
R949 VSS.n2065 VSS.t468 214.456
R950 VSS.n2054 VSS.t467 214.456
R951 VSS.n970 VSS.t632 214.456
R952 VSS.n2044 VSS.t631 214.456
R953 VSS.n2002 VSS.t476 214.456
R954 VSS.n2001 VSS.t475 214.456
R955 VSS.n990 VSS.t456 214.456
R956 VSS.n1960 VSS.t455 214.456
R957 VSS.n2060 VSS.t375 214.456
R958 VSS.n2060 VSS.t374 214.456
R959 VSS.n2061 VSS.t669 214.456
R960 VSS.n2061 VSS.t668 214.456
R961 VSS.n2399 VSS.t667 214.456
R962 VSS.n2399 VSS.t666 214.456
R963 VSS.n2468 VSS.t641 214.456
R964 VSS.n2468 VSS.t640 214.456
R965 VSS.n2604 VSS.t606 214.456
R966 VSS.n2604 VSS.t581 214.456
R967 VSS.n2596 VSS.t580 214.456
R968 VSS.n2582 VSS.t605 214.456
R969 VSS.n2578 VSS.t473 214.456
R970 VSS.n224 VSS.t472 214.456
R971 VSS.n2578 VSS.t448 214.456
R972 VSS.n224 VSS.t447 214.456
R973 VSS.n225 VSS.t575 214.456
R974 VSS.n227 VSS.t644 214.456
R975 VSS.n2540 VSS.t574 214.456
R976 VSS.n244 VSS.t430 214.456
R977 VSS.n2518 VSS.t438 214.456
R978 VSS.n2598 VSS.t503 214.456
R979 VSS.n2598 VSS.t502 214.456
R980 VSS.n2599 VSS.t479 214.456
R981 VSS.n2599 VSS.t478 214.456
R982 VSS.n2717 VSS.t405 214.456
R983 VSS.n101 VSS.t404 214.456
R984 VSS.n2821 VSS.t526 214.456
R985 VSS.n98 VSS.t525 214.456
R986 VSS.n84 VSS.t609 214.456
R987 VSS.n90 VSS.t608 214.456
R988 VSS.n2847 VSS.t436 214.456
R989 VSS.n2853 VSS.t435 214.456
R990 VSS.n117 VSS.n114 214.409
R991 VSS.n2696 VSS.n2695 213.911
R992 VSS.n8 VSS.n7 212.78
R993 VSS.n1529 VSS.n1470 212.317
R994 VSS.t431 VSS.t570 211.531
R995 VSS.t764 VSS 210.728
R996 VSS.n1481 VSS.n1480 207.965
R997 VSS.n2028 VSS.n2027 207.965
R998 VSS.n2141 VSS.n891 206.909
R999 VSS.n1569 VSS.n1568 205.971
R1000 VSS.n882 VSS.n881 205.899
R1001 VSS.n2159 VSS.n885 205.899
R1002 VSS.n2166 VSS.n2165 205.481
R1003 VSS.n1434 VSS.n1433 205.481
R1004 VSS.n2246 VSS.n2245 205.385
R1005 VSS.n2187 VSS.n2185 204.692
R1006 VSS.n887 VSS.n886 204.692
R1007 VSS.n988 VSS.n986 204.457
R1008 VSS.n988 VSS.n987 204.457
R1009 VSS.n2014 VSS.n2013 204.457
R1010 VSS.n2707 VSS.n103 204.457
R1011 VSS.n791 VSS.n790 204.201
R1012 VSS.n1005 VSS.n1004 204.201
R1013 VSS.n993 VSS.n992 204.201
R1014 VSS.n864 VSS.n863 202.724
R1015 VSS.n2220 VSS.n2219 202.724
R1016 VSS.n2145 VSS.n2142 202.724
R1017 VSS.n1553 VSS.n1448 202.724
R1018 VSS.n1460 VSS.n1459 202.724
R1019 VSS VSS.t272 202.299
R1020 VSS.t214 VSS.t52 202.299
R1021 VSS.t159 VSS.t765 202.299
R1022 VSS.t342 VSS.t834 202.299
R1023 VSS.n2240 VSS.n851 201.458
R1024 VSS.n1437 VSS.n1436 201.458
R1025 VSS.n873 VSS.n872 201.129
R1026 VSS.n2255 VSS.n846 201.129
R1027 VSS.n2250 VSS.n2249 201.129
R1028 VSS.n1578 VSS.n1435 201.129
R1029 VSS.n164 VSS.n163 200.692
R1030 VSS.n437 VSS.n436 200.692
R1031 VSS.n1853 VSS.n1852 200.692
R1032 VSS.n627 VSS.n626 200.692
R1033 VSS.n1600 VSS.n1599 200.692
R1034 VSS.n1502 VSS.n1482 200.516
R1035 VSS.n1115 VSS.n1114 200.516
R1036 VSS.n2257 VSS.n845 200.508
R1037 VSS.n2232 VSS.n855 200.508
R1038 VSS.n853 VSS.n852 200.508
R1039 VSS.n2151 VSS.n889 200.508
R1040 VSS.n1422 VSS.n1421 200.508
R1041 VSS.n1563 VSS.n1442 200.508
R1042 VSS.n1445 VSS.n1444 200.508
R1043 VSS.n2192 VSS.n870 200.231
R1044 VSS.n2844 VSS.n73 200.231
R1045 VSS.n2836 VSS.n79 200.231
R1046 VSS.n1489 VSS.n1488 200.127
R1047 VSS.n1652 VSS.n1121 200.127
R1048 VSS.n88 VSS.n82 200.105
R1049 VSS.n143 VSS.n142 199.739
R1050 VSS.n1750 VSS.n1747 199.739
R1051 VSS.n1740 VSS.n1687 199.739
R1052 VSS.n1726 VSS.n1693 199.739
R1053 VSS.n1695 VSS.n1694 199.739
R1054 VSS.n1047 VSS.n1046 199.739
R1055 VSS.n1054 VSS.n1053 199.739
R1056 VSS.n1874 VSS.n1072 199.739
R1057 VSS.n584 VSS.n582 199.739
R1058 VSS.n584 VSS.n583 199.739
R1059 VSS.n2140 VSS.n894 199.739
R1060 VSS.n1527 VSS.n1472 199.739
R1061 VSS.n1107 VSS.n1095 199.739
R1062 VSS.n1786 VSS.n1785 199.739
R1063 VSS.n1794 VSS.n1793 199.739
R1064 VSS.n1818 VSS.n1808 199.739
R1065 VSS.n768 VSS.n767 199.662
R1066 VSS.n712 VSS.n577 199.53
R1067 VSS.n712 VSS.n579 199.53
R1068 VSS.n2160 VSS.n884 199.53
R1069 VSS.n1535 VSS.n1467 199.53
R1070 VSS.n2109 VSS.n920 199.53
R1071 VSS.n1664 VSS.n1113 199.53
R1072 VSS.n1014 VSS.n1013 199.53
R1073 VSS.n2038 VSS.n2035 199.53
R1074 VSS.t240 VSS 198.519
R1075 VSS.t731 VSS 198.519
R1076 VSS.t747 VSS 198.519
R1077 VSS.t354 VSS 198.519
R1078 VSS.n1158 VSS.n1157 197.476
R1079 VSS.n2592 VSS.n2591 196.831
R1080 VSS.n1592 VSS.n1420 196.589
R1081 VSS.n2101 VSS.n923 196.589
R1082 VSS.n1146 VSS.n1145 196.442
R1083 VSS.n2144 VSS.n2143 196.442
R1084 VSS.n1571 VSS.n1439 196.442
R1085 VSS.n925 VSS.n924 196.442
R1086 VSS.n955 VSS.n943 196.442
R1087 VSS VSS.t469 195.036
R1088 VSS.n2790 VSS.n2789 195
R1089 VSS.n2791 VSS.n2790 195
R1090 VSS.n2764 VSS.n2763 195
R1091 VSS.n2765 VSS.n2764 195
R1092 VSS.n2769 VSS.n2768 195
R1093 VSS.n2768 VSS.n2767 195
R1094 VSS.n2747 VSS.n2746 195
R1095 VSS.n2746 VSS.n2745 195
R1096 VSS.n2752 VSS.n2751 195
R1097 VSS.n2753 VSS.n2752 195
R1098 VSS.n2781 VSS.n2780 195
R1099 VSS.n2782 VSS.n2781 195
R1100 VSS.n2756 VSS.n2731 195
R1101 VSS.n2757 VSS.n2756 195
R1102 VSS.n2786 VSS.n2785 195
R1103 VSS.n2785 VSS.n2784 195
R1104 VSS.t170 VSS.t139 193.87
R1105 VSS.t891 VSS.t953 193.87
R1106 VSS.n162 VSS.n161 190.399
R1107 VSS.n294 VSS.n292 190.399
R1108 VSS.n1851 VSS.n1850 190.399
R1109 VSS.n625 VSS.n624 190.399
R1110 VSS.n1417 VSS.n1414 190.399
R1111 VSS.n1010 VSS.n1009 189.268
R1112 VSS.n969 VSS.n968 189.201
R1113 VSS.t806 VSS.t80 185.441
R1114 VSS.t824 VSS.t44 185.441
R1115 VSS.t864 VSS.t853 177.012
R1116 VSS.t242 VSS.t129 177.012
R1117 VSS.t930 VSS.t836 177.012
R1118 VSS VSS.t959 177.012
R1119 VSS.n2683 VSS 174.232
R1120 VSS.t74 VSS.t85 168.583
R1121 VSS.t754 VSS.t838 168.583
R1122 VSS.t123 VSS 163.831
R1123 VSS.n2813 VSS.t237 162.471
R1124 VSS.n2808 VSS.t734 162.471
R1125 VSS.n2804 VSS.t745 162.471
R1126 VSS.n2799 VSS.t357 162.471
R1127 VSS.n2839 VSS.t768 162.471
R1128 VSS.n9 VSS.t222 162.022
R1129 VSS.n57 VSS.t323 162.022
R1130 VSS.n52 VSS.t338 162.022
R1131 VSS.n47 VSS.t33 162.022
R1132 VSS.n42 VSS.t789 162.022
R1133 VSS.n37 VSS.t770 162.022
R1134 VSS.n32 VSS.t27 162.022
R1135 VSS.n27 VSS.t921 162.022
R1136 VSS.n22 VSS.t919 162.022
R1137 VSS.n58 VSS.t11 162.022
R1138 VSS.n12 VSS.t320 162.022
R1139 VSS.n13 VSS.t316 162.022
R1140 VSS.n14 VSS.t261 162.022
R1141 VSS.n15 VSS.t964 162.022
R1142 VSS.n16 VSS.t306 162.022
R1143 VSS.n17 VSS.t192 162.022
R1144 VSS.n18 VSS.t197 162.022
R1145 VSS.n1 VSS.t751 162.022
R1146 VSS.n2844 VSS.t363 160.046
R1147 VSS.n2836 VSS.t721 160.046
R1148 VSS.n9 VSS.t9 160.017
R1149 VSS.n57 VSS.t318 160.017
R1150 VSS.n52 VSS.t314 160.017
R1151 VSS.n47 VSS.t260 160.017
R1152 VSS.n42 VSS.t963 160.017
R1153 VSS.n37 VSS.t304 160.017
R1154 VSS.n32 VSS.t193 160.017
R1155 VSS.n27 VSS.t195 160.017
R1156 VSS.n22 VSS.t753 160.017
R1157 VSS.n2719 VSS.t241 160.017
R1158 VSS.n2806 VSS.t732 160.017
R1159 VSS.n2795 VSS.t748 160.017
R1160 VSS.n97 VSS.t355 160.017
R1161 VSS.n58 VSS.t223 160.017
R1162 VSS.n12 VSS.t324 160.017
R1163 VSS.n13 VSS.t339 160.017
R1164 VSS.n14 VSS.t31 160.017
R1165 VSS.n15 VSS.t787 160.017
R1166 VSS.n16 VSS.t769 160.017
R1167 VSS.n17 VSS.t29 160.017
R1168 VSS.n18 VSS.t922 160.017
R1169 VSS.n1 VSS.t920 160.017
R1170 VSS.n2837 VSS.t926 160.017
R1171 VSS.n80 VSS.t723 160.017
R1172 VSS.n74 VSS.t505 158.534
R1173 VSS.n2096 VSS.t766 154.131
R1174 VSS VSS.n2682 152.518
R1175 VSS.n782 VSS.t211 152.381
R1176 VSS.n939 VSS.t336 152.381
R1177 VSS.n947 VSS.t82 152.381
R1178 VSS.n163 VSS.n146 152
R1179 VSS.n626 VSS.n613 152
R1180 VSS.n1601 VSS.n1600 152
R1181 VSS.n1852 VSS.n1784 152
R1182 VSS.n438 VSS.n437 152
R1183 VSS.n774 VSS.t897 150.101
R1184 VSS.n947 VSS.t330 150.101
R1185 VSS VSS.n2864 144.951
R1186 VSS.n2114 VSS.t215 144.886
R1187 VSS.n1658 VSS.t130 144.886
R1188 VSS.t881 VSS.t873 143.296
R1189 VSS.n1486 VSS 143.296
R1190 VSS.t474 VSS 143.296
R1191 VSS.n2498 VSS.t601 141.022
R1192 VSS.t203 VSS 135.415
R1193 VSS.t822 VSS.t109 134.867
R1194 VSS.t244 VSS.t127 134.867
R1195 VSS.t773 VSS.t165 134.867
R1196 VSS.t68 VSS.t327 134.867
R1197 VSS.n65 VSS.t331 133.507
R1198 VSS.t115 VSS.t72 126.438
R1199 VSS.n2579 VSS.t349 124.688
R1200 VSS.n1744 VSS.t1070 121.927
R1201 VSS.n1790 VSS.t1056 121.927
R1202 VSS.n1051 VSS.t1059 121.927
R1203 VSS.n1035 VSS.t1063 121.927
R1204 VSS.n944 VSS.t982 121.927
R1205 VSS VSS.t353 121.481
R1206 VSS VSS.t881 118.008
R1207 VSS.t683 VSS.t636 118.008
R1208 VSS.t288 VSS.t898 118.008
R1209 VSS.t862 VSS.t708 118.008
R1210 VSS.n2066 VSS.t1008 116.734
R1211 VSS.n1371 VSS.t1075 116.734
R1212 VSS.n1951 VSS.n1950 114.377
R1213 VSS.n1175 VSS.n1174 110.349
R1214 VSS.n1099 VSS.n1098 110.349
R1215 VSS.t250 VSS.t278 109.579
R1216 VSS.n1443 VSS.t286 109.579
R1217 VSS.t143 VSS.t212 109.579
R1218 VSS.t168 VSS.t810 109.579
R1219 VSS.t118 VSS.t83 109.579
R1220 VSS.n1174 VSS.t867 108.505
R1221 VSS.n1950 VSS.t19 108.505
R1222 VSS.n1098 VSS.t951 108.505
R1223 VSS VSS.t236 106.942
R1224 VSS.t77 VSS.t200 102.992
R1225 VSS.t75 VSS.t957 102.992
R1226 VSS.n506 VSS.t1072 102.353
R1227 VSS.n1238 VSS.t1068 102.353
R1228 VSS.n2405 VSS.t1036 102.353
R1229 VSS.n790 VSS.t255 101.43
R1230 VSS.n1004 VSS.t859 101.43
R1231 VSS.n992 VSS.t60 101.43
R1232 VSS.t394 VSS.t740 101.15
R1233 VSS.t344 VSS.t268 101.15
R1234 VSS.n818 VSS.t999 99.7825
R1235 VSS.n2058 VSS.t983 99.7825
R1236 VSS.t804 VSS.t101 92.7208
R1237 VSS.t262 VSS 92.7208
R1238 VSS.t270 VSS.t944 92.7208
R1239 VSS.t825 VSS.t778 92.7208
R1240 VSS.t337 VSS.t912 92.7208
R1241 VSS VSS.t117 92.7208
R1242 VSS.n2791 VSS.t744 85.9264
R1243 VSS.t925 VSS.t793 84.2917
R1244 VSS.t257 VSS.t604 84.2917
R1245 VSS.n2760 VSS 83.8426
R1246 VSS.t570 VSS 83.54
R1247 VSS.t601 VSS 83.54
R1248 VSS.t198 VSS.t718 75.8626
R1249 VSS VSS.t299 75.4142
R1250 VSS VSS.t20 75.4142
R1251 VSS VSS.t856 75.4142
R1252 VSS.t817 VSS 75.4142
R1253 VSS.t826 VSS 75.4142
R1254 VSS.t832 VSS 75.4142
R1255 VSS VSS.t762 75.4142
R1256 VSS VSS.t776 75.4142
R1257 VSS VSS.t844 75.4142
R1258 VSS.n577 VSS.t860 74.8666
R1259 VSS.n579 VSS.t795 74.8666
R1260 VSS.n884 VSS.t187 74.8666
R1261 VSS.n1420 VSS.t251 74.8666
R1262 VSS.n1467 VSS.t249 74.8666
R1263 VSS.n920 VSS.t140 74.8666
R1264 VSS.n923 VSS.t15 74.8666
R1265 VSS.n1113 VSS.t892 74.8666
R1266 VSS.n1013 VSS.t185 74.8666
R1267 VSS.n2035 VSS.t229 74.8666
R1268 VSS.n986 VSS.t861 72.8576
R1269 VSS.n987 VSS.t831 72.8576
R1270 VSS.n2013 VSS.t742 72.8576
R1271 VSS.n103 VSS.t958 72.8576
R1272 VSS.n82 VSS.t928 72.8576
R1273 VSS.n2683 VSS 72.0437
R1274 VSS.n2691 VSS.n2690 70.7128
R1275 VSS.n2692 VSS.n2691 70.7128
R1276 VSS.t208 VSS.t779 67.4452
R1277 VSS.t141 VSS.t153 67.4335
R1278 VSS.t871 VSS.t294 67.4335
R1279 VSS.t176 VSS.t743 67.4335
R1280 VSS.n2690 VSS.t904 59.664
R1281 VSS.t179 VSS.t847 59.0043
R1282 VSS.n870 VSS.t150 58.5719
R1283 VSS.n1157 VSS.t322 58.5719
R1284 VSS.n73 VSS.t202 58.5719
R1285 VSS.n79 VSS.t960 58.5719
R1286 VSS.t6 VSS.n2692 58.1908
R1287 VSS.t6 VSS.n4 58.1908
R1288 VSS VSS.t431 57.4818
R1289 VSS VSS.n2498 57.4818
R1290 VSS.n2682 VSS 57.4818
R1291 VSS.n2865 VSS.t203 57.2177
R1292 VSS.t200 VSS.t75 57.2177
R1293 VSS.n2856 VSS.n65 57.2177
R1294 VSS.n2776 VSS.n2731 54.2123
R1295 VSS.n2751 VSS.n2742 54.2123
R1296 VSS.n2770 VSS.n2769 54.2123
R1297 VSS.n2789 VSS.n2724 54.2123
R1298 VSS.n2685 VSS.n2684 53.1823
R1299 VSS.n2684 VSS.t906 53.1823
R1300 VSS.n2689 VSS.n2688 53.1823
R1301 VSS.n2690 VSS.n2689 53.1823
R1302 VSS.n2695 VSS.n2694 53.1823
R1303 VSS.n2694 VSS.n4 53.1823
R1304 VSS.n118 VSS.n117 53.1823
R1305 VSS.n2692 VSS.n118 53.1823
R1306 VSS.n767 VSS.t191 52.8576
R1307 VSS.t95 VSS.t182 50.5752
R1308 VSS VSS.t262 50.5752
R1309 VSS.t121 VSS.t362 50.5752
R1310 VSS.t673 VSS.t720 50.5752
R1311 VSS.n2687 VSS.n120 48.7505
R1312 VSS.n122 VSS.n120 48.7505
R1313 VSS.n121 VSS.n119 48.7505
R1314 VSS.n122 VSS.n119 48.7505
R1315 VSS.n1465 VSS.t715 48.5719
R1316 VSS.t236 VSS.n2759 47.9103
R1317 VSS.n1473 VSS.t939 47.1434
R1318 VSS.n2036 VSS.t719 47.1434
R1319 VSS.n2709 VSS 43.9579
R1320 VSS.n2864 VSS.t331 41.9598
R1321 VSS.n767 VSS.t308 40.0005
R1322 VSS.n577 VSS.t333 40.0005
R1323 VSS.n579 VSS.t25 40.0005
R1324 VSS.n872 VSS.t102 40.0005
R1325 VSS.n872 VSS.t114 40.0005
R1326 VSS.n846 VSS.t678 40.0005
R1327 VSS.n846 VSS.t696 40.0005
R1328 VSS.n2249 VSS.t688 40.0005
R1329 VSS.n2249 VSS.t700 40.0005
R1330 VSS.n845 VSS.t676 40.0005
R1331 VSS.n845 VSS.t684 40.0005
R1332 VSS.n863 VSS.t886 40.0005
R1333 VSS.n863 VSS.t911 40.0005
R1334 VSS.n2219 VSS.t809 40.0005
R1335 VSS.n2219 VSS.t690 40.0005
R1336 VSS.n855 VSS.t702 40.0005
R1337 VSS.n855 VSS.t686 40.0005
R1338 VSS.n852 VSS.t698 40.0005
R1339 VSS.n852 VSS.t682 40.0005
R1340 VSS.n851 VSS.t692 40.0005
R1341 VSS.n851 VSS.t706 40.0005
R1342 VSS.n2245 VSS.t680 40.0005
R1343 VSS.n881 VSS.t106 40.0005
R1344 VSS.n2165 VSS.t104 40.0005
R1345 VSS.n2165 VSS.t86 40.0005
R1346 VSS.n2185 VSS.t96 40.0005
R1347 VSS.n2185 VSS.t108 40.0005
R1348 VSS.n884 VSS.t792 40.0005
R1349 VSS.n885 VSS.t110 40.0005
R1350 VSS.n885 VSS.t94 40.0005
R1351 VSS.n886 VSS.t88 40.0005
R1352 VSS.n886 VSS.t98 40.0005
R1353 VSS.n889 VSS.t90 40.0005
R1354 VSS.n889 VSS.t100 40.0005
R1355 VSS.n2142 VSS.t882 40.0005
R1356 VSS.n2142 VSS.t116 40.0005
R1357 VSS.n891 VSS.t880 40.0005
R1358 VSS.n891 VSS.t890 40.0005
R1359 VSS.n1421 VSS.t281 40.0005
R1360 VSS.n1421 VSS.t293 40.0005
R1361 VSS.n1420 VSS.t785 40.0005
R1362 VSS.n1433 VSS.t275 40.0005
R1363 VSS.n1433 VSS.t289 40.0005
R1364 VSS.n1435 VSS.t269 40.0005
R1365 VSS.n1435 VSS.t285 40.0005
R1366 VSS.n1436 VSS.t283 40.0005
R1367 VSS.n1568 VSS.t263 40.0005
R1368 VSS.n1568 VSS.t277 40.0005
R1369 VSS.n1442 VSS.t291 40.0005
R1370 VSS.n1442 VSS.t273 40.0005
R1371 VSS.n1444 VSS.t287 40.0005
R1372 VSS.n1444 VSS.t267 40.0005
R1373 VSS.n1448 VSS.t271 40.0005
R1374 VSS.n1448 VSS.t144 40.0005
R1375 VSS.n1459 VSS.t841 40.0005
R1376 VSS.n1459 VSS.t884 40.0005
R1377 VSS.n1467 VSS.t949 40.0005
R1378 VSS.n920 VSS.t739 40.0005
R1379 VSS.n923 VSS.t956 40.0005
R1380 VSS.n1113 VSS.t799 40.0005
R1381 VSS.n1013 VSS.t70 40.0005
R1382 VSS.n2035 VSS.t199 40.0005
R1383 VSS.n1174 VSS.t966 38.7697
R1384 VSS.n1482 VSS.t312 38.7697
R1385 VSS.n1114 VSS.t837 38.7697
R1386 VSS.n1950 VSS.t328 38.7697
R1387 VSS.n1098 VSS.t870 38.7697
R1388 VSS.n1095 VSS.t177 38.5719
R1389 VSS.n1095 VSS.t709 38.5719
R1390 VSS.n582 VSS.t247 38.5719
R1391 VSS.n582 VSS.t220 38.5719
R1392 VSS.n583 VSS.t933 38.5719
R1393 VSS.n583 VSS.t40 38.5719
R1394 VSS.n2245 VSS.t704 38.5719
R1395 VSS.n881 VSS.t92 38.5719
R1396 VSS.n2143 VSS.t874 38.5719
R1397 VSS.n2143 VSS.t73 38.5719
R1398 VSS.n1436 VSS.t265 38.5719
R1399 VSS.n1439 VSS.t900 38.5719
R1400 VSS.n1439 VSS.t711 38.5719
R1401 VSS.n1470 VSS.t17 38.5719
R1402 VSS.n1470 VSS.t937 38.5719
R1403 VSS.n1472 VSS.t167 38.5719
R1404 VSS.n1472 VSS.t839 38.5719
R1405 VSS.n924 VSS.t50 38.5719
R1406 VSS.n924 VSS.t48 38.5719
R1407 VSS.n943 VSS.t158 38.5719
R1408 VSS.n943 VSS.t935 38.5719
R1409 VSS.n1009 VSS.t66 38.5719
R1410 VSS.n1009 VSS.t876 38.5719
R1411 VSS.n968 VSS.t120 38.5719
R1412 VSS.n968 VSS.t5 38.5719
R1413 VSS.n1473 VSS.t755 35.4291
R1414 VSS.n2036 VSS.t848 35.4291
R1415 VSS.t135 VSS.t931 35.3567
R1416 VSS.t931 VSS.t12 35.3567
R1417 VSS.t224 VSS.t137 35.3567
R1418 VSS.t137 VSS.t226 35.3567
R1419 VSS.t226 VSS.t904 35.3567
R1420 VSS.n2154 VSS.n2153 34.6358
R1421 VSS.n2677 VSS.n123 34.6358
R1422 VSS.n1742 VSS.n1741 34.6358
R1423 VSS.n1725 VSS.n1724 34.6358
R1424 VSS.n1905 VSS.n1904 34.6358
R1425 VSS.n1886 VSS.n1067 34.6358
R1426 VSS.n749 VSS.n748 34.6358
R1427 VSS.n714 VSS.n713 34.6358
R1428 VSS.n714 VSS.n575 34.6358
R1429 VSS.n718 VSS.n575 34.6358
R1430 VSS.n707 VSS.n580 34.6358
R1431 VSS.n711 VSS.n580 34.6358
R1432 VSS.n2184 VSS.n873 34.6358
R1433 VSS.n2158 VSS.n2157 34.6358
R1434 VSS.n2150 VSS.n890 34.6358
R1435 VSS.n1556 VSS.n1555 34.6358
R1436 VSS.n1552 VSS.n1449 34.6358
R1437 VSS.n1539 VSS.n1463 34.6358
R1438 VSS.n1534 VSS.n1533 34.6358
R1439 VSS.n1533 VSS.n1468 34.6358
R1440 VSS.n1521 VSS.n1477 34.6358
R1441 VSS.n2113 VSS.n916 34.6358
R1442 VSS.n2107 VSS.n921 34.6358
R1443 VSS.n2095 VSS.n927 34.6358
R1444 VSS.n1936 VSS.n1027 34.6358
R1445 VSS.n1937 VSS.n1936 34.6358
R1446 VSS.n1938 VSS.n1937 34.6358
R1447 VSS.n1991 VSS.n1990 34.6358
R1448 VSS.n1995 VSS.n1994 34.6358
R1449 VSS.n1996 VSS.n1995 34.6358
R1450 VSS.n2033 VSS.n974 34.6358
R1451 VSS.n2034 VSS.n2033 34.6358
R1452 VSS.n2042 VSS.n972 34.6358
R1453 VSS.n1106 VSS.n1096 34.6358
R1454 VSS.n1932 VSS.n1028 34.6358
R1455 VSS.n1842 VSS.n1841 34.6358
R1456 VSS.n1823 VSS.n1822 34.6358
R1457 VSS.n1822 VSS.n1806 34.6358
R1458 VSS.n2709 VSS.n2708 34.6358
R1459 VSS.n2706 VSS.n66 34.6358
R1460 VSS.n162 VSS.t1042 34.2973
R1461 VSS.n294 VSS.t1004 34.2973
R1462 VSS.n1851 VSS.t1050 34.2973
R1463 VSS.n625 VSS.t984 34.2973
R1464 VSS.n1417 VSS.t992 34.2973
R1465 VSS.n1571 VSS.n1570 33.8829
R1466 VSS.n2097 VSS.n925 33.8829
R1467 VSS.t107 VSS.t802 33.717
R1468 VSS.t942 VSS.t883 33.717
R1469 VSS.t16 VSS.t756 33.717
R1470 VSS VSS.t79 33.717
R1471 VSS.t335 VSS.t216 33.717
R1472 VSS.t724 VSS.t869 33.717
R1473 VSS.n142 VSS.t780 33.462
R1474 VSS.n142 VSS.t209 33.462
R1475 VSS.n1747 VSS.t857 33.462
R1476 VSS.n1747 VSS.t772 33.462
R1477 VSS.n1687 VSS.t21 33.462
R1478 VSS.n1687 VSS.t23 33.462
R1479 VSS.n1693 VSS.t962 33.462
R1480 VSS.n1693 VSS.t124 33.462
R1481 VSS.n1694 VSS.t300 33.462
R1482 VSS.n1694 VSS.t302 33.462
R1483 VSS.n1046 VSS.t818 33.462
R1484 VSS.n1046 VSS.t820 33.462
R1485 VSS.n1053 VSS.t827 33.462
R1486 VSS.n1053 VSS.t797 33.462
R1487 VSS.n1072 VSS.t833 33.462
R1488 VSS.n1072 VSS.t326 33.462
R1489 VSS.n1145 VSS.t852 33.462
R1490 VSS.n1145 VSS.t347 33.462
R1491 VSS.n894 VSS.t235 33.462
R1492 VSS.n894 VSS.t46 33.462
R1493 VSS.n1785 VSS.t763 33.462
R1494 VSS.n1785 VSS.t947 33.462
R1495 VSS.n1793 VSS.t777 33.462
R1496 VSS.n1793 VSS.t829 33.462
R1497 VSS.n1808 VSS.t845 33.462
R1498 VSS.n1808 VSS.t207 33.462
R1499 VSS.n109 VSS.t905 32.8043
R1500 VSS.n106 VSS.t907 32.8043
R1501 VSS.n1465 VSS.t761 32.5719
R1502 VSS.n721 VSS.n720 32.377
R1503 VSS.n1656 VSS.n1119 32.377
R1504 VSS.n2025 VSS.n977 32.377
R1505 VSS.n1101 VSS.n1028 32.377
R1506 VSS.n1576 VSS.n1575 32.377
R1507 VSS.n1099 VSS.n1096 31.624
R1508 VSS.n720 VSS.n719 31.2476
R1509 VSS.n1491 VSS.n1490 31.2476
R1510 VSS.n1657 VSS.n1656 31.2476
R1511 VSS.n2026 VSS.n2025 31.2476
R1512 VSS.n712 VSS.n711 30.8711
R1513 VSS.n1535 VSS.n1534 30.8711
R1514 VSS.n1665 VSS.n1664 30.8711
R1515 VSS.n1949 VSS.n1014 30.8711
R1516 VSS.n2778 VSS.n2731 30.8711
R1517 VSS.n2751 VSS.n2750 30.8711
R1518 VSS.n2769 VSS.n2736 30.8711
R1519 VSS.n2789 VSS.n2788 30.8711
R1520 VSS.n1432 VSS.n1422 30.4946
R1521 VSS.n1522 VSS.n1521 30.4946
R1522 VSS.n1666 VSS.n1665 30.4946
R1523 VSS.n2698 VSS.t7 30.3424
R1524 VSS.n2168 VSS.n2167 30.1181
R1525 VSS.n1579 VSS.n1578 30.1181
R1526 VSS.n1462 VSS.n1461 30.1181
R1527 VSS.n1029 VSS.n1027 30.1181
R1528 VSS.n2863 VSS.n8 29.8168
R1529 VSS.n2166 VSS.n2164 29.7417
R1530 VSS.n1496 VSS.n1495 29.3652
R1531 VSS.n2188 VSS.n2187 28.9887
R1532 VSS.n2760 VSS.n5 28.4645
R1533 VSS.n2146 VSS.n2145 27.8593
R1534 VSS.n1553 VSS.n1552 27.8593
R1535 VSS.n707 VSS.n706 27.4829
R1536 VSS.n1529 VSS.n1468 27.4829
R1537 VSS.n1502 VSS.n1501 27.4829
R1538 VSS.n2109 VSS.n2108 27.4829
R1539 VSS.n2103 VSS.n921 27.4829
R1540 VSS.n1112 VSS.n1093 27.4829
R1541 VSS.n1659 VSS.n1115 27.4829
R1542 VSS.n1952 VSS.n1951 27.4829
R1543 VSS.n1952 VSS.n1011 27.4829
R1544 VSS.n2146 VSS.n2141 27.1064
R1545 VSS.n2830 VSS.n2829 26.9246
R1546 VSS.n1523 VSS.n1474 26.7299
R1547 VSS.n174 VSS.n173 26.6009
R1548 VSS.n1990 VSS.n1989 26.314
R1549 VSS.n109 VSS.n108 26.1653
R1550 VSS.n111 VSS.n110 26.1653
R1551 VSS.n106 VSS.n105 26.1653
R1552 VSS.n790 VSS.t310 25.9346
R1553 VSS.n1004 VSS.t58 25.9346
R1554 VSS.n992 VSS.t148 25.9346
R1555 VSS.n1560 VSS.n1559 25.7355
R1556 VSS.n1720 VSS.n1719 25.7355
R1557 VSS.n2012 VSS.n983 25.7355
R1558 VSS.n2043 VSS.n2042 25.7355
R1559 VSS.n1817 VSS.n1816 25.7355
R1560 VSS.n2677 VSS.n2676 25.6926
R1561 VSS.n1758 VSS.n1742 25.6926
R1562 VSS.n1739 VSS.n1689 25.6926
R1563 VSS.n1730 VSS.n1691 25.6926
R1564 VSS.n1904 VSS.n1048 25.6926
R1565 VSS.n1886 VSS.n1885 25.6926
R1566 VSS.n1878 VSS.n1070 25.6926
R1567 VSS.n1841 VSS.n1787 25.6926
R1568 VSS.n2854 VSS.n66 25.6926
R1569 VSS.n748 VSS.n722 25.6005
R1570 VSS.n1575 VSS.n1437 25.6005
R1571 VSS.n870 VSS.t233 25.4291
R1572 VSS.n1157 VSS.t231 25.4291
R1573 VSS.n73 VSS.t122 25.4291
R1574 VSS.n79 VSS.t674 25.4291
R1575 VSS.t252 VSS.t521 25.2879
R1576 VSS.t791 VSS.t93 25.2879
R1577 VSS.t178 VSS.t259 25.2879
R1578 VSS.n1434 VSS.n1432 25.224
R1579 VSS.n1579 VSS.n1434 25.224
R1580 VSS.n2813 VSS.n2812 25.224
R1581 VSS.n2812 VSS.n2719 25.224
R1582 VSS.n2808 VSS.n2807 25.224
R1583 VSS.n2807 VSS.n2806 25.224
R1584 VSS.n2804 VSS.n2803 25.224
R1585 VSS.n2803 VSS.n2795 25.224
R1586 VSS.n2799 VSS.n2798 25.224
R1587 VSS.n2798 VSS.n97 25.224
R1588 VSS.n59 VSS.n9 25.224
R1589 VSS.n59 VSS.n58 25.224
R1590 VSS.n57 VSS.n56 25.224
R1591 VSS.n56 VSS.n12 25.224
R1592 VSS.n52 VSS.n51 25.224
R1593 VSS.n51 VSS.n13 25.224
R1594 VSS.n47 VSS.n46 25.224
R1595 VSS.n46 VSS.n14 25.224
R1596 VSS.n42 VSS.n41 25.224
R1597 VSS.n41 VSS.n15 25.224
R1598 VSS.n37 VSS.n36 25.224
R1599 VSS.n36 VSS.n16 25.224
R1600 VSS.n32 VSS.n31 25.224
R1601 VSS.n31 VSS.n17 25.224
R1602 VSS.n27 VSS.n26 25.224
R1603 VSS.n26 VSS.n18 25.224
R1604 VSS.n22 VSS.n21 25.224
R1605 VSS.n21 VSS.n1 25.224
R1606 VSS.n2839 VSS.n2838 25.224
R1607 VSS.n2838 VSS.n2837 25.224
R1608 VSS.n2835 VSS.n80 25.224
R1609 VSS.n169 VSS.n168 24.9894
R1610 VSS.n1847 VSS.n1846 24.9894
R1611 VSS.n691 VSS.n690 24.968
R1612 VSS.n573 VSS.t781 24.9236
R1613 VSS.n573 VSS.t783 24.9236
R1614 VSS.n572 VSS.t132 24.9236
R1615 VSS.n572 VSS.t1 24.9236
R1616 VSS.n2186 VSS.t183 24.9236
R1617 VSS.n2186 VSS.t803 24.9236
R1618 VSS.n1413 VSS.t56 24.9236
R1619 VSS.n1413 VSS.t903 24.9236
R1620 VSS.n1447 VSS.t945 24.9236
R1621 VSS.n1447 VSS.t213 24.9236
R1622 VSS.n1480 VSS.t913 24.9236
R1623 VSS.n1480 VSS.t854 24.9236
R1624 VSS.n1482 VSS.t865 24.9236
R1625 VSS.n1488 VSS.t142 24.9236
R1626 VSS.n1488 VSS.t872 24.9236
R1627 VSS.n1487 VSS.t154 24.9236
R1628 VSS.n1487 VSS.t295 24.9236
R1629 VSS.n918 VSS.t171 24.9236
R1630 VSS.n918 VSS.t351 24.9236
R1631 VSS.n1114 VSS.t954 24.9236
R1632 VSS.n1118 VSS.t245 24.9236
R1633 VSS.n1118 VSS.t774 24.9236
R1634 VSS.n1121 VSS.t126 24.9236
R1635 VSS.n1121 VSS.t128 24.9236
R1636 VSS.n976 VSS.t341 24.9236
R1637 VSS.n976 VSS.t181 24.9236
R1638 VSS.n2027 VSS.t835 24.9236
R1639 VSS.n2027 VSS.t84 24.9236
R1640 VSS.n1100 VSS.t727 24.9236
R1641 VSS.n1100 VSS.t725 24.9236
R1642 VSS.n2591 VSS.t843 24.9236
R1643 VSS.n2591 VSS.t918 24.9236
R1644 VSS.n7 VSS.t78 24.9236
R1645 VSS.n7 VSS.t76 24.9236
R1646 VSS VSS.t77 24.7946
R1647 VSS.n1593 VSS.n1592 24.4711
R1648 VSS.n2102 VSS.n2101 24.4711
R1649 VSS.n1481 VSS.n1477 24.4711
R1650 VSS.n2097 VSS.n2096 24.4711
R1651 VSS.n2096 VSS.n2095 24.4711
R1652 VSS.n2028 VSS.n974 24.4711
R1653 VSS.n2843 VSS.n74 24.0946
R1654 VSS.n1497 VSS.n1485 23.7181
R1655 VSS.n2681 VSS.n123 23.7181
R1656 VSS.n1927 VSS.n1031 23.7181
R1657 VSS.n1751 VSS.n1746 23.7181
R1658 VSS.n1910 VSS.n1909 23.7181
R1659 VSS.n1897 VSS.n1896 23.7181
R1660 VSS.n1873 VSS.n1872 23.7181
R1661 VSS.n1387 VSS.n1137 23.7181
R1662 VSS.n1378 VSS.n1137 23.7181
R1663 VSS.n2206 VSS.n866 23.7181
R1664 VSS.n2207 VSS.n2206 23.7181
R1665 VSS.n1540 VSS.n1539 23.7181
R1666 VSS.n1501 VSS.n1485 23.7181
R1667 VSS.n2114 VSS.n915 23.7181
R1668 VSS.n2114 VSS.n2113 23.7181
R1669 VSS.n1659 VSS.n1658 23.7181
R1670 VSS.n1996 VSS.n984 23.7181
R1671 VSS.n1834 VSS.n1833 23.7181
R1672 VSS.n941 VSS.n940 23.4338
R1673 VSS.n2151 VSS.n2150 23.3417
R1674 VSS.n1556 VSS.n1445 23.3417
R1675 VSS.n705 VSS.n584 22.9652
R1676 VSS.n706 VSS.n705 22.9652
R1677 VSS.n1529 VSS.n1528 22.9652
R1678 VSS.n1528 VSS.n1527 22.9652
R1679 VSS.n1491 VSS.n1489 22.9652
R1680 VSS.n2103 VSS.n2102 22.9652
R1681 VSS.n1108 VSS.n1093 22.9652
R1682 VSS.n1108 VSS.n1107 22.9652
R1683 VSS.n1653 VSS.n1652 22.9652
R1684 VSS.n1956 VSS.n1011 22.9652
R1685 VSS.n1957 VSS.n1956 22.9652
R1686 VSS.n2038 VSS.n2037 22.9652
R1687 VSS.t353 VSS.n64 22.8805
R1688 VSS.n2683 VSS.t135 22.8347
R1689 VSS.n1540 VSS.n1462 22.5887
R1690 VSS.n986 VSS.t219 22.3257
R1691 VSS.n987 VSS.t156 22.3257
R1692 VSS.n2013 VSS.t924 22.3257
R1693 VSS.n103 VSS.t332 22.3257
R1694 VSS.n82 VSS.t713 22.3257
R1695 VSS.t779 VSS 22.2266
R1696 VSS.n173 VSS.n143 22.2123
R1697 VSS.n169 VSS.n143 22.2123
R1698 VSS.n1750 VSS.n1031 22.2123
R1699 VSS.n1751 VSS.n1750 22.2123
R1700 VSS.n1741 VSS.n1740 22.2123
R1701 VSS.n1740 VSS.n1739 22.2123
R1702 VSS.n1726 VSS.n1691 22.2123
R1703 VSS.n1724 VSS.n1695 22.2123
R1704 VSS.n1726 VSS.n1725 22.2123
R1705 VSS.n1720 VSS.n1695 22.2123
R1706 VSS.n1909 VSS.n1047 22.2123
R1707 VSS.n1905 VSS.n1047 22.2123
R1708 VSS.n1896 VSS.n1054 22.2123
R1709 VSS.n1067 VSS.n1054 22.2123
R1710 VSS.n1874 VSS.n1070 22.2123
R1711 VSS.n1874 VSS.n1873 22.2123
R1712 VSS.n719 VSS.n718 22.2123
R1713 VSS.n1490 VSS.n915 22.2123
R1714 VSS.n2108 VSS.n2107 22.2123
R1715 VSS.n2029 VSS.n2026 22.2123
R1716 VSS.n1846 VSS.n1786 22.2123
R1717 VSS.n1842 VSS.n1786 22.2123
R1718 VSS.n1833 VSS.n1794 22.2123
R1719 VSS.n1823 VSS.n1794 22.2123
R1720 VSS.n1818 VSS.n1806 22.2123
R1721 VSS.n1818 VSS.n1817 22.2123
R1722 VSS.n691 VSS.n584 21.4593
R1723 VSS.n1527 VSS.n1526 21.4593
R1724 VSS.n1495 VSS.n1489 21.4593
R1725 VSS.n1951 VSS.n1949 21.4593
R1726 VSS.n1107 VSS.n1106 21.4593
R1727 VSS.n2844 VSS.n2843 21.4593
R1728 VSS.n2836 VSS.n2835 21.4593
R1729 VSS.n1597 VSS.n1418 20.8482
R1730 VSS.n2168 VSS.n2166 20.7064
R1731 VSS.n2187 VSS.n2184 20.7064
R1732 VSS.n2808 VSS.n2719 20.3299
R1733 VSS.n2799 VSS.n2795 20.3299
R1734 VSS.n5 VSS.t403 20.292
R1735 VSS.t38 VSS.n2865 19.6304
R1736 VSS.n2814 VSS.n2813 19.2926
R1737 VSS.t957 VSS 19.0729
R1738 VSS.n58 VSS.n57 18.824
R1739 VSS.n52 VSS.n12 18.824
R1740 VSS.n47 VSS.n13 18.824
R1741 VSS.n42 VSS.n14 18.824
R1742 VSS.n37 VSS.n15 18.824
R1743 VSS.n32 VSS.n16 18.824
R1744 VSS.n27 VSS.n17 18.824
R1745 VSS.n22 VSS.n18 18.824
R1746 VSS.n388 VSS.n387 18.2791
R1747 VSS.n796 VSS.n795 18.2791
R1748 VSS.n1169 VSS.n1168 18.2791
R1749 VSS.n91 VSS.n80 17.7867
R1750 VSS.n339 VSS.n321 17.7007
R1751 VSS.t12 VSS.n122 17.6786
R1752 VSS.n122 VSS.t224 17.6786
R1753 VSS.n196 VSS.n195 17.4137
R1754 VSS.n2192 VSS.n869 17.3181
R1755 VSS.n2805 VSS.n2804 17.3181
R1756 VSS.n2569 VSS.n2568 17.195
R1757 VSS.n2307 VSS.n2306 16.9936
R1758 VSS.n434 VSS.n295 16.9545
R1759 VSS.n1503 VSS.n1502 16.9417
R1760 VSS.n1663 VSS.n1115 16.9417
R1761 VSS.t851 VSS.t491 16.8587
R1762 VSS.t902 VSS.t449 16.8587
R1763 VSS.t57 VSS.t454 16.8587
R1764 VSS.t940 VSS.t434 16.8587
R1765 VSS.n454 VSS.n286 16.8353
R1766 VSS.n449 VSS.n287 16.7924
R1767 VSS.n2580 VSS.n2579 16.763
R1768 VSS.n2164 VSS.n882 16.1887
R1769 VSS.n2188 VSS.n869 16.1887
R1770 VSS.n1593 VSS.n1418 16.1887
R1771 VSS.n2806 VSS.n2805 15.8123
R1772 VSS.n2829 VSS.n97 15.8123
R1773 VSS.n63 VSS.n9 15.8123
R1774 VSS.n2870 VSS.n1 15.8123
R1775 VSS.n2681 VSS.n124 15.3963
R1776 VSS.n1184 VSS.n893 15.3963
R1777 VSS.n2497 VSS.n2496 15.3963
R1778 VSS.n2497 VSS.n268 14.8179
R1779 VSS.n2000 VSS.n984 14.8179
R1780 VSS.n1927 VSS.n1032 14.775
R1781 VSS.n731 VSS.n730 14.775
R1782 VSS.n2201 VSS.n866 14.775
R1783 VSS.n1619 VSS.n1618 14.775
R1784 VSS.n1642 VSS.n1641 14.775
R1785 VSS.n1872 VSS.n1871 14.775
R1786 VSS.n2829 VSS.n2828 14.775
R1787 VSS.n2846 VSS.n2845 14.775
R1788 VSS.n2635 VSS.n2634 14.2735
R1789 VSS.n2051 VSS.n2050 14.065
R1790 VSS.n814 VSS.n813 14.0503
R1791 VSS.n2267 VSS.n2264 14.0503
R1792 VSS.n2603 VSS.n2600 14.0503
R1793 VSS.n1523 VSS.n1522 13.9299
R1794 VSS.n1666 VSS.n1112 13.9299
R1795 VSS.n2064 VSS.n2063 13.8859
R1796 VSS.n2839 VSS.n74 13.5534
R1797 VSS.n500 VSS.n478 12.8005
R1798 VSS.n1232 VSS.n1208 12.8005
R1799 VSS.n952 VSS.n951 12.8005
R1800 VSS.n2469 VSS.n2398 12.8005
R1801 VSS.n2859 VSS.n63 12.8005
R1802 VSS.n2863 VSS.n6 12.8005
R1803 VSS.n2859 VSS.n6 12.8005
R1804 VSS.n1652 VSS.n1651 12.5161
R1805 VSS.n2307 VSS.n550 12.1384
R1806 VSS.n1570 VSS.n1569 11.9309
R1807 VSS.n1559 VSS.n1445 11.2946
R1808 VSS.n1658 VSS.n1657 11.2946
R1809 VSS.n2712 VSS.n2711 11.2844
R1810 VSS.n2787 VSS.n2723 11.0382
R1811 VSS.n2723 VSS.n2 11.0382
R1812 VSS.n2726 VSS.n2722 11.0382
R1813 VSS.n2722 VSS.n2 11.0382
R1814 VSS.n2762 VSS.n2739 11.0382
R1815 VSS.n2766 VSS.n2739 11.0382
R1816 VSS.n2738 VSS.n2737 11.0382
R1817 VSS.n2766 VSS.n2738 11.0382
R1818 VSS.n2748 VSS.n2741 11.0382
R1819 VSS.n2744 VSS.n2741 11.0382
R1820 VSS.n2743 VSS.n2740 11.0382
R1821 VSS.n2744 VSS.n2740 11.0382
R1822 VSS.n2779 VSS.n2729 11.0382
R1823 VSS.n2755 VSS.n2729 11.0382
R1824 VSS.n2730 VSS.n2728 11.0382
R1825 VSS.n2755 VSS.n2728 11.0382
R1826 VSS.n2353 VSS.n526 10.9091
R1827 VSS.n2209 VSS.n2208 10.8805
R1828 VSS.n1378 VSS.n1377 10.5983
R1829 VSS.n713 VSS.n712 10.5417
R1830 VSS.n2160 VSS.n882 10.5417
R1831 VSS.n1664 VSS.n1663 10.5417
R1832 VSS.n1938 VSS.n1014 10.5417
R1833 VSS.n2038 VSS.n2034 10.5417
R1834 VSS.n2778 VSS.n2777 10.4476
R1835 VSS.n2750 VSS.n2749 10.4476
R1836 VSS.n2771 VSS.n2736 10.4476
R1837 VSS.n2788 VSS.n2725 10.4476
R1838 VSS.n2140 VSS.n893 10.1652
R1839 VSS.n2141 VSS.n2140 10.1652
R1840 VSS.n1592 VSS.n1591 10.1652
R1841 VSS.n1503 VSS.n1481 10.1652
R1842 VSS.n2101 VSS.n2100 10.1652
R1843 VSS.n2029 VSS.n2028 10.1652
R1844 VSS.n2837 VSS.n2836 10.1652
R1845 VSS.n738 VSS.n722 9.88085
R1846 VSS.n1705 VSS.n1702 9.7205
R1847 VSS.n302 VSS.n301 9.7205
R1848 VSS.n190 VSS.n189 9.71789
R1849 VSS.n1811 VSS.n1810 9.71789
R1850 VSS.n2712 VSS.n101 9.70901
R1851 VSS.n2822 VSS.n2821 9.70901
R1852 VSS.n85 VSS.n84 9.70901
R1853 VSS.n1535 VSS.n1466 9.41227
R1854 VSS.n1991 VSS.n988 9.41227
R1855 VSS.n2015 VSS.n2014 9.41227
R1856 VSS.n2707 VSS.n2706 9.41227
R1857 VSS.n483 VSS.n478 9.3031
R1858 VSS.n1214 VSS.n1208 9.3031
R1859 VSS.n1387 VSS.n1134 9.3031
R1860 VSS.n1619 VSS.n1397 9.3031
R1861 VSS.n1641 VSS.n1640 9.3031
R1862 VSS.n2469 VSS.n2393 9.3031
R1863 VSS.n679 VSS.n678 9.3005
R1864 VSS.n676 VSS.n675 9.3005
R1865 VSS.n674 VSS.n597 9.3005
R1866 VSS.n673 VSS.n672 9.3005
R1867 VSS.n671 VSS.n670 9.3005
R1868 VSS.n669 VSS.n599 9.3005
R1869 VSS.n667 VSS.n666 9.3005
R1870 VSS.n677 VSS.n595 9.3005
R1871 VSS.n684 VSS.n683 9.3005
R1872 VSS.n685 VSS.n593 9.3005
R1873 VSS.n687 VSS.n686 9.3005
R1874 VSS.n690 VSS.n591 9.3005
R1875 VSS.n585 VSS.n584 9.3005
R1876 VSS.n706 VSS.n581 9.3005
R1877 VSS.n740 VSS.n722 9.3005
R1878 VSS.n734 VSS.n733 9.3005
R1879 VSS.n732 VSS.n731 9.3005
R1880 VSS.n736 VSS.n724 9.3005
R1881 VSS.n739 VSS.n738 9.3005
R1882 VSS.n748 VSS.n747 9.3005
R1883 VSS.n750 VSS.n749 9.3005
R1884 VSS.n720 VSS.n570 9.3005
R1885 VSS.n719 VSS.n574 9.3005
R1886 VSS.n718 VSS.n717 9.3005
R1887 VSS.n716 VSS.n575 9.3005
R1888 VSS.n715 VSS.n714 9.3005
R1889 VSS.n713 VSS.n576 9.3005
R1890 VSS.n712 VSS.n578 9.3005
R1891 VSS.n711 VSS.n710 9.3005
R1892 VSS.n709 VSS.n580 9.3005
R1893 VSS.n708 VSS.n707 9.3005
R1894 VSS.n705 VSS.n704 9.3005
R1895 VSS.n692 VSS.n691 9.3005
R1896 VSS.n665 VSS.n600 9.3005
R1897 VSS.n657 VSS.n656 9.3005
R1898 VSS.n654 VSS.n605 9.3005
R1899 VSS.n653 VSS.n652 9.3005
R1900 VSS.n646 VSS.n645 9.3005
R1901 VSS.n488 VSS.n478 9.3005
R1902 VSS.n490 VSS.n478 9.3005
R1903 VSS.n2357 VSS.n522 9.3005
R1904 VSS.n2356 VSS.n2355 9.3005
R1905 VSS.n2353 VSS.n2352 9.3005
R1906 VSS.n528 VSS.n527 9.3005
R1907 VSS.n622 VSS.n621 9.3005
R1908 VSS.n623 VSS.n612 9.3005
R1909 VSS.n629 VSS.n628 9.3005
R1910 VSS.n630 VSS.n611 9.3005
R1911 VSS.n632 VSS.n631 9.3005
R1912 VSS.n634 VSS.n610 9.3005
R1913 VSS.n636 VSS.n635 9.3005
R1914 VSS.n638 VSS.n637 9.3005
R1915 VSS.n639 VSS.n608 9.3005
R1916 VSS.n641 VSS.n640 9.3005
R1917 VSS.n643 VSS.n642 9.3005
R1918 VSS.n502 VSS.n501 9.3005
R1919 VSS.n504 VSS.n503 9.3005
R1920 VSS.n505 VSS.n474 9.3005
R1921 VSS.n509 VSS.n508 9.3005
R1922 VSS.n512 VSS.n511 9.3005
R1923 VSS.n514 VSS.n468 9.3005
R1924 VSS.n515 VSS.n469 9.3005
R1925 VSS.n2377 VSS.n2376 9.3005
R1926 VSS.n2375 VSS.n2374 9.3005
R1927 VSS.n2373 VSS.n2372 9.3005
R1928 VSS.n2371 VSS.n518 9.3005
R1929 VSS.n2370 VSS.n2369 9.3005
R1930 VSS.n2368 VSS.n2367 9.3005
R1931 VSS.n2366 VSS.n520 9.3005
R1932 VSS.n2365 VSS.n2364 9.3005
R1933 VSS.n2363 VSS.n2362 9.3005
R1934 VSS.n2359 VSS.n2358 9.3005
R1935 VSS.n2312 VSS.n2311 9.3005
R1936 VSS.n2314 VSS.n2313 9.3005
R1937 VSS.n2316 VSS.n547 9.3005
R1938 VSS.n2318 VSS.n2317 9.3005
R1939 VSS.n2320 VSS.n2319 9.3005
R1940 VSS.n2321 VSS.n545 9.3005
R1941 VSS.n2323 VSS.n2322 9.3005
R1942 VSS.n2324 VSS.n544 9.3005
R1943 VSS.n2333 VSS.n2332 9.3005
R1944 VSS.n2336 VSS.n2335 9.3005
R1945 VSS.n2310 VSS.n2309 9.3005
R1946 VSS.n2308 VSS.n2307 9.3005
R1947 VSS.n2304 VSS.n2303 9.3005
R1948 VSS.n775 VSS.n774 9.3005
R1949 VSS.n771 VSS.n770 9.3005
R1950 VSS.n781 VSS.n780 9.3005
R1951 VSS.n783 VSS.n769 9.3005
R1952 VSS.n787 VSS.n786 9.3005
R1953 VSS.n788 VSS.n768 9.3005
R1954 VSS.n789 VSS 9.3005
R1955 VSS.n793 VSS.n792 9.3005
R1956 VSS.n795 VSS.n794 9.3005
R1957 VSS.n796 VSS.n765 9.3005
R1958 VSS.n799 VSS.n798 9.3005
R1959 VSS.n800 VSS.n764 9.3005
R1960 VSS.n802 VSS.n801 9.3005
R1961 VSS.n803 VSS.n762 9.3005
R1962 VSS.n832 VSS.n831 9.3005
R1963 VSS.n830 VSS.n829 9.3005
R1964 VSS.n822 VSS.n805 9.3005
R1965 VSS.n821 VSS.n820 9.3005
R1966 VSS.n819 VSS.n807 9.3005
R1967 VSS.n817 VSS.n816 9.3005
R1968 VSS.n815 VSS.n814 9.3005
R1969 VSS.n1221 VSS.n1208 9.3005
R1970 VSS.n1217 VSS.n1208 9.3005
R1971 VSS.n1234 VSS.n1233 9.3005
R1972 VSS.n1236 VSS.n1235 9.3005
R1973 VSS.n1237 VSS.n1204 9.3005
R1974 VSS.n1241 VSS.n1240 9.3005
R1975 VSS.n1244 VSS.n1243 9.3005
R1976 VSS.n1246 VSS.n1201 9.3005
R1977 VSS.n1248 VSS.n1247 9.3005
R1978 VSS.n1261 VSS.n1260 9.3005
R1979 VSS.n1263 VSS.n1262 9.3005
R1980 VSS.n1265 VSS.n1264 9.3005
R1981 VSS.n1266 VSS.n1192 9.3005
R1982 VSS.n1269 VSS.n1268 9.3005
R1983 VSS.n1270 VSS.n1191 9.3005
R1984 VSS.n1272 VSS.n1271 9.3005
R1985 VSS.n1273 VSS.n1190 9.3005
R1986 VSS.n1276 VSS.n1275 9.3005
R1987 VSS.n1331 VSS.n1330 9.3005
R1988 VSS.n1329 VSS.n1189 9.3005
R1989 VSS.n1328 VSS.n1327 9.3005
R1990 VSS.n1327 VSS.n1326 9.3005
R1991 VSS.n1290 VSS.n1281 9.3005
R1992 VSS.n1290 VSS.n1289 9.3005
R1993 VSS.n1317 VSS.n1316 9.3005
R1994 VSS.n1314 VSS.n1286 9.3005
R1995 VSS.n1313 VSS.n1312 9.3005
R1996 VSS.n1311 VSS.n1292 9.3005
R1997 VSS.n1310 VSS.n1309 9.3005
R1998 VSS.n1308 VSS.n1293 9.3005
R1999 VSS.n1306 VSS.n1305 9.3005
R2000 VSS.n1304 VSS.n1294 9.3005
R2001 VSS.n1303 VSS.n1302 9.3005
R2002 VSS.n1300 VSS.n1295 9.3005
R2003 VSS.n2140 VSS.n2139 9.3005
R2004 VSS.n2148 VSS.n890 9.3005
R2005 VSS.n2153 VSS.n888 9.3005
R2006 VSS.n2192 VSS.n2191 9.3005
R2007 VSS.n2202 VSS.n2201 9.3005
R2008 VSS.n2204 VSS.n865 9.3005
R2009 VSS.n2212 VSS.n2211 9.3005
R2010 VSS.n2218 VSS.n2217 9.3005
R2011 VSS.n2222 VSS.n2221 9.3005
R2012 VSS.n857 VSS.n856 9.3005
R2013 VSS.n2231 VSS.n2230 9.3005
R2014 VSS.n2233 VSS.n854 9.3005
R2015 VSS.n2236 VSS.n2235 9.3005
R2016 VSS.n2238 VSS.n2237 9.3005
R2017 VSS.n2239 VSS.n850 9.3005
R2018 VSS.n2242 VSS.n2241 9.3005
R2019 VSS.n2244 VSS.n2243 9.3005
R2020 VSS.n2247 VSS.n848 9.3005
R2021 VSS.n2252 VSS.n2251 9.3005
R2022 VSS.n2253 VSS.n847 9.3005
R2023 VSS.n2255 VSS.n2254 9.3005
R2024 VSS.n2256 VSS.n843 9.3005
R2025 VSS.n2287 VSS.n2286 9.3005
R2026 VSS.n2285 VSS.n2284 9.3005
R2027 VSS.n2277 VSS.n2276 9.3005
R2028 VSS.n2274 VSS.n2273 9.3005
R2029 VSS.n2272 VSS.n2271 9.3005
R2030 VSS.n2270 VSS.n2261 9.3005
R2031 VSS.n2267 VSS.n2266 9.3005
R2032 VSS.n2206 VSS.n2205 9.3005
R2033 VSS.n2203 VSS.n866 9.3005
R2034 VSS.n2197 VSS.n867 9.3005
R2035 VSS.n2196 VSS.n2195 9.3005
R2036 VSS.n2194 VSS.n2193 9.3005
R2037 VSS.n2190 VSS.n869 9.3005
R2038 VSS.n2189 VSS.n2188 9.3005
R2039 VSS.n2187 VSS.n871 9.3005
R2040 VSS.n2184 VSS.n2183 9.3005
R2041 VSS.n2173 VSS.n873 9.3005
R2042 VSS.n2169 VSS.n2168 9.3005
R2043 VSS.n2166 VSS.n880 9.3005
R2044 VSS.n2164 VSS.n2163 9.3005
R2045 VSS.n2162 VSS.n882 9.3005
R2046 VSS.n2161 VSS.n2160 9.3005
R2047 VSS.n2158 VSS.n883 9.3005
R2048 VSS.n2157 VSS.n2156 9.3005
R2049 VSS.n2155 VSS.n2154 9.3005
R2050 VSS.n2150 VSS.n2149 9.3005
R2051 VSS.n2147 VSS.n2146 9.3005
R2052 VSS.n2141 VSS.n892 9.3005
R2053 VSS.n1180 VSS.n893 9.3005
R2054 VSS.n1388 VSS.n1387 9.3005
R2055 VSS.n1387 VSS.n1385 9.3005
R2056 VSS.n1380 VSS.n1137 9.3005
R2057 VSS.n1379 VSS.n1378 9.3005
R2058 VSS.n1376 VSS.n1375 9.3005
R2059 VSS.n1374 VSS.n1373 9.3005
R2060 VSS.n1372 VSS.n1143 9.3005
R2061 VSS.n1371 VSS.n1370 9.3005
R2062 VSS.n1369 VSS.n1368 9.3005
R2063 VSS.n1367 VSS.n1366 9.3005
R2064 VSS.n1365 VSS.n1146 9.3005
R2065 VSS.n1364 VSS.n1363 9.3005
R2066 VSS.n1361 VSS.n1360 9.3005
R2067 VSS.n1359 VSS.n1147 9.3005
R2068 VSS.n1159 VSS.n1148 9.3005
R2069 VSS.n1168 VSS.n1167 9.3005
R2070 VSS.n1185 VSS.n1184 9.3005
R2071 VSS.n1187 VSS.n1186 9.3005
R2072 VSS.n1337 VSS.n1178 9.3005
R2073 VSS.n1339 VSS.n1338 9.3005
R2074 VSS.n1340 VSS.n1176 9.3005
R2075 VSS.n1342 VSS.n1341 9.3005
R2076 VSS.n1343 VSS.n1173 9.3005
R2077 VSS.n1345 VSS.n1344 9.3005
R2078 VSS.n1346 VSS.n1172 9.3005
R2079 VSS.n1348 VSS.n1347 9.3005
R2080 VSS.n1350 VSS.n1349 9.3005
R2081 VSS.n1169 VSS.n1156 9.3005
R2082 VSS.n1620 VSS.n1619 9.3005
R2083 VSS.n1619 VSS.n1401 9.3005
R2084 VSS.n1618 VSS.n1617 9.3005
R2085 VSS.n1616 VSS.n1615 9.3005
R2086 VSS.n1610 VSS.n1609 9.3005
R2087 VSS.n1608 VSS.n1412 9.3005
R2088 VSS.n1606 VSS.n1605 9.3005
R2089 VSS.n1604 VSS.n1603 9.3005
R2090 VSS.n1416 VSS.n1415 9.3005
R2091 VSS.n1597 VSS.n1596 9.3005
R2092 VSS.n1595 VSS.n1418 9.3005
R2093 VSS.n1594 VSS.n1593 9.3005
R2094 VSS.n1591 VSS.n1590 9.3005
R2095 VSS.n1432 VSS.n1431 9.3005
R2096 VSS.n1434 VSS.n1428 9.3005
R2097 VSS.n1580 VSS.n1579 9.3005
R2098 VSS.n1577 VSS.n1429 9.3005
R2099 VSS.n1575 VSS.n1574 9.3005
R2100 VSS.n1573 VSS.n1572 9.3005
R2101 VSS.n1570 VSS.n1438 9.3005
R2102 VSS.n1567 VSS.n1566 9.3005
R2103 VSS.n1565 VSS.n1564 9.3005
R2104 VSS.n1560 VSS.n1441 9.3005
R2105 VSS.n1559 VSS.n1558 9.3005
R2106 VSS.n1557 VSS.n1556 9.3005
R2107 VSS.n1555 VSS.n1446 9.3005
R2108 VSS.n1552 VSS.n1551 9.3005
R2109 VSS.n1451 VSS.n1449 9.3005
R2110 VSS.n1462 VSS.n1458 9.3005
R2111 VSS.n1541 VSS.n1540 9.3005
R2112 VSS.n1539 VSS.n1538 9.3005
R2113 VSS.n1537 VSS.n1463 9.3005
R2114 VSS.n1536 VSS.n1535 9.3005
R2115 VSS.n1534 VSS.n1464 9.3005
R2116 VSS.n1533 VSS.n1532 9.3005
R2117 VSS.n1531 VSS.n1468 9.3005
R2118 VSS.n1530 VSS.n1529 9.3005
R2119 VSS.n1528 VSS.n1469 9.3005
R2120 VSS.n1527 VSS.n1471 9.3005
R2121 VSS.n1526 VSS.n1525 9.3005
R2122 VSS.n1524 VSS.n1523 9.3005
R2123 VSS.n1522 VSS.n1476 9.3005
R2124 VSS.n1521 VSS.n1520 9.3005
R2125 VSS.n1505 VSS.n1477 9.3005
R2126 VSS.n1504 VSS.n1503 9.3005
R2127 VSS.n1502 VSS.n1479 9.3005
R2128 VSS.n1501 VSS.n1500 9.3005
R2129 VSS.n1498 VSS.n1497 9.3005
R2130 VSS.n1495 VSS.n1494 9.3005
R2131 VSS.n1493 VSS.n1489 9.3005
R2132 VSS.n1492 VSS.n1491 9.3005
R2133 VSS.n1490 VSS.n911 9.3005
R2134 VSS.n915 VSS.n912 9.3005
R2135 VSS.n2115 VSS.n2114 9.3005
R2136 VSS.n2113 VSS.n2112 9.3005
R2137 VSS.n2111 VSS.n916 9.3005
R2138 VSS.n2110 VSS.n2109 9.3005
R2139 VSS.n2108 VSS.n917 9.3005
R2140 VSS.n2107 VSS.n2106 9.3005
R2141 VSS.n2105 VSS.n921 9.3005
R2142 VSS.n2104 VSS.n2103 9.3005
R2143 VSS.n2102 VSS.n922 9.3005
R2144 VSS.n2100 VSS.n2099 9.3005
R2145 VSS.n2098 VSS.n2097 9.3005
R2146 VSS.n2096 VSS.n926 9.3005
R2147 VSS.n2095 VSS.n2094 9.3005
R2148 VSS.n929 VSS.n927 9.3005
R2149 VSS.n941 VSS.n937 9.3005
R2150 VSS.n957 VSS.n956 9.3005
R2151 VSS.n954 VSS.n938 9.3005
R2152 VSS.n952 VSS.n946 9.3005
R2153 VSS.n1641 VSS.n1127 9.3005
R2154 VSS.n1641 VSS.n1126 9.3005
R2155 VSS.n1643 VSS.n1642 9.3005
R2156 VSS.n1645 VSS.n1644 9.3005
R2157 VSS.n1649 VSS.n1648 9.3005
R2158 VSS.n1651 VSS.n1650 9.3005
R2159 VSS.n1652 VSS.n1120 9.3005
R2160 VSS.n1654 VSS.n1653 9.3005
R2161 VSS.n1656 VSS.n1655 9.3005
R2162 VSS.n1657 VSS.n1117 9.3005
R2163 VSS.n1658 VSS.n1116 9.3005
R2164 VSS.n1660 VSS.n1659 9.3005
R2165 VSS.n1661 VSS.n1115 9.3005
R2166 VSS.n1663 VSS.n1662 9.3005
R2167 VSS.n1664 VSS.n1089 9.3005
R2168 VSS.n1665 VSS.n1090 9.3005
R2169 VSS.n1667 VSS.n1666 9.3005
R2170 VSS.n1112 VSS.n1111 9.3005
R2171 VSS.n1110 VSS.n1093 9.3005
R2172 VSS.n1109 VSS.n1108 9.3005
R2173 VSS.n1934 VSS.n1027 9.3005
R2174 VSS.n1936 VSS.n1935 9.3005
R2175 VSS.n1937 VSS.n1022 9.3005
R2176 VSS.n1939 VSS.n1938 9.3005
R2177 VSS.n1015 VSS.n1014 9.3005
R2178 VSS.n1949 VSS.n1948 9.3005
R2179 VSS.n1951 VSS.n1012 9.3005
R2180 VSS.n1953 VSS.n1952 9.3005
R2181 VSS.n1954 VSS.n1011 9.3005
R2182 VSS.n1956 VSS.n1955 9.3005
R2183 VSS.n1958 VSS.n1008 9.3005
R2184 VSS.n1962 VSS.n1961 9.3005
R2185 VSS.n1963 VSS.n1007 9.3005
R2186 VSS.n1965 VSS.n1964 9.3005
R2187 VSS.n1966 VSS.n1006 9.3005
R2188 VSS.n1968 VSS.n1967 9.3005
R2189 VSS.n1970 VSS.n1969 9.3005
R2190 VSS.n1973 VSS.n1972 9.3005
R2191 VSS.n1984 VSS.n1983 9.3005
R2192 VSS.n1985 VSS.n991 9.3005
R2193 VSS.n1987 VSS.n1986 9.3005
R2194 VSS.n1989 VSS.n1988 9.3005
R2195 VSS.n1990 VSS.n989 9.3005
R2196 VSS.n1992 VSS.n1991 9.3005
R2197 VSS.n1994 VSS.n1993 9.3005
R2198 VSS.n1995 VSS.n985 9.3005
R2199 VSS.n1997 VSS.n1996 9.3005
R2200 VSS.n1998 VSS.n984 9.3005
R2201 VSS.n2000 VSS.n1999 9.3005
R2202 VSS.n2005 VSS.n2004 9.3005
R2203 VSS.n2006 VSS.n983 9.3005
R2204 VSS.n2012 VSS.n2011 9.3005
R2205 VSS.n2016 VSS.n2015 9.3005
R2206 VSS.n2025 VSS.n2024 9.3005
R2207 VSS.n2026 VSS.n975 9.3005
R2208 VSS.n2030 VSS.n2029 9.3005
R2209 VSS.n2031 VSS.n974 9.3005
R2210 VSS.n2033 VSS.n2032 9.3005
R2211 VSS.n2034 VSS.n973 9.3005
R2212 VSS.n2039 VSS.n2038 9.3005
R2213 VSS.n2040 VSS.n972 9.3005
R2214 VSS.n2042 VSS.n2041 9.3005
R2215 VSS.n2043 VSS.n971 9.3005
R2216 VSS.n2048 VSS.n2047 9.3005
R2217 VSS.n2050 VSS.n2049 9.3005
R2218 VSS.n2052 VSS.n966 9.3005
R2219 VSS.n2082 VSS.n2081 9.3005
R2220 VSS.n2080 VSS.n2079 9.3005
R2221 VSS.n2072 VSS.n2071 9.3005
R2222 VSS.n2070 VSS.n2057 9.3005
R2223 VSS.n2069 VSS.n2068 9.3005
R2224 VSS.n2067 VSS.n2066 9.3005
R2225 VSS.n2064 VSS.n2059 9.3005
R2226 VSS.n1107 VSS.n1094 9.3005
R2227 VSS.n1106 VSS.n1105 9.3005
R2228 VSS.n1104 VSS.n1096 9.3005
R2229 VSS.n1103 VSS.n1102 9.3005
R2230 VSS.n1097 VSS.n1028 9.3005
R2231 VSS.n1933 VSS.n1932 9.3005
R2232 VSS.n1814 VSS.n1813 9.3005
R2233 VSS.n1816 VSS.n1815 9.3005
R2234 VSS.n1708 VSS.n1707 9.3005
R2235 VSS.n1719 VSS.n1718 9.3005
R2236 VSS.n1721 VSS.n1720 9.3005
R2237 VSS.n1722 VSS.n1695 9.3005
R2238 VSS.n1724 VSS.n1723 9.3005
R2239 VSS.n1725 VSS.n1692 9.3005
R2240 VSS.n1727 VSS.n1726 9.3005
R2241 VSS.n1728 VSS.n1691 9.3005
R2242 VSS.n1730 VSS.n1729 9.3005
R2243 VSS.n1732 VSS.n1690 9.3005
R2244 VSS.n1736 VSS.n1735 9.3005
R2245 VSS.n1737 VSS.n1689 9.3005
R2246 VSS.n1739 VSS.n1738 9.3005
R2247 VSS.n1740 VSS.n1688 9.3005
R2248 VSS.n1741 VSS.n1683 9.3005
R2249 VSS.n1742 VSS.n1684 9.3005
R2250 VSS.n1759 VSS.n1758 9.3005
R2251 VSS.n1756 VSS.n1755 9.3005
R2252 VSS.n1754 VSS.n1743 9.3005
R2253 VSS.n1752 VSS.n1751 9.3005
R2254 VSS.n1750 VSS.n1749 9.3005
R2255 VSS.n1748 VSS.n1031 9.3005
R2256 VSS.n1927 VSS.n1926 9.3005
R2257 VSS.n1925 VSS.n1032 9.3005
R2258 VSS.n1924 VSS.n1923 9.3005
R2259 VSS.n1922 VSS.n1921 9.3005
R2260 VSS.n1910 VSS.n1037 9.3005
R2261 VSS.n1910 VSS.n1045 9.3005
R2262 VSS.n1911 VSS.n1910 9.3005
R2263 VSS.n1909 VSS.n1908 9.3005
R2264 VSS.n1907 VSS.n1047 9.3005
R2265 VSS.n1906 VSS.n1905 9.3005
R2266 VSS.n1904 VSS.n1903 9.3005
R2267 VSS.n1902 VSS.n1048 9.3005
R2268 VSS.n1901 VSS.n1900 9.3005
R2269 VSS.n1899 VSS.n1049 9.3005
R2270 VSS.n1896 VSS.n1895 9.3005
R2271 VSS.n1060 VSS.n1054 9.3005
R2272 VSS.n1067 VSS.n1066 9.3005
R2273 VSS.n1887 VSS.n1886 9.3005
R2274 VSS.n1885 VSS.n1884 9.3005
R2275 VSS.n1883 VSS.n1882 9.3005
R2276 VSS.n1881 VSS.n1069 9.3005
R2277 VSS.n1878 VSS.n1877 9.3005
R2278 VSS.n1876 VSS.n1070 9.3005
R2279 VSS.n1875 VSS.n1874 9.3005
R2280 VSS.n1873 VSS.n1071 9.3005
R2281 VSS.n1872 VSS.n1074 9.3005
R2282 VSS.n1871 VSS.n1870 9.3005
R2283 VSS.n1869 VSS.n1868 9.3005
R2284 VSS.n1867 VSS.n1076 9.3005
R2285 VSS.n1866 VSS.n1865 9.3005
R2286 VSS.n1780 VSS.n1077 9.3005
R2287 VSS.n1849 VSS.n1782 9.3005
R2288 VSS.n1855 VSS.n1854 9.3005
R2289 VSS.n1847 VSS.n1783 9.3005
R2290 VSS.n1846 VSS.n1845 9.3005
R2291 VSS.n1844 VSS.n1786 9.3005
R2292 VSS.n1843 VSS.n1842 9.3005
R2293 VSS.n1841 VSS.n1840 9.3005
R2294 VSS.n1839 VSS.n1787 9.3005
R2295 VSS.n1838 VSS.n1837 9.3005
R2296 VSS.n1836 VSS.n1788 9.3005
R2297 VSS.n1834 VSS.n1791 9.3005
R2298 VSS.n1833 VSS.n1832 9.3005
R2299 VSS.n1805 VSS.n1794 9.3005
R2300 VSS.n1824 VSS.n1823 9.3005
R2301 VSS.n1822 VSS.n1821 9.3005
R2302 VSS.n1820 VSS.n1806 9.3005
R2303 VSS.n1819 VSS.n1818 9.3005
R2304 VSS.n1817 VSS.n1807 9.3005
R2305 VSS.n2603 VSS.n2602 9.3005
R2306 VSS.n2606 VSS.n2597 9.3005
R2307 VSS.n2608 VSS.n2607 9.3005
R2308 VSS.n2610 VSS.n2609 9.3005
R2309 VSS.n2613 VSS.n2612 9.3005
R2310 VSS.n2595 VSS.n2590 9.3005
R2311 VSS.n2593 VSS.n2589 9.3005
R2312 VSS.n2584 VSS.n2583 9.3005
R2313 VSS.n2628 VSS.n2627 9.3005
R2314 VSS.n2629 VSS.n2581 9.3005
R2315 VSS.n2631 VSS.n2630 9.3005
R2316 VSS.n2633 VSS.n2632 9.3005
R2317 VSS.n2470 VSS.n2469 9.3005
R2318 VSS.n2469 VSS.n2467 9.3005
R2319 VSS.n2505 VSS.n2504 9.3005
R2320 VSS.n2506 VSS.n2505 9.3005
R2321 VSS.n2515 VSS.n250 9.3005
R2322 VSS.n2515 VSS.n2514 9.3005
R2323 VSS.n2517 VSS.n249 9.3005
R2324 VSS.n2520 VSS.n2519 9.3005
R2325 VSS.n2521 VSS.n248 9.3005
R2326 VSS.n2523 VSS.n2522 9.3005
R2327 VSS.n2524 VSS.n247 9.3005
R2328 VSS.n2526 VSS.n2525 9.3005
R2329 VSS.n2528 VSS.n2527 9.3005
R2330 VSS.n2529 VSS.n245 9.3005
R2331 VSS.n2532 VSS.n2531 9.3005
R2332 VSS.n2534 VSS.n2533 9.3005
R2333 VSS.n2542 VSS.n2541 9.3005
R2334 VSS.n2539 VSS.n2538 9.3005
R2335 VSS.n2551 VSS.n231 9.3005
R2336 VSS.n2553 VSS.n2552 9.3005
R2337 VSS.n2554 VSS.n230 9.3005
R2338 VSS.n2556 VSS.n2555 9.3005
R2339 VSS.n2558 VSS.n2557 9.3005
R2340 VSS.n2559 VSS.n228 9.3005
R2341 VSS.n2562 VSS.n2561 9.3005
R2342 VSS.n2564 VSS.n2563 9.3005
R2343 VSS.n2566 VSS.n2565 9.3005
R2344 VSS.n2568 VSS.n2567 9.3005
R2345 VSS.n2570 VSS.n2569 9.3005
R2346 VSS.n2572 VSS.n2571 9.3005
R2347 VSS.n2573 VSS.n220 9.3005
R2348 VSS.n2574 VSS.n221 9.3005
R2349 VSS.n2648 VSS.n2647 9.3005
R2350 VSS.n2646 VSS.n2645 9.3005
R2351 VSS.n2644 VSS.n2575 9.3005
R2352 VSS.n2643 VSS.n2642 9.3005
R2353 VSS.n2640 VSS.n2576 9.3005
R2354 VSS.n2639 VSS.n2638 9.3005
R2355 VSS.n2637 VSS.n2577 9.3005
R2356 VSS.n2636 VSS.n2635 9.3005
R2357 VSS.n2461 VSS.n2460 9.3005
R2358 VSS.n2458 VSS.n2403 9.3005
R2359 VSS.n2457 VSS.n2456 9.3005
R2360 VSS.n2455 VSS.n2404 9.3005
R2361 VSS.n2453 VSS.n2452 9.3005
R2362 VSS.n2450 VSS.n2449 9.3005
R2363 VSS.n2416 VSS.n2410 9.3005
R2364 VSS.n2421 VSS.n2418 9.3005
R2365 VSS.n2439 VSS.n2438 9.3005
R2366 VSS.n2436 VSS.n2419 9.3005
R2367 VSS.n2435 VSS.n2434 9.3005
R2368 VSS.n2433 VSS.n2422 9.3005
R2369 VSS.n2432 VSS.n2431 9.3005
R2370 VSS.n2430 VSS.n2423 9.3005
R2371 VSS.n2429 VSS.n2428 9.3005
R2372 VSS.n2427 VSS.n2426 9.3005
R2373 VSS.n2501 VSS.n266 9.3005
R2374 VSS.n2503 VSS.n2502 9.3005
R2375 VSS.n2871 VSS.n2870 9.3005
R2376 VSS.n19 VSS.n1 9.3005
R2377 VSS.n2861 VSS.n6 9.3005
R2378 VSS.n2860 VSS.n2859 9.3005
R2379 VSS.n63 VSS.n62 9.3005
R2380 VSS.n61 VSS.n9 9.3005
R2381 VSS.n60 VSS.n59 9.3005
R2382 VSS.n58 VSS.n10 9.3005
R2383 VSS.n57 VSS.n11 9.3005
R2384 VSS.n56 VSS.n55 9.3005
R2385 VSS.n54 VSS.n12 9.3005
R2386 VSS.n53 VSS.n52 9.3005
R2387 VSS.n51 VSS.n50 9.3005
R2388 VSS.n49 VSS.n13 9.3005
R2389 VSS.n48 VSS.n47 9.3005
R2390 VSS.n46 VSS.n45 9.3005
R2391 VSS.n44 VSS.n14 9.3005
R2392 VSS.n43 VSS.n42 9.3005
R2393 VSS.n41 VSS.n40 9.3005
R2394 VSS.n39 VSS.n15 9.3005
R2395 VSS.n38 VSS.n37 9.3005
R2396 VSS.n36 VSS.n35 9.3005
R2397 VSS.n34 VSS.n16 9.3005
R2398 VSS.n33 VSS.n32 9.3005
R2399 VSS.n31 VSS.n30 9.3005
R2400 VSS.n29 VSS.n17 9.3005
R2401 VSS.n28 VSS.n27 9.3005
R2402 VSS.n26 VSS.n25 9.3005
R2403 VSS.n24 VSS.n18 9.3005
R2404 VSS.n23 VSS.n22 9.3005
R2405 VSS.n21 VSS.n20 9.3005
R2406 VSS.n2863 VSS.n2862 9.3005
R2407 VSS.n87 VSS.n86 9.3005
R2408 VSS.n89 VSS.n81 9.3005
R2409 VSS.n92 VSS.n91 9.3005
R2410 VSS.n2710 VSS.n2709 9.3005
R2411 VSS.n2708 VSS.n102 9.3005
R2412 VSS.n2706 VSS.n2705 9.3005
R2413 VSS.n2704 VSS.n66 9.3005
R2414 VSS.n2854 VSS.n67 9.3005
R2415 VSS.n2852 VSS.n2851 9.3005
R2416 VSS.n2850 VSS.n2849 9.3005
R2417 VSS.n2846 VSS.n69 9.3005
R2418 VSS.n2845 VSS.n71 9.3005
R2419 VSS.n2844 VSS.n72 9.3005
R2420 VSS.n2843 VSS.n2842 9.3005
R2421 VSS.n2841 VSS.n74 9.3005
R2422 VSS.n2840 VSS.n2839 9.3005
R2423 VSS.n2838 VSS.n76 9.3005
R2424 VSS.n2837 VSS.n77 9.3005
R2425 VSS.n2836 VSS.n78 9.3005
R2426 VSS.n2835 VSS.n2834 9.3005
R2427 VSS.n93 VSS.n80 9.3005
R2428 VSS.n2831 VSS.n2830 9.3005
R2429 VSS.n2824 VSS.n2823 9.3005
R2430 VSS.n2826 VSS.n2825 9.3005
R2431 VSS.n2828 VSS.n2827 9.3005
R2432 VSS.n2829 VSS.n94 9.3005
R2433 VSS.n2714 VSS.n2713 9.3005
R2434 VSS.n2715 VSS.n100 9.3005
R2435 VSS.n2815 VSS.n2814 9.3005
R2436 VSS.n2813 VSS.n2718 9.3005
R2437 VSS.n2812 VSS.n2811 9.3005
R2438 VSS.n2810 VSS.n2719 9.3005
R2439 VSS.n2809 VSS.n2808 9.3005
R2440 VSS.n2807 VSS.n2720 9.3005
R2441 VSS.n2806 VSS.n2721 9.3005
R2442 VSS.n2805 VSS.n2793 9.3005
R2443 VSS.n2804 VSS.n2794 9.3005
R2444 VSS.n2803 VSS.n2802 9.3005
R2445 VSS.n2801 VSS.n2795 9.3005
R2446 VSS.n2800 VSS.n2799 9.3005
R2447 VSS.n2798 VSS.n2797 9.3005
R2448 VSS.n2796 VSS.n97 9.3005
R2449 VSS.n306 VSS.n305 9.3005
R2450 VSS.n308 VSS.n286 9.3005
R2451 VSS.n455 VSS.n454 9.3005
R2452 VSS.n452 VSS.n285 9.3005
R2453 VSS.n449 VSS.n448 9.3005
R2454 VSS.n447 VSS.n287 9.3005
R2455 VSS.n446 VSS.n445 9.3005
R2456 VSS.n444 VSS.n288 9.3005
R2457 VSS.n443 VSS.n442 9.3005
R2458 VSS.n441 VSS.n290 9.3005
R2459 VSS.n440 VSS.n439 9.3005
R2460 VSS.n293 VSS.n291 9.3005
R2461 VSS.n434 VSS.n433 9.3005
R2462 VSS.n432 VSS.n295 9.3005
R2463 VSS.n421 VSS.n296 9.3005
R2464 VSS.n424 VSS.n423 9.3005
R2465 VSS.n422 VSS.n275 9.3005
R2466 VSS.n2484 VSS.n274 9.3005
R2467 VSS.n2486 VSS.n2485 9.3005
R2468 VSS.n2487 VSS.n273 9.3005
R2469 VSS.n2489 VSS.n2488 9.3005
R2470 VSS.n2491 VSS.n2490 9.3005
R2471 VSS.n2492 VSS.n271 9.3005
R2472 VSS.n2494 VSS.n2493 9.3005
R2473 VSS.n2496 VSS.n2495 9.3005
R2474 VSS.n2497 VSS.n269 9.3005
R2475 VSS.n324 VSS.n268 9.3005
R2476 VSS.n329 VSS.n328 9.3005
R2477 VSS.n331 VSS.n321 9.3005
R2478 VSS.n339 VSS.n338 9.3005
R2479 VSS.n341 VSS.n319 9.3005
R2480 VSS.n404 VSS.n403 9.3005
R2481 VSS.n402 VSS.n320 9.3005
R2482 VSS.n401 VSS.n400 9.3005
R2483 VSS.n399 VSS.n342 9.3005
R2484 VSS.n398 VSS.n397 9.3005
R2485 VSS.n396 VSS.n343 9.3005
R2486 VSS.n394 VSS.n393 9.3005
R2487 VSS.n392 VSS.n344 9.3005
R2488 VSS.n391 VSS.n390 9.3005
R2489 VSS.n388 VSS 9.3005
R2490 VSS.n387 VSS.n386 9.3005
R2491 VSS.n385 VSS.n384 9.3005
R2492 VSS.n383 VSS.n382 9.3005
R2493 VSS.n349 VSS.n347 9.3005
R2494 VSS.n374 VSS.n373 9.3005
R2495 VSS.n372 VSS.n358 9.3005
R2496 VSS.n371 VSS.n370 9.3005
R2497 VSS.n369 VSS.n359 9.3005
R2498 VSS.n368 VSS.n367 9.3005
R2499 VSS.n366 VSS.n360 9.3005
R2500 VSS.n365 VSS.n364 9.3005
R2501 VSS.n363 VSS.n124 9.3005
R2502 VSS.n2681 VSS.n2680 9.3005
R2503 VSS.n2679 VSS.n123 9.3005
R2504 VSS.n2678 VSS.n2677 9.3005
R2505 VSS.n2676 VSS.n2675 9.3005
R2506 VSS.n151 VSS.n126 9.3005
R2507 VSS.n153 VSS.n152 9.3005
R2508 VSS.n156 VSS.n147 9.3005
R2509 VSS.n159 VSS.n158 9.3005
R2510 VSS.n160 VSS.n145 9.3005
R2511 VSS.n166 VSS.n165 9.3005
R2512 VSS.n168 VSS.n167 9.3005
R2513 VSS.n170 VSS.n169 9.3005
R2514 VSS.n171 VSS.n143 9.3005
R2515 VSS.n173 VSS.n172 9.3005
R2516 VSS.n174 VSS.n141 9.3005
R2517 VSS.n177 VSS.n176 9.3005
R2518 VSS.n178 VSS.n140 9.3005
R2519 VSS.n180 VSS.n179 9.3005
R2520 VSS.n181 VSS.n137 9.3005
R2521 VSS.n208 VSS.n207 9.3005
R2522 VSS.n206 VSS.n205 9.3005
R2523 VSS.n203 VSS.n182 9.3005
R2524 VSS.n202 VSS.n201 9.3005
R2525 VSS.n200 VSS.n185 9.3005
R2526 VSS.n199 VSS.n198 9.3005
R2527 VSS.n197 VSS.n196 9.3005
R2528 VSS.n195 VSS.n194 9.3005
R2529 VSS.n193 VSS.n192 9.3005
R2530 VSS.n2193 VSS.n2192 9.12791
R2531 VSS.n2154 VSS.n887 9.03579
R2532 VSS.n2152 VSS.n2151 9.03579
R2533 VSS.n1572 VSS.n1437 9.03579
R2534 VSS.n2247 VSS.n2246 8.9684
R2535 VSS.n2773 VSS.n2772 8.44328
R2536 VSS.t234 VSS.t887 8.42962
R2537 VSS.t879 VSS.t45 8.42962
R2538 VSS.t494 VSS.t290 8.42962
R2539 VSS.n2734 VSS.n2733 8.33966
R2540 VSS.n2109 VSS.n919 8.28285
R2541 VSS.n176 VSS.n140 8.23546
R2542 VSS.n180 VSS.n140 8.23546
R2543 VSS.n181 VSS.n180 8.23546
R2544 VSS.n207 VSS.n181 8.23546
R2545 VSS.n207 VSS.n206 8.23546
R2546 VSS.n206 VSS.n182 8.23546
R2547 VSS.n201 VSS.n200 8.23546
R2548 VSS.n200 VSS.n199 8.23546
R2549 VSS.n384 VSS.n383 8.23546
R2550 VSS.n383 VSS.n347 8.23546
R2551 VSS.n373 VSS.n347 8.23546
R2552 VSS.n373 VSS.n372 8.23546
R2553 VSS.n372 VSS.n371 8.23546
R2554 VSS.n371 VSS.n359 8.23546
R2555 VSS.n367 VSS.n366 8.23546
R2556 VSS.n366 VSS.n365 8.23546
R2557 VSS.n403 VSS.n341 8.23546
R2558 VSS.n403 VSS.n402 8.23546
R2559 VSS.n402 VSS.n401 8.23546
R2560 VSS.n401 VSS.n342 8.23546
R2561 VSS.n397 VSS.n342 8.23546
R2562 VSS.n397 VSS.n396 8.23546
R2563 VSS.n394 VSS.n344 8.23546
R2564 VSS.n390 VSS.n344 8.23546
R2565 VSS.n798 VSS.n764 8.23546
R2566 VSS.n802 VSS.n764 8.23546
R2567 VSS.n774 VSS.n770 8.23546
R2568 VSS.n781 VSS.n770 8.23546
R2569 VSS.n789 VSS.n768 8.23546
R2570 VSS.n792 VSS.n789 8.23546
R2571 VSS.n1331 VSS.n1189 8.23546
R2572 VSS.n2255 VSS.n847 8.23546
R2573 VSS.n2256 VSS.n2255 8.23546
R2574 VSS.n2286 VSS.n2285 8.23546
R2575 VSS.n2221 VSS.n2218 8.23546
R2576 VSS.n2231 VSS.n856 8.23546
R2577 VSS.n2235 VSS.n2233 8.23546
R2578 VSS.n2239 VSS.n2238 8.23546
R2579 VSS.n1367 VSS.n1146 8.23546
R2580 VSS.n1363 VSS.n1146 8.23546
R2581 VSS.n1361 VSS.n1147 8.23546
R2582 VSS.n1349 VSS.n1348 8.23546
R2583 VSS.n1348 VSS.n1172 8.23546
R2584 VSS.n1344 VSS.n1343 8.23546
R2585 VSS.n1343 VSS.n1342 8.23546
R2586 VSS.n1342 VSS.n1176 8.23546
R2587 VSS.n1338 VSS.n1337 8.23546
R2588 VSS.n1337 VSS.n1187 8.23546
R2589 VSS.n1961 VSS.n1007 8.23546
R2590 VSS.n1965 VSS.n1007 8.23546
R2591 VSS.n1966 VSS.n1965 8.23546
R2592 VSS.n1967 VSS.n1966 8.23546
R2593 VSS.n1972 VSS.n1970 8.23546
R2594 VSS.n1985 VSS.n1984 8.23546
R2595 VSS.n1986 VSS.n1985 8.23546
R2596 VSS.n2630 VSS.n2629 8.23546
R2597 VSS.n2629 VSS.n2628 8.23546
R2598 VSS.n2628 VSS.n2583 8.23546
R2599 VSS.n2612 VSS.n2595 8.23546
R2600 VSS.n2502 VSS.n2501 8.23546
R2601 VSS.n423 VSS.n421 8.23546
R2602 VSS.n423 VSS.n422 8.23546
R2603 VSS.n422 VSS.n274 8.23546
R2604 VSS.n2486 VSS.n274 8.23546
R2605 VSS.n2487 VSS.n2486 8.23546
R2606 VSS.n2488 VSS.n2487 8.23546
R2607 VSS.n2492 VSS.n2491 8.23546
R2608 VSS.n2493 VSS.n2492 8.23546
R2609 VSS.n783 VSS.n782 8.14595
R2610 VSS.n2593 VSS.n2592 8.05644
R2611 VSS.n2775 VSS.n2774 7.97888
R2612 VSS.n2773 VSS.n2735 7.97601
R2613 VSS.n2160 VSS.n2159 7.90638
R2614 VSS.n1526 VSS.n1474 7.90638
R2615 VSS.n2037 VSS.n972 7.90638
R2616 VSS.n1159 VSS.n1158 7.78791
R2617 VSS.n1959 VSS.n1010 7.72113
R2618 VSS.n176 VSS.n175 7.6984
R2619 VSS.n199 VSS.n187 7.6984
R2620 VSS.n384 VSS.n345 7.6984
R2621 VSS.n365 VSS.n362 7.6984
R2622 VSS.n341 VSS.n340 7.6984
R2623 VSS.n390 VSS.n389 7.6984
R2624 VSS.n798 VSS.n797 7.6984
R2625 VSS.n786 VSS.n784 7.6984
R2626 VSS.n2251 VSS.n2248 7.6984
R2627 VSS.n2211 VSS.n2210 7.6984
R2628 VSS.n2211 VSS.n864 7.6984
R2629 VSS.n2241 VSS.n849 7.6984
R2630 VSS.n1160 VSS.n1159 7.6984
R2631 VSS.n1187 VSS.n1179 7.6984
R2632 VSS.n1961 VSS.n1960 7.6984
R2633 VSS.n1986 VSS.n990 7.6984
R2634 VSS.n2565 VSS.n225 7.6984
R2635 VSS.n2630 VSS.n2582 7.6984
R2636 VSS.n421 VSS.n420 7.6984
R2637 VSS.n2493 VSS.n270 7.6984
R2638 VSS.n2053 VSS.n969 7.6005
R2639 VSS.n1344 VSS.n1175 7.51938
R2640 VSS.n792 VSS.n791 7.34036
R2641 VSS.n1970 VSS.n1005 7.34036
R2642 VSS.n2257 VSS.n2256 7.25085
R2643 VSS.n1171 VSS.n1170 7.25085
R2644 VSS.n2777 VSS.n2775 7.16724
R2645 VSS.n2749 VSS.n2735 7.16724
R2646 VSS.n2772 VSS.n2771 7.16724
R2647 VSS.n2733 VSS.n2725 7.16724
R2648 VSS.n2250 VSS.n847 7.16134
R2649 VSS.n2845 VSS.n2844 7.15344
R2650 VSS.n2311 VSS.n2310 7.11268
R2651 VSS.n2565 VSS.n2564 7.11268
R2652 VSS.n2594 VSS.n2593 6.98232
R2653 VSS.n803 VSS.n802 6.88949
R2654 VSS.n1368 VSS.n1367 6.88949
R2655 VSS.n2221 VSS.n2220 6.62428
R2656 VSS.n1290 VSS.n1280 6.61527
R2657 VSS.n2515 VSS.n252 6.61527
R2658 VSS.n108 VSS.t138 6.6005
R2659 VSS.n108 VSS.t227 6.6005
R2660 VSS.n110 VSS.t13 6.6005
R2661 VSS.n110 VSS.t225 6.6005
R2662 VSS.n105 VSS.t136 6.6005
R2663 VSS.n105 VSS.t932 6.6005
R2664 VSS.n1327 VSS.n1280 6.57117
R2665 VSS.n1612 VSS.n1411 6.57117
R2666 VSS.n1614 VSS.n1612 6.57117
R2667 VSS.n2505 VSS.n252 6.57117
R2668 VSS.n2285 VSS.n2258 6.53477
R2669 VSS.n2833 VSS.n2832 6.50373
R2670 VSS.n1994 VSS.n988 6.4005
R2671 VSS.n2014 VSS.n2012 6.4005
R2672 VSS.n2708 VSS.n2707 6.4005
R2673 VSS.n152 VSS.n151 6.26433
R2674 VSS.n152 VSS.n147 6.26433
R2675 VSS.n1756 VSS.n1743 6.26433
R2676 VSS.n1735 VSS.n1732 6.26433
R2677 VSS.n1923 VSS.n1922 6.26433
R2678 VSS.n1900 VSS.n1899 6.26433
R2679 VSS.n1882 VSS.n1881 6.26433
R2680 VSS.n2197 VSS.n2196 6.26433
R2681 VSS.n1609 VSS.n1608 6.26433
R2682 VSS.n1648 VSS.n1645 6.26433
R2683 VSS.n1868 VSS.n1867 6.26433
R2684 VSS.n1867 VSS.n1866 6.26433
R2685 VSS.n1837 VSS.n1836 6.26433
R2686 VSS.n2715 VSS.n2714 6.26433
R2687 VSS.n2825 VSS.n2824 6.26433
R2688 VSS.n445 VSS.n444 6.26433
R2689 VSS.n444 VSS.n443 6.26433
R2690 VSS.n955 VSS.n954 6.12816
R2691 VSS.n736 VSS.n735 6.06007
R2692 VSS.n645 VSS.n643 6.02861
R2693 VSS.n667 VSS.n600 6.02861
R2694 VSS.n2376 VSS.n2375 6.02861
R2695 VSS.n1262 VSS.n1261 6.02861
R2696 VSS.n2438 VSS.n2421 6.02861
R2697 VSS.n2157 VSS.n887 6.02403
R2698 VSS.n2145 VSS.n2144 6.02403
R2699 VSS.n192 VSS.n188 5.98311
R2700 VSS.n328 VSS.n325 5.98311
R2701 VSS.n1707 VSS.n1697 5.98311
R2702 VSS.n1564 VSS.n1440 5.98311
R2703 VSS.n2004 VSS.n2001 5.98311
R2704 VSS.n2047 VSS.n2044 5.98311
R2705 VSS.n1813 VSS.n1809 5.98311
R2706 VSS.n453 VSS.n452 5.98311
R2707 VSS.n305 VSS.n304 5.98311
R2708 VSS.n151 VSS.n125 5.85582
R2709 VSS.n1757 VSS.n1756 5.85582
R2710 VSS.n1732 VSS.n1731 5.85582
R2711 VSS.n1923 VSS.n1034 5.85582
R2712 VSS.n1900 VSS.n1050 5.85582
R2713 VSS.n1882 VSS.n1068 5.85582
R2714 VSS.n737 VSS.n736 5.85582
R2715 VSS.n2196 VSS.n868 5.85582
R2716 VSS.n1615 VSS.n1403 5.85582
R2717 VSS.n956 VSS.n942 5.85582
R2718 VSS.n1645 VSS.n1123 5.85582
R2719 VSS.n2081 VSS.n2054 5.85582
R2720 VSS.n1868 VSS.n1075 5.85582
R2721 VSS.n1837 VSS.n1789 5.85582
R2722 VSS.n2714 VSS.n101 5.85582
R2723 VSS.n2825 VSS.n98 5.85582
R2724 VSS.n2853 VSS.n2852 5.85582
R2725 VSS.n2849 VSS.n68 5.85582
R2726 VSS.n90 VSS.n89 5.85582
R2727 VSS.n445 VSS.n289 5.85582
R2728 VSS.n159 VSS.n147 5.65809
R2729 VSS.n1866 VSS.n1077 5.65809
R2730 VSS.n443 VSS.n290 5.65809
R2731 VSS.n774 VSS.n552 5.63966
R2732 VSS.n2310 VSS.n550 5.63966
R2733 VSS.n1278 VSS.n1189 5.63966
R2734 VSS.n2502 VSS.n264 5.63966
R2735 VSS.n680 VSS.n595 5.5878
R2736 VSS.n2232 VSS.n2231 5.55015
R2737 VSS.n2360 VSS.n2359 5.48621
R2738 VSS.n632 VSS.n611 5.48128
R2739 VSS.n2081 VSS.n2080 5.37524
R2740 VSS.n1497 VSS.n1496 5.27109
R2741 VSS.n1607 VSS.n1606 5.24958
R2742 VSS.n478 VSS.n476 5.13108
R2743 VSS.n478 VSS.n477 5.13108
R2744 VSS.n730 VSS.n727 5.13108
R2745 VSS.n730 VSS.n729 5.13108
R2746 VSS.n500 VSS.n479 5.13108
R2747 VSS.n500 VSS.n499 5.13108
R2748 VSS.n813 VSS.n810 5.13108
R2749 VSS.n813 VSS.n812 5.13108
R2750 VSS.n1208 VSS.n1206 5.13108
R2751 VSS.n1208 VSS.n1207 5.13108
R2752 VSS.n1232 VSS.n1209 5.13108
R2753 VSS.n1232 VSS.n1231 5.13108
R2754 VSS.n1387 VSS.n1138 5.13108
R2755 VSS.n1387 VSS.n1386 5.13108
R2756 VSS.n2264 VSS.n2262 5.13108
R2757 VSS.n2264 VSS.n2263 5.13108
R2758 VSS.n1619 VSS.n1400 5.13108
R2759 VSS.n1619 VSS.n1402 5.13108
R2760 VSS.n951 VSS.n948 5.13108
R2761 VSS.n951 VSS.n949 5.13108
R2762 VSS.n1641 VSS.n1125 5.13108
R2763 VSS.n1641 VSS.n1128 5.13108
R2764 VSS.n2063 VSS.n2060 5.13108
R2765 VSS.n2063 VSS.n2061 5.13108
R2766 VSS.n2469 VSS.n2399 5.13108
R2767 VSS.n2469 VSS.n2468 5.13108
R2768 VSS.n2600 VSS.n2598 5.13108
R2769 VSS.n2600 VSS.n2599 5.13108
R2770 VSS.n2398 VSS.n2396 5.13108
R2771 VSS.n2398 VSS.n2397 5.13108
R2772 VSS.n2241 VSS.n2240 4.92358
R2773 VSS.n163 VSS.n162 4.85762
R2774 VSS.n437 VSS.n294 4.85762
R2775 VSS.n1852 VSS.n1851 4.85762
R2776 VSS.n626 VSS.n625 4.85762
R2777 VSS.n1600 VSS.n1417 4.85762
R2778 VSS.n192 VSS.n191 4.8005
R2779 VSS.n328 VSS.n327 4.8005
R2780 VSS.n1707 VSS.n1706 4.8005
R2781 VSS.n2004 VSS.n2003 4.8005
R2782 VSS.n1813 VSS.n1812 4.8005
R2783 VSS.n452 VSS.n451 4.8005
R2784 VSS.n305 VSS.n303 4.8005
R2785 VSS.n2832 VSS.n94 4.788
R2786 VSS.n1299 VSS.n1298 4.72533
R2787 VSS.n2536 VSS.n2535 4.72533
R2788 VSS.n635 VSS.n634 4.67352
R2789 VSS.n639 VSS.n638 4.67352
R2790 VSS.n640 VSS.n639 4.67352
R2791 VSS.n654 VSS.n653 4.67352
R2792 VSS.n656 VSS.n654 4.67352
R2793 VSS.n670 VSS.n669 4.67352
R2794 VSS.n674 VSS.n673 4.67352
R2795 VSS.n675 VSS.n674 4.67352
R2796 VSS.n515 VSS.n514 4.67352
R2797 VSS.n2372 VSS.n2371 4.67352
R2798 VSS.n2371 VSS.n2370 4.67352
R2799 VSS.n2367 VSS.n2366 4.67352
R2800 VSS.n2366 VSS.n2365 4.67352
R2801 VSS.n1247 VSS.n1246 4.67352
R2802 VSS.n1266 VSS.n1265 4.67352
R2803 VSS.n1268 VSS.n1266 4.67352
R2804 VSS.n1272 VSS.n1191 4.67352
R2805 VSS.n1273 VSS.n1272 4.67352
R2806 VSS.n1314 VSS.n1313 4.67352
R2807 VSS.n1313 VSS.n1292 4.67352
R2808 VSS.n1309 VSS.n1292 4.67352
R2809 VSS.n1309 VSS.n1308 4.67352
R2810 VSS.n1306 VSS.n1294 4.67352
R2811 VSS.n2333 VSS.n544 4.67352
R2812 VSS.n2322 VSS.n544 4.67352
R2813 VSS.n2322 VSS.n2321 4.67352
R2814 VSS.n2321 VSS.n2320 4.67352
R2815 VSS.n2317 VSS.n2316 4.67352
R2816 VSS.n2519 VSS.n248 4.67352
R2817 VSS.n2523 VSS.n248 4.67352
R2818 VSS.n2524 VSS.n2523 4.67352
R2819 VSS.n2525 VSS.n2524 4.67352
R2820 VSS.n2529 VSS.n2528 4.67352
R2821 VSS.n2539 VSS.n231 4.67352
R2822 VSS.n2553 VSS.n231 4.67352
R2823 VSS.n2554 VSS.n2553 4.67352
R2824 VSS.n2555 VSS.n2554 4.67352
R2825 VSS.n2559 VSS.n2558 4.67352
R2826 VSS.n2573 VSS.n2572 4.67352
R2827 VSS.n2574 VSS.n2573 4.67352
R2828 VSS.n2647 VSS.n2574 4.67352
R2829 VSS.n2647 VSS.n2646 4.67352
R2830 VSS.n2646 VSS.n2575 4.67352
R2831 VSS.n2642 VSS.n2575 4.67352
R2832 VSS.n2640 VSS.n2639 4.67352
R2833 VSS.n2639 VSS.n2577 4.67352
R2834 VSS.n2450 VSS.n2410 4.67352
R2835 VSS.n2436 VSS.n2435 4.67352
R2836 VSS.n2435 VSS.n2422 4.67352
R2837 VSS.n2431 VSS.n2430 4.67352
R2838 VSS.n2430 VSS.n2429 4.67352
R2839 VSS.n1291 VSS.n1290 4.63943
R2840 VSS.n1298 VSS.n543 4.63943
R2841 VSS.n2516 VSS.n2515 4.63943
R2842 VSS.n2537 VSS.n2536 4.63943
R2843 VSS.n952 VSS.n945 4.62124
R2844 VSS.n1834 VSS.n1792 4.62124
R2845 VSS.n2304 VSS.n553 4.62124
R2846 VSS.n1298 VSS.n1297 4.62124
R2847 VSS.n1612 VSS.n1611 4.62124
R2848 VSS.n2536 VSS.n243 4.62124
R2849 VSS.n1327 VSS.n1278 4.6085
R2850 VSS.n2505 VSS.n264 4.6085
R2851 VSS.n1300 VSS.n1299 4.60638
R2852 VSS.n2535 VSS.n2534 4.60638
R2853 VSS.n1316 VSS.n1291 4.55559
R2854 VSS.n2335 VSS.n543 4.55559
R2855 VSS.n2517 VSS.n2516 4.55559
R2856 VSS.n2541 VSS.n2537 4.55559
R2857 VSS.n2167 VSS.n873 4.51815
R2858 VSS.n2159 VSS.n2158 4.51815
R2859 VSS.n1578 VSS.n1577 4.51815
R2860 VSS.n1554 VSS.n1553 4.51815
R2861 VSS.n1932 VSS.n1029 4.51815
R2862 VSS.n2674 VSS.n2673 4.51401
R2863 VSS.n157 VSS.n132 4.51401
R2864 VSS.n211 VSS.n136 4.51401
R2865 VSS.n204 VSS.n135 4.51401
R2866 VSS.n2657 VSS.n218 4.51401
R2867 VSS.n223 VSS.n222 4.51401
R2868 VSS.n1801 VSS.n1798 4.51401
R2869 VSS.n1826 VSS.n1825 4.51401
R2870 VSS.n2010 VSS.n2009 4.51401
R2871 VSS.n2023 VSS.n2022 4.51401
R2872 VSS.n301 VSS.n300 4.51401
R2873 VSS.n457 VSS.n456 4.51401
R2874 VSS.n2473 VSS.n2393 4.51401
R2875 VSS.n2464 VSS.n2463 4.51401
R2876 VSS.n1711 VSS.n1702 4.51401
R2877 VSS.n1715 VSS.n1696 4.51401
R2878 VSS.n2412 VSS.n2408 4.51401
R2879 VSS.n2441 VSS.n2440 4.51401
R2880 VSS.n2124 VSS.n909 4.51401
R2881 VSS.n914 VSS.n913 4.51401
R2882 VSS.n1623 VSS.n1397 4.51401
R2883 VSS.n1410 VSS.n1409 4.51401
R2884 VSS.n930 VSS.n928 4.51401
R2885 VSS.n959 VSS.n958 4.51401
R2886 VSS.n1391 VSS.n1134 4.51401
R2887 VSS.n1382 VSS.n1381 4.51401
R2888 VSS.n2290 VSS.n841 4.51401
R2889 VSS.n2283 VSS.n2282 4.51401
R2890 VSS.n2216 VSS.n2215 4.51401
R2891 VSS.n2229 VSS.n2228 4.51401
R2892 VSS.n330 VSS.n323 4.51401
R2893 VSS.n406 VSS.n405 4.51401
R2894 VSS.n2509 VSS.n259 4.51401
R2895 VSS VSS.n2513 4.51401
R2896 VSS.n353 VSS.n346 4.51401
R2897 VSS.n376 VSS.n375 4.51401
R2898 VSS.n2545 VSS.n238 4.51401
R2899 VSS.n2550 VSS.n2549 4.51401
R2900 VSS.n1254 VSS.n1199 4.51401
R2901 VSS.n1259 VSS.n1258 4.51401
R2902 VSS.n1224 VSS.n1214 4.51401
R2903 VSS.n1229 VSS.n1228 4.51401
R2904 VSS.n835 VSS.n760 4.51401
R2905 VSS.n828 VSS.n827 4.51401
R2906 VSS.n555 VSS.n554 4.51401
R2907 VSS.n779 VSS.n778 4.51401
R2908 VSS.n1282 VSS.n1277 4.51401
R2909 VSS.n1318 VSS 4.51401
R2910 VSS.n2386 VSS.n466 4.51401
R2911 VSS.n471 VSS.n470 4.51401
R2912 VSS.n485 VSS.n483 4.51401
R2913 VSS.n497 VSS.n496 4.51401
R2914 VSS.n753 VSS.n568 4.51401
R2915 VSS.n746 VSS.n745 4.51401
R2916 VSS.n698 VSS.n589 4.51401
R2917 VSS.n703 VSS.n702 4.51401
R2918 VSS.n651 VSS.n650 4.51401
R2919 VSS.n664 VSS.n663 4.51401
R2920 VSS.n529 VSS.n524 4.51401
R2921 VSS.n620 VSS.n619 4.51401
R2922 VSS.n2339 VSS.n540 4.51401
R2923 VSS.n2329 VSS.n2325 4.51401
R2924 VSS.n2176 VSS.n2170 4.51401
R2925 VSS.n2180 VSS.n875 4.51401
R2926 VSS.n1512 VSS.n1475 4.51401
R2927 VSS.n1517 VSS.n1506 4.51401
R2928 VSS.n1976 VSS.n1001 4.51401
R2929 VSS.n1980 VSS.n995 4.51401
R2930 VSS.n1894 VSS.n1893 4.51401
R2931 VSS.n1889 VSS.n1888 4.51401
R2932 VSS.n1452 VSS.n1450 4.51401
R2933 VSS.n1543 VSS.n1542 4.51401
R2934 VSS.n1942 VSS.n1020 4.51401
R2935 VSS.n1947 VSS.n1946 4.51401
R2936 VSS.n1038 VSS.n1033 4.51401
R2937 VSS.n1913 VSS.n1912 4.51401
R2938 VSS.n1183 VSS.n1182 4.51401
R2939 VSS.n2133 VSS 4.51401
R2940 VSS.n1358 VSS.n1357 4.51401
R2941 VSS.n1352 VSS.n1351 4.51401
R2942 VSS.n1424 VSS.n1419 4.51401
R2943 VSS.n1582 VSS.n1581 4.51401
R2944 VSS.n1676 VSS.n1087 4.51401
R2945 VSS.n1092 VSS.n1091 4.51401
R2946 VSS.n1768 VSS.n1681 4.51401
R2947 VSS.n1686 VSS.n1685 4.51401
R2948 VSS.n1640 VSS.n1639 4.51401
R2949 VSS.n1630 VSS.n1124 4.51401
R2950 VSS.n2085 VSS.n964 4.51401
R2951 VSS.n2078 VSS.n2077 4.51401
R2952 VSS.n1080 VSS.n1078 4.51401
R2953 VSS.n1857 VSS.n1856 4.51401
R2954 VSS.n2626 VSS.n2625 4.51401
R2955 VSS.n2617 VSS.n2614 4.51401
R2956 VSS.n431 VSS.n430 4.51401
R2957 VSS.n2483 VSS.n2482 4.51401
R2958 VSS.n2832 VSS.n2831 4.50726
R2959 VSS.n618 VSS.n616 4.5005
R2960 VSS.n648 VSS.n647 4.5005
R2961 VSS.n659 VSS.n658 4.5005
R2962 VSS.n602 VSS.n601 4.5005
R2963 VSS.n697 VSS.n696 4.5005
R2964 VSS.n695 VSS.n694 4.5005
R2965 VSS.n592 VSS.n586 4.5005
R2966 VSS.n752 VSS.n751 4.5005
R2967 VSS.n741 VSS.n571 4.5005
R2968 VSS.n744 VSS.n723 4.5005
R2969 VSS.n487 VSS.n486 4.5005
R2970 VSS.n492 VSS.n491 4.5005
R2971 VSS.n489 VSS.n480 4.5005
R2972 VSS.n2385 VSS.n2384 4.5005
R2973 VSS.n2383 VSS.n2382 4.5005
R2974 VSS.n2379 VSS.n2378 4.5005
R2975 VSS.n2351 VSS.n2350 4.5005
R2976 VSS.n615 VSS.n530 4.5005
R2977 VSS.n1288 VSS.n1285 4.5005
R2978 VSS.n2302 VSS.n2301 4.5005
R2979 VSS.n773 VSS.n556 4.5005
R2980 VSS.n777 VSS.n776 4.5005
R2981 VSS.n834 VSS.n833 4.5005
R2982 VSS.n823 VSS.n763 4.5005
R2983 VSS.n826 VSS.n806 4.5005
R2984 VSS.n1223 VSS.n1222 4.5005
R2985 VSS.n1220 VSS.n1219 4.5005
R2986 VSS.n1216 VSS.n1210 4.5005
R2987 VSS.n1253 VSS.n1252 4.5005
R2988 VSS.n1251 VSS.n1250 4.5005
R2989 VSS.n1196 VSS.n1195 4.5005
R2990 VSS.n1325 VSS.n1324 4.5005
R2991 VSS.n1287 VSS.n1283 4.5005
R2992 VSS.n2338 VSS.n2337 4.5005
R2993 VSS.n2326 VSS.n542 4.5005
R2994 VSS.n2331 VSS.n2330 4.5005
R2995 VSS.n1181 VSS.n895 4.5005
R2996 VSS.n2138 VSS.n2137 4.5005
R2997 VSS.n898 VSS.n896 4.5005
R2998 VSS.n2175 VSS.n2174 4.5005
R2999 VSS.n2171 VSS.n874 4.5005
R3000 VSS.n2182 VSS.n2181 4.5005
R3001 VSS.n2213 VSS.n861 4.5005
R3002 VSS.n2224 VSS.n2223 4.5005
R3003 VSS.n862 VSS.n858 4.5005
R3004 VSS.n2289 VSS.n2288 4.5005
R3005 VSS.n2278 VSS.n844 4.5005
R3006 VSS.n2281 VSS.n2259 4.5005
R3007 VSS.n1390 VSS.n1389 4.5005
R3008 VSS.n1139 VSS.n1136 4.5005
R3009 VSS.n1384 VSS.n1383 4.5005
R3010 VSS.n1161 VSS.n1149 4.5005
R3011 VSS.n1165 VSS.n1164 4.5005
R3012 VSS.n1166 VSS.n1155 4.5005
R3013 VSS.n936 VSS.n934 4.5005
R3014 VSS.n1622 VSS.n1621 4.5005
R3015 VSS.n1404 VSS.n1399 4.5005
R3016 VSS.n1408 VSS.n1407 4.5005
R3017 VSS.n1550 VSS.n1549 4.5005
R3018 VSS.n1456 VSS.n1453 4.5005
R3019 VSS.n1457 VSS.n1455 4.5005
R3020 VSS.n1511 VSS.n1510 4.5005
R3021 VSS.n1508 VSS.n1478 4.5005
R3022 VSS.n1519 VSS.n1518 4.5005
R3023 VSS.n2123 VSS.n2122 4.5005
R3024 VSS.n2121 VSS.n2120 4.5005
R3025 VSS.n2117 VSS.n2116 4.5005
R3026 VSS.n2093 VSS.n2092 4.5005
R3027 VSS.n935 VSS.n931 4.5005
R3028 VSS.n1589 VSS.n1588 4.5005
R3029 VSS.n1425 VSS.n1423 4.5005
R3030 VSS.n1430 VSS.n1427 4.5005
R3031 VSS.n2076 VSS.n2056 4.5005
R3032 VSS.n1130 VSS.n1129 4.5005
R3033 VSS.n1635 VSS.n1634 4.5005
R3034 VSS.n1629 VSS.n1628 4.5005
R3035 VSS.n1675 VSS.n1674 4.5005
R3036 VSS.n1673 VSS.n1672 4.5005
R3037 VSS.n1669 VSS.n1668 4.5005
R3038 VSS.n1941 VSS.n1940 4.5005
R3039 VSS.n1026 VSS.n1025 4.5005
R3040 VSS.n1023 VSS.n1016 4.5005
R3041 VSS.n1975 VSS.n1974 4.5005
R3042 VSS.n1002 VSS.n994 4.5005
R3043 VSS.n1982 VSS.n1981 4.5005
R3044 VSS.n2007 VSS.n982 4.5005
R3045 VSS.n2018 VSS.n2017 4.5005
R3046 VSS.n979 VSS.n978 4.5005
R3047 VSS.n2084 VSS.n2083 4.5005
R3048 VSS.n2073 VSS.n967 4.5005
R3049 VSS.n1804 VSS.n1796 4.5005
R3050 VSS.n1710 VSS.n1709 4.5005
R3051 VSS.n1703 VSS.n1698 4.5005
R3052 VSS.n1717 VSS.n1716 4.5005
R3053 VSS.n1767 VSS.n1766 4.5005
R3054 VSS.n1765 VSS.n1764 4.5005
R3055 VSS.n1761 VSS.n1760 4.5005
R3056 VSS.n1920 VSS.n1919 4.5005
R3057 VSS.n1043 VSS.n1039 4.5005
R3058 VSS.n1044 VSS.n1042 4.5005
R3059 VSS.n1059 VSS.n1055 4.5005
R3060 VSS.n1064 VSS.n1063 4.5005
R3061 VSS.n1065 VSS.n1058 4.5005
R3062 VSS.n1800 VSS.n1799 4.5005
R3063 VSS.n1831 VSS.n1830 4.5005
R3064 VSS.n1864 VSS.n1863 4.5005
R3065 VSS.n1081 VSS.n1079 4.5005
R3066 VSS.n1781 VSS.n1779 4.5005
R3067 VSS.n2588 VSS.n2585 4.5005
R3068 VSS.n2621 VSS.n2620 4.5005
R3069 VSS.n2619 VSS.n2618 4.5005
R3070 VSS.n2472 VSS.n2471 4.5005
R3071 VSS.n2400 VSS.n2395 4.5005
R3072 VSS.n2466 VSS.n2465 4.5005
R3073 VSS.n2448 VSS.n2447 4.5005
R3074 VSS.n2413 VSS.n2411 4.5005
R3075 VSS.n2417 VSS.n2415 4.5005
R3076 VSS.n2508 VSS.n2507 4.5005
R3077 VSS.n262 VSS.n261 4.5005
R3078 VSS.n254 VSS.n253 4.5005
R3079 VSS.n2544 VSS.n2543 4.5005
R3080 VSS.n242 VSS.n241 4.5005
R3081 VSS.n233 VSS.n232 4.5005
R3082 VSS.n2656 VSS.n2655 4.5005
R3083 VSS.n2654 VSS.n2653 4.5005
R3084 VSS.n2650 VSS.n2649 4.5005
R3085 VSS.n184 VSS.n183 4.5005
R3086 VSS.n299 VSS.n297 4.5005
R3087 VSS.n310 VSS.n309 4.5005
R3088 VSS.n307 VSS.n284 4.5005
R3089 VSS.n333 VSS.n332 4.5005
R3090 VSS.n337 VSS.n336 4.5005
R3091 VSS.n322 VSS.n318 4.5005
R3092 VSS.n352 VSS.n348 4.5005
R3093 VSS.n381 VSS.n380 4.5005
R3094 VSS.n357 VSS.n351 4.5005
R3095 VSS.n148 VSS.n127 4.5005
R3096 VSS.n150 VSS.n149 4.5005
R3097 VSS.n155 VSS.n154 4.5005
R3098 VSS.n210 VSS.n209 4.5005
R3099 VSS.n139 VSS.n138 4.5005
R3100 VSS.n429 VSS.n428 4.5005
R3101 VSS.n427 VSS.n426 4.5005
R3102 VSS.n419 VSS.n276 4.5005
R3103 VSS.n2687 VSS.n2686 4.4805
R3104 VSS.n2046 VSS.n2045 4.38311
R3105 VSS.n634 VSS.n633 4.36875
R3106 VSS.n640 VSS.n607 4.36875
R3107 VSS.n656 VSS.n655 4.36875
R3108 VSS.n669 VSS.n668 4.36875
R3109 VSS.n675 VSS.n596 4.36875
R3110 VSS.n514 VSS.n513 4.36875
R3111 VSS.n516 VSS.n515 4.36875
R3112 VSS.n2372 VSS.n517 4.36875
R3113 VSS.n2365 VSS.n521 4.36875
R3114 VSS.n1246 VSS.n1245 4.36875
R3115 VSS.n1247 VSS.n1194 4.36875
R3116 VSS.n1265 VSS.n1193 4.36875
R3117 VSS.n1274 VSS.n1273 4.36875
R3118 VSS.n1315 VSS.n1314 4.36875
R3119 VSS.n1302 VSS.n1301 4.36875
R3120 VSS.n2334 VSS.n2333 4.36875
R3121 VSS.n2314 VSS.n548 4.36875
R3122 VSS.n2519 VSS.n2518 4.36875
R3123 VSS.n2531 VSS.n244 4.36875
R3124 VSS.n2540 VSS.n2539 4.36875
R3125 VSS.n2561 VSS.n227 4.36875
R3126 VSS.n2572 VSS.n224 4.36875
R3127 VSS.n2578 VSS.n2577 4.36875
R3128 VSS.n2451 VSS.n2450 4.36875
R3129 VSS.n2420 VSS.n2410 4.36875
R3130 VSS.n2437 VSS.n2436 4.36875
R3131 VSS.n2429 VSS.n2425 4.36875
R3132 VSS.n1745 VSS.n1743 4.28986
R3133 VSS.n1922 VSS.n1036 4.28986
R3134 VSS.n1899 VSS.n1898 4.28986
R3135 VSS.n1615 VSS.n1614 4.28986
R3136 VSS.n1609 VSS.n1411 4.28986
R3137 VSS.n954 VSS.n953 4.28986
R3138 VSS.n1836 VSS.n1835 4.28986
R3139 VSS.n1591 VSS.n1422 4.14168
R3140 VSS.n186 VSS.n182 4.11798
R3141 VSS.n201 VSS.n186 4.11798
R3142 VSS.n361 VSS.n359 4.11798
R3143 VSS.n367 VSS.n361 4.11798
R3144 VSS.n396 VSS.n395 4.11798
R3145 VSS.n395 VSS.n394 4.11798
R3146 VSS.n786 VSS.n785 4.11798
R3147 VSS.n785 VSS.n768 4.11798
R3148 VSS.n2235 VSS.n2234 4.11798
R3149 VSS.n1363 VSS.n1362 4.11798
R3150 VSS.n1362 VSS.n1361 4.11798
R3151 VSS.n1177 VSS.n1176 4.11798
R3152 VSS.n1338 VSS.n1177 4.11798
R3153 VSS.n1972 VSS.n1971 4.11798
R3154 VSS.n2488 VSS.n272 4.11798
R3155 VSS.n2491 VSS.n272 4.11798
R3156 VSS.n2305 VSS.n2304 4.09013
R3157 VSS.n1746 VSS.n1745 4.07323
R3158 VSS.n1910 VSS.n1036 4.07323
R3159 VSS.n1898 VSS.n1897 4.07323
R3160 VSS.n953 VSS.n952 4.07323
R3161 VSS.n1835 VSS.n1834 4.07323
R3162 VSS.n2276 VSS.n2275 4.03876
R3163 VSS.n2612 VSS.n2611 4.03876
R3164 VSS.n2732 VSS 4.02175
R3165 VSS.n1331 VSS.n1188 3.97459
R3166 VSS.n2501 VSS.n265 3.97459
R3167 VSS.n687 VSS.n593 3.96548
R3168 VSS.n505 VSS.n504 3.96548
R3169 VSS.n508 VSS.n505 3.96548
R3170 VSS.n831 VSS.n830 3.96548
R3171 VSS.n830 VSS.n805 3.96548
R3172 VSS.n820 VSS.n819 3.96548
R3173 VSS.n1237 VSS.n1236 3.96548
R3174 VSS.n1240 VSS.n1237 3.96548
R3175 VSS.n2271 VSS.n2270 3.96548
R3176 VSS.n1373 VSS.n1372 3.96548
R3177 VSS.n1372 VSS.n1371 3.96548
R3178 VSS.n2607 VSS.n2606 3.96548
R3179 VSS.n2458 VSS.n2457 3.96548
R3180 VSS.n2457 VSS.n2404 3.96548
R3181 VSS.n1485 VSS.n1483 3.90948
R3182 VSS.n1485 VSS.n1484 3.90948
R3183 VSS.n2777 VSS.n2776 3.78485
R3184 VSS.n2749 VSS.n2742 3.78485
R3185 VSS.n2771 VSS.n2770 3.78485
R3186 VSS.n2725 VSS.n2724 3.78485
R3187 VSS.n2238 VSS.n853 3.75994
R3188 VSS.n682 VSS.n593 3.7069
R3189 VSS.n2355 VSS.n525 3.7069
R3190 VSS.n2355 VSS.n2354 3.7069
R3191 VSS.n504 VSS.n475 3.7069
R3192 VSS.n831 VSS.n804 3.7069
R3193 VSS.n817 VSS.n809 3.7069
R3194 VSS.n1236 VSS.n1205 3.7069
R3195 VSS.n2271 VSS.n2260 3.7069
R3196 VSS.n1373 VSS.n1142 3.7069
R3197 VSS.n1371 VSS.n1144 3.7069
R3198 VSS.n2607 VSS.n2596 3.7069
R3199 VSS.n2459 VSS.n2458 3.7069
R3200 VSS.n161 VSS.n160 3.50735
R3201 VSS.n1603 VSS.n1414 3.50735
R3202 VSS.n1850 VSS.n1849 3.50735
R3203 VSS.n439 VSS.n292 3.50735
R3204 VSS.n2071 VSS.n2070 3.44377
R3205 VSS.n2070 VSS.n2069 3.44377
R3206 VSS.n222 VSS.n215 3.43925
R3207 VSS.n2658 VSS.n2657 3.43925
R3208 VSS.n1827 VSS.n1826 3.43925
R3209 VSS.n1802 VSS.n1801 3.43925
R3210 VSS.n2022 VSS.n2021 3.43925
R3211 VSS.n2009 VSS.n2008 3.43925
R3212 VSS.n2464 VSS.n460 3.43925
R3213 VSS.n2474 VSS.n2473 3.43925
R3214 VSS.n1715 VSS.n1714 3.43925
R3215 VSS.n1712 VSS.n1711 3.43925
R3216 VSS.n2442 VSS.n2441 3.43925
R3217 VSS.n2444 VSS.n2412 3.43925
R3218 VSS.n913 VSS.n906 3.43925
R3219 VSS.n2125 VSS.n2124 3.43925
R3220 VSS.n1409 VSS.n1395 3.43925
R3221 VSS.n1624 VSS.n1623 3.43925
R3222 VSS.n960 VSS.n959 3.43925
R3223 VSS.n2089 VSS.n930 3.43925
R3224 VSS.n1382 VSS.n1132 3.43925
R3225 VSS.n1392 VSS.n1391 3.43925
R3226 VSS.n2282 VSS.n838 3.43925
R3227 VSS.n2291 VSS.n2290 3.43925
R3228 VSS.n2228 VSS.n2227 3.43925
R3229 VSS.n2215 VSS.n2214 3.43925
R3230 VSS.n2513 VSS.n2512 3.43925
R3231 VSS.n2510 VSS.n2509 3.43925
R3232 VSS.n2549 VSS.n2548 3.43925
R3233 VSS.n2546 VSS.n2545 3.43925
R3234 VSS.n1258 VSS.n1257 3.43925
R3235 VSS.n1255 VSS.n1254 3.43925
R3236 VSS.n1228 VSS.n1227 3.43925
R3237 VSS.n1225 VSS.n1224 3.43925
R3238 VSS.n827 VSS.n758 3.43925
R3239 VSS.n836 VSS.n835 3.43925
R3240 VSS.n778 VSS.n559 3.43925
R3241 VSS.n2298 VSS.n555 3.43925
R3242 VSS.n1319 VSS.n1318 3.43925
R3243 VSS.n1321 VSS.n1282 3.43925
R3244 VSS.n470 VSS.n463 3.43925
R3245 VSS.n2387 VSS.n2386 3.43925
R3246 VSS.n496 VSS.n495 3.43925
R3247 VSS.n485 VSS.n484 3.43925
R3248 VSS.n745 VSS.n566 3.43925
R3249 VSS.n754 VSS.n753 3.43925
R3250 VSS.n702 VSS.n701 3.43925
R3251 VSS.n699 VSS.n698 3.43925
R3252 VSS.n663 VSS.n662 3.43925
R3253 VSS.n650 VSS.n649 3.43925
R3254 VSS.n619 VSS.n532 3.43925
R3255 VSS.n2347 VSS.n529 3.43925
R3256 VSS.n2329 VSS.n537 3.43925
R3257 VSS.n2340 VSS.n2339 3.43925
R3258 VSS.n2180 VSS.n2179 3.43925
R3259 VSS.n2177 VSS.n2176 3.43925
R3260 VSS.n1517 VSS.n1516 3.43925
R3261 VSS.n1513 VSS.n1512 3.43925
R3262 VSS.n1980 VSS.n1979 3.43925
R3263 VSS.n1977 VSS.n1976 3.43925
R3264 VSS.n1890 VSS.n1889 3.43925
R3265 VSS.n1893 VSS.n1892 3.43925
R3266 VSS.n1544 VSS.n1543 3.43925
R3267 VSS.n1546 VSS.n1452 3.43925
R3268 VSS.n1946 VSS.n1945 3.43925
R3269 VSS.n1943 VSS.n1942 3.43925
R3270 VSS.n1914 VSS.n1913 3.43925
R3271 VSS.n1916 VSS.n1038 3.43925
R3272 VSS.n1353 VSS.n1352 3.43925
R3273 VSS.n1357 VSS.n1356 3.43925
R3274 VSS.n1583 VSS.n1582 3.43925
R3275 VSS.n1585 VSS.n1424 3.43925
R3276 VSS.n1091 VSS.n1085 3.43925
R3277 VSS.n1677 VSS.n1676 3.43925
R3278 VSS.n1685 VSS.n1679 3.43925
R3279 VSS.n1769 VSS.n1768 3.43925
R3280 VSS.n2077 VSS.n961 3.43925
R3281 VSS.n2086 VSS.n2085 3.43925
R3282 VSS.n1858 VSS.n1857 3.43925
R3283 VSS.n1860 VSS.n1080 3.43925
R3284 VSS.n458 VSS.n457 3.41839
R3285 VSS.n300 VSS.n282 3.41839
R3286 VSS.n2482 VSS.n2481 3.41636
R3287 VSS.n430 VSS.n279 3.41636
R3288 VSS.n407 VSS.n406 3.41624
R3289 VSS.n323 VSS.n317 3.41624
R3290 VSS.n377 VSS.n376 3.41605
R3291 VSS.n355 VSS.n353 3.41605
R3292 VSS.n2665 VSS.n211 3.4105
R3293 VSS.n219 VSS.n217 3.4105
R3294 VSS.n2652 VSS.n2651 3.4105
R3295 VSS.n1797 VSS.n1795 3.4105
R3296 VSS.n1829 VSS.n1828 3.4105
R3297 VSS.n981 VSS.n980 3.4105
R3298 VSS.n2020 VSS.n2019 3.4105
R3299 VSS.n312 VSS.n311 3.4105
R3300 VSS.n298 VSS.n283 3.4105
R3301 VSS.n2394 VSS.n2392 3.4105
R3302 VSS.n2402 VSS.n2401 3.4105
R3303 VSS.n1704 VSS.n1701 3.4105
R3304 VSS.n1700 VSS.n1699 3.4105
R3305 VSS.n2446 VSS.n2445 3.4105
R3306 VSS.n2443 VSS.n2414 3.4105
R3307 VSS.n910 VSS.n908 3.4105
R3308 VSS.n2119 VSS.n2118 3.4105
R3309 VSS.n1398 VSS.n1396 3.4105
R3310 VSS.n1406 VSS.n1405 3.4105
R3311 VSS.n2091 VSS.n2090 3.4105
R3312 VSS.n933 VSS.n932 3.4105
R3313 VSS.n1135 VSS.n1133 3.4105
R3314 VSS.n1141 VSS.n1140 3.4105
R3315 VSS.n842 VSS.n840 3.4105
R3316 VSS.n2280 VSS.n2279 3.4105
R3317 VSS.n860 VSS.n859 3.4105
R3318 VSS.n2226 VSS.n2225 3.4105
R3319 VSS.n334 VSS.n315 3.4105
R3320 VSS.n335 VSS.n316 3.4105
R3321 VSS.n263 VSS.n258 3.4105
R3322 VSS.n260 VSS.n255 3.4105
R3323 VSS.n354 VSS.n350 3.4105
R3324 VSS.n379 VSS.n378 3.4105
R3325 VSS.n239 VSS.n237 3.4105
R3326 VSS.n240 VSS.n234 3.4105
R3327 VSS.n1200 VSS.n1198 3.4105
R3328 VSS.n1249 VSS.n1197 3.4105
R3329 VSS.n1215 VSS.n1213 3.4105
R3330 VSS.n1218 VSS.n1211 3.4105
R3331 VSS.n761 VSS.n759 3.4105
R3332 VSS.n825 VSS.n824 3.4105
R3333 VSS.n2300 VSS.n2299 3.4105
R3334 VSS.n772 VSS.n557 3.4105
R3335 VSS.n1323 VSS.n1322 3.4105
R3336 VSS.n1320 VSS.n1284 3.4105
R3337 VSS.n467 VSS.n465 3.4105
R3338 VSS.n2381 VSS.n2380 3.4105
R3339 VSS.n482 VSS.n481 3.4105
R3340 VSS.n494 VSS.n493 3.4105
R3341 VSS.n569 VSS.n567 3.4105
R3342 VSS.n743 VSS.n742 3.4105
R3343 VSS.n590 VSS.n588 3.4105
R3344 VSS.n693 VSS.n587 3.4105
R3345 VSS.n604 VSS.n603 3.4105
R3346 VSS.n661 VSS.n660 3.4105
R3347 VSS.n2349 VSS.n2348 3.4105
R3348 VSS.n617 VSS.n531 3.4105
R3349 VSS.n541 VSS.n539 3.4105
R3350 VSS.n2328 VSS.n2327 3.4105
R3351 VSS.n2172 VSS.n879 3.4105
R3352 VSS.n877 VSS.n876 3.4105
R3353 VSS.n1514 VSS.n1509 3.4105
R3354 VSS.n1515 VSS.n1507 3.4105
R3355 VSS.n1003 VSS.n1000 3.4105
R3356 VSS.n997 VSS.n996 3.4105
R3357 VSS.n1061 VSS.n1056 3.4105
R3358 VSS.n1062 VSS.n1057 3.4105
R3359 VSS.n1548 VSS.n1547 3.4105
R3360 VSS.n1545 VSS.n1454 3.4105
R3361 VSS.n1021 VSS.n1019 3.4105
R3362 VSS.n1024 VSS.n1017 3.4105
R3363 VSS.n1918 VSS.n1917 3.4105
R3364 VSS.n1041 VSS.n1040 3.4105
R3365 VSS.n2134 VSS.n2132 3.4105
R3366 VSS.n2132 VSS.n902 3.4105
R3367 VSS.n2134 VSS.n2133 3.4105
R3368 VSS.n1182 VSS.n902 3.4105
R3369 VSS.n901 VSS.n897 3.4105
R3370 VSS.n2136 VSS.n2135 3.4105
R3371 VSS.n1162 VSS.n1150 3.4105
R3372 VSS.n1163 VSS.n1154 3.4105
R3373 VSS.n1587 VSS.n1586 3.4105
R3374 VSS.n1584 VSS.n1426 3.4105
R3375 VSS.n1088 VSS.n1086 3.4105
R3376 VSS.n1671 VSS.n1670 3.4105
R3377 VSS.n1682 VSS.n1680 3.4105
R3378 VSS.n1763 VSS.n1762 3.4105
R3379 VSS.n1631 VSS.n1626 3.4105
R3380 VSS.n1638 VSS.n1626 3.4105
R3381 VSS.n1631 VSS.n1630 3.4105
R3382 VSS.n1639 VSS.n1638 3.4105
R3383 VSS.n1637 VSS.n1636 3.4105
R3384 VSS.n1633 VSS.n1632 3.4105
R3385 VSS.n965 VSS.n963 3.4105
R3386 VSS.n2075 VSS.n2074 3.4105
R3387 VSS.n1862 VSS.n1861 3.4105
R3388 VSS.n1778 VSS.n1082 3.4105
R3389 VSS.n2616 VSS.n213 3.4105
R3390 VSS.n2624 VSS.n213 3.4105
R3391 VSS.n2617 VSS.n2616 3.4105
R3392 VSS.n2625 VSS.n2624 3.4105
R3393 VSS.n2623 VSS.n2622 3.4105
R3394 VSS.n2615 VSS.n2587 3.4105
R3395 VSS.n418 VSS.n417 3.4105
R3396 VSS.n425 VSS.n277 3.4105
R3397 VSS.n2667 VSS.n132 3.4105
R3398 VSS.n2673 VSS.n2672 3.4105
R3399 VSS.n2670 VSS.n130 3.4105
R3400 VSS.n2669 VSS.n131 3.4105
R3401 VSS.n2665 VSS.n135 3.4105
R3402 VSS.n2665 VSS.n134 3.4105
R3403 VSS.n2665 VSS.n133 3.4105
R3404 VSS.n88 VSS.n87 3.40476
R3405 VSS.n2240 VSS.n2239 3.31239
R3406 VSS.n1971 VSS.n993 3.22288
R3407 VSS.n2071 VSS.n2055 3.21921
R3408 VSS.n2066 VSS.n2065 3.21921
R3409 VSS.n165 VSS.n146 3.2005
R3410 VSS.n1601 VSS.n1416 3.2005
R3411 VSS.n1854 VSS.n1784 3.2005
R3412 VSS.n438 VSS.n293 3.2005
R3413 VSS.n1735 VSS.n1734 3.13241
R3414 VSS.n1881 VSS.n1880 3.13241
R3415 VSS.n734 VSS.n725 3.13241
R3416 VSS.n2198 VSS.n2197 3.13241
R3417 VSS.n2716 VSS.n2715 3.13241
R3418 VSS.n2824 VSS.n2820 3.13241
R3419 VSS.n2849 VSS.n2848 3.13241
R3420 VSS.n87 VSS.n83 3.13241
R3421 VSS.n2697 VSS.n2696 3.1005
R3422 VSS.n527 VSS.n526 3.09945
R3423 VSS.n1275 VSS.n1188 3.05276
R3424 VSS.n2426 VSS.n265 3.05276
R3425 VSS.n730 VSS.n728 3.04861
R3426 VSS.n813 VSS.n811 3.04861
R3427 VSS.n1232 VSS.n1230 3.04861
R3428 VSS.n2265 VSS.n2264 3.04861
R3429 VSS.n951 VSS.n950 3.04861
R3430 VSS.n2063 VSS.n2062 3.04861
R3431 VSS.n1897 VSS.n1052 3.04861
R3432 VSS.n2601 VSS.n2600 3.04861
R3433 VSS.n500 VSS.n498 3.04861
R3434 VSS.n1753 VSS.n1746 3.04861
R3435 VSS.n2462 VSS.n2398 3.04861
R3436 VSS.n1102 VSS.n1099 3.01226
R3437 VSS.n1564 VSS.n1563 2.92224
R3438 VSS.n2304 VSS.n552 2.92166
R3439 VSS.n508 VSS.n507 2.88804
R3440 VSS.n1240 VSS.n1239 2.88804
R3441 VSS.n2406 VSS.n2404 2.88804
R3442 VSS.n89 VSS.n88 2.86007
R3443 VSS.n507 VSS.n506 2.79323
R3444 VSS.n1239 VSS.n1238 2.79323
R3445 VSS.n2406 VSS.n2405 2.79323
R3446 VSS.n2275 VSS.n2274 2.77203
R3447 VSS.n2611 VSS.n2610 2.77203
R3448 VSS.n1734 VSS.n1733 2.7239
R3449 VSS.n1880 VSS.n1879 2.7239
R3450 VSS.n726 VSS.n725 2.7239
R3451 VSS.n2199 VSS.n2198 2.7239
R3452 VSS.n1646 VSS.n1122 2.7239
R3453 VSS.n2717 VSS.n2716 2.7239
R3454 VSS.n2821 VSS.n2820 2.7239
R3455 VSS.n2848 VSS.n2847 2.7239
R3456 VSS.n84 VSS.n83 2.7239
R3457 VSS.n2233 VSS.n2232 2.68581
R3458 VSS.n2703 VSS.n2702 2.63717
R3459 VSS.n164 VSS.n144 2.63064
R3460 VSS.n1599 VSS.n1598 2.63064
R3461 VSS.n1853 VSS.n1848 2.63064
R3462 VSS.n436 VSS.n435 2.63064
R3463 VSS.n624 VSS.n623 2.55412
R3464 VSS.n2207 VSS.n865 2.50679
R3465 VSS.n1958 VSS.n1957 2.50679
R3466 VSS.n2634 VSS.n2633 2.50679
R3467 VSS.n2306 VSS.n2305 2.38348
R3468 VSS.n635 VSS.n609 2.33701
R3469 VSS.n638 VSS.n609 2.33701
R3470 VSS.n653 VSS.n606 2.33701
R3471 VSS.n670 VSS.n598 2.33701
R3472 VSS.n673 VSS.n598 2.33701
R3473 VSS.n2370 VSS.n519 2.33701
R3474 VSS.n2367 VSS.n519 2.33701
R3475 VSS.n1268 VSS.n1267 2.33701
R3476 VSS.n1267 VSS.n1191 2.33701
R3477 VSS.n1308 VSS.n1307 2.33701
R3478 VSS.n1307 VSS.n1306 2.33701
R3479 VSS.n1296 VSS.n1294 2.33701
R3480 VSS.n1302 VSS.n1296 2.33701
R3481 VSS.n2320 VSS.n546 2.33701
R3482 VSS.n2317 VSS.n546 2.33701
R3483 VSS.n2316 VSS.n2315 2.33701
R3484 VSS.n2315 VSS.n2314 2.33701
R3485 VSS.n2525 VSS.n246 2.33701
R3486 VSS.n2528 VSS.n246 2.33701
R3487 VSS.n2530 VSS.n2529 2.33701
R3488 VSS.n2531 VSS.n2530 2.33701
R3489 VSS.n2555 VSS.n229 2.33701
R3490 VSS.n2558 VSS.n229 2.33701
R3491 VSS.n2560 VSS.n2559 2.33701
R3492 VSS.n2561 VSS.n2560 2.33701
R3493 VSS.n2642 VSS.n2641 2.33701
R3494 VSS.n2641 VSS.n2640 2.33701
R3495 VSS.n2424 VSS.n2422 2.33701
R3496 VSS.n2431 VSS.n2424 2.33701
R3497 VSS.n628 VSS.n613 2.33067
R3498 VSS.n749 VSS.n721 2.25932
R3499 VSS.n2153 VSS.n2152 2.25932
R3500 VSS.n1577 VSS.n1576 2.25932
R3501 VSS.n1555 VSS.n1554 2.25932
R3502 VSS.n1460 VSS.n1449 2.25932
R3503 VSS.n1461 VSS.n1460 2.25932
R3504 VSS.n919 VSS.n916 2.25932
R3505 VSS.n1653 VSS.n1119 2.25932
R3506 VSS.n2015 VSS.n977 2.25932
R3507 VSS.n1102 VSS.n1101 2.25932
R3508 VSS.n510 VSS.n473 2.25312
R3509 VSS.n1242 VSS.n1203 2.25312
R3510 VSS.n2454 VSS.n2407 2.25312
R3511 VSS.n1499 VSS.n1485 2.25293
R3512 VSS.n473 VSS.n472 2.2228
R3513 VSS.n1203 VSS.n1202 2.2228
R3514 VSS.n2409 VSS.n2407 2.2228
R3515 VSS.n1647 VSS.n1646 2.17922
R3516 VSS.n2873 VSS.n2872 2.14347
R3517 VSS.n1614 VSS.n1613 2.13383
R3518 VSS.n1280 VSS.n1279 2.11085
R3519 VSS.n252 VSS.n251 2.11085
R3520 VSS.n819 VSS.n818 2.06919
R3521 VSS.n644 VSS.n606 2.03225
R3522 VSS.n688 VSS.n687 1.98299
R3523 VSS.n808 VSS.n805 1.98299
R3524 VSS.n820 VSS.n808 1.98299
R3525 VSS.n2270 VSS.n2269 1.98299
R3526 VSS.n2606 VSS.n2605 1.98299
R3527 VSS.n2052 VSS.n2051 1.97497
R3528 VSS.n627 VSS.n614 1.91571
R3529 VSS.n818 VSS.n817 1.8968
R3530 VSS.n940 VSS.n939 1.88285
R3531 VSS.n1563 VSS.n1562 1.87876
R3532 VSS.n2069 VSS.n2058 1.79699
R3533 VSS.n2246 VSS.n2244 1.75824
R3534 VSS.n2819 VSS.n2818 1.753
R3535 VSS.n2817 VSS.n2816 1.753
R3536 VSS.n1569 VSS.n1567 1.7528
R3537 VSS.n689 VSS.n688 1.72441
R3538 VSS.n2269 VSS.n2268 1.72441
R3539 VSS.n2605 VSS.n2604 1.72441
R3540 VSS.n2668 VSS.n129 1.70468
R3541 VSS.n2671 VSS.n129 1.70468
R3542 VSS.n377 VSS.n356 1.70348
R3543 VSS.n356 VSS.n355 1.70348
R3544 VSS.n408 VSS.n407 1.70338
R3545 VSS.n408 VSS.n317 1.70338
R3546 VSS.n2481 VSS.n2480 1.70332
R3547 VSS.n2480 VSS.n279 1.70332
R3548 VSS.n459 VSS.n458 1.70231
R3549 VSS.n459 VSS.n282 1.70231
R3550 VSS.n2276 VSS.n2258 1.7012
R3551 VSS.n1891 VSS.n1890 1.69188
R3552 VSS.n1892 VSS.n1891 1.69188
R3553 VSS.n1979 VSS.n1978 1.69188
R3554 VSS.n1978 VSS.n1977 1.69188
R3555 VSS.n1516 VSS.n998 1.69188
R3556 VSS.n1513 VSS.n998 1.69188
R3557 VSS.n2179 VSS.n2178 1.69188
R3558 VSS.n2178 VSS.n2177 1.69188
R3559 VSS.n2341 VSS.n537 1.69188
R3560 VSS.n2341 VSS.n2340 1.69188
R3561 VSS.n662 VSS.n536 1.69188
R3562 VSS.n649 VSS.n536 1.69188
R3563 VSS.n2548 VSS.n2547 1.69188
R3564 VSS.n2547 VSS.n2546 1.69188
R3565 VSS.n1915 VSS.n1914 1.69188
R3566 VSS.n1916 VSS.n1915 1.69188
R3567 VSS.n1945 VSS.n1944 1.69188
R3568 VSS.n1944 VSS.n1943 1.69188
R3569 VSS.n1544 VSS.n903 1.69188
R3570 VSS.n1546 VSS.n903 1.69188
R3571 VSS.n1319 VSS.n533 1.69188
R3572 VSS.n1321 VSS.n533 1.69188
R3573 VSS.n2346 VSS.n532 1.69188
R3574 VSS.n2347 VSS.n2346 1.69188
R3575 VSS.n2512 VSS.n2511 1.69188
R3576 VSS.n2511 VSS.n2510 1.69188
R3577 VSS.n2132 VSS.n899 1.69188
R3578 VSS.n1770 VSS.n1679 1.69188
R3579 VSS.n1770 VSS.n1769 1.69188
R3580 VSS.n1678 VSS.n1085 1.69188
R3581 VSS.n1678 VSS.n1677 1.69188
R3582 VSS.n1583 VSS.n1084 1.69188
R3583 VSS.n1585 VSS.n1084 1.69188
R3584 VSS.n1355 VSS.n1353 1.69188
R3585 VSS.n1356 VSS.n1355 1.69188
R3586 VSS.n1257 VSS.n1256 1.69188
R3587 VSS.n1256 VSS.n1255 1.69188
R3588 VSS.n2388 VSS.n463 1.69188
R3589 VSS.n2388 VSS.n2387 1.69188
R3590 VSS.n2442 VSS.n280 1.69188
R3591 VSS.n2444 VSS.n280 1.69188
R3592 VSS.n1714 VSS.n1713 1.69188
R3593 VSS.n1713 VSS.n1712 1.69188
R3594 VSS.n1625 VSS.n1395 1.69188
R3595 VSS.n1625 VSS.n1624 1.69188
R3596 VSS.n1393 VSS.n1132 1.69188
R3597 VSS.n1393 VSS.n1392 1.69188
R3598 VSS.n1227 VSS.n1226 1.69188
R3599 VSS.n1226 VSS.n1225 1.69188
R3600 VSS.n495 VSS.n461 1.69188
R3601 VSS.n484 VSS.n461 1.69188
R3602 VSS.n2475 VSS.n460 1.69188
R3603 VSS.n2475 VSS.n2474 1.69188
R3604 VSS.n1627 VSS.n1626 1.69188
R3605 VSS.n1859 VSS.n1858 1.69188
R3606 VSS.n1860 VSS.n1859 1.69188
R3607 VSS.n2021 VSS.n907 1.69188
R3608 VSS.n2008 VSS.n907 1.69188
R3609 VSS.n2126 VSS.n906 1.69188
R3610 VSS.n2126 VSS.n2125 1.69188
R3611 VSS.n2227 VSS.n560 1.69188
R3612 VSS.n2214 VSS.n560 1.69188
R3613 VSS.n2297 VSS.n559 1.69188
R3614 VSS.n2298 VSS.n2297 1.69188
R3615 VSS.n701 VSS.n700 1.69188
R3616 VSS.n700 VSS.n699 1.69188
R3617 VSS.n2659 VSS.n215 1.69188
R3618 VSS.n2659 VSS.n2658 1.69188
R3619 VSS.n1827 VSS.n1803 1.69188
R3620 VSS.n1803 VSS.n1802 1.69188
R3621 VSS.n2087 VSS.n961 1.69188
R3622 VSS.n2087 VSS.n2086 1.69188
R3623 VSS.n2088 VSS.n960 1.69188
R3624 VSS.n2089 VSS.n2088 1.69188
R3625 VSS.n2292 VSS.n838 1.69188
R3626 VSS.n2292 VSS.n2291 1.69188
R3627 VSS.n837 VSS.n758 1.69188
R3628 VSS.n837 VSS.n836 1.69188
R3629 VSS.n755 VSS.n566 1.69188
R3630 VSS.n755 VSS.n754 1.69188
R3631 VSS.n2586 VSS.n213 1.69188
R3632 VSS.n2066 VSS.n2058 1.64728
R3633 VSS.n2220 VSS.n856 1.61169
R3634 VSS VSS.n8 1.54822
R3635 VSS.n680 VSS.n679 1.47352
R3636 VSS.n2362 VSS.n2361 1.34658
R3637 VSS.n2305 VSS.n551 1.3283
R3638 VSS.n512 VSS.n472 1.29527
R3639 VSS.n1244 VSS.n1202 1.29527
R3640 VSS.n2452 VSS.n2409 1.29527
R3641 VSS.n2595 VSS.n2594 1.25365
R3642 VSS.n2360 VSS.n522 1.25033
R3643 VSS.n75 VSS.n0 1.21169
R3644 VSS.n1377 VSS.n1376 1.20723
R3645 VSS.n191 VSS.n190 1.18311
R3646 VSS.n327 VSS.n326 1.18311
R3647 VSS.n1706 VSS.n1705 1.18311
R3648 VSS.n1562 VSS.n1561 1.18311
R3649 VSS.n2003 VSS.n2002 1.18311
R3650 VSS.n2045 VSS.n970 1.18311
R3651 VSS.n1812 VSS.n1811 1.18311
R3652 VSS.n451 VSS.n450 1.18311
R3653 VSS.n303 VSS.n302 1.18311
R3654 VSS.n165 VSS.n164 1.14023
R3655 VSS.n1599 VSS.n1416 1.14023
R3656 VSS.n1854 VSS.n1853 1.14023
R3657 VSS.n436 VSS.n293 1.14023
R3658 VSS.n1466 VSS.n1463 1.12991
R3659 VSS.n683 VSS.n681 1.12954
R3660 VSS.n278 VSS 1.12383
R3661 VSS.n409 VSS 1.11689
R3662 VSS.n212 VSS 1.11689
R3663 VSS.n411 VSS 1.07702
R3664 VSS.n2251 VSS.n2250 1.07463
R3665 VSS.n107 VSS.n104 0.993972
R3666 VSS.n2286 VSS.n2257 0.985115
R3667 VSS.n1648 VSS.n1647 0.953691
R3668 VSS.n1745 VSS.n1744 0.952566
R3669 VSS.n1036 VSS.n1035 0.952566
R3670 VSS.n1898 VSS.n1051 0.952566
R3671 VSS.n953 VSS.n944 0.952566
R3672 VSS.n1835 VSS.n1790 0.952566
R3673 VSS.n952 VSS.n947 0.899674
R3674 VSS.n1967 VSS.n1005 0.895605
R3675 VSS.n1984 VSS.n993 0.895605
R3676 VSS.n507 VSS.n473 0.892621
R3677 VSS.n1239 VSS.n1203 0.892621
R3678 VSS.n2407 VSS.n2406 0.892621
R3679 VSS.n2665 VSS.n2664 0.853
R3680 VSS.n2700 VSS.n2699 0.842928
R3681 VSS.n160 VSS.n146 0.833377
R3682 VSS.n1849 VSS.n1784 0.833377
R3683 VSS.n439 VSS.n438 0.833377
R3684 VSS.n628 VSS.n627 0.830425
R3685 VSS.n622 VSS.n526 0.798505
R3686 VSS.n2686 VSS.n113 0.777453
R3687 VSS.n2818 VSS.n2817 0.761313
R3688 VSS.n2144 VSS.n890 0.753441
R3689 VSS.n1572 VSS.n1571 0.753441
R3690 VSS.n2100 VSS.n925 0.753441
R3691 VSS.n1175 VSS.n1172 0.716584
R3692 VSS.n623 VSS.n613 0.606984
R3693 VSS.n175 VSS.n174 0.537563
R3694 VSS.n196 VSS.n187 0.537563
R3695 VSS.n387 VSS.n345 0.537563
R3696 VSS.n362 VSS.n124 0.537563
R3697 VSS.n340 VSS.n339 0.537563
R3698 VSS.n389 VSS.n388 0.537563
R3699 VSS.n797 VSS.n796 0.537563
R3700 VSS.n784 VSS.n783 0.537563
R3701 VSS.n795 VSS.n766 0.537563
R3702 VSS.n2248 VSS.n2247 0.537563
R3703 VSS.n2218 VSS.n864 0.537563
R3704 VSS.n2244 VSS.n849 0.537563
R3705 VSS.n1168 VSS.n1160 0.537563
R3706 VSS.n1170 VSS.n1169 0.537563
R3707 VSS.n1184 VSS.n1179 0.537563
R3708 VSS.n1989 VSS.n990 0.537563
R3709 VSS.n2568 VSS.n225 0.537563
R3710 VSS.n420 VSS.n295 0.537563
R3711 VSS.n2496 VSS.n270 0.537563
R3712 VSS.n161 VSS.n159 0.526527
R3713 VSS.n1606 VSS.n1414 0.526527
R3714 VSS.n1603 VSS.n1602 0.526527
R3715 VSS.n1850 VSS.n1077 0.526527
R3716 VSS.n292 VSS.n290 0.526527
R3717 VSS.n1394 VSS.n904 0.500125
R3718 VSS.n1772 VSS.n1083 0.500125
R3719 VSS.n2391 VSS.n2390 0.500125
R3720 VSS.n1212 VSS.n534 0.500125
R3721 VSS.n1152 VSS.n1131 0.500125
R3722 VSS.n2478 VSS.n2476 0.500125
R3723 VSS.n2732 VSS.n99 0.482665
R3724 VSS.n2774 VSS.n2773 0.467019
R3725 VSS.n2872 VSS 0.448179
R3726 VSS.n1158 VSS.n1147 0.448052
R3727 VSS.n1349 VSS.n1171 0.448052
R3728 VSS.n2582 VSS.n2580 0.448052
R3729 VSS.n195 VSS.n188 0.417891
R3730 VSS.n325 VSS.n268 0.417891
R3731 VSS.n326 VSS.n321 0.417891
R3732 VSS.n1719 VSS.n1697 0.417891
R3733 VSS.n1567 VSS.n1440 0.417891
R3734 VSS.n1561 VSS.n1560 0.417891
R3735 VSS.n2001 VSS.n2000 0.417891
R3736 VSS.n2002 VSS.n983 0.417891
R3737 VSS.n2044 VSS.n2043 0.417891
R3738 VSS.n2047 VSS.n2046 0.417891
R3739 VSS.n2050 VSS.n970 0.417891
R3740 VSS.n1816 VSS.n1809 0.417891
R3741 VSS.n454 VSS.n453 0.417891
R3742 VSS.n450 VSS.n449 0.417891
R3743 VSS.n304 VSS.n286 0.417891
R3744 VSS.n2697 VSS.n113 0.410656
R3745 VSS.n2676 VSS.n125 0.409011
R3746 VSS.n1758 VSS.n1757 0.409011
R3747 VSS.n1731 VSS.n1730 0.409011
R3748 VSS.n1733 VSS.n1689 0.409011
R3749 VSS.n1034 VSS.n1032 0.409011
R3750 VSS.n1050 VSS.n1048 0.409011
R3751 VSS.n1885 VSS.n1068 0.409011
R3752 VSS.n1879 VSS.n1878 0.409011
R3753 VSS.n738 VSS.n737 0.409011
R3754 VSS.n731 VSS.n726 0.409011
R3755 VSS.n2193 VSS.n868 0.409011
R3756 VSS.n1618 VSS.n1403 0.409011
R3757 VSS.n1608 VSS.n1607 0.409011
R3758 VSS.n942 VSS.n941 0.409011
R3759 VSS.n1642 VSS.n1123 0.409011
R3760 VSS.n1651 VSS.n1122 0.409011
R3761 VSS.n1871 VSS.n1075 0.409011
R3762 VSS.n1789 VSS.n1787 0.409011
R3763 VSS.n2814 VSS.n2717 0.409011
R3764 VSS.n2828 VSS.n98 0.409011
R3765 VSS.n2854 VSS.n2853 0.409011
R3766 VSS.n2852 VSS.n68 0.409011
R3767 VSS.n2847 VSS.n2846 0.409011
R3768 VSS.n91 VSS.n90 0.409011
R3769 VSS.n289 VSS.n287 0.409011
R3770 VSS.n624 VSS.n622 0.383542
R3771 VSS.n561 VSS.n538 0.3805
R3772 VSS.n2343 VSS.n2342 0.3805
R3773 VSS.n562 VSS.n236 0.3805
R3774 VSS.n1774 VSS.n999 0.3805
R3775 VSS.n2129 VSS.n878 0.3805
R3776 VSS.n235 VSS.n214 0.3805
R3777 VSS.n2477 VSS.n256 0.3805
R3778 VSS.n462 VSS.n257 0.3805
R3779 VSS.n2345 VSS.n2344 0.3805
R3780 VSS.n1151 VSS.n900 0.3805
R3781 VSS.n2131 VSS.n2130 0.3805
R3782 VSS.n1773 VSS.n1018 0.3805
R3783 VSS.n2479 VSS.n2478 0.3805
R3784 VSS.n2390 VSS.n2389 0.3805
R3785 VSS.n534 VSS.n464 0.3805
R3786 VSS.n1153 VSS.n1152 0.3805
R3787 VSS.n1354 VSS.n904 0.3805
R3788 VSS.n1772 VSS.n1771 0.3805
R3789 VSS.n2661 VSS.n2660 0.3805
R3790 VSS.n563 VSS.n216 0.3805
R3791 VSS.n558 VSS.n535 0.3805
R3792 VSS.n2296 VSS.n2295 0.3805
R3793 VSS.n2128 VSS.n2127 0.3805
R3794 VSS.n1777 VSS.n1776 0.3805
R3795 VSS.n2294 VSS.n2293 0.3805
R3796 VSS.n757 VSS.n756 0.3805
R3797 VSS.n565 VSS.n564 0.3805
R3798 VSS.n2663 VSS.n2662 0.3805
R3799 VSS.n1775 VSS.n962 0.3805
R3800 VSS.n905 VSS.n839 0.3805
R3801 VSS.n939 VSS.n927 0.376971
R3802 VSS VSS.n2873 0.366908
R3803 VSS.n2702 VSS.n2701 0.358995
R3804 VSS.n791 VSS.n766 0.358542
R3805 VSS.n2210 VSS.n2209 0.358542
R3806 VSS.n2234 VSS.n853 0.358542
R3807 VSS.n1959 VSS.n1958 0.358542
R3808 VSS.n2201 VSS.n2200 0.340926
R3809 VSS.n1602 VSS.n1601 0.307349
R3810 VSS.n633 VSS.n632 0.305262
R3811 VSS.n643 VSS.n607 0.305262
R3812 VSS.n645 VSS.n644 0.305262
R3813 VSS.n655 VSS.n600 0.305262
R3814 VSS.n668 VSS.n667 0.305262
R3815 VSS.n679 VSS.n596 0.305262
R3816 VSS.n513 VSS.n512 0.305262
R3817 VSS.n2376 VSS.n516 0.305262
R3818 VSS.n2375 VSS.n517 0.305262
R3819 VSS.n2362 VSS.n521 0.305262
R3820 VSS.n1245 VSS.n1244 0.305262
R3821 VSS.n1261 VSS.n1194 0.305262
R3822 VSS.n1262 VSS.n1193 0.305262
R3823 VSS.n1275 VSS.n1274 0.305262
R3824 VSS.n1316 VSS.n1315 0.305262
R3825 VSS.n1301 VSS.n1300 0.305262
R3826 VSS.n2335 VSS.n2334 0.305262
R3827 VSS.n2311 VSS.n548 0.305262
R3828 VSS.n2518 VSS.n2517 0.305262
R3829 VSS.n2534 VSS.n244 0.305262
R3830 VSS.n2541 VSS.n2540 0.305262
R3831 VSS.n2564 VSS.n227 0.305262
R3832 VSS.n2569 VSS.n224 0.305262
R3833 VSS.n2635 VSS.n2578 0.305262
R3834 VSS.n2452 VSS.n2451 0.305262
R3835 VSS.n2421 VSS.n2420 0.305262
R3836 VSS.n2438 VSS.n2437 0.305262
R3837 VSS.n2426 VSS.n2425 0.305262
R3838 VSS.n2700 VSS.n104 0.298799
R3839 VSS.n510 VSS.n509 0.298074
R3840 VSS.n1242 VSS.n1241 0.298074
R3841 VSS.n2455 VSS.n2454 0.298074
R3842 VSS.n413 VSS.n412 0.278782
R3843 VSS.n168 VSS.n144 0.263514
R3844 VSS.n1598 VSS.n1597 0.263514
R3845 VSS.n1848 VSS.n1847 0.263514
R3846 VSS.n435 VSS.n434 0.263514
R3847 VSS VSS.n0 0.260439
R3848 VSS.n683 VSS.n682 0.259086
R3849 VSS.n690 VSS.n689 0.259086
R3850 VSS.n525 VSS.n522 0.259086
R3851 VSS.n2354 VSS.n2353 0.259086
R3852 VSS.n501 VSS.n475 0.259086
R3853 VSS.n804 VSS.n803 0.259086
R3854 VSS.n814 VSS.n809 0.259086
R3855 VSS.n1233 VSS.n1205 0.259086
R3856 VSS.n2274 VSS.n2260 0.259086
R3857 VSS.n2268 VSS.n2267 0.259086
R3858 VSS.n1376 VSS.n1142 0.259086
R3859 VSS.n1368 VSS.n1144 0.259086
R3860 VSS.n2610 VSS.n2596 0.259086
R3861 VSS.n2604 VSS.n2603 0.259086
R3862 VSS.n2460 VSS.n2459 0.259086
R3863 VSS.n2696 VSS.n114 0.2565
R3864 VSS.n1754 VSS.n1753 0.239726
R3865 VSS.n1052 VSS.n1049 0.239381
R3866 VSS VSS.n1499 0.237784
R3867 VSS.n2701 VSS.n2700 0.23574
R3868 VSS.n2080 VSS.n2055 0.225061
R3869 VSS.n2065 VSS.n2064 0.225061
R3870 VSS.n2666 VSS.n104 0.224703
R3871 VSS.n459 VSS.n281 0.218753
R3872 VSS.n735 VSS.n734 0.204755
R3873 VSS.n2053 VSS.n2052 0.204755
R3874 VSS.n2054 VSS.n2053 0.204755
R3875 VSS.n1499 VSS 0.200023
R3876 VSS VSS.n510 0.199635
R3877 VSS VSS.n1242 0.199635
R3878 VSS.n2454 VSS 0.199635
R3879 VSS.n410 VSS.n281 0.196532
R3880 VSS.n416 VSS.n415 0.196532
R3881 VSS.n412 VSS.n212 0.195539
R3882 VSS.n614 VSS.n611 0.192021
R3883 VSS.n2667 VSS.n2666 0.184476
R3884 VSS.n2734 VSS.n2732 0.1838
R3885 VSS.n1792 VSS.n1788 0.180304
R3886 VSS.n950 VSS 0.17983
R3887 VSS.n2062 VSS 0.17983
R3888 VSS.n2209 VSS.n865 0.179521
R3889 VSS.n1960 VSS.n1959 0.179521
R3890 VSS.n2592 VSS.n2583 0.179521
R3891 VSS.n728 VSS 0.179485
R3892 VSS.n811 VSS 0.179485
R3893 VSS VSS.n2265 0.179485
R3894 VSS VSS.n2601 0.179485
R3895 VSS.n2672 VSS.n128 0.175416
R3896 VSS.n113 VSS.n112 0.173577
R3897 VSS.n416 VSS.n314 0.169759
R3898 VSS.n1978 VSS.n998 0.1603
R3899 VSS.n1944 VSS.n903 0.1603
R3900 VSS.n1678 VSS.n1084 0.1603
R3901 VSS.n1626 VSS.n1625 0.1603
R3902 VSS.n2126 VSS.n907 0.1603
R3903 VSS.n2088 VSS.n2087 0.1603
R3904 VSS.n2178 VSS.n878 0.159712
R3905 VSS.n2132 VSS.n2131 0.159712
R3906 VSS.n1355 VSS.n1354 0.159712
R3907 VSS.n1394 VSS.n1393 0.159712
R3908 VSS.n2127 VSS.n560 0.159712
R3909 VSS.n2292 VSS.n839 0.159712
R3910 VSS.n1297 VSS 0.158169
R3911 VSS.n553 VSS 0.158169
R3912 VSS VSS.n243 0.158169
R3913 VSS VSS.n945 0.156867
R3914 VSS.n1798 VSS.n1792 0.151658
R3915 VSS.n498 VSS.n497 0.143372
R3916 VSS.n2463 VSS.n2462 0.143372
R3917 VSS.n1230 VSS.n1229 0.143027
R3918 VSS.n728 VSS 0.14207
R3919 VSS.n1230 VSS 0.14207
R3920 VSS.n811 VSS 0.14207
R3921 VSS.n2265 VSS 0.14207
R3922 VSS VSS.n1052 0.14207
R3923 VSS.n2601 VSS 0.14207
R3924 VSS.n498 VSS 0.141725
R3925 VSS.n950 VSS 0.141725
R3926 VSS.n2062 VSS 0.141725
R3927 VSS.n1753 VSS 0.141725
R3928 VSS.n2462 VSS 0.141725
R3929 VSS.n2547 VSS.n235 0.137387
R3930 VSS.n2511 VSS.n256 0.137387
R3931 VSS.n2479 VSS.n280 0.137387
R3932 VSS.n2476 VSS.n2475 0.137387
R3933 VSS.n2660 VSS.n2659 0.137387
R3934 VSS.n2663 VSS.n213 0.137387
R3935 VSS.n956 VSS.n955 0.13667
R3936 VSS.n1891 VSS.n999 0.126812
R3937 VSS.n1915 VSS.n1018 0.126812
R3938 VSS.n1771 VSS.n1770 0.126812
R3939 VSS.n1713 VSS.n1083 0.126812
R3940 VSS.n1859 VSS.n1777 0.126812
R3941 VSS.n1803 VSS.n962 0.126812
R3942 VSS.n2361 VSS.n2360 0.126617
R3943 VSS.n2341 VSS.n538 0.125637
R3944 VSS.n900 VSS.n533 0.125637
R3945 VSS.n1256 VSS.n1153 0.125637
R3946 VSS.n1226 VSS.n1131 0.125637
R3947 VSS.n2297 VSS.n2296 0.125637
R3948 VSS.n2293 VSS.n837 0.125637
R3949 VSS.n2831 VSS.n95 0.1255
R3950 VSS.n2702 VSS.n0 0.122556
R3951 VSS.n681 VSS.n680 0.120632
R3952 VSS.n1611 VSS 0.120408
R3953 VSS.n503 VSS.n502 0.120292
R3954 VSS.n503 VSS.n474 0.120292
R3955 VSS.n509 VSS.n474 0.120292
R3956 VSS.n2374 VSS.n2373 0.120292
R3957 VSS.n2373 VSS.n518 0.120292
R3958 VSS.n2369 VSS.n518 0.120292
R3959 VSS.n2369 VSS.n2368 0.120292
R3960 VSS.n2368 VSS.n520 0.120292
R3961 VSS.n2364 VSS.n520 0.120292
R3962 VSS.n2364 VSS.n2363 0.120292
R3963 VSS.n2357 VSS.n2356 0.120292
R3964 VSS.n629 VSS.n612 0.120292
R3965 VSS.n630 VSS.n629 0.120292
R3966 VSS.n631 VSS.n610 0.120292
R3967 VSS.n636 VSS.n610 0.120292
R3968 VSS.n637 VSS.n636 0.120292
R3969 VSS.n637 VSS.n608 0.120292
R3970 VSS.n641 VSS.n608 0.120292
R3971 VSS.n642 VSS.n641 0.120292
R3972 VSS.n652 VSS.n646 0.120292
R3973 VSS.n666 VSS.n599 0.120292
R3974 VSS.n671 VSS.n599 0.120292
R3975 VSS.n672 VSS.n671 0.120292
R3976 VSS.n672 VSS.n597 0.120292
R3977 VSS.n676 VSS.n597 0.120292
R3978 VSS.n678 VSS.n676 0.120292
R3979 VSS.n685 VSS.n684 0.120292
R3980 VSS.n686 VSS.n685 0.120292
R3981 VSS.n704 VSS.n581 0.120292
R3982 VSS.n708 VSS.n581 0.120292
R3983 VSS.n709 VSS.n708 0.120292
R3984 VSS.n710 VSS.n709 0.120292
R3985 VSS.n710 VSS.n578 0.120292
R3986 VSS.n578 VSS.n576 0.120292
R3987 VSS.n715 VSS.n576 0.120292
R3988 VSS.n716 VSS.n715 0.120292
R3989 VSS.n717 VSS.n716 0.120292
R3990 VSS.n717 VSS.n574 0.120292
R3991 VSS.n739 VSS.n724 0.120292
R3992 VSS.n733 VSS.n724 0.120292
R3993 VSS.n1235 VSS.n1234 0.120292
R3994 VSS.n1235 VSS.n1204 0.120292
R3995 VSS.n1241 VSS.n1204 0.120292
R3996 VSS.n1264 VSS.n1263 0.120292
R3997 VSS.n1264 VSS.n1192 0.120292
R3998 VSS.n1269 VSS.n1192 0.120292
R3999 VSS.n1270 VSS.n1269 0.120292
R4000 VSS.n1271 VSS.n1270 0.120292
R4001 VSS.n1271 VSS.n1190 0.120292
R4002 VSS.n1276 VSS.n1190 0.120292
R4003 VSS.n1317 VSS.n1286 0.120292
R4004 VSS.n1312 VSS.n1286 0.120292
R4005 VSS.n1312 VSS.n1311 0.120292
R4006 VSS.n1311 VSS.n1310 0.120292
R4007 VSS.n1310 VSS.n1293 0.120292
R4008 VSS.n1305 VSS.n1293 0.120292
R4009 VSS.n1305 VSS.n1304 0.120292
R4010 VSS.n1304 VSS.n1303 0.120292
R4011 VSS.n1303 VSS.n1295 0.120292
R4012 VSS.n2324 VSS.n2323 0.120292
R4013 VSS.n2323 VSS.n545 0.120292
R4014 VSS.n2319 VSS.n545 0.120292
R4015 VSS.n2319 VSS.n2318 0.120292
R4016 VSS.n2318 VSS.n547 0.120292
R4017 VSS.n2313 VSS.n547 0.120292
R4018 VSS.n2313 VSS.n2312 0.120292
R4019 VSS.n787 VSS.n769 0.120292
R4020 VSS.n788 VSS.n787 0.120292
R4021 VSS VSS.n788 0.120292
R4022 VSS.n794 VSS.n793 0.120292
R4023 VSS.n799 VSS.n765 0.120292
R4024 VSS.n800 VSS.n799 0.120292
R4025 VSS.n822 VSS.n821 0.120292
R4026 VSS.n821 VSS.n807 0.120292
R4027 VSS.n816 VSS.n807 0.120292
R4028 VSS.n816 VSS.n815 0.120292
R4029 VSS.n1375 VSS.n1374 0.120292
R4030 VSS.n1374 VSS.n1143 0.120292
R4031 VSS.n1370 VSS.n1143 0.120292
R4032 VSS.n1370 VSS.n1369 0.120292
R4033 VSS.n1365 VSS.n1364 0.120292
R4034 VSS.n1360 VSS.n1359 0.120292
R4035 VSS.n1347 VSS.n1346 0.120292
R4036 VSS.n1346 VSS.n1345 0.120292
R4037 VSS.n1345 VSS.n1173 0.120292
R4038 VSS.n1341 VSS.n1173 0.120292
R4039 VSS.n1341 VSS.n1340 0.120292
R4040 VSS.n1340 VSS.n1339 0.120292
R4041 VSS.n1186 VSS.n1185 0.120292
R4042 VSS.n2149 VSS.n2148 0.120292
R4043 VSS.n2149 VSS.n888 0.120292
R4044 VSS.n2155 VSS.n888 0.120292
R4045 VSS.n2156 VSS.n2155 0.120292
R4046 VSS.n2156 VSS.n883 0.120292
R4047 VSS.n2161 VSS.n883 0.120292
R4048 VSS.n2162 VSS.n2161 0.120292
R4049 VSS.n2163 VSS.n2162 0.120292
R4050 VSS.n2163 VSS.n880 0.120292
R4051 VSS.n2169 VSS.n880 0.120292
R4052 VSS.n2189 VSS.n871 0.120292
R4053 VSS.n2195 VSS.n2194 0.120292
R4054 VSS.n2195 VSS.n867 0.120292
R4055 VSS.n2202 VSS.n867 0.120292
R4056 VSS.n2230 VSS.n854 0.120292
R4057 VSS.n2236 VSS.n854 0.120292
R4058 VSS.n2237 VSS.n2236 0.120292
R4059 VSS.n2237 VSS.n850 0.120292
R4060 VSS.n2242 VSS.n850 0.120292
R4061 VSS.n2243 VSS.n2242 0.120292
R4062 VSS.n2252 VSS.n848 0.120292
R4063 VSS.n2253 VSS.n2252 0.120292
R4064 VSS.n2254 VSS.n2253 0.120292
R4065 VSS.n2273 VSS.n2272 0.120292
R4066 VSS.n2272 VSS.n2261 0.120292
R4067 VSS.n2266 VSS.n2261 0.120292
R4068 VSS.n1617 VSS.n1616 0.120292
R4069 VSS.n1610 VSS.n1412 0.120292
R4070 VSS.n1605 VSS.n1412 0.120292
R4071 VSS.n1605 VSS.n1604 0.120292
R4072 VSS.n1604 VSS.n1415 0.120292
R4073 VSS.n1596 VSS.n1415 0.120292
R4074 VSS.n1595 VSS.n1594 0.120292
R4075 VSS.n1580 VSS.n1429 0.120292
R4076 VSS.n1574 VSS.n1429 0.120292
R4077 VSS.n1574 VSS.n1573 0.120292
R4078 VSS.n1573 VSS.n1438 0.120292
R4079 VSS.n1566 VSS.n1565 0.120292
R4080 VSS.n1565 VSS.n1441 0.120292
R4081 VSS.n1557 VSS.n1446 0.120292
R4082 VSS.n1537 VSS.n1536 0.120292
R4083 VSS.n1536 VSS.n1464 0.120292
R4084 VSS.n1532 VSS.n1464 0.120292
R4085 VSS.n1532 VSS.n1531 0.120292
R4086 VSS.n1531 VSS.n1530 0.120292
R4087 VSS.n1530 VSS.n1469 0.120292
R4088 VSS.n1505 VSS.n1504 0.120292
R4089 VSS.n1504 VSS.n1479 0.120292
R4090 VSS.n1494 VSS.n1493 0.120292
R4091 VSS.n1493 VSS.n1492 0.120292
R4092 VSS.n2112 VSS.n2111 0.120292
R4093 VSS.n2111 VSS.n2110 0.120292
R4094 VSS.n2110 VSS.n917 0.120292
R4095 VSS.n2106 VSS.n917 0.120292
R4096 VSS.n2106 VSS.n2105 0.120292
R4097 VSS.n2105 VSS.n2104 0.120292
R4098 VSS.n2104 VSS.n922 0.120292
R4099 VSS.n2099 VSS.n922 0.120292
R4100 VSS.n2099 VSS.n2098 0.120292
R4101 VSS.n957 VSS.n938 0.120292
R4102 VSS.n1644 VSS.n1643 0.120292
R4103 VSS.n1654 VSS.n1120 0.120292
R4104 VSS.n1655 VSS.n1654 0.120292
R4105 VSS.n1655 VSS.n1117 0.120292
R4106 VSS.n1117 VSS.n1116 0.120292
R4107 VSS.n1662 VSS.n1661 0.120292
R4108 VSS.n1109 VSS.n1094 0.120292
R4109 VSS.n1105 VSS.n1094 0.120292
R4110 VSS.n1104 VSS.n1103 0.120292
R4111 VSS.n1103 VSS.n1097 0.120292
R4112 VSS.n1948 VSS.n1012 0.120292
R4113 VSS.n1953 VSS.n1012 0.120292
R4114 VSS.n1955 VSS.n1954 0.120292
R4115 VSS.n1962 VSS.n1008 0.120292
R4116 VSS.n1964 VSS.n1006 0.120292
R4117 VSS.n1968 VSS.n1006 0.120292
R4118 VSS.n1969 VSS.n1968 0.120292
R4119 VSS.n1987 VSS.n991 0.120292
R4120 VSS.n1988 VSS.n1987 0.120292
R4121 VSS.n1992 VSS.n989 0.120292
R4122 VSS.n1993 VSS.n1992 0.120292
R4123 VSS.n1993 VSS.n985 0.120292
R4124 VSS.n1997 VSS.n985 0.120292
R4125 VSS.n2030 VSS.n975 0.120292
R4126 VSS.n2031 VSS.n2030 0.120292
R4127 VSS.n2032 VSS.n2031 0.120292
R4128 VSS.n2032 VSS.n973 0.120292
R4129 VSS.n2039 VSS.n973 0.120292
R4130 VSS.n2040 VSS.n2039 0.120292
R4131 VSS.n2041 VSS.n2040 0.120292
R4132 VSS.n2048 VSS.n971 0.120292
R4133 VSS.n2049 VSS.n2048 0.120292
R4134 VSS.n2072 VSS.n2057 0.120292
R4135 VSS.n2068 VSS.n2057 0.120292
R4136 VSS.n2068 VSS.n2067 0.120292
R4137 VSS.n2067 VSS.n2059 0.120292
R4138 VSS.n1723 VSS.n1722 0.120292
R4139 VSS.n1727 VSS.n1692 0.120292
R4140 VSS.n1728 VSS.n1727 0.120292
R4141 VSS.n1729 VSS.n1690 0.120292
R4142 VSS.n1736 VSS.n1690 0.120292
R4143 VSS.n1737 VSS.n1736 0.120292
R4144 VSS.n1755 VSS.n1754 0.120292
R4145 VSS.n1749 VSS.n1748 0.120292
R4146 VSS.n1925 VSS.n1924 0.120292
R4147 VSS.n1907 VSS.n1906 0.120292
R4148 VSS.n1902 VSS.n1901 0.120292
R4149 VSS.n1901 VSS.n1049 0.120292
R4150 VSS.n1884 VSS.n1883 0.120292
R4151 VSS.n1883 VSS.n1069 0.120292
R4152 VSS.n1877 VSS.n1069 0.120292
R4153 VSS.n1875 VSS.n1071 0.120292
R4154 VSS.n1870 VSS.n1869 0.120292
R4155 VSS.n1869 VSS.n1076 0.120292
R4156 VSS.n1855 VSS.n1783 0.120292
R4157 VSS.n1844 VSS.n1843 0.120292
R4158 VSS.n1839 VSS.n1838 0.120292
R4159 VSS.n1838 VSS.n1788 0.120292
R4160 VSS.n1819 VSS.n1807 0.120292
R4161 VSS.n1815 VSS.n1814 0.120292
R4162 VSS.n1814 VSS.n1810 0.120292
R4163 VSS.n2461 VSS.n2403 0.120292
R4164 VSS.n2456 VSS.n2403 0.120292
R4165 VSS.n2456 VSS.n2455 0.120292
R4166 VSS.n2439 VSS.n2419 0.120292
R4167 VSS.n2434 VSS.n2419 0.120292
R4168 VSS.n2434 VSS.n2433 0.120292
R4169 VSS.n2433 VSS.n2432 0.120292
R4170 VSS.n2432 VSS.n2423 0.120292
R4171 VSS.n2428 VSS.n2423 0.120292
R4172 VSS.n2428 VSS.n2427 0.120292
R4173 VSS.n2520 VSS.n249 0.120292
R4174 VSS.n2521 VSS.n2520 0.120292
R4175 VSS.n2522 VSS.n2521 0.120292
R4176 VSS.n2522 VSS.n247 0.120292
R4177 VSS.n2526 VSS.n247 0.120292
R4178 VSS.n2527 VSS.n2526 0.120292
R4179 VSS.n2527 VSS.n245 0.120292
R4180 VSS.n2532 VSS.n245 0.120292
R4181 VSS.n2533 VSS.n2532 0.120292
R4182 VSS.n2552 VSS.n2551 0.120292
R4183 VSS.n2552 VSS.n230 0.120292
R4184 VSS.n2556 VSS.n230 0.120292
R4185 VSS.n2557 VSS.n2556 0.120292
R4186 VSS.n2557 VSS.n228 0.120292
R4187 VSS.n2562 VSS.n228 0.120292
R4188 VSS.n2563 VSS.n2562 0.120292
R4189 VSS.n2571 VSS.n2570 0.120292
R4190 VSS.n2645 VSS.n2644 0.120292
R4191 VSS.n2644 VSS.n2643 0.120292
R4192 VSS.n2643 VSS.n2576 0.120292
R4193 VSS.n2638 VSS.n2576 0.120292
R4194 VSS.n2638 VSS.n2637 0.120292
R4195 VSS.n2637 VSS.n2636 0.120292
R4196 VSS.n2632 VSS.n2631 0.120292
R4197 VSS.n2631 VSS.n2581 0.120292
R4198 VSS.n2627 VSS.n2581 0.120292
R4199 VSS.n2609 VSS.n2608 0.120292
R4200 VSS.n2608 VSS.n2597 0.120292
R4201 VSS.n2602 VSS.n2597 0.120292
R4202 VSS.n2710 VSS.n102 0.120292
R4203 VSS.n2705 VSS.n102 0.120292
R4204 VSS.n2705 VSS.n2704 0.120292
R4205 VSS.n2850 VSS.n69 0.120292
R4206 VSS.n2840 VSS.n76 0.120292
R4207 VSS.n77 VSS.n76 0.120292
R4208 VSS.n2834 VSS.n78 0.120292
R4209 VSS.n92 VSS.n81 0.120292
R4210 VSS.n86 VSS.n81 0.120292
R4211 VSS.n86 VSS.n85 0.120292
R4212 VSS.n2713 VSS.n2712 0.120292
R4213 VSS.n2713 VSS.n100 0.120292
R4214 VSS.n2811 VSS.n2718 0.120292
R4215 VSS.n2811 VSS.n2810 0.120292
R4216 VSS.n2809 VSS.n2720 0.120292
R4217 VSS.n2721 VSS.n2720 0.120292
R4218 VSS.n2802 VSS.n2794 0.120292
R4219 VSS.n2802 VSS.n2801 0.120292
R4220 VSS.n2800 VSS.n2797 0.120292
R4221 VSS.n2797 VSS.n2796 0.120292
R4222 VSS.n2827 VSS.n2826 0.120292
R4223 VSS.n2823 VSS.n2822 0.120292
R4224 VSS.n455 VSS.n285 0.120292
R4225 VSS.n448 VSS.n285 0.120292
R4226 VSS.n447 VSS.n446 0.120292
R4227 VSS.n446 VSS.n288 0.120292
R4228 VSS.n442 VSS.n288 0.120292
R4229 VSS.n442 VSS.n441 0.120292
R4230 VSS.n441 VSS.n440 0.120292
R4231 VSS.n440 VSS.n291 0.120292
R4232 VSS.n433 VSS.n291 0.120292
R4233 VSS.n2485 VSS.n2484 0.120292
R4234 VSS.n2485 VSS.n273 0.120292
R4235 VSS.n2489 VSS.n273 0.120292
R4236 VSS.n2490 VSS.n2489 0.120292
R4237 VSS.n2490 VSS.n271 0.120292
R4238 VSS.n2494 VSS.n271 0.120292
R4239 VSS.n2495 VSS.n2494 0.120292
R4240 VSS.n329 VSS.n324 0.120292
R4241 VSS.n404 VSS.n320 0.120292
R4242 VSS.n400 VSS.n320 0.120292
R4243 VSS.n400 VSS.n399 0.120292
R4244 VSS.n399 VSS.n398 0.120292
R4245 VSS.n398 VSS.n343 0.120292
R4246 VSS.n393 VSS.n343 0.120292
R4247 VSS.n393 VSS.n392 0.120292
R4248 VSS.n392 VSS.n391 0.120292
R4249 VSS.n391 VSS 0.120292
R4250 VSS.n386 VSS.n385 0.120292
R4251 VSS.n374 VSS.n358 0.120292
R4252 VSS.n370 VSS.n358 0.120292
R4253 VSS.n370 VSS.n369 0.120292
R4254 VSS.n369 VSS.n368 0.120292
R4255 VSS.n368 VSS.n360 0.120292
R4256 VSS.n364 VSS.n360 0.120292
R4257 VSS.n364 VSS.n363 0.120292
R4258 VSS.n2679 VSS.n2678 0.120292
R4259 VSS.n158 VSS.n145 0.120292
R4260 VSS.n166 VSS.n145 0.120292
R4261 VSS.n167 VSS.n166 0.120292
R4262 VSS.n172 VSS.n171 0.120292
R4263 VSS.n177 VSS.n141 0.120292
R4264 VSS.n178 VSS.n177 0.120292
R4265 VSS.n179 VSS.n178 0.120292
R4266 VSS.n203 VSS.n202 0.120292
R4267 VSS.n202 VSS.n185 0.120292
R4268 VSS.n198 VSS.n185 0.120292
R4269 VSS.n198 VSS.n197 0.120292
R4270 VSS.n194 VSS.n193 0.120292
R4271 VSS.n193 VSS.n189 0.120292
R4272 VSS.n2130 VSS.n904 0.120125
R4273 VSS.n2130 VSS.n2129 0.120125
R4274 VSS.n2129 VSS.n2128 0.120125
R4275 VSS.n2128 VSS.n905 0.120125
R4276 VSS.n1773 VSS.n1772 0.120125
R4277 VSS.n1774 VSS.n1773 0.120125
R4278 VSS.n1776 VSS.n1774 0.120125
R4279 VSS.n1776 VSS.n1775 0.120125
R4280 VSS.n2390 VSS.n462 0.120125
R4281 VSS.n562 VSS.n462 0.120125
R4282 VSS.n563 VSS.n562 0.120125
R4283 VSS.n564 VSS.n563 0.120125
R4284 VSS.n2344 VSS.n534 0.120125
R4285 VSS.n2344 VSS.n2343 0.120125
R4286 VSS.n2343 VSS.n535 0.120125
R4287 VSS.n756 VSS.n535 0.120125
R4288 VSS.n1152 VSS.n1151 0.120125
R4289 VSS.n1151 VSS.n561 0.120125
R4290 VSS.n2295 VSS.n561 0.120125
R4291 VSS.n2295 VSS.n2294 0.120125
R4292 VSS.n2478 VSS.n2477 0.120125
R4293 VSS.n2477 VSS.n214 0.120125
R4294 VSS.n2661 VSS.n214 0.120125
R4295 VSS.n2662 VSS.n2661 0.120125
R4296 VSS.n2701 VSS 0.114397
R4297 VSS.n2774 VSS.n2734 0.113648
R4298 VSS.n60 VSS.n10 0.111077
R4299 VSS.n55 VSS.n54 0.111077
R4300 VSS.n50 VSS.n49 0.111077
R4301 VSS.n45 VSS.n44 0.111077
R4302 VSS.n40 VSS.n39 0.111077
R4303 VSS.n35 VSS.n34 0.111077
R4304 VSS.n30 VSS.n29 0.111077
R4305 VSS.n25 VSS.n24 0.111077
R4306 VSS.n20 VSS.n19 0.111077
R4307 VSS.n554 VSS.n553 0.109992
R4308 VSS.n414 VSS.n128 0.10744
R4309 VSS.n536 VSS.n236 0.103312
R4310 VSS.n2346 VSS.n257 0.103312
R4311 VSS.n2389 VSS.n2388 0.103312
R4312 VSS.n2391 VSS.n461 0.103312
R4313 VSS.n700 VSS.n216 0.103312
R4314 VSS.n755 VSS.n565 0.103312
R4315 VSS.n1351 VSS.n1350 0.102062
R4316 VSS.n1581 VSS.n1580 0.102062
R4317 VSS.n1111 VSS.n1092 0.102062
R4318 VSS.n1755 VSS.n1686 0.102062
R4319 VSS.n2484 VSS.n2483 0.102062
R4320 VSS.n2374 VSS 0.0981562
R4321 VSS.n2358 VSS 0.0981562
R4322 VSS.n646 VSS 0.0981562
R4323 VSS.n666 VSS 0.0981562
R4324 VSS VSS.n677 0.0981562
R4325 VSS.n1263 VSS 0.0981562
R4326 VSS.n1330 VSS 0.0981562
R4327 VSS.n2309 VSS 0.0981562
R4328 VSS VSS.n765 0.0981562
R4329 VSS VSS.n1365 0.0981562
R4330 VSS.n2148 VSS 0.0981562
R4331 VSS.n2212 VSS 0.0981562
R4332 VSS VSS.n848 0.0981562
R4333 VSS.n1525 VSS 0.0981562
R4334 VSS.n1650 VSS 0.0981562
R4335 VSS VSS.n1109 0.0981562
R4336 VSS.n1964 VSS 0.0981562
R4337 VSS.n2006 VSS 0.0981562
R4338 VSS VSS.n2439 0.0981562
R4339 VSS VSS.n266 0.0981562
R4340 VSS.n2566 VSS 0.0981562
R4341 VSS.n2632 VSS 0.0981562
R4342 VSS VSS.n2850 0.0981562
R4343 VSS VSS.n269 0.0981562
R4344 VSS.n386 VSS 0.0981562
R4345 VSS.n2680 VSS 0.0981562
R4346 VSS.n194 VSS 0.0981562
R4347 VSS.n704 VSS.n703 0.0968542
R4348 VSS.n780 VSS.n779 0.0968542
R4349 VSS.n2230 VSS.n2229 0.0968542
R4350 VSS VSS.n1537 0.0968542
R4351 VSS.n1661 VSS 0.0968542
R4352 VSS.n1856 VSS.n1855 0.0968542
R4353 VSS.n2645 VSS.n223 0.0968542
R4354 VSS.n158 VSS.n157 0.0968542
R4355 VSS.n1722 VSS 0.0955521
R4356 VSS VSS.n1688 0.0955521
R4357 VSS.n1749 VSS 0.0955521
R4358 VSS VSS.n1907 0.0955521
R4359 VSS VSS.n1875 0.0955521
R4360 VSS VSS.n1844 0.0955521
R4361 VSS VSS.n1819 0.0955521
R4362 VSS.n171 VSS 0.0955521
R4363 VSS.n2673 VSS.n127 0.0950946
R4364 VSS.n154 VSS.n132 0.0950946
R4365 VSS.n211 VSS.n210 0.0950946
R4366 VSS.n183 VSS.n135 0.0950946
R4367 VSS.n2657 VSS.n2656 0.0950946
R4368 VSS.n2650 VSS.n222 0.0950946
R4369 VSS.n1801 VSS.n1800 0.0950946
R4370 VSS.n1826 VSS.n1796 0.0950946
R4371 VSS.n2009 VSS.n2007 0.0950946
R4372 VSS.n2022 VSS.n979 0.0950946
R4373 VSS.n300 VSS.n297 0.0950946
R4374 VSS.n457 VSS.n284 0.0950946
R4375 VSS.n2473 VSS.n2472 0.0950946
R4376 VSS.n2465 VSS.n2464 0.0950946
R4377 VSS.n1711 VSS.n1710 0.0950946
R4378 VSS.n1716 VSS.n1715 0.0950946
R4379 VSS.n2447 VSS.n2412 0.0950946
R4380 VSS.n2441 VSS.n2415 0.0950946
R4381 VSS.n2124 VSS.n2123 0.0950946
R4382 VSS.n2117 VSS.n913 0.0950946
R4383 VSS.n1623 VSS.n1622 0.0950946
R4384 VSS.n1409 VSS.n1408 0.0950946
R4385 VSS.n2092 VSS.n930 0.0950946
R4386 VSS.n959 VSS.n934 0.0950946
R4387 VSS.n1391 VSS.n1390 0.0950946
R4388 VSS.n1383 VSS.n1382 0.0950946
R4389 VSS.n2290 VSS.n2289 0.0950946
R4390 VSS.n2282 VSS.n2281 0.0950946
R4391 VSS.n2215 VSS.n2213 0.0950946
R4392 VSS.n2228 VSS.n858 0.0950946
R4393 VSS.n333 VSS.n323 0.0950946
R4394 VSS.n406 VSS.n318 0.0950946
R4395 VSS.n2509 VSS.n2508 0.0950946
R4396 VSS.n2513 VSS.n254 0.0950946
R4397 VSS.n353 VSS.n352 0.0950946
R4398 VSS.n376 VSS.n351 0.0950946
R4399 VSS.n2545 VSS.n2544 0.0950946
R4400 VSS.n2549 VSS.n233 0.0950946
R4401 VSS.n1254 VSS.n1253 0.0950946
R4402 VSS.n1258 VSS.n1196 0.0950946
R4403 VSS.n1224 VSS.n1223 0.0950946
R4404 VSS.n1228 VSS.n1210 0.0950946
R4405 VSS.n835 VSS.n834 0.0950946
R4406 VSS.n827 VSS.n826 0.0950946
R4407 VSS.n2301 VSS.n555 0.0950946
R4408 VSS.n778 VSS.n777 0.0950946
R4409 VSS.n1324 VSS.n1282 0.0950946
R4410 VSS.n1318 VSS.n1285 0.0950946
R4411 VSS.n2386 VSS.n2385 0.0950946
R4412 VSS.n2379 VSS.n470 0.0950946
R4413 VSS.n486 VSS.n485 0.0950946
R4414 VSS.n496 VSS.n480 0.0950946
R4415 VSS.n753 VSS.n752 0.0950946
R4416 VSS.n745 VSS.n744 0.0950946
R4417 VSS.n698 VSS.n697 0.0950946
R4418 VSS.n702 VSS.n586 0.0950946
R4419 VSS.n650 VSS.n648 0.0950946
R4420 VSS.n663 VSS.n602 0.0950946
R4421 VSS.n2350 VSS.n529 0.0950946
R4422 VSS.n619 VSS.n618 0.0950946
R4423 VSS.n2339 VSS.n2338 0.0950946
R4424 VSS.n2330 VSS.n2329 0.0950946
R4425 VSS.n2176 VSS.n2175 0.0950946
R4426 VSS.n2181 VSS.n2180 0.0950946
R4427 VSS.n1512 VSS.n1511 0.0950946
R4428 VSS.n1518 VSS.n1517 0.0950946
R4429 VSS.n1976 VSS.n1975 0.0950946
R4430 VSS.n1981 VSS.n1980 0.0950946
R4431 VSS.n1893 VSS.n1055 0.0950946
R4432 VSS.n1889 VSS.n1058 0.0950946
R4433 VSS.n1549 VSS.n1452 0.0950946
R4434 VSS.n1543 VSS.n1455 0.0950946
R4435 VSS.n1942 VSS.n1941 0.0950946
R4436 VSS.n1946 VSS.n1016 0.0950946
R4437 VSS.n1919 VSS.n1038 0.0950946
R4438 VSS.n1913 VSS.n1042 0.0950946
R4439 VSS.n1182 VSS.n1181 0.0950946
R4440 VSS.n2133 VSS.n898 0.0950946
R4441 VSS.n1357 VSS.n1149 0.0950946
R4442 VSS.n1352 VSS.n1155 0.0950946
R4443 VSS.n1588 VSS.n1424 0.0950946
R4444 VSS.n1582 VSS.n1427 0.0950946
R4445 VSS.n1676 VSS.n1675 0.0950946
R4446 VSS.n1669 VSS.n1091 0.0950946
R4447 VSS.n1768 VSS.n1767 0.0950946
R4448 VSS.n1761 VSS.n1685 0.0950946
R4449 VSS.n1639 VSS.n1130 0.0950946
R4450 VSS.n1630 VSS.n1629 0.0950946
R4451 VSS.n2085 VSS.n2084 0.0950946
R4452 VSS.n2077 VSS.n2076 0.0950946
R4453 VSS.n1863 VSS.n1080 0.0950946
R4454 VSS.n1857 VSS.n1779 0.0950946
R4455 VSS.n2625 VSS.n2585 0.0950946
R4456 VSS.n2618 VSS.n2617 0.0950946
R4457 VSS.n430 VSS.n429 0.0950946
R4458 VSS.n2482 VSS.n276 0.0950946
R4459 VSS.n2711 VSS 0.09425
R4460 VSS.n574 VSS.n568 0.0916458
R4461 VSS.n2254 VSS.n841 0.0916458
R4462 VSS.n928 VSS.n926 0.0916458
R4463 VSS.n2627 VSS.n2626 0.0916458
R4464 VSS.n179 VSS.n136 0.0916458
R4465 VSS.n2342 VSS.n536 0.0915625
R4466 VSS.n2346 VSS.n2345 0.0915625
R4467 VSS.n2388 VSS.n464 0.0915625
R4468 VSS.n1212 VSS.n461 0.0915625
R4469 VSS.n700 VSS.n558 0.0915625
R4470 VSS.n757 VSS.n755 0.0915625
R4471 VSS.n2699 VSS 0.0907344
R4472 VSS VSS.n60 0.0906442
R4473 VSS.n55 VSS 0.0906442
R4474 VSS.n50 VSS 0.0906442
R4475 VSS.n45 VSS 0.0906442
R4476 VSS.n40 VSS 0.0906442
R4477 VSS.n35 VSS 0.0906442
R4478 VSS.n30 VSS 0.0906442
R4479 VSS.n25 VSS 0.0906442
R4480 VSS.n20 VSS 0.0906442
R4481 VSS.n782 VSS.n781 0.0900105
R4482 VSS.n2633 VSS.n2580 0.0900105
R4483 VSS.n413 VSS.n410 0.0898892
R4484 VSS.n415 VSS.n414 0.0898892
R4485 VSS.n2818 VSS 0.0881354
R4486 VSS.n2356 VSS.n524 0.0864375
R4487 VSS.n1328 VSS.n1277 0.0864375
R4488 VSS.n1450 VSS.n1446 0.0864375
R4489 VSS.n1924 VSS.n1033 0.0864375
R4490 VSS.n2504 VSS.n259 0.0864375
R4491 VSS.n330 VSS.n329 0.0864375
R4492 VSS.n2384 VSS.n2383 0.0838333
R4493 VSS.n616 VSS.n615 0.0838333
R4494 VSS.n651 VSS.n647 0.0838333
R4495 VSS.n664 VSS.n601 0.0838333
R4496 VSS.n723 VSS.n571 0.0838333
R4497 VSS.n1252 VSS.n1251 0.0838333
R4498 VSS.n1288 VSS.n1287 0.0838333
R4499 VSS.n2331 VSS.n2325 0.0838333
R4500 VSS.n806 VSS.n763 0.0838333
R4501 VSS.n1165 VSS.n1161 0.0838333
R4502 VSS.n2138 VSS.n896 0.0838333
R4503 VSS.n2174 VSS.n2170 0.0838333
R4504 VSS.n2182 VSS.n875 0.0838333
R4505 VSS.n2223 VSS.n861 0.0838333
R4506 VSS.n2259 VSS.n844 0.0838333
R4507 VSS.n1589 VSS.n1423 0.0838333
R4508 VSS.n1457 VSS.n1456 0.0838333
R4509 VSS.n1510 VSS.n1475 0.0838333
R4510 VSS.n1519 VSS.n1506 0.0838333
R4511 VSS.n2122 VSS.n2121 0.0838333
R4512 VSS.n1674 VSS.n1673 0.0838333
R4513 VSS.n1026 VSS.n1023 0.0838333
R4514 VSS.n1982 VSS.n995 0.0838333
R4515 VSS.n2017 VSS.n982 0.0838333
R4516 VSS.n1044 VSS.n1043 0.0838333
R4517 VSS.n1864 VSS.n1079 0.0838333
R4518 VSS.n2448 VSS.n2411 0.0838333
R4519 VSS.n261 VSS.n253 0.0838333
R4520 VSS.n2550 VSS.n232 0.0838333
R4521 VSS.n2655 VSS.n2654 0.0838333
R4522 VSS.n2620 VSS.n2619 0.0838333
R4523 VSS.n428 VSS.n427 0.0838333
R4524 VSS.n337 VSS.n322 0.0838333
R4525 VSS.n348 VSS.n346 0.0838333
R4526 VSS.n375 VSS.n357 0.0838333
R4527 VSS.n150 VSS.n148 0.0838333
R4528 VSS.n184 VSS.n139 0.0838333
R4529 VSS.n905 VSS 0.0827875
R4530 VSS.n1775 VSS 0.0827875
R4531 VSS.n564 VSS 0.0827875
R4532 VSS.n756 VSS 0.0827875
R4533 VSS.n2294 VSS 0.0827875
R4534 VSS.n2662 VSS 0.0827875
R4535 VSS VSS.n945 0.082648
R4536 VSS.n1611 VSS 0.082648
R4537 VSS.n1804 VSS 0.0773229
R4538 VSS.n468 VSS.n466 0.0760208
R4539 VSS.n1201 VSS.n1199 0.0760208
R4540 VSS.n1358 VSS.n1148 0.0760208
R4541 VSS.n1590 VSS.n1419 0.0760208
R4542 VSS.n1089 VSS.n1087 0.0760208
R4543 VSS.n1683 VSS.n1681 0.0760208
R4544 VSS.n2449 VSS.n2408 0.0760208
R4545 VSS.n431 VSS.n296 0.0760208
R4546 VSS.n2698 VSS.n2697 0.0747188
R4547 VSS.n2823 VSS.n2819 0.0721146
R4548 VSS.n491 VSS.n490 0.0708125
R4549 VSS.n2351 VSS.n528 0.0708125
R4550 VSS.n591 VSS.n589 0.0708125
R4551 VSS.n1220 VSS.n1217 0.0708125
R4552 VSS.n1325 VSS.n1281 0.0708125
R4553 VSS.n2303 VSS.n554 0.0708125
R4554 VSS.n1385 VSS.n1136 0.0708125
R4555 VSS.n2139 VSS.n895 0.0708125
R4556 VSS.n2217 VSS.n2216 0.0708125
R4557 VSS.n1401 VSS.n1399 0.0708125
R4558 VSS.n1550 VSS.n1451 0.0708125
R4559 VSS.n911 VSS.n909 0.0708125
R4560 VSS.n1634 VSS.n1126 0.0708125
R4561 VSS.n1940 VSS.n1939 0.0708125
R4562 VSS.n1718 VSS.n1698 0.0708125
R4563 VSS.n1920 VSS.n1037 0.0708125
R4564 VSS.n1865 VSS.n1078 0.0708125
R4565 VSS.n2467 VSS.n2395 0.0708125
R4566 VSS.n2507 VSS.n250 0.0708125
R4567 VSS.n220 VSS.n218 0.0708125
R4568 VSS.n2842 VSS.n75 0.0708125
R4569 VSS.n309 VSS.n308 0.0708125
R4570 VSS.n2674 VSS.n126 0.0708125
R4571 VSS.n2337 VSS 0.0695104
R4572 VSS.n2543 VSS 0.0695104
R4573 VSS.n2342 VSS.n2341 0.0692375
R4574 VSS.n2345 VSS.n533 0.0692375
R4575 VSS.n1256 VSS.n464 0.0692375
R4576 VSS.n1226 VSS.n1212 0.0692375
R4577 VSS.n2297 VSS.n558 0.0692375
R4578 VSS.n837 VSS.n757 0.0692375
R4579 VSS.n2200 VSS.n2199 0.0685851
R4580 VSS.n1297 VSS.n540 0.068325
R4581 VSS.n243 VSS.n238 0.068325
R4582 VSS.n149 VSS.n130 0.0680676
R4583 VSS.n149 VSS.n131 0.0680676
R4584 VSS.n138 VSS.n134 0.0680676
R4585 VSS.n138 VSS.n133 0.0680676
R4586 VSS.n2653 VSS.n219 0.0680676
R4587 VSS.n2653 VSS.n2652 0.0680676
R4588 VSS.n1830 VSS.n1795 0.0680676
R4589 VSS.n1830 VSS.n1829 0.0680676
R4590 VSS.n2018 VSS.n981 0.0680676
R4591 VSS.n2019 VSS.n2018 0.0680676
R4592 VSS.n311 VSS.n310 0.0680676
R4593 VSS.n310 VSS.n298 0.0680676
R4594 VSS.n2400 VSS.n2394 0.0680676
R4595 VSS.n2402 VSS.n2400 0.0680676
R4596 VSS.n1704 VSS.n1703 0.0680676
R4597 VSS.n1703 VSS.n1699 0.0680676
R4598 VSS.n2446 VSS.n2413 0.0680676
R4599 VSS.n2414 VSS.n2413 0.0680676
R4600 VSS.n2120 VSS.n910 0.0680676
R4601 VSS.n2120 VSS.n2119 0.0680676
R4602 VSS.n1404 VSS.n1398 0.0680676
R4603 VSS.n1406 VSS.n1404 0.0680676
R4604 VSS.n2091 VSS.n931 0.0680676
R4605 VSS.n933 VSS.n931 0.0680676
R4606 VSS.n1139 VSS.n1135 0.0680676
R4607 VSS.n1141 VSS.n1139 0.0680676
R4608 VSS.n2278 VSS.n842 0.0680676
R4609 VSS.n2280 VSS.n2278 0.0680676
R4610 VSS.n2224 VSS.n860 0.0680676
R4611 VSS.n2225 VSS.n2224 0.0680676
R4612 VSS.n336 VSS.n334 0.0680676
R4613 VSS.n336 VSS.n335 0.0680676
R4614 VSS.n263 VSS.n262 0.0680676
R4615 VSS.n262 VSS.n260 0.0680676
R4616 VSS.n380 VSS.n350 0.0680676
R4617 VSS.n380 VSS.n379 0.0680676
R4618 VSS.n241 VSS.n239 0.0680676
R4619 VSS.n241 VSS.n240 0.0680676
R4620 VSS.n1250 VSS.n1200 0.0680676
R4621 VSS.n1250 VSS.n1249 0.0680676
R4622 VSS.n1219 VSS.n1215 0.0680676
R4623 VSS.n1219 VSS.n1218 0.0680676
R4624 VSS.n823 VSS.n761 0.0680676
R4625 VSS.n825 VSS.n823 0.0680676
R4626 VSS.n2300 VSS.n556 0.0680676
R4627 VSS.n772 VSS.n556 0.0680676
R4628 VSS.n1323 VSS.n1283 0.0680676
R4629 VSS.n1284 VSS.n1283 0.0680676
R4630 VSS.n2382 VSS.n467 0.0680676
R4631 VSS.n2382 VSS.n2381 0.0680676
R4632 VSS.n492 VSS.n482 0.0680676
R4633 VSS.n493 VSS.n492 0.0680676
R4634 VSS.n741 VSS.n569 0.0680676
R4635 VSS.n743 VSS.n741 0.0680676
R4636 VSS.n694 VSS.n590 0.0680676
R4637 VSS.n694 VSS.n693 0.0680676
R4638 VSS.n659 VSS.n604 0.0680676
R4639 VSS.n660 VSS.n659 0.0680676
R4640 VSS.n2349 VSS.n530 0.0680676
R4641 VSS.n617 VSS.n530 0.0680676
R4642 VSS.n2326 VSS.n541 0.0680676
R4643 VSS.n2328 VSS.n2326 0.0680676
R4644 VSS.n2172 VSS.n2171 0.0680676
R4645 VSS.n2171 VSS.n876 0.0680676
R4646 VSS.n1509 VSS.n1508 0.0680676
R4647 VSS.n1508 VSS.n1507 0.0680676
R4648 VSS.n1003 VSS.n1002 0.0680676
R4649 VSS.n1002 VSS.n996 0.0680676
R4650 VSS.n1063 VSS.n1061 0.0680676
R4651 VSS.n1063 VSS.n1062 0.0680676
R4652 VSS.n1548 VSS.n1453 0.0680676
R4653 VSS.n1454 VSS.n1453 0.0680676
R4654 VSS.n1025 VSS.n1021 0.0680676
R4655 VSS.n1025 VSS.n1024 0.0680676
R4656 VSS.n1918 VSS.n1039 0.0680676
R4657 VSS.n1041 VSS.n1039 0.0680676
R4658 VSS.n2137 VSS.n897 0.0680676
R4659 VSS.n2137 VSS.n2136 0.0680676
R4660 VSS.n1164 VSS.n1162 0.0680676
R4661 VSS.n1164 VSS.n1163 0.0680676
R4662 VSS.n1587 VSS.n1425 0.0680676
R4663 VSS.n1426 VSS.n1425 0.0680676
R4664 VSS.n1672 VSS.n1088 0.0680676
R4665 VSS.n1672 VSS.n1671 0.0680676
R4666 VSS.n1764 VSS.n1682 0.0680676
R4667 VSS.n1764 VSS.n1763 0.0680676
R4668 VSS.n1636 VSS.n1635 0.0680676
R4669 VSS.n1635 VSS.n1633 0.0680676
R4670 VSS.n2073 VSS.n965 0.0680676
R4671 VSS.n2075 VSS.n2073 0.0680676
R4672 VSS.n1862 VSS.n1081 0.0680676
R4673 VSS.n1778 VSS.n1081 0.0680676
R4674 VSS.n2622 VSS.n2621 0.0680676
R4675 VSS.n2621 VSS.n2587 0.0680676
R4676 VSS.n426 VSS.n418 0.0680676
R4677 VSS.n426 VSS.n425 0.0680676
R4678 VSS.n1059 VSS 0.0669062
R4679 VSS.n2378 VSS.n2377 0.0656042
R4680 VSS.n658 VSS.n657 0.0656042
R4681 VSS.n751 VSS.n750 0.0656042
R4682 VSS.n1260 VSS.n1195 0.0656042
R4683 VSS.n2332 VSS.n542 0.0656042
R4684 VSS.n833 VSS.n832 0.0656042
R4685 VSS.n829 VSS.n828 0.0656042
R4686 VSS.n1166 VSS.n1156 0.0656042
R4687 VSS.n2183 VSS.n874 0.0656042
R4688 VSS.n2288 VSS.n2287 0.0656042
R4689 VSS.n2284 VSS.n2283 0.0656042
R4690 VSS.n1430 VSS.n1428 0.0656042
R4691 VSS.n1520 VSS.n1478 0.0656042
R4692 VSS.n2093 VSS.n929 0.0656042
R4693 VSS.n958 VSS.n937 0.0656042
R4694 VSS.n1668 VSS.n1667 0.0656042
R4695 VSS.n1983 VSS.n994 0.0656042
R4696 VSS.n2083 VSS.n2082 0.0656042
R4697 VSS.n2079 VSS.n2078 0.0656042
R4698 VSS.n1066 VSS.n1064 0.0656042
R4699 VSS.n1825 VSS.n1805 0.0656042
R4700 VSS.n2418 VSS.n2417 0.0656042
R4701 VSS.n2538 VSS.n242 0.0656042
R4702 VSS.n2589 VSS.n2588 0.0656042
R4703 VSS.n419 VSS.n275 0.0656042
R4704 VSS.n381 VSS.n349 0.0656042
R4705 VSS.n209 VSS.n208 0.0656042
R4706 VSS.n205 VSS.n204 0.0656042
R4707 VSS.n2775 VSS 0.064875
R4708 VSS.n2735 VSS 0.064875
R4709 VSS.n2772 VSS 0.064875
R4710 VSS.n2733 VSS 0.064875
R4711 VSS.n487 VSS 0.0643021
R4712 VSS.n1222 VSS 0.0643021
R4713 VSS.n1389 VSS 0.0643021
R4714 VSS.n1621 VSS 0.0643021
R4715 VSS.n1129 VSS 0.0643021
R4716 VSS VSS.n1020 0.0643021
R4717 VSS.n1709 VSS 0.0643021
R4718 VSS.n2471 VSS 0.0643021
R4719 VSS VSS.n299 0.0643021
R4720 VSS.n2816 VSS.n100 0.0616979
R4721 VSS.n502 VSS 0.0603958
R4722 VSS.n511 VSS 0.0603958
R4723 VSS VSS.n2357 0.0603958
R4724 VSS.n621 VSS.n620 0.0603958
R4725 VSS.n620 VSS.n612 0.0603958
R4726 VSS.n631 VSS 0.0603958
R4727 VSS.n684 VSS 0.0603958
R4728 VSS.n592 VSS.n585 0.0603958
R4729 VSS.n747 VSS 0.0603958
R4730 VSS VSS.n739 0.0603958
R4731 VSS.n733 VSS 0.0603958
R4732 VSS VSS.n732 0.0603958
R4733 VSS.n1234 VSS 0.0603958
R4734 VSS.n1243 VSS 0.0603958
R4735 VSS VSS.n1329 0.0603958
R4736 VSS VSS.n1328 0.0603958
R4737 VSS VSS.n1317 0.0603958
R4738 VSS VSS.n2308 0.0603958
R4739 VSS.n776 VSS.n775 0.0603958
R4740 VSS.n776 VSS.n771 0.0603958
R4741 VSS VSS.n769 0.0603958
R4742 VSS.n793 VSS 0.0603958
R4743 VSS.n801 VSS 0.0603958
R4744 VSS VSS.n1379 0.0603958
R4745 VSS.n1375 VSS 0.0603958
R4746 VSS.n1366 VSS 0.0603958
R4747 VSS.n1364 VSS 0.0603958
R4748 VSS.n1360 VSS 0.0603958
R4749 VSS.n1347 VSS 0.0603958
R4750 VSS.n1178 VSS 0.0603958
R4751 VSS.n1186 VSS 0.0603958
R4752 VSS.n892 VSS 0.0603958
R4753 VSS.n2147 VSS 0.0603958
R4754 VSS VSS.n2189 0.0603958
R4755 VSS.n2190 VSS 0.0603958
R4756 VSS VSS.n2190 0.0603958
R4757 VSS.n2191 VSS 0.0603958
R4758 VSS.n2194 VSS 0.0603958
R4759 VSS.n2203 VSS 0.0603958
R4760 VSS.n2205 VSS 0.0603958
R4761 VSS VSS.n2204 0.0603958
R4762 VSS.n2222 VSS.n862 0.0603958
R4763 VSS.n862 VSS.n857 0.0603958
R4764 VSS.n2277 VSS 0.0603958
R4765 VSS.n2273 VSS 0.0603958
R4766 VSS VSS.n1610 0.0603958
R4767 VSS VSS.n1595 0.0603958
R4768 VSS.n1566 VSS 0.0603958
R4769 VSS.n1558 VSS 0.0603958
R4770 VSS VSS.n1557 0.0603958
R4771 VSS.n1542 VSS.n1458 0.0603958
R4772 VSS.n1542 VSS.n1541 0.0603958
R4773 VSS.n1538 VSS 0.0603958
R4774 VSS VSS.n1469 0.0603958
R4775 VSS.n1471 VSS 0.0603958
R4776 VSS VSS.n1524 0.0603958
R4777 VSS VSS.n1479 0.0603958
R4778 VSS.n1500 VSS 0.0603958
R4779 VSS VSS.n1498 0.0603958
R4780 VSS.n1494 VSS 0.0603958
R4781 VSS.n2116 VSS.n912 0.0603958
R4782 VSS.n2116 VSS.n2115 0.0603958
R4783 VSS.n2112 VSS 0.0603958
R4784 VSS.n926 VSS 0.0603958
R4785 VSS.n946 VSS 0.0603958
R4786 VSS.n1649 VSS 0.0603958
R4787 VSS VSS.n1120 0.0603958
R4788 VSS.n1116 VSS 0.0603958
R4789 VSS.n1660 VSS 0.0603958
R4790 VSS.n1111 VSS 0.0603958
R4791 VSS VSS.n1110 0.0603958
R4792 VSS VSS.n1104 0.0603958
R4793 VSS.n1097 VSS 0.0603958
R4794 VSS.n1933 VSS 0.0603958
R4795 VSS.n1934 VSS 0.0603958
R4796 VSS.n1935 VSS 0.0603958
R4797 VSS.n1947 VSS.n1015 0.0603958
R4798 VSS.n1948 VSS.n1947 0.0603958
R4799 VSS VSS.n1953 0.0603958
R4800 VSS.n1954 VSS 0.0603958
R4801 VSS VSS.n1008 0.0603958
R4802 VSS.n1963 VSS 0.0603958
R4803 VSS VSS.n989 0.0603958
R4804 VSS.n1998 VSS 0.0603958
R4805 VSS.n1999 VSS 0.0603958
R4806 VSS.n2005 VSS 0.0603958
R4807 VSS.n2011 VSS 0.0603958
R4808 VSS.n2016 VSS.n978 0.0603958
R4809 VSS.n2024 VSS.n978 0.0603958
R4810 VSS VSS.n975 0.0603958
R4811 VSS VSS.n971 0.0603958
R4812 VSS.n1723 VSS 0.0603958
R4813 VSS VSS.n1692 0.0603958
R4814 VSS.n1729 VSS 0.0603958
R4815 VSS.n1738 VSS 0.0603958
R4816 VSS VSS.n1759 0.0603958
R4817 VSS VSS.n1752 0.0603958
R4818 VSS.n1748 VSS 0.0603958
R4819 VSS.n1926 VSS 0.0603958
R4820 VSS VSS.n1925 0.0603958
R4821 VSS.n1912 VSS.n1045 0.0603958
R4822 VSS.n1912 VSS.n1911 0.0603958
R4823 VSS.n1908 VSS 0.0603958
R4824 VSS.n1906 VSS 0.0603958
R4825 VSS.n1903 VSS 0.0603958
R4826 VSS VSS.n1902 0.0603958
R4827 VSS.n1895 VSS 0.0603958
R4828 VSS.n1884 VSS 0.0603958
R4829 VSS VSS.n1876 0.0603958
R4830 VSS VSS.n1071 0.0603958
R4831 VSS.n1074 VSS 0.0603958
R4832 VSS.n1870 VSS 0.0603958
R4833 VSS.n1781 VSS.n1780 0.0603958
R4834 VSS.n1782 VSS.n1781 0.0603958
R4835 VSS.n1845 VSS 0.0603958
R4836 VSS.n1843 VSS 0.0603958
R4837 VSS.n1840 VSS 0.0603958
R4838 VSS VSS.n1839 0.0603958
R4839 VSS.n1832 VSS 0.0603958
R4840 VSS.n1824 VSS 0.0603958
R4841 VSS.n1821 VSS 0.0603958
R4842 VSS VSS.n1820 0.0603958
R4843 VSS VSS.n1807 0.0603958
R4844 VSS.n1815 VSS 0.0603958
R4845 VSS VSS.n2461 0.0603958
R4846 VSS VSS.n2453 0.0603958
R4847 VSS.n2503 VSS 0.0603958
R4848 VSS.n2504 VSS 0.0603958
R4849 VSS VSS.n249 0.0603958
R4850 VSS.n2567 VSS 0.0603958
R4851 VSS.n2570 VSS 0.0603958
R4852 VSS.n2649 VSS.n221 0.0603958
R4853 VSS.n2649 VSS.n2648 0.0603958
R4854 VSS.n2609 VSS 0.0603958
R4855 VSS.n2704 VSS 0.0603958
R4856 VSS.n2851 VSS 0.0603958
R4857 VSS.n71 VSS 0.0603958
R4858 VSS.n72 VSS 0.0603958
R4859 VSS.n2842 VSS 0.0603958
R4860 VSS VSS.n2841 0.0603958
R4861 VSS VSS.n2840 0.0603958
R4862 VSS.n78 VSS 0.0603958
R4863 VSS.n2834 VSS 0.0603958
R4864 VSS VSS.n92 0.0603958
R4865 VSS.n2718 VSS 0.0603958
R4866 VSS VSS.n2809 0.0603958
R4867 VSS.n2793 VSS 0.0603958
R4868 VSS.n2794 VSS 0.0603958
R4869 VSS VSS.n2800 0.0603958
R4870 VSS VSS.n94 0.0603958
R4871 VSS.n2827 VSS 0.0603958
R4872 VSS VSS.n447 0.0603958
R4873 VSS VSS.n432 0.0603958
R4874 VSS.n324 VSS 0.0603958
R4875 VSS.n338 VSS 0.0603958
R4876 VSS.n405 VSS.n319 0.0603958
R4877 VSS.n405 VSS.n404 0.0603958
R4878 VSS VSS.n2679 0.0603958
R4879 VSS.n2675 VSS 0.0603958
R4880 VSS.n155 VSS.n153 0.0603958
R4881 VSS.n156 VSS.n155 0.0603958
R4882 VSS.n170 VSS 0.0603958
R4883 VSS.n172 VSS 0.0603958
R4884 VSS VSS.n141 0.0603958
R4885 VSS VSS.n2833 0.0590938
R4886 VSS.n2816 VSS.n2815 0.0590938
R4887 VSS.n2547 VSS.n236 0.0574875
R4888 VSS.n2511 VSS.n257 0.0574875
R4889 VSS.n2389 VSS.n280 0.0574875
R4890 VSS.n2475 VSS.n2391 0.0574875
R4891 VSS.n2659 VSS.n216 0.0574875
R4892 VSS.n565 VSS.n213 0.0574875
R4893 VSS.n2651 VSS.n217 0.0574697
R4894 VSS.n1828 VSS.n1797 0.0574697
R4895 VSS.n2020 VSS.n980 0.0574697
R4896 VSS.n2401 VSS.n2392 0.0574697
R4897 VSS.n1701 VSS.n1700 0.0574697
R4898 VSS.n2445 VSS.n2443 0.0574697
R4899 VSS.n2118 VSS.n908 0.0574697
R4900 VSS.n1405 VSS.n1396 0.0574697
R4901 VSS.n2090 VSS.n932 0.0574697
R4902 VSS.n1140 VSS.n1133 0.0574697
R4903 VSS.n2279 VSS.n840 0.0574697
R4904 VSS.n2226 VSS.n859 0.0574697
R4905 VSS.n258 VSS.n255 0.0574697
R4906 VSS.n237 VSS.n234 0.0574697
R4907 VSS.n1198 VSS.n1197 0.0574697
R4908 VSS.n1213 VSS.n1211 0.0574697
R4909 VSS.n824 VSS.n759 0.0574697
R4910 VSS.n2299 VSS.n557 0.0574697
R4911 VSS.n1322 VSS.n1320 0.0574697
R4912 VSS.n2380 VSS.n465 0.0574697
R4913 VSS.n494 VSS.n481 0.0574697
R4914 VSS.n742 VSS.n567 0.0574697
R4915 VSS.n588 VSS.n587 0.0574697
R4916 VSS.n661 VSS.n603 0.0574697
R4917 VSS.n2348 VSS.n531 0.0574697
R4918 VSS.n2327 VSS.n539 0.0574697
R4919 VSS.n879 VSS.n877 0.0574697
R4920 VSS.n1515 VSS.n1514 0.0574697
R4921 VSS.n1000 VSS.n997 0.0574697
R4922 VSS.n1057 VSS.n1056 0.0574697
R4923 VSS.n1547 VSS.n1545 0.0574697
R4924 VSS.n1019 VSS.n1017 0.0574697
R4925 VSS.n1917 VSS.n1040 0.0574697
R4926 VSS.n902 VSS.n901 0.0574697
R4927 VSS.n2135 VSS.n2134 0.0574697
R4928 VSS.n1154 VSS.n1150 0.0574697
R4929 VSS.n1586 VSS.n1584 0.0574697
R4930 VSS.n1670 VSS.n1086 0.0574697
R4931 VSS.n1762 VSS.n1680 0.0574697
R4932 VSS.n1638 VSS.n1637 0.0574697
R4933 VSS.n1632 VSS.n1631 0.0574697
R4934 VSS.n2074 VSS.n963 0.0574697
R4935 VSS.n1861 VSS.n1082 0.0574697
R4936 VSS.n2624 VSS.n2623 0.0574697
R4937 VSS.n2616 VSS.n2615 0.0574697
R4938 VSS.n2862 VSS 0.0557885
R4939 VSS VSS.n2861 0.0557885
R4940 VSS VSS.n2860 0.0557885
R4941 VSS.n62 VSS 0.0557885
R4942 VSS VSS.n61 0.0557885
R4943 VSS.n11 VSS 0.0557885
R4944 VSS VSS.n53 0.0557885
R4945 VSS VSS.n48 0.0557885
R4946 VSS VSS.n43 0.0557885
R4947 VSS VSS.n38 0.0557885
R4948 VSS VSS.n33 0.0557885
R4949 VSS VSS.n28 0.0557885
R4950 VSS VSS.n23 0.0557885
R4951 VSS.n2871 VSS 0.0557885
R4952 VSS.n2378 VSS.n469 0.0551875
R4953 VSS.n658 VSS.n605 0.0551875
R4954 VSS.n751 VSS.n570 0.0551875
R4955 VSS.n746 VSS.n740 0.0551875
R4956 VSS.n1248 VSS.n1195 0.0551875
R4957 VSS.n2336 VSS.n542 0.0551875
R4958 VSS.n833 VSS.n762 0.0551875
R4959 VSS.n828 VSS.n822 0.0551875
R4960 VSS.n2173 VSS.n874 0.0551875
R4961 VSS.n2288 VSS.n843 0.0551875
R4962 VSS.n2283 VSS.n2277 0.0551875
R4963 VSS.n1431 VSS.n1430 0.0551875
R4964 VSS.n1478 VSS.n1476 0.0551875
R4965 VSS.n2094 VSS.n2093 0.0551875
R4966 VSS.n958 VSS.n957 0.0551875
R4967 VSS.n1668 VSS.n1090 0.0551875
R4968 VSS.n1973 VSS.n994 0.0551875
R4969 VSS.n2083 VSS.n966 0.0551875
R4970 VSS.n2078 VSS.n2072 0.0551875
R4971 VSS.n1064 VSS.n1060 0.0551875
R4972 VSS.n1825 VSS.n1824 0.0551875
R4973 VSS.n2417 VSS.n2416 0.0551875
R4974 VSS.n2542 VSS.n242 0.0551875
R4975 VSS.n2588 VSS.n2584 0.0551875
R4976 VSS.n2614 VSS.n2613 0.0551875
R4977 VSS.n424 VSS.n419 0.0551875
R4978 VSS.n382 VSS.n381 0.0551875
R4979 VSS.n209 VSS.n137 0.0551875
R4980 VSS.n204 VSS.n203 0.0551875
R4981 VSS VSS.n99 0.0527529
R4982 VSS VSS.n1001 0.0525833
R4983 VSS.n1766 VSS 0.0525833
R4984 VSS.n2817 VSS.n99 0.0519696
R4985 VSS.n2873 VSS 0.0518289
R4986 VSS.n491 VSS.n488 0.0499792
R4987 VSS.n686 VSS.n589 0.0499792
R4988 VSS.n1221 VSS.n1220 0.0499792
R4989 VSS.n1388 VSS.n1136 0.0499792
R4990 VSS.n2216 VSS.n2212 0.0499792
R4991 VSS.n1620 VSS.n1399 0.0499792
R4992 VSS.n1551 VSS.n1550 0.0499792
R4993 VSS.n1492 VSS.n909 0.0499792
R4994 VSS.n1634 VSS.n1127 0.0499792
R4995 VSS.n1940 VSS.n1022 0.0499792
R4996 VSS.n1708 VSS.n1698 0.0499792
R4997 VSS.n1921 VSS.n1920 0.0499792
R4998 VSS.n1078 VSS.n1076 0.0499792
R4999 VSS.n2470 VSS.n2395 0.0499792
R5000 VSS.n2571 VSS.n218 0.0499792
R5001 VSS.n75 VSS.n72 0.0499792
R5002 VSS.n309 VSS.n306 0.0499792
R5003 VSS.n2675 VSS.n2674 0.0499792
R5004 VSS.n2826 VSS.n2819 0.0486771
R5005 VSS.n489 VSS 0.047375
R5006 VSS.n1216 VSS 0.047375
R5007 VSS.n1384 VSS 0.047375
R5008 VSS.n1407 VSS 0.047375
R5009 VSS.n1628 VSS 0.047375
R5010 VSS.n1717 VSS 0.047375
R5011 VSS.n2466 VSS 0.047375
R5012 VSS.n307 VSS 0.047375
R5013 VSS.n314 VSS 0.0469438
R5014 VSS VSS.n2703 0.0460729
R5015 VSS.n511 VSS.n466 0.0447708
R5016 VSS.n1243 VSS.n1199 0.0447708
R5017 VSS.n1359 VSS.n1358 0.0447708
R5018 VSS.n1594 VSS.n1419 0.0447708
R5019 VSS.n1662 VSS.n1087 0.0447708
R5020 VSS.n1688 VSS.n1681 0.0447708
R5021 VSS.n2453 VSS.n2408 0.0447708
R5022 VSS.n432 VSS.n431 0.0447708
R5023 VSS.n936 VSS 0.0421667
R5024 VSS.n2056 VSS 0.0421667
R5025 VSS.n1065 VSS 0.0421667
R5026 VSS.n1888 VSS 0.0421667
R5027 VSS.n111 VSS.n109 0.0414836
R5028 VSS.n130 VSS.n127 0.0410405
R5029 VSS.n154 VSS.n131 0.0410405
R5030 VSS.n210 VSS.n134 0.0410405
R5031 VSS.n183 VSS.n133 0.0410405
R5032 VSS.n2656 VSS.n219 0.0410405
R5033 VSS.n2652 VSS.n2650 0.0410405
R5034 VSS.n1800 VSS.n1795 0.0410405
R5035 VSS.n1829 VSS.n1796 0.0410405
R5036 VSS.n2007 VSS.n981 0.0410405
R5037 VSS.n2019 VSS.n979 0.0410405
R5038 VSS.n311 VSS.n297 0.0410405
R5039 VSS.n298 VSS.n284 0.0410405
R5040 VSS.n2472 VSS.n2394 0.0410405
R5041 VSS.n2465 VSS.n2402 0.0410405
R5042 VSS.n1710 VSS.n1704 0.0410405
R5043 VSS.n1716 VSS.n1699 0.0410405
R5044 VSS.n2447 VSS.n2446 0.0410405
R5045 VSS.n2415 VSS.n2414 0.0410405
R5046 VSS.n2123 VSS.n910 0.0410405
R5047 VSS.n2119 VSS.n2117 0.0410405
R5048 VSS.n1622 VSS.n1398 0.0410405
R5049 VSS.n1408 VSS.n1406 0.0410405
R5050 VSS.n2092 VSS.n2091 0.0410405
R5051 VSS.n934 VSS.n933 0.0410405
R5052 VSS.n1390 VSS.n1135 0.0410405
R5053 VSS.n1383 VSS.n1141 0.0410405
R5054 VSS.n2289 VSS.n842 0.0410405
R5055 VSS.n2281 VSS.n2280 0.0410405
R5056 VSS.n2213 VSS.n860 0.0410405
R5057 VSS.n2225 VSS.n858 0.0410405
R5058 VSS.n334 VSS.n333 0.0410405
R5059 VSS.n335 VSS.n318 0.0410405
R5060 VSS.n2508 VSS.n263 0.0410405
R5061 VSS.n260 VSS.n254 0.0410405
R5062 VSS.n352 VSS.n350 0.0410405
R5063 VSS.n379 VSS.n351 0.0410405
R5064 VSS.n2544 VSS.n239 0.0410405
R5065 VSS.n240 VSS.n233 0.0410405
R5066 VSS.n1253 VSS.n1200 0.0410405
R5067 VSS.n1249 VSS.n1196 0.0410405
R5068 VSS.n1223 VSS.n1215 0.0410405
R5069 VSS.n1218 VSS.n1210 0.0410405
R5070 VSS.n834 VSS.n761 0.0410405
R5071 VSS.n826 VSS.n825 0.0410405
R5072 VSS.n2301 VSS.n2300 0.0410405
R5073 VSS.n777 VSS.n772 0.0410405
R5074 VSS.n1324 VSS.n1323 0.0410405
R5075 VSS.n1285 VSS.n1284 0.0410405
R5076 VSS.n2385 VSS.n467 0.0410405
R5077 VSS.n2381 VSS.n2379 0.0410405
R5078 VSS.n486 VSS.n482 0.0410405
R5079 VSS.n493 VSS.n480 0.0410405
R5080 VSS.n752 VSS.n569 0.0410405
R5081 VSS.n744 VSS.n743 0.0410405
R5082 VSS.n697 VSS.n590 0.0410405
R5083 VSS.n693 VSS.n586 0.0410405
R5084 VSS.n648 VSS.n604 0.0410405
R5085 VSS.n660 VSS.n602 0.0410405
R5086 VSS.n2350 VSS.n2349 0.0410405
R5087 VSS.n618 VSS.n617 0.0410405
R5088 VSS.n2338 VSS.n541 0.0410405
R5089 VSS.n2330 VSS.n2328 0.0410405
R5090 VSS.n2175 VSS.n2172 0.0410405
R5091 VSS.n2181 VSS.n876 0.0410405
R5092 VSS.n1511 VSS.n1509 0.0410405
R5093 VSS.n1518 VSS.n1507 0.0410405
R5094 VSS.n1975 VSS.n1003 0.0410405
R5095 VSS.n1981 VSS.n996 0.0410405
R5096 VSS.n1061 VSS.n1055 0.0410405
R5097 VSS.n1062 VSS.n1058 0.0410405
R5098 VSS.n1549 VSS.n1548 0.0410405
R5099 VSS.n1455 VSS.n1454 0.0410405
R5100 VSS.n1941 VSS.n1021 0.0410405
R5101 VSS.n1024 VSS.n1016 0.0410405
R5102 VSS.n1919 VSS.n1918 0.0410405
R5103 VSS.n1042 VSS.n1041 0.0410405
R5104 VSS.n1181 VSS.n897 0.0410405
R5105 VSS.n2136 VSS.n898 0.0410405
R5106 VSS.n1162 VSS.n1149 0.0410405
R5107 VSS.n1163 VSS.n1155 0.0410405
R5108 VSS.n1588 VSS.n1587 0.0410405
R5109 VSS.n1427 VSS.n1426 0.0410405
R5110 VSS.n1675 VSS.n1088 0.0410405
R5111 VSS.n1671 VSS.n1669 0.0410405
R5112 VSS.n1767 VSS.n1682 0.0410405
R5113 VSS.n1763 VSS.n1761 0.0410405
R5114 VSS.n1636 VSS.n1130 0.0410405
R5115 VSS.n1633 VSS.n1629 0.0410405
R5116 VSS.n2084 VSS.n965 0.0410405
R5117 VSS.n2076 VSS.n2075 0.0410405
R5118 VSS.n1863 VSS.n1862 0.0410405
R5119 VSS.n1779 VSS.n1778 0.0410405
R5120 VSS.n2622 VSS.n2585 0.0410405
R5121 VSS.n2618 VSS.n2587 0.0410405
R5122 VSS.n429 VSS.n418 0.0410405
R5123 VSS.n425 VSS.n276 0.0410405
R5124 VSS.n412 VSS.n411 0.0393869
R5125 VSS VSS.n592 0.0382604
R5126 VSS.n497 VSS 0.0369583
R5127 VSS VSS.n695 0.0369583
R5128 VSS.n1229 VSS 0.0369583
R5129 VSS.n773 VSS 0.0369583
R5130 VSS.n1381 VSS 0.0369583
R5131 VSS.n1410 VSS 0.0369583
R5132 VSS VSS.n914 0.0369583
R5133 VSS VSS.n1124 0.0369583
R5134 VSS.n2023 VSS 0.0369583
R5135 VSS VSS.n1696 0.0369583
R5136 VSS.n2463 VSS 0.0369583
R5137 VSS.n456 VSS 0.0369583
R5138 VSS.n2699 VSS.n2698 0.0352656
R5139 VSS.n2178 VSS.n538 0.0351625
R5140 VSS.n2132 VSS.n900 0.0351625
R5141 VSS.n1355 VSS.n1153 0.0351625
R5142 VSS.n1393 VSS.n1131 0.0351625
R5143 VSS.n2296 VSS.n560 0.0351625
R5144 VSS.n2293 VSS.n2292 0.0351625
R5145 VSS.n314 VSS.n313 0.0349852
R5146 VSS.n488 VSS.n487 0.0343542
R5147 VSS.n2352 VSS.n524 0.0343542
R5148 VSS.n1222 VSS.n1221 0.0343542
R5149 VSS.n1326 VSS.n1277 0.0343542
R5150 VSS.n1389 VSS.n1388 0.0343542
R5151 VSS.n1379 VSS 0.0343542
R5152 VSS.n1183 VSS.n1180 0.0343542
R5153 VSS.n1621 VSS.n1620 0.0343542
R5154 VSS.n1616 VSS 0.0343542
R5155 VSS.n1551 VSS.n1450 0.0343542
R5156 VSS.n1129 VSS.n1127 0.0343542
R5157 VSS.n1644 VSS 0.0343542
R5158 VSS.n1022 VSS.n1020 0.0343542
R5159 VSS.n1955 VSS 0.0343542
R5160 VSS.n1999 VSS 0.0343542
R5161 VSS.n1709 VSS.n1708 0.0343542
R5162 VSS.n1921 VSS.n1033 0.0343542
R5163 VSS.n2471 VSS.n2470 0.0343542
R5164 VSS.n2506 VSS.n259 0.0343542
R5165 VSS VSS.n67 0.0343542
R5166 VSS.n306 VSS.n299 0.0343542
R5167 VSS.n331 VSS.n330 0.0343542
R5168 VSS.n2678 VSS 0.0343542
R5169 VSS.n1978 VSS.n999 0.0339875
R5170 VSS.n1944 VSS.n1018 0.0339875
R5171 VSS.n1771 VSS.n1678 0.0339875
R5172 VSS.n1626 VSS.n1083 0.0339875
R5173 VSS.n1777 VSS.n907 0.0339875
R5174 VSS.n2087 VSS.n962 0.0339875
R5175 VSS.n2358 VSS 0.0330521
R5176 VSS.n677 VSS 0.0330521
R5177 VSS.n1330 VSS 0.0330521
R5178 VSS.n2309 VSS 0.0330521
R5179 VSS VSS.n1166 0.0330521
R5180 VSS VSS.n1178 0.0330521
R5181 VSS VSS.n2203 0.0330521
R5182 VSS.n1558 VSS 0.0330521
R5183 VSS VSS.n1933 0.0330521
R5184 VSS VSS.n1998 0.0330521
R5185 VSS.n1926 VSS 0.0330521
R5186 VSS VSS.n1074 0.0330521
R5187 VSS.n1799 VSS 0.0330521
R5188 VSS.n266 VSS 0.0330521
R5189 VSS VSS.n2566 0.0330521
R5190 VSS VSS.n71 0.0330521
R5191 VSS VSS.n2793 0.0330521
R5192 VSS VSS.n269 0.0330521
R5193 VSS.n2680 VSS 0.0330521
R5194 VSS.n1329 VSS 0.03175
R5195 VSS.n801 VSS 0.03175
R5196 VSS VSS.n760 0.03175
R5197 VSS.n1380 VSS 0.03175
R5198 VSS.n2191 VSS 0.03175
R5199 VSS.n2205 VSS 0.03175
R5200 VSS VSS.n1934 0.03175
R5201 VSS.n1974 VSS 0.03175
R5202 VSS VSS.n964 0.03175
R5203 VSS VSS.n1765 0.03175
R5204 VSS VSS.n1684 0.03175
R5205 VSS.n1903 VSS 0.03175
R5206 VSS.n1887 VSS 0.03175
R5207 VSS.n1840 VSS 0.03175
R5208 VSS.n1821 VSS 0.03175
R5209 VSS VSS.n2503 0.03175
R5210 VSS.n2613 VSS 0.03175
R5211 VSS VSS.n95 0.03175
R5212 VSS.n107 VSS.n106 0.0308279
R5213 VSS.n2862 VSS 0.0305481
R5214 VSS.n2861 VSS 0.0305481
R5215 VSS.n2860 VSS 0.0305481
R5216 VSS.n62 VSS 0.0305481
R5217 VSS VSS.n2871 0.0305481
R5218 VSS.n1892 VSS.n1056 0.0292489
R5219 VSS.n1890 VSS.n1057 0.0292489
R5220 VSS.n1977 VSS.n1000 0.0292489
R5221 VSS.n1979 VSS.n997 0.0292489
R5222 VSS.n1514 VSS.n1513 0.0292489
R5223 VSS.n1516 VSS.n1515 0.0292489
R5224 VSS.n2177 VSS.n879 0.0292489
R5225 VSS.n2179 VSS.n877 0.0292489
R5226 VSS.n2340 VSS.n539 0.0292489
R5227 VSS.n2327 VSS.n537 0.0292489
R5228 VSS.n649 VSS.n603 0.0292489
R5229 VSS.n662 VSS.n661 0.0292489
R5230 VSS.n2546 VSS.n237 0.0292489
R5231 VSS.n2548 VSS.n234 0.0292489
R5232 VSS.n1917 VSS.n1916 0.0292489
R5233 VSS.n1914 VSS.n1040 0.0292489
R5234 VSS.n1943 VSS.n1019 0.0292489
R5235 VSS.n1945 VSS.n1017 0.0292489
R5236 VSS.n1547 VSS.n1546 0.0292489
R5237 VSS.n1545 VSS.n1544 0.0292489
R5238 VSS.n1322 VSS.n1321 0.0292489
R5239 VSS.n1320 VSS.n1319 0.0292489
R5240 VSS.n2348 VSS.n2347 0.0292489
R5241 VSS.n532 VSS.n531 0.0292489
R5242 VSS.n2510 VSS.n258 0.0292489
R5243 VSS.n2512 VSS.n255 0.0292489
R5244 VSS.n2135 VSS.n899 0.0292489
R5245 VSS.n901 VSS.n899 0.0292489
R5246 VSS.n1769 VSS.n1680 0.0292489
R5247 VSS.n1762 VSS.n1679 0.0292489
R5248 VSS.n1677 VSS.n1086 0.0292489
R5249 VSS.n1670 VSS.n1085 0.0292489
R5250 VSS.n1586 VSS.n1585 0.0292489
R5251 VSS.n1584 VSS.n1583 0.0292489
R5252 VSS.n1356 VSS.n1150 0.0292489
R5253 VSS.n1353 VSS.n1154 0.0292489
R5254 VSS.n1255 VSS.n1198 0.0292489
R5255 VSS.n1257 VSS.n1197 0.0292489
R5256 VSS.n2387 VSS.n465 0.0292489
R5257 VSS.n2380 VSS.n463 0.0292489
R5258 VSS.n2445 VSS.n2444 0.0292489
R5259 VSS.n2443 VSS.n2442 0.0292489
R5260 VSS.n1712 VSS.n1701 0.0292489
R5261 VSS.n1714 VSS.n1700 0.0292489
R5262 VSS.n1624 VSS.n1396 0.0292489
R5263 VSS.n1405 VSS.n1395 0.0292489
R5264 VSS.n1392 VSS.n1133 0.0292489
R5265 VSS.n1140 VSS.n1132 0.0292489
R5266 VSS.n1225 VSS.n1213 0.0292489
R5267 VSS.n1227 VSS.n1211 0.0292489
R5268 VSS.n484 VSS.n481 0.0292489
R5269 VSS.n495 VSS.n494 0.0292489
R5270 VSS.n2474 VSS.n2392 0.0292489
R5271 VSS.n2401 VSS.n460 0.0292489
R5272 VSS.n1632 VSS.n1627 0.0292489
R5273 VSS.n1637 VSS.n1627 0.0292489
R5274 VSS.n1861 VSS.n1860 0.0292489
R5275 VSS.n1858 VSS.n1082 0.0292489
R5276 VSS.n2008 VSS.n980 0.0292489
R5277 VSS.n2021 VSS.n2020 0.0292489
R5278 VSS.n2125 VSS.n908 0.0292489
R5279 VSS.n2118 VSS.n906 0.0292489
R5280 VSS.n2214 VSS.n859 0.0292489
R5281 VSS.n2227 VSS.n2226 0.0292489
R5282 VSS.n2299 VSS.n2298 0.0292489
R5283 VSS.n559 VSS.n557 0.0292489
R5284 VSS.n699 VSS.n588 0.0292489
R5285 VSS.n701 VSS.n587 0.0292489
R5286 VSS.n2658 VSS.n217 0.0292489
R5287 VSS.n2651 VSS.n215 0.0292489
R5288 VSS.n1802 VSS.n1797 0.0292489
R5289 VSS.n1828 VSS.n1827 0.0292489
R5290 VSS.n2086 VSS.n963 0.0292489
R5291 VSS.n2074 VSS.n961 0.0292489
R5292 VSS.n2090 VSS.n2089 0.0292489
R5293 VSS.n960 VSS.n932 0.0292489
R5294 VSS.n2291 VSS.n840 0.0292489
R5295 VSS.n2279 VSS.n838 0.0292489
R5296 VSS.n836 VSS.n759 0.0292489
R5297 VSS.n824 VSS.n758 0.0292489
R5298 VSS.n754 VSS.n567 0.0292489
R5299 VSS.n742 VSS.n566 0.0292489
R5300 VSS.n2615 VSS.n2586 0.0292489
R5301 VSS.n2623 VSS.n2586 0.0292489
R5302 VSS.n2383 VSS.n469 0.0291458
R5303 VSS.n647 VSS.n605 0.0291458
R5304 VSS.n570 VSS.n568 0.0291458
R5305 VSS.n1251 VSS.n1248 0.0291458
R5306 VSS.n2337 VSS.n2336 0.0291458
R5307 VSS.n762 VSS.n760 0.0291458
R5308 VSS.n1167 VSS.n1165 0.0291458
R5309 VSS.n2174 VSS.n2173 0.0291458
R5310 VSS.n843 VSS.n841 0.0291458
R5311 VSS.n1431 VSS.n1423 0.0291458
R5312 VSS.n1510 VSS.n1476 0.0291458
R5313 VSS.n2094 VSS.n928 0.0291458
R5314 VSS.n1673 VSS.n1090 0.0291458
R5315 VSS.n1974 VSS.n1973 0.0291458
R5316 VSS.n966 VSS.n964 0.0291458
R5317 VSS.n1765 VSS.n1684 0.0291458
R5318 VSS.n1060 VSS.n1059 0.0291458
R5319 VSS.n1798 VSS.n1791 0.0291458
R5320 VSS.n2416 VSS.n2411 0.0291458
R5321 VSS.n2543 VSS.n2542 0.0291458
R5322 VSS.n2626 VSS.n2584 0.0291458
R5323 VSS.n427 VSS.n424 0.0291458
R5324 VSS.n382 VSS.n348 0.0291458
R5325 VSS.n137 VSS.n136 0.0291458
R5326 VSS VSS.n2351 0.0278438
R5327 VSS VSS.n1325 0.0278438
R5328 VSS VSS.n895 0.0278438
R5329 VSS.n2010 VSS 0.0278438
R5330 VSS.n2507 VSS 0.0278438
R5331 VSS.n332 VSS 0.0278438
R5332 VSS VSS.n1183 0.0265417
R5333 VSS VSS.n1721 0.0252396
R5334 VSS.n1738 VSS 0.0252396
R5335 VSS.n1752 VSS 0.0252396
R5336 VSS.n1908 VSS 0.0252396
R5337 VSS.n1876 VSS 0.0252396
R5338 VSS.n1845 VSS 0.0252396
R5339 VSS.n1820 VSS 0.0252396
R5340 VSS VSS.n170 0.0252396
R5341 VSS.n2666 VSS.n2665 0.024993
R5342 VSS.n621 VSS.n616 0.0239375
R5343 VSS.n695 VSS.n692 0.0239375
R5344 VSS.n703 VSS.n585 0.0239375
R5345 VSS.n1289 VSS.n1288 0.0239375
R5346 VSS.n775 VSS.n773 0.0239375
R5347 VSS.n779 VSS.n771 0.0239375
R5348 VSS.n1381 VSS.n1380 0.0239375
R5349 VSS.n896 VSS.n892 0.0239375
R5350 VSS.n2223 VSS.n2222 0.0239375
R5351 VSS.n2229 VSS.n857 0.0239375
R5352 VSS.n1617 VSS.n1410 0.0239375
R5353 VSS.n1458 VSS.n1457 0.0239375
R5354 VSS.n1538 VSS 0.0239375
R5355 VSS.n2121 VSS.n912 0.0239375
R5356 VSS.n2115 VSS.n914 0.0239375
R5357 VSS.n946 VSS 0.0239375
R5358 VSS.n1643 VSS.n1124 0.0239375
R5359 VSS VSS.n1660 0.0239375
R5360 VSS.n1023 VSS.n1015 0.0239375
R5361 VSS.n2017 VSS.n2016 0.0239375
R5362 VSS.n2024 VSS.n2023 0.0239375
R5363 VSS.n1721 VSS.n1696 0.0239375
R5364 VSS.n1760 VSS 0.0239375
R5365 VSS.n1045 VSS.n1044 0.0239375
R5366 VSS.n1780 VSS.n1079 0.0239375
R5367 VSS.n1856 VSS.n1782 0.0239375
R5368 VSS.n2514 VSS.n253 0.0239375
R5369 VSS.n2654 VSS.n221 0.0239375
R5370 VSS.n2648 VSS.n223 0.0239375
R5371 VSS.n456 VSS.n455 0.0239375
R5372 VSS.n322 VSS.n319 0.0239375
R5373 VSS.n153 VSS.n150 0.0239375
R5374 VSS.n157 VSS.n156 0.0239375
R5375 VSS.n356 VSS.n235 0.0234125
R5376 VSS.n408 VSS.n256 0.0234125
R5377 VSS.n2480 VSS.n2479 0.0234125
R5378 VSS.n2476 VSS.n459 0.0234125
R5379 VSS.n2660 VSS.n129 0.0234125
R5380 VSS.n2664 VSS.n2663 0.0234125
R5381 VSS.n2363 VSS 0.0226354
R5382 VSS.n2352 VSS 0.0226354
R5383 VSS VSS.n630 0.0226354
R5384 VSS.n642 VSS 0.0226354
R5385 VSS VSS.n665 0.0226354
R5386 VSS.n678 VSS 0.0226354
R5387 VSS.n692 VSS 0.0226354
R5388 VSS.n740 VSS 0.0226354
R5389 VSS.n732 VSS 0.0226354
R5390 VSS VSS.n1276 0.0226354
R5391 VSS.n1326 VSS 0.0226354
R5392 VSS.n1289 VSS 0.0226354
R5393 VSS VSS.n1295 0.0226354
R5394 VSS.n2312 VSS 0.0226354
R5395 VSS.n2308 VSS 0.0226354
R5396 VSS.n794 VSS 0.0226354
R5397 VSS VSS.n800 0.0226354
R5398 VSS.n815 VSS 0.0226354
R5399 VSS.n1369 VSS 0.0226354
R5400 VSS.n1366 VSS 0.0226354
R5401 VSS.n1167 VSS 0.0226354
R5402 VSS.n1350 VSS 0.0226354
R5403 VSS.n1339 VSS 0.0226354
R5404 VSS.n1185 VSS 0.0226354
R5405 VSS.n1180 VSS 0.0226354
R5406 VSS VSS.n2147 0.0226354
R5407 VSS VSS.n2202 0.0226354
R5408 VSS.n2204 VSS 0.0226354
R5409 VSS.n2243 VSS 0.0226354
R5410 VSS.n2266 VSS 0.0226354
R5411 VSS.n1596 VSS 0.0226354
R5412 VSS VSS.n1438 0.0226354
R5413 VSS VSS.n1441 0.0226354
R5414 VSS.n1541 VSS 0.0226354
R5415 VSS VSS.n1471 0.0226354
R5416 VSS.n1525 VSS 0.0226354
R5417 VSS.n1498 VSS 0.0226354
R5418 VSS.n2098 VSS 0.0226354
R5419 VSS VSS.n938 0.0226354
R5420 VSS VSS.n1649 0.0226354
R5421 VSS.n1650 VSS 0.0226354
R5422 VSS.n1110 VSS 0.0226354
R5423 VSS.n1105 VSS 0.0226354
R5424 VSS.n1935 VSS 0.0226354
R5425 VSS VSS.n1962 0.0226354
R5426 VSS VSS.n1963 0.0226354
R5427 VSS.n1988 VSS 0.0226354
R5428 VSS VSS.n1997 0.0226354
R5429 VSS VSS.n2005 0.0226354
R5430 VSS VSS.n2006 0.0226354
R5431 VSS.n2041 VSS 0.0226354
R5432 VSS.n2049 VSS 0.0226354
R5433 VSS VSS.n2059 0.0226354
R5434 VSS VSS.n1737 0.0226354
R5435 VSS.n1911 VSS 0.0226354
R5436 VSS.n1877 VSS 0.0226354
R5437 VSS VSS.n1783 0.0226354
R5438 VSS VSS.n1791 0.0226354
R5439 VSS.n1810 VSS 0.0226354
R5440 VSS.n2427 VSS 0.0226354
R5441 VSS VSS.n2506 0.0226354
R5442 VSS.n2514 VSS 0.0226354
R5443 VSS.n2533 VSS 0.0226354
R5444 VSS.n2563 VSS 0.0226354
R5445 VSS.n2567 VSS 0.0226354
R5446 VSS.n2636 VSS 0.0226354
R5447 VSS VSS.n2590 0.0226354
R5448 VSS.n2602 VSS 0.0226354
R5449 VSS.n2851 VSS 0.0226354
R5450 VSS VSS.n69 0.0226354
R5451 VSS.n2841 VSS 0.0226354
R5452 VSS VSS.n77 0.0226354
R5453 VSS.n93 VSS 0.0226354
R5454 VSS.n85 VSS 0.0226354
R5455 VSS.n2815 VSS 0.0226354
R5456 VSS.n2810 VSS 0.0226354
R5457 VSS VSS.n2721 0.0226354
R5458 VSS.n2801 VSS 0.0226354
R5459 VSS.n2796 VSS 0.0226354
R5460 VSS.n2822 VSS 0.0226354
R5461 VSS.n448 VSS 0.0226354
R5462 VSS.n433 VSS 0.0226354
R5463 VSS.n2495 VSS 0.0226354
R5464 VSS VSS.n331 0.0226354
R5465 VSS.n363 VSS 0.0226354
R5466 VSS.n167 VSS 0.0226354
R5467 VSS.n197 VSS 0.0226354
R5468 VSS.n189 VSS 0.0226354
R5469 VSS.n2872 VSS 0.0219286
R5470 VSS.n414 VSS.n413 0.0218125
R5471 VSS.n780 VSS 0.0213333
R5472 VSS.n1500 VSS 0.0213333
R5473 VSS.n61 VSS 0.0209327
R5474 VSS VSS.n10 0.0209327
R5475 VSS VSS.n11 0.0209327
R5476 VSS.n54 VSS 0.0209327
R5477 VSS.n53 VSS 0.0209327
R5478 VSS.n49 VSS 0.0209327
R5479 VSS.n48 VSS 0.0209327
R5480 VSS.n44 VSS 0.0209327
R5481 VSS.n43 VSS 0.0209327
R5482 VSS.n39 VSS 0.0209327
R5483 VSS.n38 VSS 0.0209327
R5484 VSS.n34 VSS 0.0209327
R5485 VSS.n33 VSS 0.0209327
R5486 VSS.n29 VSS 0.0209327
R5487 VSS.n28 VSS 0.0209327
R5488 VSS.n24 VSS 0.0209327
R5489 VSS.n23 VSS 0.0209327
R5490 VSS.n19 VSS 0.0209327
R5491 VSS.n483 VSS 0.0200312
R5492 VSS VSS.n1214 0.0200312
R5493 VSS VSS.n1134 0.0200312
R5494 VSS VSS.n1397 0.0200312
R5495 VSS.n1640 VSS 0.0200312
R5496 VSS VSS.n1702 0.0200312
R5497 VSS VSS.n1728 0.0200312
R5498 VSS VSS.n2393 0.0200312
R5499 VSS.n301 VSS 0.0200312
R5500 VSS.n2377 VSS.n471 0.0187292
R5501 VSS.n657 VSS.n601 0.0187292
R5502 VSS.n665 VSS.n664 0.0187292
R5503 VSS.n750 VSS.n571 0.0187292
R5504 VSS.n747 VSS.n723 0.0187292
R5505 VSS.n1260 VSS.n1259 0.0187292
R5506 VSS.n2332 VSS.n2331 0.0187292
R5507 VSS.n2325 VSS.n2324 0.0187292
R5508 VSS.n832 VSS.n763 0.0187292
R5509 VSS.n829 VSS.n806 0.0187292
R5510 VSS.n1351 VSS.n1156 0.0187292
R5511 VSS.n2183 VSS.n2182 0.0187292
R5512 VSS.n875 VSS.n871 0.0187292
R5513 VSS.n2287 VSS.n844 0.0187292
R5514 VSS.n2284 VSS.n2259 0.0187292
R5515 VSS.n1581 VSS.n1428 0.0187292
R5516 VSS.n1520 VSS.n1519 0.0187292
R5517 VSS.n1506 VSS.n1505 0.0187292
R5518 VSS.n935 VSS.n929 0.0187292
R5519 VSS.n937 VSS.n936 0.0187292
R5520 VSS.n1667 VSS.n1092 0.0187292
R5521 VSS.n1983 VSS.n1982 0.0187292
R5522 VSS.n995 VSS.n991 0.0187292
R5523 VSS.n2082 VSS.n967 0.0187292
R5524 VSS.n2079 VSS.n2056 0.0187292
R5525 VSS.n1759 VSS.n1686 0.0187292
R5526 VSS.n1066 VSS.n1065 0.0187292
R5527 VSS.n1888 VSS.n1887 0.0187292
R5528 VSS.n1832 VSS.n1831 0.0187292
R5529 VSS.n1805 VSS.n1804 0.0187292
R5530 VSS.n2440 VSS.n2418 0.0187292
R5531 VSS.n2538 VSS.n232 0.0187292
R5532 VSS.n2551 VSS.n2550 0.0187292
R5533 VSS.n2620 VSS.n2589 0.0187292
R5534 VSS.n2619 VSS.n2590 0.0187292
R5535 VSS.n2483 VSS.n275 0.0187292
R5536 VSS.n357 VSS.n349 0.0187292
R5537 VSS.n375 VSS.n374 0.0187292
R5538 VSS.n208 VSS.n139 0.0187292
R5539 VSS.n205 VSS.n184 0.0187292
R5540 VSS.n281 VSS.n278 0.0183038
R5541 VSS.n410 VSS.n409 0.0182893
R5542 VSS.n1894 VSS 0.0174271
R5543 VSS VSS.n540 0.0148229
R5544 VSS VSS.n238 0.0148229
R5545 VSS.n2703 VSS.n67 0.0148229
R5546 VSS.n490 VSS.n489 0.0135208
R5547 VSS.n615 VSS.n528 0.0135208
R5548 VSS.n696 VSS.n591 0.0135208
R5549 VSS.n1217 VSS.n1216 0.0135208
R5550 VSS.n1287 VSS.n1281 0.0135208
R5551 VSS.n2303 VSS.n2302 0.0135208
R5552 VSS.n1385 VSS.n1384 0.0135208
R5553 VSS.n2139 VSS.n2138 0.0135208
R5554 VSS.n2217 VSS.n861 0.0135208
R5555 VSS.n1407 VSS.n1401 0.0135208
R5556 VSS.n1456 VSS.n1451 0.0135208
R5557 VSS.n2122 VSS.n911 0.0135208
R5558 VSS.n1628 VSS.n1126 0.0135208
R5559 VSS.n1939 VSS.n1026 0.0135208
R5560 VSS.n2011 VSS.n982 0.0135208
R5561 VSS.n1718 VSS.n1717 0.0135208
R5562 VSS.n1043 VSS.n1037 0.0135208
R5563 VSS.n1865 VSS.n1864 0.0135208
R5564 VSS.n2467 VSS.n2466 0.0135208
R5565 VSS.n261 VSS.n250 0.0135208
R5566 VSS.n2655 VSS.n220 0.0135208
R5567 VSS.n308 VSS.n307 0.0135208
R5568 VSS.n338 VSS.n337 0.0135208
R5569 VSS.n148 VSS.n126 0.0135208
R5570 VSS VSS.n2010 0.0109167
R5571 VSS.n332 VSS 0.0109167
R5572 VSS.n696 VSS 0.00961458
R5573 VSS.n2302 VSS 0.00961458
R5574 VSS.n312 VSS.n282 0.00838554
R5575 VSS.n458 VSS.n283 0.00838554
R5576 VSS.n2384 VSS.n468 0.0083125
R5577 VSS.n652 VSS.n651 0.0083125
R5578 VSS.n1252 VSS.n1201 0.0083125
R5579 VSS.n1161 VSS.n1148 0.0083125
R5580 VSS.n2170 VSS.n2169 0.0083125
R5581 VSS.n1590 VSS.n1589 0.0083125
R5582 VSS.n1524 VSS.n1475 0.0083125
R5583 VSS.n1674 VSS.n1089 0.0083125
R5584 VSS.n1969 VSS.n1001 0.0083125
R5585 VSS.n1766 VSS.n1683 0.0083125
R5586 VSS.n1895 VSS.n1894 0.0083125
R5587 VSS.n2449 VSS.n2448 0.0083125
R5588 VSS.n428 VSS.n296 0.0083125
R5589 VSS.n385 VSS.n346 0.0083125
R5590 VSS.n112 VSS.n107 0.00808197
R5591 VSS.n313 VSS.n312 0.00790157
R5592 VSS.n313 VSS.n283 0.00790157
R5593 VSS.n1891 VSS 0.00755
R5594 VSS.n1915 VSS 0.00755
R5595 VSS.n1770 VSS 0.00755
R5596 VSS.n1713 VSS 0.00755
R5597 VSS.n1859 VSS 0.00755
R5598 VSS.n1803 VSS 0.00755
R5599 VSS.n1831 VSS 0.00701042
R5600 VSS.n415 VSS.n316 0.00653911
R5601 VSS.n416 VSS.n277 0.00640857
R5602 VSS.n417 VSS.n279 0.00636298
R5603 VSS.n2481 VSS.n277 0.00636298
R5604 VSS.n378 VSS.n128 0.00631183
R5605 VSS.n317 VSS.n315 0.00624332
R5606 VSS.n407 VSS.n316 0.00624332
R5607 VSS.n355 VSS.n354 0.00604629
R5608 VSS.n378 VSS.n377 0.00604629
R5609 VSS.n2670 VSS.n2669 0.00579577
R5610 VSS VSS.n746 0.00570833
R5611 VSS.n1760 VSS 0.00570833
R5612 VSS.n1799 VSS 0.00570833
R5613 VSS.n2614 VSS 0.00570833
R5614 VSS.n417 VSS.n416 0.00533429
R5615 VSS.n409 VSS.n408 0.0052
R5616 VSS.n2480 VSS.n278 0.0052
R5617 VSS.n411 VSS.n129 0.0052
R5618 VSS.n2664 VSS.n212 0.0052
R5619 VSS.n415 VSS.n315 0.00496369
R5620 VSS.n354 VSS.n128 0.0047957
R5621 VSS VSS.n471 0.00440625
R5622 VSS.n1259 VSS 0.00440625
R5623 VSS VSS.n967 0.00440625
R5624 VSS.n2440 VSS 0.00440625
R5625 VSS.n2711 VSS.n2710 0.00440625
R5626 VSS.n2671 VSS.n2670 0.00364583
R5627 VSS.n2668 VSS.n2667 0.00364583
R5628 VSS.n2669 VSS.n2668 0.00364583
R5629 VSS.n2672 VSS.n2671 0.00364583
R5630 VSS VSS.n935 0.00310417
R5631 VSS.n2833 VSS.n93 0.00180208
R5632 VSS.n95 VSS.n94 0.00180208
R5633 VSS.n112 VSS.n111 0.00152459
R5634 VSS.n998 VSS.n878 0.0010875
R5635 VSS.n2131 VSS.n903 0.0010875
R5636 VSS.n1354 VSS.n1084 0.0010875
R5637 VSS.n1625 VSS.n1394 0.0010875
R5638 VSS.n2127 VSS.n2126 0.0010875
R5639 VSS.n2088 VSS.n839 0.0010875
R5640 x4.clknet_1_0__leaf_clk.n26 x4.clknet_1_0__leaf_clk.n24 333.392
R5641 x4.clknet_1_0__leaf_clk.n26 x4.clknet_1_0__leaf_clk.n25 301.392
R5642 x4.clknet_1_0__leaf_clk.n28 x4.clknet_1_0__leaf_clk.n27 301.392
R5643 x4.clknet_1_0__leaf_clk.n22 x4.clknet_1_0__leaf_clk.n4 301.392
R5644 x4.clknet_1_0__leaf_clk.n31 x4.clknet_1_0__leaf_clk.n23 301.392
R5645 x4.clknet_1_0__leaf_clk.n30 x4.clknet_1_0__leaf_clk.n29 301.392
R5646 x4.clknet_1_0__leaf_clk.n21 x4.clknet_1_0__leaf_clk.n5 297.863
R5647 x4.clknet_1_0__leaf_clk.n2 x4.clknet_1_0__leaf_clk.t38 294.557
R5648 x4.clknet_1_0__leaf_clk.n0 x4.clknet_1_0__leaf_clk.t36 294.557
R5649 x4.clknet_1_0__leaf_clk.n41 x4.clknet_1_0__leaf_clk.t35 294.557
R5650 x4.clknet_1_0__leaf_clk.n38 x4.clknet_1_0__leaf_clk.t33 294.557
R5651 x4.clknet_1_0__leaf_clk.n36 x4.clknet_1_0__leaf_clk.t39 294.557
R5652 x4.clknet_1_0__leaf_clk.n34 x4.clknet_1_0__leaf_clk.n33 287.303
R5653 x4.clknet_1_0__leaf_clk.n8 x4.clknet_1_0__leaf_clk.n6 248.638
R5654 x4.clknet_1_0__leaf_clk.n2 x4.clknet_1_0__leaf_clk.t40 211.01
R5655 x4.clknet_1_0__leaf_clk.n0 x4.clknet_1_0__leaf_clk.t34 211.01
R5656 x4.clknet_1_0__leaf_clk.n41 x4.clknet_1_0__leaf_clk.t37 211.01
R5657 x4.clknet_1_0__leaf_clk.n38 x4.clknet_1_0__leaf_clk.t32 211.01
R5658 x4.clknet_1_0__leaf_clk.n36 x4.clknet_1_0__leaf_clk.t41 211.01
R5659 x4.clknet_1_0__leaf_clk.n8 x4.clknet_1_0__leaf_clk.n7 203.463
R5660 x4.clknet_1_0__leaf_clk.n10 x4.clknet_1_0__leaf_clk.n9 203.463
R5661 x4.clknet_1_0__leaf_clk.n14 x4.clknet_1_0__leaf_clk.n13 203.463
R5662 x4.clknet_1_0__leaf_clk.n16 x4.clknet_1_0__leaf_clk.n15 203.463
R5663 x4.clknet_1_0__leaf_clk.n18 x4.clknet_1_0__leaf_clk.n17 203.463
R5664 x4.clknet_1_0__leaf_clk.n12 x4.clknet_1_0__leaf_clk.n11 202.456
R5665 x4.clknet_1_0__leaf_clk x4.clknet_1_0__leaf_clk.n19 199.607
R5666 x4.clknet_1_0__leaf_clk x4.clknet_1_0__leaf_clk.n2 156.207
R5667 x4.clknet_1_0__leaf_clk.n37 x4.clknet_1_0__leaf_clk.n36 153.097
R5668 x4.clknet_1_0__leaf_clk.n39 x4.clknet_1_0__leaf_clk.n38 152.296
R5669 x4.clknet_1_0__leaf_clk.n1 x4.clknet_1_0__leaf_clk.n0 152
R5670 x4.clknet_1_0__leaf_clk.n42 x4.clknet_1_0__leaf_clk.n41 152
R5671 x4.clknet_1_0__leaf_clk.n10 x4.clknet_1_0__leaf_clk.n8 45.177
R5672 x4.clknet_1_0__leaf_clk.n16 x4.clknet_1_0__leaf_clk.n14 45.177
R5673 x4.clknet_1_0__leaf_clk.n18 x4.clknet_1_0__leaf_clk.n16 45.177
R5674 x4.clknet_1_0__leaf_clk.n12 x4.clknet_1_0__leaf_clk.n10 44.0476
R5675 x4.clknet_1_0__leaf_clk.n14 x4.clknet_1_0__leaf_clk.n12 44.0476
R5676 x4.clknet_1_0__leaf_clk.n6 x4.clknet_1_0__leaf_clk.t23 40.0005
R5677 x4.clknet_1_0__leaf_clk.n6 x4.clknet_1_0__leaf_clk.t29 40.0005
R5678 x4.clknet_1_0__leaf_clk.n7 x4.clknet_1_0__leaf_clk.t21 40.0005
R5679 x4.clknet_1_0__leaf_clk.n7 x4.clknet_1_0__leaf_clk.t27 40.0005
R5680 x4.clknet_1_0__leaf_clk.n9 x4.clknet_1_0__leaf_clk.t19 40.0005
R5681 x4.clknet_1_0__leaf_clk.n9 x4.clknet_1_0__leaf_clk.t24 40.0005
R5682 x4.clknet_1_0__leaf_clk.n11 x4.clknet_1_0__leaf_clk.t31 40.0005
R5683 x4.clknet_1_0__leaf_clk.n11 x4.clknet_1_0__leaf_clk.t18 40.0005
R5684 x4.clknet_1_0__leaf_clk.n13 x4.clknet_1_0__leaf_clk.t30 40.0005
R5685 x4.clknet_1_0__leaf_clk.n13 x4.clknet_1_0__leaf_clk.t22 40.0005
R5686 x4.clknet_1_0__leaf_clk.n15 x4.clknet_1_0__leaf_clk.t28 40.0005
R5687 x4.clknet_1_0__leaf_clk.n15 x4.clknet_1_0__leaf_clk.t17 40.0005
R5688 x4.clknet_1_0__leaf_clk.n17 x4.clknet_1_0__leaf_clk.t26 40.0005
R5689 x4.clknet_1_0__leaf_clk.n17 x4.clknet_1_0__leaf_clk.t16 40.0005
R5690 x4.clknet_1_0__leaf_clk.n19 x4.clknet_1_0__leaf_clk.t20 40.0005
R5691 x4.clknet_1_0__leaf_clk.n19 x4.clknet_1_0__leaf_clk.t25 40.0005
R5692 x4.clknet_1_0__leaf_clk.n28 x4.clknet_1_0__leaf_clk.n26 32.0005
R5693 x4.clknet_1_0__leaf_clk.n32 x4.clknet_1_0__leaf_clk.n22 32.0005
R5694 x4.clknet_1_0__leaf_clk.n32 x4.clknet_1_0__leaf_clk.n31 32.0005
R5695 x4.clknet_1_0__leaf_clk.n30 x4.clknet_1_0__leaf_clk.n28 32.0005
R5696 x4.clknet_1_0__leaf_clk.n31 x4.clknet_1_0__leaf_clk.n30 31.2005
R5697 x4.clknet_1_0__leaf_clk.n35 x4.clknet_1_0__leaf_clk.n34 28.6283
R5698 x4.clknet_1_0__leaf_clk.n3 x4.clknet_1_0__leaf_clk 28.0697
R5699 x4.clknet_1_0__leaf_clk.n24 x4.clknet_1_0__leaf_clk.t7 27.5805
R5700 x4.clknet_1_0__leaf_clk.n24 x4.clknet_1_0__leaf_clk.t13 27.5805
R5701 x4.clknet_1_0__leaf_clk.n25 x4.clknet_1_0__leaf_clk.t5 27.5805
R5702 x4.clknet_1_0__leaf_clk.n25 x4.clknet_1_0__leaf_clk.t11 27.5805
R5703 x4.clknet_1_0__leaf_clk.n27 x4.clknet_1_0__leaf_clk.t3 27.5805
R5704 x4.clknet_1_0__leaf_clk.n27 x4.clknet_1_0__leaf_clk.t8 27.5805
R5705 x4.clknet_1_0__leaf_clk.n4 x4.clknet_1_0__leaf_clk.t10 27.5805
R5706 x4.clknet_1_0__leaf_clk.n4 x4.clknet_1_0__leaf_clk.t0 27.5805
R5707 x4.clknet_1_0__leaf_clk.n5 x4.clknet_1_0__leaf_clk.t4 27.5805
R5708 x4.clknet_1_0__leaf_clk.n5 x4.clknet_1_0__leaf_clk.t9 27.5805
R5709 x4.clknet_1_0__leaf_clk.n33 x4.clknet_1_0__leaf_clk.t12 27.5805
R5710 x4.clknet_1_0__leaf_clk.n33 x4.clknet_1_0__leaf_clk.t1 27.5805
R5711 x4.clknet_1_0__leaf_clk.n23 x4.clknet_1_0__leaf_clk.t14 27.5805
R5712 x4.clknet_1_0__leaf_clk.n23 x4.clknet_1_0__leaf_clk.t6 27.5805
R5713 x4.clknet_1_0__leaf_clk.n29 x4.clknet_1_0__leaf_clk.t15 27.5805
R5714 x4.clknet_1_0__leaf_clk.n29 x4.clknet_1_0__leaf_clk.t2 27.5805
R5715 x4.clknet_1_0__leaf_clk.n43 x4.clknet_1_0__leaf_clk.n42 27.3319
R5716 x4.clknet_1_0__leaf_clk.n40 x4.clknet_1_0__leaf_clk.n39 21.4985
R5717 x4.clknet_1_0__leaf_clk.n3 x4.clknet_1_0__leaf_clk.n1 21.401
R5718 x4.clknet_1_0__leaf_clk.n34 x4.clknet_1_0__leaf_clk.n32 14.0898
R5719 x4.clknet_1_0__leaf_clk.n20 x4.clknet_1_0__leaf_clk.n18 13.177
R5720 x4.clknet_1_0__leaf_clk.n40 x4.clknet_1_0__leaf_clk.n37 11.0654
R5721 x4.clknet_1_0__leaf_clk.n22 x4.clknet_1_0__leaf_clk.n21 10.4484
R5722 x4.clknet_1_0__leaf_clk.n43 x4.clknet_1_0__leaf_clk.n40 7.18319
R5723 x4.clknet_1_0__leaf_clk.n35 x4.clknet_1_0__leaf_clk.n3 5.63649
R5724 x4.clknet_1_0__leaf_clk x4.clknet_1_0__leaf_clk.n20 3.13183
R5725 x4.clknet_1_0__leaf_clk.n37 x4.clknet_1_0__leaf_clk 3.10907
R5726 x4.clknet_1_0__leaf_clk x4.clknet_1_0__leaf_clk.n43 2.66671
R5727 x4.clknet_1_0__leaf_clk x4.clknet_1_0__leaf_clk.n35 2.66671
R5728 x4.clknet_1_0__leaf_clk.n42 x4.clknet_1_0__leaf_clk 2.01193
R5729 x4.clknet_1_0__leaf_clk.n21 x4.clknet_1_0__leaf_clk 1.75844
R5730 x4.clknet_1_0__leaf_clk.n39 x4.clknet_1_0__leaf_clk 1.67435
R5731 x4.clknet_1_0__leaf_clk.n1 x4.clknet_1_0__leaf_clk 1.37896
R5732 x4.clknet_1_0__leaf_clk.n20 x4.clknet_1_0__leaf_clk 0.604792
R5733 ring_out.n0 ring_out.t10 844.321
R5734 ring_out.n0 ring_out.t12 354.322
R5735 ring_out.n3 ring_out.n1 243.68
R5736 ring_out.n8 ring_out.t14 212.081
R5737 ring_out.n7 ring_out.t11 212.081
R5738 ring_out.n5 ring_out.n4 206.249
R5739 ring_out.n3 ring_out.n2 205.28
R5740 ring_out.n9 ring_out.n8 184.806
R5741 ring_out.n8 ring_out.t13 139.78
R5742 ring_out.n7 ring_out.t15 139.78
R5743 ring_out.n8 ring_out.n7 61.346
R5744 ring_out.n1 ring_out.t3 26.5955
R5745 ring_out.n1 ring_out.t2 26.5955
R5746 ring_out.n2 ring_out.t0 26.5955
R5747 ring_out.n2 ring_out.t4 26.5955
R5748 ring_out.n11 ring_out.t6 26.3998
R5749 ring_out ring_out.n3 24.9955
R5750 ring_out.n4 ring_out.t1 24.9236
R5751 ring_out.n4 ring_out.t5 24.9236
R5752 ring_out.n11 ring_out.t7 23.5483
R5753 ring_out.n10 ring_out.n9 21.363
R5754 ring_out ring_out.n5 14.8576
R5755 ring_out.n12 ring_out.t9 12.9758
R5756 ring_out.n6 ring_out 10.9719
R5757 ring_out.n12 ring_out.t8 10.8618
R5758 ring_out.n10 ring_out.n6 9.53262
R5759 ring_out.n6 ring_out 4.57193
R5760 ring_out.n13 ring_out.n11 3.06895
R5761 ring_out.n9 ring_out 2.32777
R5762 ring_out.n13 ring_out.n12 2.14822
R5763 ring_out ring_out.n13 1.12636
R5764 ring_out.n5 ring_out 0.686214
R5765 ring_out ring_out.n10 0.631142
R5766 ring_out ring_out.n0 0.534429
R5767 a_21119_n968.n0 a_21119_n968.t9 1681.78
R5768 a_21119_n968.n2 a_21119_n968.t14 1681.21
R5769 a_21119_n968.n1 a_21119_n968.t6 1681.21
R5770 a_21119_n968.n0 a_21119_n968.t7 1681.21
R5771 a_21119_n968.n13 a_21119_n968.t12 1681.21
R5772 a_21119_n968.n11 a_21119_n968.t13 1681.21
R5773 a_21119_n968.n9 a_21119_n968.t8 1681.21
R5774 a_21119_n968.n7 a_21119_n968.t10 1681.21
R5775 a_21119_n968.n3 a_21119_n968.t2 703.317
R5776 a_21119_n968.n7 a_21119_n968.t17 702.768
R5777 a_21119_n968.n5 a_21119_n968.t16 702.747
R5778 a_21119_n968.n4 a_21119_n968.t3 702.747
R5779 a_21119_n968.n3 a_21119_n968.t15 702.747
R5780 a_21119_n968.n12 a_21119_n968.t5 702.747
R5781 a_21119_n968.n10 a_21119_n968.t4 702.747
R5782 a_21119_n968.n8 a_21119_n968.t11 702.747
R5783 a_21119_n968.n6 a_21119_n968.t1 30.088
R5784 a_21119_n968.t0 a_21119_n968.n15 26.0464
R5785 a_21119_n968.n15 a_21119_n968.n2 20.0759
R5786 a_21119_n968.n6 a_21119_n968.n5 0.875353
R5787 a_21119_n968.n1 a_21119_n968.n0 0.576859
R5788 a_21119_n968.n2 a_21119_n968.n1 0.576859
R5789 a_21119_n968.n4 a_21119_n968.n3 0.570292
R5790 a_21119_n968.n5 a_21119_n968.n4 0.570292
R5791 a_21119_n968.n15 a_21119_n968.n14 0.267403
R5792 a_21119_n968.n14 a_21119_n968.n6 0.10833
R5793 a_21119_n968.n14 a_21119_n968.n13 0.0744583
R5794 a_21119_n968.n8 a_21119_n968.n7 0.0205
R5795 a_21119_n968.n9 a_21119_n968.n8 0.0205
R5796 a_21119_n968.n10 a_21119_n968.n9 0.0205
R5797 a_21119_n968.n11 a_21119_n968.n10 0.0205
R5798 a_21119_n968.n12 a_21119_n968.n11 0.0205
R5799 a_21119_n968.n13 a_21119_n968.n12 0.0205
R5800 x3.x2.GP4.n2 x3.x2.GP4.t4 450.938
R5801 x3.x2.GP4.n2 x3.x2.GP4.t5 445.666
R5802 x3.x2.GP4.n5 x3.x2.GP4.n4 208.965
R5803 x3.x1.x14.Y x3.x2.GP4.n0 96.8352
R5804 x3.x2.GP4.n4 x3.x2.GP4.t1 26.5955
R5805 x3.x2.GP4.n4 x3.x2.GP4.t0 26.5955
R5806 x3.x2.GP4.n0 x3.x2.GP4.t2 24.9236
R5807 x3.x2.GP4.n0 x3.x2.GP4.t3 24.9236
R5808 x3.x1.gpo3 x3.x2.x4.GP 16.5032
R5809 x3.x1.x14.Y x3.x2.GP4.n3 10.2405
R5810 x3.x2.GP4.n3 x3.x1.gpo3 7.76481
R5811 x3.x2.GP4.n1 x3.x1.x14.Y 6.1445
R5812 x3.x2.GP4.n1 x3.x1.x14.Y 4.65505
R5813 x3.x2.x4.GP x3.x2.GP4.n2 2.95993
R5814 x3.x2.GP4.n5 x3.x1.x14.Y 2.0485
R5815 x3.x1.x14.Y x3.x2.GP4.n5 1.55202
R5816 x3.x2.GP4.n3 x3.x2.GP4.n1 1.0245
R5817 x4._11_ x4._11_.n0 623.909
R5818 x4._11_.n24 x4._11_.t5 334.723
R5819 x4._11_.n5 x4._11_.t17 334.723
R5820 x4._11_.n18 x4._11_.t19 261.887
R5821 x4._11_.n14 x4._11_.t20 256.07
R5822 x4._11_.n8 x4._11_.t9 241.536
R5823 x4._11_.n3 x4._11_.t10 241.536
R5824 x4._11_.n1 x4._11_.t7 231.835
R5825 x4._11_.n21 x4._11_.t21 230.363
R5826 x4._11_ x4._11_.n30 216.464
R5827 x4._11_.n24 x4._11_.t12 206.19
R5828 x4._11_.n5 x4._11_.t14 206.19
R5829 x4._11_.n11 x4._11_.t15 183.505
R5830 x4._11_.n8 x4._11_.t6 169.237
R5831 x4._11_.n3 x4._11_.t8 169.237
R5832 x4._11_.n21 x4._11_.t4 158.064
R5833 x4._11_ x4._11_.n3 157.555
R5834 x4._11_ x4._11_.n8 157.166
R5835 x4._11_.n1 x4._11_.t11 157.07
R5836 x4._11_.n18 x4._11_.t13 155.847
R5837 x4._11_.n22 x4._11_.n21 154.048
R5838 x4._11_.n12 x4._11_.n11 153.863
R5839 x4._11_.n19 x4._11_.n18 153.13
R5840 x4._11_.n25 x4._11_.n24 152
R5841 x4._11_.n15 x4._11_.n14 152
R5842 x4._11_.n6 x4._11_.n5 152
R5843 x4._11_.n2 x4._11_.n1 152
R5844 x4._11_.n14 x4._11_.t18 150.03
R5845 x4._11_.n11 x4._11_.t16 114.532
R5846 x4._11_.n27 x4._11_.n26 41.0809
R5847 x4._11_.n30 x4._11_.t2 38.5719
R5848 x4._11_.n30 x4._11_.t3 38.5719
R5849 x4._11_.n0 x4._11_.t0 26.5955
R5850 x4._11_.n0 x4._11_.t1 26.5955
R5851 x4._11_.n17 x4._11_.n16 25.2401
R5852 x4._11_.n20 x4._11_.n19 22.3199
R5853 x4._11_.n10 x4._11_.n9 21.8442
R5854 x4._11_.n10 x4._11_.n7 20.8523
R5855 x4._11_.n28 x4._11_.n27 13.7699
R5856 x4._11_.n28 x4._11_.n2 12.7179
R5857 x4._11_.n4 x4._11_ 12.3175
R5858 x4._11_.n9 x4._11_ 11.4531
R5859 x4._11_.n7 x4._11_.n4 11.4418
R5860 x4._11_.n23 x4._11_.n20 10.8618
R5861 x4._11_.n7 x4._11_.n6 10.3976
R5862 x4._11_.n25 x4._11_ 9.6005
R5863 x4._11_.n29 x4._11_ 9.6005
R5864 x4._11_ x4._11_.n22 9.39918
R5865 x4._11_.n13 x4._11_.n12 9.3005
R5866 x4._11_.n29 x4._11_.n28 9.3005
R5867 x4._11_.n23 x4._11_ 8.80957
R5868 x4._11_.n6 x4._11_ 8.22907
R5869 x4._11_.n15 x4._11_ 7.6805
R5870 x4._11_.n16 x4._11_.n15 4.6085
R5871 x4._11_.n16 x4._11_ 4.58918
R5872 x4._11_.n22 x4._11_ 4.3525
R5873 x4._11_.n4 x4._11_ 4.10616
R5874 x4._11_.n9 x4._11_ 3.81804
R5875 x4._11_.n26 x4._11_ 3.62717
R5876 x4._11_.n19 x4._11_ 3.2005
R5877 x4._11_ x4._11_.n29 3.2005
R5878 x4._11_.n17 x4._11_.n13 2.49494
R5879 x4._11_.n2 x4._11_ 2.3045
R5880 x4._11_.n12 x4._11_ 1.97868
R5881 x4._11_.n13 x4._11_.n10 1.71582
R5882 x4._11_.n27 x4._11_.n23 1.38649
R5883 x4._11_.n26 x4._11_.n25 1.2805
R5884 x4._11_.n20 x4._11_.n17 1.24753
R5885 drv_out.n7 drv_out.t24 184.768
R5886 drv_out.n6 drv_out.t20 184.768
R5887 drv_out.n5 drv_out.t26 184.768
R5888 drv_out.n4 drv_out.t22 184.768
R5889 drv_out.n8 drv_out.n7 171.375
R5890 drv_out.n7 drv_out.t25 146.208
R5891 drv_out.n6 drv_out.t21 146.208
R5892 drv_out.n5 drv_out.t27 146.208
R5893 drv_out.n4 drv_out.t23 146.208
R5894 drv_out.n7 drv_out.n6 40.6397
R5895 drv_out.n6 drv_out.n5 40.6397
R5896 drv_out.n5 drv_out.n4 40.6397
R5897 drv_out.n0 drv_out.t2 26.3998
R5898 drv_out.n21 drv_out.n20 26.0838
R5899 drv_out.n21 drv_out.n17 26.0838
R5900 drv_out.n21 drv_out.n19 26.0838
R5901 drv_out.n21 drv_out.n18 26.0838
R5902 drv_out.n16 drv_out.n12 24.902
R5903 drv_out.n16 drv_out.n14 24.902
R5904 drv_out.n16 drv_out.n13 24.902
R5905 drv_out.n16 drv_out.n15 24.902
R5906 drv_out.n0 drv_out.t3 23.5483
R5907 drv_out.n1 drv_out.t1 12.9758
R5908 drv_out drv_out.n8 12.3171
R5909 drv_out.n1 drv_out.t0 10.8618
R5910 drv_out.n20 drv_out.t16 6.6005
R5911 drv_out.n20 drv_out.t13 6.6005
R5912 drv_out.n17 drv_out.t17 6.6005
R5913 drv_out.n17 drv_out.t18 6.6005
R5914 drv_out.n19 drv_out.t15 6.6005
R5915 drv_out.n19 drv_out.t14 6.6005
R5916 drv_out.n18 drv_out.t12 6.6005
R5917 drv_out.n18 drv_out.t19 6.6005
R5918 drv_out.n11 drv_out 5.69273
R5919 drv_out.n12 drv_out.t4 3.61217
R5920 drv_out.n12 drv_out.t6 3.61217
R5921 drv_out.n14 drv_out.t10 3.61217
R5922 drv_out.n14 drv_out.t9 3.61217
R5923 drv_out.n13 drv_out.t8 3.61217
R5924 drv_out.n13 drv_out.t7 3.61217
R5925 drv_out.n15 drv_out.t11 3.61217
R5926 drv_out.n15 drv_out.t5 3.61217
R5927 drv_out.n2 drv_out.n0 3.06895
R5928 drv_out.n11 drv_out 2.87193
R5929 drv_out.n8 drv_out 2.23542
R5930 drv_out.n2 drv_out.n1 2.14822
R5931 drv_out.n10 drv_out 1.7806
R5932 drv_out drv_out.n10 1.54574
R5933 drv_out.n9 drv_out 1.25273
R5934 drv_out.n3 drv_out.n2 1.12636
R5935 drv_out drv_out.n22 0.461707
R5936 drv_out.n9 drv_out 0.316378
R5937 drv_out drv_out.n11 0.188041
R5938 drv_out drv_out.n3 0.138152
R5939 drv_out.n22 drv_out.n16 0.0921193
R5940 drv_out.n22 drv_out.n21 0.069392
R5941 drv_out.n3 drv_out 0.0655
R5942 drv_out.n10 drv_out.n9 0.0596216
R5943 mux_out.n6 mux_out.t1 23.6581
R5944 mux_out.n12 mux_out.t13 23.6581
R5945 mux_out.n19 mux_out.t5 23.6581
R5946 mux_out.n1 mux_out.t14 23.6581
R5947 mux_out.n5 mux_out.t0 23.3739
R5948 mux_out.n11 mux_out.t12 23.3739
R5949 mux_out.n18 mux_out.t4 23.3739
R5950 mux_out.n0 mux_out.t15 23.3739
R5951 mux_out.n6 mux_out.t6 10.7528
R5952 mux_out.n12 mux_out.t10 10.7528
R5953 mux_out.n19 mux_out.t9 10.7528
R5954 mux_out.n1 mux_out.t2 10.7528
R5955 mux_out.n8 mux_out.t7 10.6417
R5956 mux_out.n14 mux_out.t11 10.6417
R5957 mux_out.n21 mux_out.t8 10.6417
R5958 mux_out.n3 mux_out.t3 10.6417
R5959 mux_out.n7 mux_out.n6 1.30064
R5960 mux_out.n13 mux_out.n12 1.30064
R5961 mux_out.n20 mux_out.n19 1.30064
R5962 mux_out.n2 mux_out.n1 1.30064
R5963 mux_out mux_out.n4 0.983856
R5964 mux_out.n23 mux_out.n22 0.946356
R5965 mux_out.n16 mux_out.n15 0.927606
R5966 mux_out.n10 mux_out.n9 0.925106
R5967 mux_out.n17 mux_out 0.748625
R5968 mux_out.n7 mux_out.n5 0.726502
R5969 mux_out.n13 mux_out.n11 0.726502
R5970 mux_out.n20 mux_out.n18 0.726502
R5971 mux_out.n2 mux_out.n0 0.726502
R5972 mux_out.n24 mux_out.n17 0.54425
R5973 mux_out.n8 mux_out.n7 0.512491
R5974 mux_out.n14 mux_out.n13 0.512491
R5975 mux_out.n21 mux_out.n20 0.512491
R5976 mux_out.n3 mux_out.n2 0.512491
R5977 mux_out.n9 mux_out.n8 0.359663
R5978 mux_out.n15 mux_out.n14 0.359663
R5979 mux_out.n22 mux_out.n21 0.359663
R5980 mux_out.n4 mux_out.n3 0.359663
R5981 mux_out.n9 mux_out.n5 0.216071
R5982 mux_out.n15 mux_out.n11 0.216071
R5983 mux_out.n22 mux_out.n18 0.216071
R5984 mux_out.n4 mux_out.n0 0.216071
R5985 mux_out.n17 mux_out 0.20175
R5986 mux_out.n24 mux_out 0.17925
R5987 mux_out.n24 mux_out 0.063
R5988 mux_out.n10 mux_out 0.05925
R5989 mux_out.n16 mux_out 0.05675
R5990 mux_out mux_out.n16 0.0561931
R5991 mux_out mux_out.n10 0.0561872
R5992 mux_out.n23 mux_out 0.038
R5993 mux_out mux_out.n23 0.0376287
R5994 mux_out mux_out.n24 0.004875
R5995 x4.clknet_1_1__leaf_clk.n29 x4.clknet_1_1__leaf_clk.n27 333.392
R5996 x4.clknet_1_1__leaf_clk.n29 x4.clknet_1_1__leaf_clk.n28 301.392
R5997 x4.clknet_1_1__leaf_clk.n31 x4.clknet_1_1__leaf_clk.n30 301.392
R5998 x4.clknet_1_1__leaf_clk.n33 x4.clknet_1_1__leaf_clk.n32 301.392
R5999 x4.clknet_1_1__leaf_clk.n35 x4.clknet_1_1__leaf_clk.n34 301.392
R6000 x4.clknet_1_1__leaf_clk.n37 x4.clknet_1_1__leaf_clk.n36 301.392
R6001 x4.clknet_1_1__leaf_clk.n39 x4.clknet_1_1__leaf_clk.n38 301.392
R6002 x4.clknet_1_1__leaf_clk.n40 x4.clknet_1_1__leaf_clk.n26 297.863
R6003 x4.clknet_1_1__leaf_clk.n18 x4.clknet_1_1__leaf_clk.t38 294.557
R6004 x4.clknet_1_1__leaf_clk.n15 x4.clknet_1_1__leaf_clk.t40 294.557
R6005 x4.clknet_1_1__leaf_clk.n13 x4.clknet_1_1__leaf_clk.t34 294.557
R6006 x4.clknet_1_1__leaf_clk.n11 x4.clknet_1_1__leaf_clk.t36 294.557
R6007 x4.clknet_1_1__leaf_clk.n10 x4.clknet_1_1__leaf_clk.t32 294.557
R6008 x4.clknet_1_1__leaf_clk.n2 x4.clknet_1_1__leaf_clk.n0 248.638
R6009 x4.clknet_1_1__leaf_clk.n18 x4.clknet_1_1__leaf_clk.t41 211.01
R6010 x4.clknet_1_1__leaf_clk.n15 x4.clknet_1_1__leaf_clk.t39 211.01
R6011 x4.clknet_1_1__leaf_clk.n13 x4.clknet_1_1__leaf_clk.t37 211.01
R6012 x4.clknet_1_1__leaf_clk.n11 x4.clknet_1_1__leaf_clk.t35 211.01
R6013 x4.clknet_1_1__leaf_clk.n10 x4.clknet_1_1__leaf_clk.t33 211.01
R6014 x4.clknet_1_1__leaf_clk.n2 x4.clknet_1_1__leaf_clk.n1 203.463
R6015 x4.clknet_1_1__leaf_clk.n4 x4.clknet_1_1__leaf_clk.n3 203.463
R6016 x4.clknet_1_1__leaf_clk.n8 x4.clknet_1_1__leaf_clk.n7 203.463
R6017 x4.clknet_1_1__leaf_clk.n25 x4.clknet_1_1__leaf_clk.n24 203.463
R6018 x4.clknet_1_1__leaf_clk.n6 x4.clknet_1_1__leaf_clk.n5 202.456
R6019 x4.clknet_1_1__leaf_clk x4.clknet_1_1__leaf_clk.n42 199.607
R6020 x4.clknet_1_1__leaf_clk.n22 x4.clknet_1_1__leaf_clk.n9 188.201
R6021 x4.clknet_1_1__leaf_clk x4.clknet_1_1__leaf_clk.n13 156.207
R6022 x4.clknet_1_1__leaf_clk x4.clknet_1_1__leaf_clk.n10 156.207
R6023 x4.clknet_1_1__leaf_clk.n19 x4.clknet_1_1__leaf_clk.n18 153.097
R6024 x4.clknet_1_1__leaf_clk.n16 x4.clknet_1_1__leaf_clk.n15 152.296
R6025 x4.clknet_1_1__leaf_clk.n12 x4.clknet_1_1__leaf_clk.n11 152.296
R6026 x4.clknet_1_1__leaf_clk.n4 x4.clknet_1_1__leaf_clk.n2 45.177
R6027 x4.clknet_1_1__leaf_clk.n23 x4.clknet_1_1__leaf_clk.n8 45.177
R6028 x4.clknet_1_1__leaf_clk.n25 x4.clknet_1_1__leaf_clk.n23 45.177
R6029 x4.clknet_1_1__leaf_clk.n6 x4.clknet_1_1__leaf_clk.n4 44.0476
R6030 x4.clknet_1_1__leaf_clk.n8 x4.clknet_1_1__leaf_clk.n6 44.0476
R6031 x4.clknet_1_1__leaf_clk.n0 x4.clknet_1_1__leaf_clk.t18 40.0005
R6032 x4.clknet_1_1__leaf_clk.n0 x4.clknet_1_1__leaf_clk.t20 40.0005
R6033 x4.clknet_1_1__leaf_clk.n1 x4.clknet_1_1__leaf_clk.t21 40.0005
R6034 x4.clknet_1_1__leaf_clk.n1 x4.clknet_1_1__leaf_clk.t28 40.0005
R6035 x4.clknet_1_1__leaf_clk.n3 x4.clknet_1_1__leaf_clk.t23 40.0005
R6036 x4.clknet_1_1__leaf_clk.n3 x4.clknet_1_1__leaf_clk.t30 40.0005
R6037 x4.clknet_1_1__leaf_clk.n5 x4.clknet_1_1__leaf_clk.t26 40.0005
R6038 x4.clknet_1_1__leaf_clk.n5 x4.clknet_1_1__leaf_clk.t16 40.0005
R6039 x4.clknet_1_1__leaf_clk.n7 x4.clknet_1_1__leaf_clk.t27 40.0005
R6040 x4.clknet_1_1__leaf_clk.n7 x4.clknet_1_1__leaf_clk.t17 40.0005
R6041 x4.clknet_1_1__leaf_clk.n9 x4.clknet_1_1__leaf_clk.t29 40.0005
R6042 x4.clknet_1_1__leaf_clk.n9 x4.clknet_1_1__leaf_clk.t19 40.0005
R6043 x4.clknet_1_1__leaf_clk.n24 x4.clknet_1_1__leaf_clk.t31 40.0005
R6044 x4.clknet_1_1__leaf_clk.n24 x4.clknet_1_1__leaf_clk.t22 40.0005
R6045 x4.clknet_1_1__leaf_clk.n42 x4.clknet_1_1__leaf_clk.t24 40.0005
R6046 x4.clknet_1_1__leaf_clk.n42 x4.clknet_1_1__leaf_clk.t25 40.0005
R6047 x4.clknet_1_1__leaf_clk.n21 x4.clknet_1_1__leaf_clk 34.5053
R6048 x4.clknet_1_1__leaf_clk.n14 x4.clknet_1_1__leaf_clk 33.8485
R6049 x4.clknet_1_1__leaf_clk.n31 x4.clknet_1_1__leaf_clk.n29 32.0005
R6050 x4.clknet_1_1__leaf_clk.n33 x4.clknet_1_1__leaf_clk.n31 32.0005
R6051 x4.clknet_1_1__leaf_clk.n37 x4.clknet_1_1__leaf_clk.n35 32.0005
R6052 x4.clknet_1_1__leaf_clk.n39 x4.clknet_1_1__leaf_clk.n37 32.0005
R6053 x4.clknet_1_1__leaf_clk.n35 x4.clknet_1_1__leaf_clk.n33 31.2005
R6054 x4.clknet_1_1__leaf_clk.n27 x4.clknet_1_1__leaf_clk.t2 27.5805
R6055 x4.clknet_1_1__leaf_clk.n27 x4.clknet_1_1__leaf_clk.t4 27.5805
R6056 x4.clknet_1_1__leaf_clk.n28 x4.clknet_1_1__leaf_clk.t5 27.5805
R6057 x4.clknet_1_1__leaf_clk.n28 x4.clknet_1_1__leaf_clk.t12 27.5805
R6058 x4.clknet_1_1__leaf_clk.n30 x4.clknet_1_1__leaf_clk.t7 27.5805
R6059 x4.clknet_1_1__leaf_clk.n30 x4.clknet_1_1__leaf_clk.t14 27.5805
R6060 x4.clknet_1_1__leaf_clk.n32 x4.clknet_1_1__leaf_clk.t10 27.5805
R6061 x4.clknet_1_1__leaf_clk.n32 x4.clknet_1_1__leaf_clk.t0 27.5805
R6062 x4.clknet_1_1__leaf_clk.n34 x4.clknet_1_1__leaf_clk.t11 27.5805
R6063 x4.clknet_1_1__leaf_clk.n34 x4.clknet_1_1__leaf_clk.t1 27.5805
R6064 x4.clknet_1_1__leaf_clk.n36 x4.clknet_1_1__leaf_clk.t13 27.5805
R6065 x4.clknet_1_1__leaf_clk.n36 x4.clknet_1_1__leaf_clk.t3 27.5805
R6066 x4.clknet_1_1__leaf_clk.n26 x4.clknet_1_1__leaf_clk.t8 27.5805
R6067 x4.clknet_1_1__leaf_clk.n26 x4.clknet_1_1__leaf_clk.t9 27.5805
R6068 x4.clknet_1_1__leaf_clk.n38 x4.clknet_1_1__leaf_clk.t15 27.5805
R6069 x4.clknet_1_1__leaf_clk.n38 x4.clknet_1_1__leaf_clk.t6 27.5805
R6070 x4.clknet_1_1__leaf_clk.n23 x4.clknet_1_1__leaf_clk.n22 15.262
R6071 x4.clknet_1_1__leaf_clk.n20 x4.clknet_1_1__leaf_clk.n19 13.8005
R6072 x4.clknet_1_1__leaf_clk.n41 x4.clknet_1_1__leaf_clk.n25 13.177
R6073 x4.clknet_1_1__leaf_clk.n14 x4.clknet_1_1__leaf_clk.n12 11.6482
R6074 x4.clknet_1_1__leaf_clk.n22 x4.clknet_1_1__leaf_clk.n21 10.8268
R6075 x4.clknet_1_1__leaf_clk.n40 x4.clknet_1_1__leaf_clk.n39 10.4484
R6076 x4.clknet_1_1__leaf_clk.n17 x4.clknet_1_1__leaf_clk.n16 9.3005
R6077 x4.clknet_1_1__leaf_clk.n20 x4.clknet_1_1__leaf_clk.n17 8.37704
R6078 x4.clknet_1_1__leaf_clk.n21 x4.clknet_1_1__leaf_clk 5.19349
R6079 x4.clknet_1_1__leaf_clk.n17 x4.clknet_1_1__leaf_clk.n14 3.99105
R6080 x4.clknet_1_1__leaf_clk.n41 x4.clknet_1_1__leaf_clk 3.13183
R6081 x4.clknet_1_1__leaf_clk.n19 x4.clknet_1_1__leaf_clk 3.10907
R6082 x4.clknet_1_1__leaf_clk x4.clknet_1_1__leaf_clk.n40 1.75844
R6083 x4.clknet_1_1__leaf_clk.n16 x4.clknet_1_1__leaf_clk 1.67435
R6084 x4.clknet_1_1__leaf_clk.n12 x4.clknet_1_1__leaf_clk 1.67435
R6085 x4.clknet_1_1__leaf_clk x4.clknet_1_1__leaf_clk.n20 0.693495
R6086 x4.clknet_1_1__leaf_clk x4.clknet_1_1__leaf_clk.n41 0.604792
R6087 x4.clknet_0_clk.n28 x4.clknet_0_clk.n26 333.392
R6088 x4.clknet_0_clk.n28 x4.clknet_0_clk.n27 301.392
R6089 x4.clknet_0_clk.n30 x4.clknet_0_clk.n29 301.392
R6090 x4.clknet_0_clk.n32 x4.clknet_0_clk.n31 301.392
R6091 x4.clknet_0_clk.n34 x4.clknet_0_clk.n33 301.392
R6092 x4.clknet_0_clk.n36 x4.clknet_0_clk.n35 301.392
R6093 x4.clknet_0_clk.n38 x4.clknet_0_clk.n37 301.392
R6094 x4.clknet_0_clk.n39 x4.clknet_0_clk.n25 297.863
R6095 x4.clknet_0_clk.n2 x4.clknet_0_clk.n0 248.638
R6096 x4.clknet_0_clk.n2 x4.clknet_0_clk.n1 203.463
R6097 x4.clknet_0_clk.n4 x4.clknet_0_clk.n3 203.463
R6098 x4.clknet_0_clk.n8 x4.clknet_0_clk.n7 203.463
R6099 x4.clknet_0_clk.n24 x4.clknet_0_clk.n23 203.463
R6100 x4.clknet_0_clk.n6 x4.clknet_0_clk.n5 202.456
R6101 x4.clknet_0_clk x4.clknet_0_clk.n41 199.607
R6102 x4.clknet_0_clk.n21 x4.clknet_0_clk.n9 188.201
R6103 x4.clknet_0_clk.n18 x4.clknet_0_clk.t32 184.768
R6104 x4.clknet_0_clk.n17 x4.clknet_0_clk.t40 184.768
R6105 x4.clknet_0_clk.n16 x4.clknet_0_clk.t34 184.768
R6106 x4.clknet_0_clk.n15 x4.clknet_0_clk.t43 184.768
R6107 x4.clknet_0_clk.n10 x4.clknet_0_clk.t36 184.768
R6108 x4.clknet_0_clk.n11 x4.clknet_0_clk.t42 184.768
R6109 x4.clknet_0_clk.n12 x4.clknet_0_clk.t38 184.768
R6110 x4.clknet_0_clk.n13 x4.clknet_0_clk.t45 184.768
R6111 x4.clknet_0_clk x4.clknet_0_clk.n18 173.609
R6112 x4.clknet_0_clk.n14 x4.clknet_0_clk.n13 171.375
R6113 x4.clknet_0_clk.n18 x4.clknet_0_clk.t33 146.208
R6114 x4.clknet_0_clk.n17 x4.clknet_0_clk.t41 146.208
R6115 x4.clknet_0_clk.n16 x4.clknet_0_clk.t35 146.208
R6116 x4.clknet_0_clk.n15 x4.clknet_0_clk.t46 146.208
R6117 x4.clknet_0_clk.n10 x4.clknet_0_clk.t37 146.208
R6118 x4.clknet_0_clk.n11 x4.clknet_0_clk.t44 146.208
R6119 x4.clknet_0_clk.n12 x4.clknet_0_clk.t39 146.208
R6120 x4.clknet_0_clk.n13 x4.clknet_0_clk.t47 146.208
R6121 x4.clknet_0_clk.n4 x4.clknet_0_clk.n2 45.177
R6122 x4.clknet_0_clk.n22 x4.clknet_0_clk.n8 45.177
R6123 x4.clknet_0_clk.n24 x4.clknet_0_clk.n22 45.177
R6124 x4.clknet_0_clk.n6 x4.clknet_0_clk.n4 44.0476
R6125 x4.clknet_0_clk.n8 x4.clknet_0_clk.n6 44.0476
R6126 x4.clknet_0_clk.n18 x4.clknet_0_clk.n17 40.6397
R6127 x4.clknet_0_clk.n17 x4.clknet_0_clk.n16 40.6397
R6128 x4.clknet_0_clk.n16 x4.clknet_0_clk.n15 40.6397
R6129 x4.clknet_0_clk.n11 x4.clknet_0_clk.n10 40.6397
R6130 x4.clknet_0_clk.n12 x4.clknet_0_clk.n11 40.6397
R6131 x4.clknet_0_clk.n13 x4.clknet_0_clk.n12 40.6397
R6132 x4.clknet_0_clk.n0 x4.clknet_0_clk.t31 40.0005
R6133 x4.clknet_0_clk.n0 x4.clknet_0_clk.t18 40.0005
R6134 x4.clknet_0_clk.n1 x4.clknet_0_clk.t23 40.0005
R6135 x4.clknet_0_clk.n1 x4.clknet_0_clk.t17 40.0005
R6136 x4.clknet_0_clk.n3 x4.clknet_0_clk.t22 40.0005
R6137 x4.clknet_0_clk.n3 x4.clknet_0_clk.t28 40.0005
R6138 x4.clknet_0_clk.n5 x4.clknet_0_clk.t20 40.0005
R6139 x4.clknet_0_clk.n5 x4.clknet_0_clk.t26 40.0005
R6140 x4.clknet_0_clk.n7 x4.clknet_0_clk.t19 40.0005
R6141 x4.clknet_0_clk.n7 x4.clknet_0_clk.t25 40.0005
R6142 x4.clknet_0_clk.n9 x4.clknet_0_clk.t16 40.0005
R6143 x4.clknet_0_clk.n9 x4.clknet_0_clk.t24 40.0005
R6144 x4.clknet_0_clk.n23 x4.clknet_0_clk.t30 40.0005
R6145 x4.clknet_0_clk.n23 x4.clknet_0_clk.t21 40.0005
R6146 x4.clknet_0_clk.n41 x4.clknet_0_clk.t27 40.0005
R6147 x4.clknet_0_clk.n41 x4.clknet_0_clk.t29 40.0005
R6148 x4.clknet_0_clk.n30 x4.clknet_0_clk.n28 32.0005
R6149 x4.clknet_0_clk.n32 x4.clknet_0_clk.n30 32.0005
R6150 x4.clknet_0_clk.n36 x4.clknet_0_clk.n34 32.0005
R6151 x4.clknet_0_clk.n38 x4.clknet_0_clk.n36 32.0005
R6152 x4.clknet_0_clk.n34 x4.clknet_0_clk.n32 31.2005
R6153 x4.clknet_0_clk.n25 x4.clknet_0_clk.t12 27.5805
R6154 x4.clknet_0_clk.n25 x4.clknet_0_clk.t14 27.5805
R6155 x4.clknet_0_clk.n26 x4.clknet_0_clk.t0 27.5805
R6156 x4.clknet_0_clk.n26 x4.clknet_0_clk.t3 27.5805
R6157 x4.clknet_0_clk.n27 x4.clknet_0_clk.t8 27.5805
R6158 x4.clknet_0_clk.n27 x4.clknet_0_clk.t2 27.5805
R6159 x4.clknet_0_clk.n29 x4.clknet_0_clk.t7 27.5805
R6160 x4.clknet_0_clk.n29 x4.clknet_0_clk.t13 27.5805
R6161 x4.clknet_0_clk.n31 x4.clknet_0_clk.t5 27.5805
R6162 x4.clknet_0_clk.n31 x4.clknet_0_clk.t11 27.5805
R6163 x4.clknet_0_clk.n33 x4.clknet_0_clk.t4 27.5805
R6164 x4.clknet_0_clk.n33 x4.clknet_0_clk.t10 27.5805
R6165 x4.clknet_0_clk.n35 x4.clknet_0_clk.t1 27.5805
R6166 x4.clknet_0_clk.n35 x4.clknet_0_clk.t9 27.5805
R6167 x4.clknet_0_clk.n37 x4.clknet_0_clk.t15 27.5805
R6168 x4.clknet_0_clk.n37 x4.clknet_0_clk.t6 27.5805
R6169 x4.clknet_0_clk x4.clknet_0_clk.n14 25.9814
R6170 x4.clknet_0_clk.n22 x4.clknet_0_clk.n21 15.262
R6171 x4.clknet_0_clk.n20 x4.clknet_0_clk.n19 14.7771
R6172 x4.clknet_0_clk.n40 x4.clknet_0_clk.n24 13.177
R6173 x4.clknet_0_clk.n39 x4.clknet_0_clk.n38 10.4484
R6174 x4.clknet_0_clk.n19 x4.clknet_0_clk 10.3624
R6175 x4.clknet_0_clk.n21 x4.clknet_0_clk.n20 9.3005
R6176 x4.clknet_0_clk.n19 x4.clknet_0_clk 3.45447
R6177 x4.clknet_0_clk.n40 x4.clknet_0_clk 3.13183
R6178 x4.clknet_0_clk.n14 x4.clknet_0_clk 2.23542
R6179 x4.clknet_0_clk x4.clknet_0_clk.n39 1.75844
R6180 x4.clknet_0_clk.n20 x4.clknet_0_clk 1.5927
R6181 x4.clknet_0_clk x4.clknet_0_clk.n40 0.604792
R6182 x4.net2.n14 x4.net2.t0 315.034
R6183 x4.net2.t1 x4.net2.n14 265.769
R6184 x4.net2 x4.net2.t1 262.318
R6185 x4.net2.n4 x4.net2.t5 260.322
R6186 x4.net2.n9 x4.net2.t11 241.536
R6187 x4.net2.n0 x4.net2.t10 212.081
R6188 x4.net2.n1 x4.net2.t9 212.081
R6189 x4.net2.n6 x4.net2.t2 183.505
R6190 x4.net2.n4 x4.net2.t7 175.169
R6191 x4.net2.n9 x4.net2.t8 169.237
R6192 x4.net2.n10 x4.net2.n9 159.952
R6193 x4.net2.n7 x4.net2.n6 153.863
R6194 x4.net2.n3 x4.net2.n2 152.698
R6195 x4.net2.n5 x4.net2.n4 152
R6196 x4.net2.n0 x4.net2.t6 139.78
R6197 x4.net2.n1 x4.net2.t4 139.78
R6198 x4.net2.n6 x4.net2.t3 114.532
R6199 x4.net2.n2 x4.net2.n0 37.246
R6200 x4.net2.n8 x4.net2.n5 34.4715
R6201 x4.net2.n2 x4.net2.n1 24.1005
R6202 x4.net2.n12 x4.net2.n3 18.9449
R6203 x4.net2.n13 x4.net2.n12 14.916
R6204 x4.net2.n11 x4.net2.n10 13.8005
R6205 x4.net2 x4.net2.n7 10.8927
R6206 x4.net2.n14 x4.net2.n13 8.72777
R6207 x4.net2.n8 x4.net2 6.07742
R6208 x4.net2.n10 x4.net2 3.33963
R6209 x4.net2.n10 x4.net2 3.29747
R6210 x4.net2 x4.net2.n13 3.29747
R6211 x4.net2.n11 x4.net2.n8 3.19006
R6212 x4.net2.n3 x4.net2 1.97868
R6213 x4.net2.n7 x4.net2 1.97868
R6214 x4.net2.n5 x4.net2 1.55726
R6215 x4.net2.n12 x4.net2.n11 1.38649
R6216 select1.n10 select1.t6 327.99
R6217 select1.n3 select1.t8 293.969
R6218 select1.n6 select1.t3 256.07
R6219 select1.n0 select1.t4 212.081
R6220 select1.n1 select1.t2 212.081
R6221 select1.n10 select1.t5 199.457
R6222 select1.n2 select1.n1 182.929
R6223 select1 select1.n3 154.065
R6224 select1.n11 select1.n10 152
R6225 select1.n7 select1.n6 152
R6226 select1.n6 select1.t7 150.03
R6227 select1.n0 select1.t1 139.78
R6228 select1.n1 select1.t9 139.78
R6229 select1.n3 select1.t0 138.338
R6230 select1.n1 select1.n0 61.346
R6231 select1.n5 select1 17.455
R6232 select1.n14 select1.n13 14.6836
R6233 select1.n13 select1.n12 14.6704
R6234 select1.n4 select1 13.8328
R6235 select1.n14 select1.n2 10.6811
R6236 select1.n7 select1.n5 10.4374
R6237 select1.n9 select1.n8 8.15776
R6238 select1.n12 select1 6.61383
R6239 select1.n2 select1 6.1445
R6240 select1.n4 select1 5.16179
R6241 select1.n11 select1 4.90717
R6242 select1.n9 select1.n4 4.65206
R6243 select1.n8 select1 3.93896
R6244 select1.n12 select1.n11 2.98717
R6245 select1.n5 select1 2.16665
R6246 select1.n8 select1.n7 1.57588
R6247 select1.n13 select1.n9 0.79438
R6248 select1 select1.n14 0.248606
R6249 x4.net6.n3 x4.net6.t8 323.342
R6250 x4.net6.n0 x4.net6.t12 323.342
R6251 x4.net6.n1 x4.net6.t2 260.322
R6252 x4.net6.n8 x4.net6.t7 241.536
R6253 x4.net6.n17 x4.net6.t0 222.679
R6254 x4.net6.n12 x4.net6.t10 212.081
R6255 x4.net6.n13 x4.net6.t11 212.081
R6256 x4.net6.n3 x4.net6.t3 194.809
R6257 x4.net6.n0 x4.net6.t13 194.809
R6258 x4.net6.n5 x4.net6.t14 183.505
R6259 x4.net6.n1 x4.net6.t5 175.169
R6260 x4.net6.n8 x4.net6.t4 169.237
R6261 x4.net6 x4.net6.n3 158.133
R6262 x4.net6 x4.net6.n0 158.133
R6263 x4.net6 x4.net6.n8 157.555
R6264 x4.net6.n15 x4.net6.n14 155.52
R6265 x4.net6.n6 x4.net6.n5 153.863
R6266 x4.net6.n2 x4.net6.n1 152
R6267 x4.net6.n12 x4.net6.t6 139.78
R6268 x4.net6.n13 x4.net6.t9 139.78
R6269 x4.net6.n18 x4.net6.t1 129.078
R6270 x4.net6.n5 x4.net6.t15 114.532
R6271 x4.net6.n18 x4.net6.n17 96.7191
R6272 x4.net6.n11 x4.net6 55.2785
R6273 x4.net6.n14 x4.net6.n13 37.246
R6274 x4.net6.n14 x4.net6.n12 24.1005
R6275 x4.net6.n10 x4.net6.n9 21.4124
R6276 x4.net6.n16 x4.net6.n15 21.1949
R6277 x4.net6.n4 x4.net6.n2 20.043
R6278 x4.net6.n7 x4.net6.n6 15.2615
R6279 x4.net6.n17 x4.net6.n16 12.4213
R6280 x4.net6.n9 x4.net6 12.3175
R6281 x4.net6.n16 x4.net6.n11 8.09819
R6282 x4.net6.n11 x4.net6.n10 7.53948
R6283 x4.net6.n4 x4.net6 7.39885
R6284 x4.net6 x4.net6.n18 5.84085
R6285 x4.net6.n15 x4.net6 5.4405
R6286 x4.net6.n9 x4.net6 4.10616
R6287 x4.net6.n7 x4.net6.n4 2.60421
R6288 x4.net6.n10 x4.net6.n7 2.43577
R6289 x4.net6.n6 x4.net6 1.97868
R6290 x4.net6.n2 x4.net6 1.55726
R6291 select0.n5 select0.t1 327.99
R6292 select0.n9 select0.t8 293.969
R6293 select0.n3 select0.t3 261.887
R6294 select0.n0 select0.t7 212.081
R6295 select0.n1 select0.t9 212.081
R6296 select0.n5 select0.t0 199.457
R6297 select0.n2 select0.n1 183.185
R6298 select0.n3 select0.t6 155.847
R6299 select0 select0.n9 154.065
R6300 select0.n4 select0.n3 153.506
R6301 select0.n6 select0.n5 152
R6302 select0.n0 select0.t4 139.78
R6303 select0.n1 select0.t5 139.78
R6304 select0.n9 select0.t2 138.338
R6305 select0.n1 select0.n0 61.346
R6306 select0.n10 select0 13.4199
R6307 select0.n11 select0.n8 11.7395
R6308 select0.n12 select0.n11 11.5949
R6309 select0.n8 select0.n4 10.4004
R6310 select0.n12 select0.n2 9.68118
R6311 select0.n6 select0 9.6005
R6312 select0.n2 select0 5.8885
R6313 select0.n10 select0 5.57469
R6314 select0.n8 select0.n7 4.6505
R6315 select0.n11 select0.n10 4.6505
R6316 select0.n7 select0.n6 2.98717
R6317 select0.n4 select0 2.82403
R6318 select0.n7 select0 1.9205
R6319 select0 select0.n12 0.559212
R6320 x4.net3.t7 x4.net3.t2 395.01
R6321 x4.net3 x4.net3.t7 320.745
R6322 x4.net3.n3 x4.net3.t4 260.322
R6323 x4.net3.n0 x4.net3.t3 229.369
R6324 x4.net3.n7 x4.net3.t0 222.68
R6325 x4.net3.n3 x4.net3.t5 175.169
R6326 x4.net3.n0 x4.net3.t6 157.07
R6327 x4.net3.n4 x4.net3.n3 152
R6328 x4.net3.n1 x4.net3.n0 152
R6329 x4.net3.n8 x4.net3.t1 132.322
R6330 x4.net3.n8 x4.net3.n7 95.0273
R6331 x4.net3.n5 x4.net3 25.2581
R6332 x4.net3.n5 x4.net3 20.1696
R6333 x4.net3.n7 x4.net3.n6 12.7813
R6334 x4.net3.n1 x4.net3 12.0005
R6335 x4.net3 x4.net3.n4 11.2497
R6336 x4.net3.n6 x4.net3.n2 9.79203
R6337 x4.net3.n6 x4.net3.n5 5.9277
R6338 x4.net3.n2 x4.net3 4.53383
R6339 x4.net3 x4.net3.n8 2.70465
R6340 x4.net3.n2 x4.net3.n1 1.6005
R6341 x4.net3.n4 x4.net3 1.55726
R6342 counter7.n0 counter7.t0 368.521
R6343 counter7.n1 counter7.t1 216.155
R6344 counter7.n1 counter7 78.8791
R6345 counter7.n4 counter7.t5 26.3998
R6346 counter7.n4 counter7.t4 23.5483
R6347 counter7.n3 counter7.n2 18.2765
R6348 counter7.n5 counter7.t2 12.9758
R6349 counter7.n5 counter7.t3 10.8618
R6350 counter7 counter7.n0 10.5563
R6351 counter7.n0 counter7 5.48477
R6352 counter7.n2 counter7 4.18512
R6353 counter7.n6 counter7.n4 3.06895
R6354 counter7.n6 counter7.n5 2.14822
R6355 counter7 counter7.n6 1.27287
R6356 counter7.n3 counter7 1.27059
R6357 counter7.n2 counter7.n1 0.985115
R6358 counter7 counter7.n3 0.647091
R6359 x3.x2.GP2.n2 x3.x2.GP2.t4 450.938
R6360 x3.x2.GP2.n2 x3.x2.GP2.t5 445.666
R6361 x3.x2.GP2.n4 x3.x2.GP2.n3 195.958
R6362 x3.x2.GP2 x3.x2.GP2.n0 96.8352
R6363 x3.x2.GP2.n3 x3.x2.GP2.t1 26.5955
R6364 x3.x2.GP2.n3 x3.x2.GP2.t0 26.5955
R6365 x3.x2.GP2.n0 x3.x2.GP2.t2 24.9236
R6366 x3.x2.GP2.n0 x3.x2.GP2.t3 24.9236
R6367 x3.x2.GP2.n5 x3.x2.GP2.n4 13.0077
R6368 x3.x2.GP2.n4 x3.x2.GP2 11.995
R6369 x3.x2.GP2 x3.x2.GP2.n1 11.2645
R6370 x3.x2.GP2.n1 x3.x2.GP2 6.1445
R6371 x3.x2.GP2.n1 x3.x2.GP2 4.65505
R6372 x3.x2.GP2 x3.x2.GP2.n2 3.12839
R6373 x3.x2.GP2.n5 x3.x2.GP2 2.0485
R6374 x3.x2.GP2 x3.x2.GP2.n5 1.55202
R6375 counter3.n0 counter3.t2 368.521
R6376 counter3.n1 counter3.t3 216.155
R6377 counter3.n1 counter3 78.8791
R6378 counter3.n4 counter3.t0 26.3998
R6379 counter3.n4 counter3.t1 23.5483
R6380 counter3.n3 counter3.n2 17.5689
R6381 counter3.n5 counter3.t4 12.9693
R6382 counter3.n5 counter3.t5 10.8444
R6383 counter3 counter3.n0 10.5563
R6384 counter3.n0 counter3 5.48477
R6385 counter3.n2 counter3 4.18512
R6386 counter3.n6 counter3.n4 3.06895
R6387 counter3.n6 counter3.n5 2.14822
R6388 counter3.n3 counter3 1.28175
R6389 counter3 counter3.n6 1.25828
R6390 counter3.n2 counter3.n1 0.985115
R6391 counter3 counter3.n3 0.688
R6392 x4._16_.n12 x4._16_.t0 339.418
R6393 x4._16_ x4._16_.t1 269.426
R6394 x4._16_.n1 x4._16_.t2 264.029
R6395 x4._16_ x4._16_.n5 241.976
R6396 x4._16_.n3 x4._16_.t9 241.536
R6397 x4._16_.n5 x4._16_.t5 241.536
R6398 x4._16_.n1 x4._16_.t6 206.19
R6399 x4._16_.n4 x4._16_.n3 171.332
R6400 x4._16_.n3 x4._16_.t7 169.237
R6401 x4._16_.n5 x4._16_.t4 169.237
R6402 x4._16_.n2 x4._16_.n1 160.96
R6403 x4._16_.n9 x4._16_.n8 153.165
R6404 x4._16_.n8 x4._16_.t3 144.548
R6405 x4._16_.n8 x4._16_.t8 128.482
R6406 x4._16_.n7 x4._16_.n2 21.45
R6407 x4._16_.n7 x4._16_.n6 16.7975
R6408 x4._16_.n10 x4._16_ 15.8161
R6409 x4._16_.n11 x4._16_.n10 14.0946
R6410 x4._16_ x4._16_.n0 11.2645
R6411 x4._16_ x4._16_.n9 9.55788
R6412 x4._16_.n6 x4._16_ 6.4005
R6413 x4._16_.n0 x4._16_ 6.1445
R6414 x4._16_.n2 x4._16_ 5.4405
R6415 x4._16_.n0 x4._16_ 4.63498
R6416 x4._16_.n4 x4._16_ 4.44132
R6417 x4._16_.n11 x4._16_ 4.3525
R6418 x4._16_.n13 x4._16_.n12 4.0914
R6419 x4._16_ x4._16_.n13 3.61789
R6420 x4._16_.n9 x4._16_ 3.29747
R6421 x4._16_.n13 x4._16_.n11 2.3045
R6422 x4._16_.n12 x4._16_ 1.74382
R6423 x4._16_.n6 x4._16_.n4 1.50638
R6424 x4._16_.n10 x4._16_.n7 1.38649
R6425 enable_ring.n0 enable_ring.t0 212.081
R6426 enable_ring.n1 enable_ring.t2 212.081
R6427 enable_ring enable_ring.n2 152.512
R6428 enable_ring.n0 enable_ring.t1 139.78
R6429 enable_ring.n1 enable_ring.t3 139.78
R6430 enable_ring.n2 enable_ring.n0 30.6732
R6431 enable_ring.n2 enable_ring.n1 30.6732
R6432 enable_ring.n3 enable_ring 16.4378
R6433 enable_ring.n3 enable_ring 0.7505
R6434 enable_ring enable_ring.n3 0.0808571
R6435 x3.x2.GP1.n2 x3.x2.GP1.t4 450.938
R6436 x3.x2.GP1.n2 x3.x2.GP1.t5 445.666
R6437 x3.x2.GP1.n4 x3.x2.GP1.n3 195.832
R6438 x3.x2.GP1 x3.x2.GP1.n0 96.8352
R6439 x3.x2.GP1.n3 x3.x2.GP1.t1 26.5955
R6440 x3.x2.GP1.n3 x3.x2.GP1.t0 26.5955
R6441 x3.x2.GP1.n0 x3.x2.GP1.t3 24.9236
R6442 x3.x2.GP1.n0 x3.x2.GP1.t2 24.9236
R6443 x3.x2.GP1.n5 x3.x2.GP1.n4 13.1346
R6444 x3.x2.GP1.n4 x3.x2.GP1 12.2007
R6445 x3.x2.GP1 x3.x2.GP1.n1 11.2645
R6446 x3.x2.GP1.n1 x3.x2.GP1 6.1445
R6447 x3.x2.GP1.n1 x3.x2.GP1 4.65505
R6448 x3.x2.GP1 x3.x2.GP1.n2 3.07707
R6449 x3.x2.GP1.n5 x3.x2.GP1 2.0485
R6450 x3.x2.GP1 x3.x2.GP1.n5 1.55202
C0 x4._20_ x4.clknet_1_1__leaf_clk 0.0051f
C1 a_28031_n8709# a_28565_n8715# 0.002698f
C2 a_26593_n7906# x4._15_ 1.57e-19
C3 a_25875_n7395# a_25600_n8741# 7.28e-21
C4 x4._11_ x4.clknet_1_1__leaf_clk 0.367667f
C5 a_18409_n2290# a_18585_n1958# 0.185422f
C6 a_17857_n2290# x3.x2.GN1 0.012445f
C7 x4.net8 a_27055_n8715# 0.00311f
C8 x4.clknet_0_clk a_25709_n7109# 1.74729f
C9 x4.net7 a_28579_n7627# 5.4e-19
C10 x4.net3 a_23851_n9829# 0.002183f
C11 a_23421_n7921# x4.net6 4.71e-21
C12 a_28031_n7261# a_27755_n7261# 0.00119f
C13 a_26529_n7849# a_26798_n8741# 1e-18
C14 a_28031_n7261# x4.net7 5.71e-19
C15 a_23946_n9147# a_23778_n8893# 0.239923f
C16 a_23505_n9259# a_24371_n8991# 0.034054f
C17 x4._21_ a_25639_n9259# 0.087922f
C18 a_27055_n8715# x4._07_ 0.009837f
C19 x4.net8 x4._22_ 0.137056f
C20 a_23615_n8171# a_24371_n8991# 3.85e-19
C21 a_27124_n9259# a_26998_n8893# 0.005525f
C22 x4._04_ a_23778_n8893# 3.52e-21
C23 x4.clknet_1_0__leaf_clk x4._16_ 4.14e-20
C24 x1.sky130_fd_sc_hd__inv_2_6.A select0 2.42e-19
C25 x4.counter[9] VDD 0.449609f
C26 select0 x3.x2.GP1 8.3e-19
C27 x4._11_ a_28470_n8893# 5.04e-19
C28 a_26159_n7409# a_26375_n8171# 2.84e-21
C29 a_25709_n7109# a_25779_n7395# 0.022122f
C30 a_27807_n9829# a_28457_n9803# 0.010893f
C31 a_23675_n5233# a_23882_n5174# 0.260055f
C32 x4.net4 a_25729_n8395# 7.88e-20
C33 a_23295_n5219# x4._01_ 1.56e-19
C34 a_23391_n5219# a_23811_n5073# 0.036838f
C35 x4._17_ a_25211_n9231# 6.88e-22
C36 x4._22_ x4._07_ 0.503878f
C37 a_27194_n8171# a_27423_n8893# 0.001605f
C38 a_23682_n5329# x4._00_ 4.06e-19
C39 x4._11_ x4._03_ 0.00174f
C40 a_29133_n9803# x4._23_ 0.113094f
C41 a_28551_n9803# a_28725_n10182# 2.21e-19
C42 VDD a_24229_n5073# 0.074934f
C43 a_27223_n8741# x4.net9 0.007609f
C44 VDD a_28197_n8709# 0.31297f
C45 a_26725_n8715# x4.clknet_1_1__leaf_clk 0.002214f
C46 x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_7.A 5.04e-19
C47 x4._24_ a_28999_n7408# 0.006166f
C48 a_28399_n7627# x4._25_ 0.001476f
C49 VDD a_28638_n9147# 0.186041f
C50 x4._22_ a_28647_n9483# 1.37e-20
C51 x4.net4 x4.net8 0.001699f
C52 a_26366_n7350# x4._06_ 2.41e-19
C53 a_27807_n9829# x4._15_ 0.086673f
C54 m2_17442_n2443# select0 0.130999f
C55 a_23682_n4633# a_23682_n5329# 0.027204f
C56 a_23675_n4933# a_23675_n5233# 0.040702f
C57 a_28895_n8715# x4._09_ 0.001217f
C58 VDD x4.net1 1.47718f
C59 x4.net9 a_26457_n7849# 0.004319f
C60 a_28031_n9259# a_28565_n8893# 0.002698f
C61 x4._09_ a_28385_n9259# 0.129132f
C62 VDD x3.x2.GN2 0.602894f
C63 a_23615_n5995# x4._10_ 0.107891f
C64 VDD a_23339_n9259# 0.741952f
C65 a_23682_n4633# x4._00_ 0.208988f
C66 a_24769_n9465# x4._15_ 1.81e-19
C67 a_26159_n7409# x4._19_ 0.074331f
C68 a_25639_n9259# x4.net7 0.003261f
C69 x4._17_ x4.clknet_1_1__leaf_clk 0.044595f
C70 a_28470_n8715# a_28596_n8337# 0.005525f
C71 x4.net3 a_24075_n5995# 0.001478f
C72 x4._18_ a_24095_n8741# 3.26e-20
C73 VDD x4._13_ 0.524973f
C74 x4._16_ a_25721_n9259# 0.00109f
C75 a_25823_n8395# x4._15_ 0.004604f
C76 x4._11_ x4.clknet_0_clk 0.042991f
C77 VDD ring_out 4.36358f
C78 x4.net8 a_25793_n9259# 8.5e-20
C79 x4.net10 x4._22_ 0.074459f
C80 a_25900_n8197# x4._16_ 0.035189f
C81 x4._12_ a_24075_n5995# 0.026119f
C82 x4._16_ x4._15_ 0.656968f
C83 x4.clknet_1_0__leaf_clk a_23778_n8893# 0.003461f
C84 VDD a_26713_n7249# 0.085296f
C85 x4.net8 a_26756_n8337# 4.88e-19
C86 select1 x3.x2.GN2 0.108649f
C87 x4.net8 a_25834_n7921# 0.063158f
C88 x4._14_ a_22837_n10182# 0.001394f
C89 a_24054_n7805# a_23969_n8171# 0.037333f
C90 a_23781_n8171# a_24563_n7805# 4.04e-19
C91 a_25779_n7395# x4._20_ 1.63e-20
C92 VDD a_23610_n4907# 4.59e-19
C93 a_26191_n8709# a_26147_n9107# 1.28e-19
C94 VDD x4.counter[1] 0.343446f
C95 x4._13_ a_23421_n7921# 0.01129f
C96 a_25639_n9259# x4.net5 5.06e-20
C97 x4._11_ a_25779_n7395# 8.65e-19
C98 x4.counter[9] a_28725_n10182# 2.34e-19
C99 x4.clknet_1_1__leaf_clk x4._23_ 0.071442f
C100 a_28743_n9483# a_28457_n9803# 0.010132f
C101 VDD a_23225_n7109# 1.52032f
C102 a_24625_n8715# x4._11_ 2.49e-20
C103 a_23969_n8171# x4._11_ 0.020189f
C104 ring_out select1 0.016625f
C105 x4.net9 a_28457_n9803# 0.008597f
C106 a_25875_n7395# x4._05_ 9.72e-20
C107 x4.net4 a_23946_n9147# 0.007782f
C108 x4._01_ a_24058_n5451# 5.75e-19
C109 a_26191_n8709# a_26559_n9259# 0.012779f
C110 x4.clknet_1_0__leaf_clk x4._10_ 0.006812f
C111 x4._14_ a_24095_n8741# 1.02e-20
C112 x4.net5 a_25297_n9231# 2.72e-19
C113 a_28638_n8741# x4._23_ 0.006211f
C114 a_27223_n8741# a_27055_n8715# 0.310858f
C115 a_17857_n2290# a_17985_n1898# 0.004764f
C116 x4.net4 x4._04_ 0.689049f
C117 VDD a_26381_n9259# 9.47e-20
C118 VDD a_23295_n4755# 0.415615f
C119 x3.x2.GN3 counter7 0.005062f
C120 x4._18_ x4._06_ 3.12e-20
C121 a_26979_n9829# x4.net6 0.211407f
C122 a_28470_n8893# x4._23_ 0.011058f
C123 VDD a_25359_n7627# 0.185924f
C124 m3_18876_n6983# x3.x2.GP2 2.65e-20
C125 a_29063_n8991# x4.net7 8.32e-20
C126 drv_out counter3 1.91048f
C127 x4._17_ a_26117_n7627# 0.002375f
C128 drv_out x4.net9 4.05e-20
C129 a_28725_n10182# a_28638_n9147# 2.21e-20
C130 a_29133_n9803# x4.net11 0.01512f
C131 a_28743_n9483# x4._15_ 0.001637f
C132 a_24095_n8741# a_23994_n9687# 6.81e-19
C133 a_26545_n8715# x4.net9 1.41e-19
C134 a_26798_n8741# x4.clknet_1_1__leaf_clk 0.01748f
C135 a_25211_n9465# a_25211_n9231# 0.012876f
C136 a_24220_n9483# a_23505_n9259# 4.63e-19
C137 VDD a_24011_n8715# 0.007439f
C138 a_27223_n8741# x4._22_ 4.4e-21
C139 x4.net10 a_29103_n9829# 0.104575f
C140 VDD a_27194_n8171# 1.3575f
C141 mux_out x3.x2.GN4 0.446429f
C142 a_25875_n7395# a_26295_n7249# 0.036838f
C143 x4.net9 x4._15_ 0.08758f
C144 a_26159_n7409# a_26366_n7350# 0.260055f
C145 a_26725_n9259# a_26998_n8893# 0.074022f
C146 a_26559_n9259# a_27591_n8991# 0.048748f
C147 a_23615_n8171# a_24220_n9483# 4.07e-21
C148 x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_6.A 0.17253f
C149 x4.clknet_1_0__leaf_clk a_22879_n5451# 3.26e-19
C150 x4.clknet_0_clk x4._17_ 0.029087f
C151 x4._06_ a_26191_n8709# 0.091082f
C152 x4._05_ x4._25_ 4.6e-21
C153 x4._21_ a_25875_n7395# 9.57e-19
C154 x4.net8 a_28551_n9803# 6.89e-20
C155 a_23615_n5995# a_23697_n5995# 0.005167f
C156 m3_18862_n5953# x3.x2.GN4 7.07e-19
C157 a_24058_n4541# x4.net1 4.16e-19
C158 a_26913_n9259# x4.clknet_1_1__leaf_clk 0.011819f
C159 a_23675_n5233# a_24075_n5995# 4.04e-19
C160 x4._02_ a_24595_n8741# 7.66e-20
C161 VDD a_28579_n7627# 0.178246f
C162 x4._04_ a_25834_n7921# 3.15e-21
C163 x4._17_ a_25779_n7395# 0.0702f
C164 a_27755_n7261# a_27837_n7261# 0.005781f
C165 a_29063_n8741# x4._24_ 0.009415f
C166 VDD a_28031_n7261# 0.002272f
C167 x4.net7 a_27837_n7261# 0.003849f
C168 x4.net3 x4._01_ 0.006403f
C169 x4.net8 x4.net6 0.806426f
C170 ring_out a_19207_65# 0.105448f
C171 a_28895_n8893# x4._24_ 0.012283f
C172 a_25709_n7109# x4._06_ 1.96e-20
C173 x4._16_ a_24371_n8991# 1.37e-19
C174 VDD x1.sky130_fd_sc_hd__nand2_2_0.B 0.787508f
C175 a_24222_n8059# a_23927_n8715# 0.004484f
C176 a_24054_n7805# a_24095_n8741# 0.004197f
C177 x4.clknet_0_clk x4._23_ 2.29e-20
C178 a_28647_n9483# a_28551_n9803# 1.26e-19
C179 x4._07_ x4.net6 0.066033f
C180 VDD a_23295_n5219# 0.399249f
C181 x4._01_ x4._12_ 0.353697f
C182 x4._08_ a_28385_n8715# 0.134213f
C183 a_26147_n9107# x4._20_ 0.113204f
C184 x4._11_ a_24095_n8741# 0.033019f
C185 a_18033_n1958# x3.x2.GN2 0.017071f
C186 VDD a_29489_n9803# 0.009314f
C187 x4.net4 x4.clknet_1_0__leaf_clk 0.158995f
C188 x4._11_ a_26147_n9107# 0.046716f
C189 x4.net11 x4.clknet_1_1__leaf_clk 1.82e-20
C190 x4.counter[8] counter7 0.068429f
C191 a_25875_n7395# x4.net7 0.037726f
C192 a_23063_n8709# a_23851_n9829# 3.4e-19
C193 x4.net3 x4.net5 9.15e-21
C194 x4._22_ a_28457_n9803# 0.140356f
C195 a_25211_n9465# x4._03_ 2.93e-20
C196 x4.clknet_1_0__leaf_clk a_23697_n5995# 2.61e-19
C197 drv_out a_27055_n8715# 2.32e-21
C198 x4.counter[9] x4.net8 1.68e-20
C199 x4._18_ a_26159_n7409# 6.58e-19
C200 x4.clknet_0_clk a_26798_n8741# 3.18e-19
C201 x4._20_ a_26559_n9259# 0.004564f
C202 a_26529_n7849# a_26630_n8715# 0.001605f
C203 a_25297_n9465# x4.net5 0.001706f
C204 x4.net10 a_28551_n9803# 0.007482f
C205 a_23811_n4907# x4._12_ 7.61e-20
C206 a_27055_n8715# x4._15_ 0.0351f
C207 x4._11_ a_26559_n9259# 0.029022f
C208 a_25729_n8715# x4._18_ 3.94e-20
C209 VDD a_23502_n8715# 0.259474f
C210 a_28895_n8893# a_28979_n8893# 0.008508f
C211 a_24563_n7805# x4._18_ 1.72e-19
C212 VDD a_25639_n9259# 0.211123f
C213 VDD x3.x2.GN3 0.649844f
C214 a_23417_n8715# x4._02_ 0.114994f
C215 a_23633_n4541# a_23391_n4933# 0.008508f
C216 a_26529_n7849# a_26593_n7906# 0.266837f
C217 x4.net3 counter7 4.2e-20
C218 x4._22_ x4._15_ 0.422897f
C219 a_26159_n7409# a_26191_n8709# 0.001493f
C220 x4.net10 x4.net6 1.08e-19
C221 a_18409_n2290# x3.x2.GN1 6.43e-20
C222 x4.net8 a_28197_n8709# 5.19e-19
C223 x4._14_ a_24316_n9803# 0.003598f
C224 x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_6.A 5.04e-19
C225 a_27755_n7261# x4._25_ 1.87e-19
C226 x4.net2 a_23505_n9259# 3.95e-20
C227 x4._23_ a_28999_n7408# 6.47e-19
C228 a_23229_n8709# a_23946_n9147# 0.001879f
C229 x4.net7 x4._25_ 3.01e-19
C230 a_23670_n8741# a_23505_n9259# 3.46e-19
C231 x1.sky130_fd_sc_hd__inv_2_11.A x3.nselect2 1.41e-19
C232 a_25729_n8715# a_26191_n8709# 1.44e-19
C233 x4._04_ x4.net6 0.050232f
C234 a_28031_n9259# x4._24_ 0.03301f
C235 a_23946_n9147# a_24203_n8893# 0.036838f
C236 VDD a_25297_n9231# 0.00273f
C237 x4._11_ x4._06_ 0.020042f
C238 a_23615_n8171# x4.net2 2.26e-20
C239 x4._04_ a_23229_n8709# 0.011144f
C240 a_23615_n8171# a_23670_n8741# 0.002941f
C241 a_28031_n9259# a_27591_n8991# 0.001745f
C242 x4._04_ a_24203_n8893# 0.001409f
C243 a_28205_n9437# x4.clknet_1_1__leaf_clk 5.67e-20
C244 select1 x3.x2.GN3 0.273713f
C245 x4._11_ a_28895_n8893# 3.81e-21
C246 a_26366_n7350# a_26375_n8171# 1.55e-20
C247 a_25709_n7109# a_26159_n7409# 0.022305f
C248 a_28457_n9803# a_29103_n9829# 0.016298f
C249 a_23675_n5233# x4._01_ 0.092611f
C250 a_23682_n5329# a_23811_n5073# 0.124967f
C251 x4._17_ a_26147_n9107# 1.09e-21
C252 x3.x1.nSEL0 x3.x2.GN2 0.154394f
C253 drv_out a_19061_n2032# 3.86e-20
C254 x4.net4 x4._15_ 0.003757f
C255 x1.sky130_fd_sc_hd__nand2_2_0.B a_19207_65# 0.110771f
C256 VDD x1.sky130_fd_sc_hd__inv_2_9.A 0.639974f
C257 a_25229_n10182# x4.counter[4] 0.001146f
C258 select0 mux_out 4.1e-22
C259 x4._05_ a_27251_n7408# 0.121098f
C260 x4._08_ a_26191_n8709# 3.42e-20
C261 x4.counter[9] x4.net10 0.092658f
C262 VDD a_24058_n5451# 0.004407f
C263 counter7 x4.counter[2] 0.003115f
C264 a_28031_n8709# x4.net9 8.34e-19
C265 VDD a_28470_n8715# 0.247111f
C266 x4.net9 a_28197_n9259# 0.047741f
C267 x4._17_ a_26559_n9259# 1.69e-21
C268 x4._22_ a_29321_n9483# 3.34e-21
C269 ring_out x3.x1.nSEL0 1.86e-21
C270 VDD a_29063_n8991# 0.462064f
C271 x3.x2.GN4 counter7 3.94045f
C272 x4._08_ x4._24_ 0.423487f
C273 a_23675_n4933# a_23882_n5174# 6.88e-20
C274 a_23882_n4933# a_23682_n5329# 1.26e-19
C275 a_23811_n4907# a_23675_n5233# 5.28e-20
C276 a_27223_n8741# x4.net6 0.002597f
C277 a_25793_n9259# x4._15_ 2.18e-19
C278 x4.net9 a_28979_n8715# 1.06e-19
C279 a_23882_n4933# x4._00_ 0.00938f
C280 x4._16_ a_24220_n9483# 3.76e-19
C281 a_26366_n7350# x4._19_ 0.034076f
C282 mux_out x3.x2.GP1 0.352376f
C283 a_28197_n8709# x4.net10 5.04e-19
C284 a_28638_n8741# a_29021_n8337# 4.67e-20
C285 x4.counter[8] VDD 0.228646f
C286 a_25900_n8197# a_25834_n7921# 0.221119f
C287 a_26457_n7849# x4.net6 4.57e-19
C288 x4._18_ a_24595_n8741# 0.002375f
C289 x4._16_ a_26309_n9259# 7.06e-20
C290 x4.net10 a_28638_n9147# 1.26e-19
C291 a_18585_n1958# x3.x2.GP3 5.21e-19
C292 a_26756_n8337# x4._15_ 0.002542f
C293 a_25834_n7921# x4._15_ 5.11e-20
C294 x3.nselect2 a_18585_n1958# 6.01e-20
C295 x4._17_ x4._06_ 0.001225f
C296 x4.net8 a_26381_n9259# 5.79e-19
C297 x4.clknet_1_0__leaf_clk x4.net6 6.56e-20
C298 x4._03_ a_23505_n9259# 0.260627f
C299 a_23339_n9259# a_23946_n9147# 0.141453f
C300 m3_18862_n5953# x3.x2.GP1 3.25e-21
C301 a_23682_n4633# a_23882_n4933# 0.074815f
C302 a_26529_n7849# x4._16_ 0.113309f
C303 a_24229_n4907# x4.net2 1.04e-19
C304 a_26559_n9259# x4._23_ 3.56e-21
C305 x4.clknet_1_0__leaf_clk a_23229_n8709# 0.158653f
C306 a_26725_n9259# x4.net7 0.030766f
C307 a_26885_n10182# a_26725_n9259# 1.2e-20
C308 x4._04_ a_23339_n9259# 2.08e-19
C309 a_23615_n8171# x4._03_ 4.31e-20
C310 VDD a_27837_n7261# 0.001434f
C311 x4.clknet_1_0__leaf_clk a_24203_n8893# 6.12e-19
C312 a_24479_n7805# a_24625_n8715# 1.65e-19
C313 x4._14_ a_24125_n10182# 4.42e-19
C314 a_23781_n8171# a_25762_n7921# 1.01e-20
C315 counter7 a_23205_n10182# 2.81e-20
C316 x4.net8 a_27194_n8171# 0.001798f
C317 a_24222_n8059# a_24180_n8171# 4.62e-19
C318 VDD x4.net3 2.1402f
C319 x4._11_ a_28031_n9259# 0.012822f
C320 a_25779_n7395# a_25667_n8171# 2.76e-20
C321 x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_5.A 0.17253f
C322 a_23693_n9259# x4.net5 2.02e-19
C323 x4.counter[9] a_29645_n10182# 0.039377f
C324 x4._11_ a_26159_n7409# 2.33e-19
C325 x4._13_ x4._04_ 1.41e-19
C326 x4.net1 a_23615_n5995# 0.232539f
C327 drv_out x3.x2.GP3 0.077808f
C328 x4._08_ a_28979_n8893# 1.22e-19
C329 a_25729_n8715# x4._20_ 1.05e-19
C330 a_26630_n8715# x4.clknet_1_1__leaf_clk 0.033626f
C331 VDD a_25297_n9465# 0.002731f
C332 a_28551_n9803# a_28457_n9803# 0.062574f
C333 a_24125_n10182# a_23994_n9687# 0.002548f
C334 a_29321_n9483# a_29103_n9829# 0.007234f
C335 a_27194_n8171# x4._07_ 0.022424f
C336 a_25729_n8715# x4._11_ 0.07562f
C337 a_24563_n7805# x4._11_ 0.002344f
C338 a_26166_n7505# x4._05_ 0.181338f
C339 x4.net4 a_24371_n8991# 0.020834f
C340 VDD x4._12_ 0.307826f
C341 a_26798_n8741# a_26559_n9259# 1.62e-19
C342 a_26357_n8709# a_26725_n9259# 1.17e-19
C343 a_26191_n8709# a_27166_n9147# 3.92e-19
C344 x4._14_ a_24595_n8741# 1.74e-20
C345 x4.net9 a_26309_n9259# 8.5e-21
C346 a_29063_n8741# x4._23_ 1.75e-20
C347 a_27055_n8715# a_28031_n8709# 1.07e-19
C348 a_18033_n1958# x3.x2.GN3 0.048646f
C349 a_27223_n8741# a_28197_n8709# 2.73e-19
C350 VDD a_27124_n9259# 1.42e-19
C351 a_23421_n7921# x4.net3 0.001185f
C352 a_28457_n9803# x4.net6 5.59e-20
C353 a_28895_n8893# x4._23_ 0.006274f
C354 VDD a_25875_n7395# 0.175351f
C355 a_28385_n9259# x4.net7 2.26e-19
C356 VDD x1.sky130_fd_sc_hd__inv_2_7.Y 0.636657f
C357 a_23610_n5085# x4.net1 1.42e-19
C358 a_27251_n7408# x4.net7 0.030401f
C359 a_28551_n9803# x4._15_ 0.038186f
C360 a_26529_n7849# x4.net9 0.170073f
C361 x4._04_ a_23225_n7109# 0.00168f
C362 VDD a_24981_n8715# 0.009139f
C363 a_28031_n8709# x4._22_ 5.82e-21
C364 x4._18_ x4._19_ 0.036736f
C365 VDD a_24149_n7805# 0.003961f
C366 a_26166_n7505# a_26295_n7249# 0.110715f
C367 a_27166_n9147# a_27591_n8991# 1.28e-19
C368 a_26725_n9259# a_27423_n8893# 0.193199f
C369 a_26559_n9259# a_26913_n9259# 0.062224f
C370 x4._08_ x4._11_ 1.44e-20
C371 x4._22_ a_28197_n9259# 3.15e-20
C372 drv_out x4.net6 2.01e-20
C373 VDD x4.counter[2] 0.494839f
C374 ring_out x1.sky130_fd_sc_hd__inv_2_11.A 0.167117f
C375 x4.clknet_1_0__leaf_clk a_24229_n5073# 0.018091f
C376 x4._06_ a_26798_n8741# 0.001008f
C377 a_26545_n8715# x4.net6 0.008614f
C378 a_25709_n7109# a_26375_n8171# 2.81e-20
C379 a_25900_n8197# x4.net6 0.016498f
C380 x4.counter[8] a_28725_n10182# 6.92e-19
C381 x4._21_ a_26166_n7505# 0.001538f
C382 x4.net6 x4._15_ 0.117386f
C383 a_24053_n8337# a_23927_n8715# 0.006169f
C384 x4._10_ a_23769_n5995# 5.49e-20
C385 a_23615_n5995# a_23225_n7109# 5.68e-19
C386 VDD x3.x2.GN4 1.23321f
C387 a_23781_n8171# x4._18_ 8.49e-20
C388 x4.clknet_1_0__leaf_clk x4.net1 0.561165f
C389 a_26191_n8709# x4._19_ 9.86e-21
C390 a_27194_n8171# x4.net10 3.58e-19
C391 a_23682_n5329# x4._11_ 4.06e-19
C392 a_23882_n5174# a_24075_n5995# 2.48e-20
C393 a_24203_n8893# x4._15_ 1.6e-20
C394 VDD x4._25_ 0.22908f
C395 x4.clknet_1_0__leaf_clk a_23339_n9259# 0.293401f
C396 a_23615_n8171# a_23969_n8171# 0.062224f
C397 x4._17_ a_26159_n7409# 0.42661f
C398 x4._11_ a_24125_n10182# 3.83e-19
C399 VDD a_26542_n7627# 0.004407f
C400 x4.net2 x4._16_ 5.41e-20
C401 x4._00_ x4._11_ 0.003231f
C402 x4._16_ a_23670_n8741# 1.76e-20
C403 a_28565_n8893# x4._24_ 7.21e-19
C404 x4._13_ x4.clknet_1_0__leaf_clk 0.02176f
C405 x4._16_ a_25211_n9231# 0.113241f
C406 a_27807_n9829# x4.clknet_1_1__leaf_clk 3.39e-19
C407 x4._19_ x4._24_ 8.27e-21
C408 a_25729_n8715# x4._17_ 9.12e-21
C409 x4.net8 a_25639_n9259# 7.44e-19
C410 a_26630_n8715# x4.clknet_0_clk 4.59e-20
C411 counter7 a_28385_n9259# 2.77e-20
C412 a_25709_n7109# x4._19_ 5.98e-19
C413 a_25179_n7627# x4._05_ 4.45e-20
C414 select1 x3.x2.GN4 0.059808f
C415 a_17405_n2032# select0 0.048888f
C416 VDD a_23675_n5233# 0.446206f
C417 a_23675_n4933# a_24075_n5995# 4.52e-21
C418 x4._14_ x4._02_ 0.166596f
C419 x4.net9 a_29133_n9803# 0.005829f
C420 x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_5.A 5.04e-19
C421 x4._11_ a_24595_n8741# 0.001227f
C422 a_18585_n1958# x3.x2.GN2 5.62e-20
C423 VDD a_23205_n10182# 0.272145f
C424 x3.x1.nSEL0 x3.x2.GN3 4.01e-20
C425 x4._07_ a_25639_n9259# 1.81e-20
C426 a_28638_n9147# a_28457_n9803# 3.15e-19
C427 VDD a_23505_n4043# 5.43e-19
C428 x4.clknet_0_clk a_26593_n7906# 7.62e-19
C429 x4.clknet_1_0__leaf_clk a_23610_n4907# 0.001704f
C430 x4._11_ a_23873_n8893# 6.67e-19
C431 a_28031_n9259# x4._23_ 0.029061f
C432 x4._09_ x4.net7 2.46e-19
C433 a_23781_n8171# x4._14_ 3.24e-22
C434 a_26166_n7505# x4.net7 0.027472f
C435 x4.clknet_1_0__leaf_clk a_23225_n7109# 1.67275f
C436 ring_out a_18585_n1958# 2.55e-19
C437 x4._16_ x4.clknet_1_1__leaf_clk 0.001692f
C438 x4._18_ a_26366_n7350# 5.4e-20
C439 x4._20_ a_27166_n9147# 6.25e-20
C440 a_27194_n8171# a_27223_n8741# 0.009572f
C441 a_27181_n8337# x4.net7 1.38e-19
C442 x4.net2 counter3 0.003151f
C443 x4.net10 a_29489_n9803# 0.003077f
C444 a_29063_n8741# x4.net11 1.16e-19
C445 a_28197_n8709# x4._15_ 0.058771f
C446 x4._11_ a_27166_n9147# 0.039242f
C447 a_24769_n9465# x4._03_ 1.17e-19
C448 x4._11_ a_26375_n8171# 1.22e-19
C449 VDD a_23927_n8715# 0.228175f
C450 a_25762_n7921# x4._18_ 0.00112f
C451 a_28895_n8893# x4.net11 0.003417f
C452 a_28638_n9147# x4._15_ 0.002208f
C453 x4._05_ a_28399_n7627# 6.38e-20
C454 VDD x1.sky130_fd_sc_hd__inv_2_7.A 0.636415f
C455 drv_out x3.x2.GN2 3.92936f
C456 a_22885_n8715# x4._02_ 0.01416f
C457 x4.clknet_1_0__leaf_clk a_23295_n4755# 0.007095f
C458 VDD a_23693_n9259# 0.083158f
C459 a_26529_n7849# x4._22_ 0.019192f
C460 a_26366_n7350# a_26191_n8709# 2.08e-22
C461 x4._11_ a_29021_n9259# 9.67e-22
C462 a_26159_n7409# a_26798_n8741# 2.9e-20
C463 a_26166_n7505# a_26357_n8709# 6.46e-19
C464 a_23295_n5219# a_23615_n5995# 3.66e-19
C465 x4.net8 a_28470_n8715# 2.79e-19
C466 x4.clknet_1_0__leaf_clk a_24011_n8715# 3.7e-19
C467 ring_out x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C468 x4.net4 a_24220_n9483# 0.01239f
C469 a_24095_n8741# a_23505_n9259# 0.00183f
C470 a_28385_n8715# a_26191_n8709# 2.33e-21
C471 ring_out drv_out 2.13841f
C472 x4._08_ x4._23_ 0.030554f
C473 x4._21_ a_25600_n8741# 0.005326f
C474 a_24371_n8991# a_24203_n8893# 0.310858f
C475 x4._06_ a_25667_n8171# 4.79e-19
C476 VDD a_26725_n9259# 0.323392f
C477 x4._16_ x4._03_ 0.005745f
C478 m2_17442_n2443# a_17405_n2032# 0.01297f
C479 a_25359_n7627# a_25449_n7261# 0.004764f
C480 x4._04_ a_23502_n8715# 3.3e-20
C481 a_23615_n8171# a_24095_n8741# 4.12e-19
C482 x4._09_ a_27423_n8893# 1.4e-19
C483 a_23417_n8715# x4._11_ 2.52e-19
C484 x1.sky130_fd_sc_hd__inv_2_7.A select1 2.42e-19
C485 counter7 x4._09_ 5.27e-21
C486 a_28385_n8715# x4._24_ 4.8e-19
C487 x1.sky130_fd_sc_hd__inv_2_8.Y select0 1.18e-19
C488 x4._11_ x4._19_ 0.032711f
C489 a_25709_n7109# a_26366_n7350# 0.007109f
C490 x4.net9 x4.clknet_1_1__leaf_clk 0.461828f
C491 a_18409_n2290# x3.x2.GP2 3.07e-19
C492 a_23882_n5174# x4._01_ 0.004715f
C493 a_23295_n5219# a_23610_n5085# 7.84e-20
C494 a_23781_n8171# a_24054_n7805# 0.074434f
C495 x4.net2 x4._10_ 0.006086f
C496 x4._11_ x4._02_ 0.012298f
C497 x4._08_ a_26798_n8741# 9.82e-20
C498 a_28551_n9803# a_28197_n9259# 1.65e-19
C499 a_25179_n7627# x4.net7 2.88e-19
C500 a_28638_n8741# x4.net9 2.66e-21
C501 a_23781_n8171# x4._11_ 0.082924f
C502 VDD a_28895_n8715# 0.233266f
C503 x4.net9 a_28470_n8893# 0.023502f
C504 a_27194_n8171# a_28457_n9803# 1.15e-20
C505 x4._22_ a_29133_n9803# 6.52e-20
C506 VDD a_28385_n9259# 0.079695f
C507 a_18409_n2290# a_18537_n1898# 0.004764f
C508 VDD a_27251_n7408# 0.209324f
C509 x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_4.A 0.17253f
C510 VDD select0 2.53226f
C511 a_23811_n4907# a_23882_n5174# 1.77e-19
C512 x4.clknet_1_0__leaf_clk a_23295_n5219# 0.01132f
C513 a_23675_n4933# x4._01_ 6.79e-20
C514 a_23882_n4933# a_23811_n5073# 1.77e-19
C515 x4.clknet_0_clk x4._16_ 0.019509f
C516 x1.sky130_fd_sc_hd__inv_2_11.A x3.x2.GN3 7.01e-21
C517 a_28031_n8709# x4.net6 2.14e-19
C518 a_22879_n5451# x4.net2 0.07281f
C519 x4._09_ a_28596_n9259# 3.07e-19
C520 a_28031_n9259# x4.net11 3.07e-19
C521 VDD a_23063_n8709# 0.684183f
C522 a_23633_n4541# x4._00_ 3.7e-19
C523 a_25600_n8741# x4.net7 0.142058f
C524 x4.net2 x4.counter[0] 0.010591f
C525 a_25359_n7627# x4._15_ 2e-21
C526 a_27194_n8171# drv_out 1.27e-19
C527 x4.counter[4] x4.net5 0.001223f
C528 a_29063_n8741# a_29021_n8337# 7.84e-20
C529 a_28470_n8715# x4.net10 3.33e-19
C530 a_25834_n7921# a_26529_n7849# 5.89e-19
C531 a_25229_n10182# x4.net5 0.233889f
C532 x4._18_ a_26191_n8709# 5.99e-21
C533 x4.net10 a_29063_n8991# 0.008159f
C534 x3.x2.GN1 x3.x2.GP3 0.002437f
C535 a_27194_n8171# x4._15_ 0.047247f
C536 a_25779_n7395# x4._16_ 3.45e-20
C537 x4.net7 a_28399_n7627# 6.19e-19
C538 x1.sky130_fd_sc_hd__inv_2_13.A x3.x2.GN2 3.88e-22
C539 x4._03_ a_23778_n8893# 0.010537f
C540 a_23339_n9259# a_24371_n8991# 0.048748f
C541 VDD x1.sky130_fd_sc_hd__inv_2_6.A 0.636415f
C542 x4.net8 a_25875_n7395# 1.55e-19
C543 VDD x3.x2.GP1 1.86414f
C544 a_23675_n4933# a_23811_n4907# 0.141453f
C545 a_23682_n4633# a_23633_n4541# 6.32e-19
C546 a_24625_n8715# x4._16_ 0.059496f
C547 a_26630_n8715# a_26559_n9259# 2.14e-19
C548 select0 select1 3.46737f
C549 a_26998_n8893# x4.net7 0.005696f
C550 x4.clknet_1_0__leaf_clk a_23502_n8715# 0.032164f
C551 x4.counter[8] x4.net10 0.009948f
C552 counter7 x4.counter[4] 0.007159f
C553 x4._17_ x4._19_ 0.214371f
C554 counter7 a_25229_n10182# 2.81e-20
C555 a_24479_n7805# a_24563_n7805# 0.008508f
C556 x1.sky130_fd_sc_hd__inv_2_9.A x1.sky130_fd_sc_hd__inv_2_11.A 0.001676f
C557 x4._11_ a_26366_n7350# 3.53e-20
C558 x4._15_ a_28579_n7627# 0.001357f
C559 x4.clknet_0_clk x4.net9 0.132797f
C560 a_28031_n7261# x4._15_ 0.001194f
C561 a_29133_n9803# a_29103_n9829# 0.025037f
C562 a_27055_n8715# x4.clknet_1_1__leaf_clk 0.024694f
C563 x4.net4 x4.net2 8.49e-21
C564 a_23781_n8171# x4._17_ 9.29e-21
C565 a_25762_n7921# x4._11_ 0.002546f
C566 x4.net4 a_23670_n8741# 5.24e-19
C567 a_26295_n7249# x4._05_ 0.001005f
C568 x1.sky130_fd_sc_hd__inv_2_6.A select1 8.27e-22
C569 x4.net3 a_23946_n9147# 3.22e-20
C570 x4.net4 a_25211_n9231# 4.87e-19
C571 m2_17442_n2443# VDD 0.14037f
C572 select1 x3.x2.GP1 8.45e-19
C573 a_26357_n8709# a_26998_n8893# 7.62e-19
C574 a_26630_n8715# x4._06_ 3.32e-19
C575 x4._22_ x4.clknet_1_1__leaf_clk 0.031888f
C576 a_25709_n7109# a_26191_n8709# 3.84e-19
C577 x4.net9 a_27507_n8893# 8.89e-19
C578 x4.net2 a_23697_n5995# 6.45e-19
C579 a_18585_n1958# x3.x2.GN3 0.004288f
C580 VDD x4._09_ 0.262387f
C581 a_28031_n8709# a_28197_n8709# 0.970499f
C582 x4._04_ x4.net3 5.28e-22
C583 x3.x1.nSEL0 x3.x2.GN4 2.26e-20
C584 x3.x2.GP2 counter3 0.148166f
C585 a_28565_n8893# x4._23_ 8.32e-19
C586 a_28031_n8709# a_28638_n9147# 1.99e-20
C587 a_28197_n8709# a_28197_n9259# 0.027195f
C588 VDD a_26166_n7505# 0.321592f
C589 x4._19_ x4._23_ 2.58e-20
C590 x4._06_ a_26593_n7906# 9.69e-19
C591 a_28197_n9259# a_28638_n9147# 0.118966f
C592 a_26309_n9259# x4.net6 1.78e-19
C593 a_23851_n9829# x4.net5 0.006016f
C594 a_28638_n8741# x4._22_ 9.3e-20
C595 VDD a_24180_n8171# 3.37e-19
C596 x4.net2 a_23337_n4363# 0.00492f
C597 a_28197_n8709# a_28979_n8715# 6.32e-19
C598 a_27166_n9147# a_26913_n9259# 3.39e-19
C599 x4._22_ a_28470_n8893# 0.004398f
C600 x4.net3 a_23615_n5995# 0.079675f
C601 a_23941_n3056# x4.net1 0.10983f
C602 a_25721_n9259# a_25639_n9259# 0.005167f
C603 x4.clknet_1_0__leaf_clk a_24058_n5451# 0.002447f
C604 a_26529_n7849# x4.net6 0.09145f
C605 x3.x1.nSEL1 a_17857_n2290# 0.073392f
C606 x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_4.A 5.04e-19
C607 x4.counter[8] a_29645_n10182# 0.111116f
C608 m2_17442_n2443# select1 0.183786f
C609 x4._21_ a_26295_n7249# 1.21e-19
C610 a_17579_n1926# x3.x2.GN2 8.86e-19
C611 a_24813_n8395# a_24595_n8741# 0.007234f
C612 drv_out x3.x2.GN3 0.243642f
C613 a_26979_n9829# a_26725_n9259# 0.002313f
C614 a_24054_n7805# x4._18_ 5.13e-20
C615 a_25900_n8197# a_25639_n9259# 7.94e-19
C616 x4._14_ a_23994_n9687# 0.089653f
C617 x4._12_ a_23615_n5995# 0.001375f
C618 x4._01_ a_24075_n5995# 0.014882f
C619 a_25639_n9259# x4._15_ 0.080244f
C620 x4._04_ a_24981_n8715# 2.55e-19
C621 x4._17_ a_26366_n7350# 0.032936f
C622 x4._16_ a_24095_n8741# 7.03e-19
C623 a_28979_n8893# x4._24_ 8.56e-19
C624 x4._11_ x4._18_ 0.035586f
C625 x4._16_ a_26147_n9107# 1.3e-19
C626 a_25762_n7921# x4._17_ 0.002503f
C627 a_24479_n7805# a_24595_n8741# 0.001534f
C628 VDD x1.sky130_fd_sc_hd__inv_2_5.A 0.636362f
C629 x4._05_ a_27755_n7261# 1.27e-19
C630 x4._05_ x4.net7 0.232588f
C631 a_22885_n8715# x4._14_ 6.31e-19
C632 a_27549_n9259# a_27423_n8893# 0.006169f
C633 a_24222_n8059# x4.net5 1.47e-21
C634 a_25297_n9231# x4._15_ 7.85e-19
C635 a_27377_n9437# x4.net7 0.001525f
C636 a_27055_n8715# x4.clknet_0_clk 0.013741f
C637 enable_counter x4.net1 0.067291f
C638 a_18033_n1958# select0 0.143958f
C639 x4.net4 x4._03_ 0.031989f
C640 VDD a_23882_n5174# 0.271061f
C641 x4._08_ a_29021_n8337# 7.43e-19
C642 x4._12_ a_23610_n5085# 0.001666f
C643 a_22962_n5131# a_22879_n5451# 2.42e-19
C644 VDD x4.counter[4] 0.454642f
C645 counter3 a_22837_n10182# 2.11e-19
C646 x4.net1 a_23769_n5995# 0.002601f
C647 x4.net5 a_24329_n9259# 6.03e-19
C648 x4._16_ a_26559_n9259# 1.25e-20
C649 x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__inv_2_11.A 0.025028f
C650 x3.x2.GN1 x3.x2.GN2 0.065153f
C651 x4._11_ a_26191_n8709# 1.58e-19
C652 VDD a_25229_n10182# 0.316408f
C653 x4.net11 a_29021_n9259# 3e-19
C654 a_25834_n7921# x4.clknet_1_1__leaf_clk 0.007927f
C655 x4.clknet_1_0__leaf_clk x4.net3 0.373279f
C656 x4.clknet_0_clk x4._22_ 0.003156f
C657 VDD a_25179_n7627# 0.252612f
C658 x4.net8 a_26725_n9259# 0.003497f
C659 a_26630_n8715# a_26159_n7409# 8.34e-21
C660 a_24054_n7805# x4._14_ 5.19e-22
C661 a_26295_n7249# x4.net7 0.035198f
C662 a_25823_n8395# x4._06_ 6.56e-20
C663 a_26357_n8709# x4._05_ 2.65e-21
C664 a_24220_n9483# a_23339_n9259# 3.11e-19
C665 x4.net1 a_23505_n4363# 0.073427f
C666 x4._11_ x4._24_ 4.57e-19
C667 a_28385_n8715# x4._23_ 0.014354f
C668 ring_out x3.x2.GN1 4.6809f
C669 x4._20_ a_27591_n8991# 3.47e-20
C670 a_27194_n8171# a_28031_n8709# 0.016172f
C671 x4._21_ x4.net7 0.326643f
C672 a_24125_n10182# a_23505_n9259# 7.04e-21
C673 x4._07_ a_26725_n9259# 0.195848f
C674 a_18033_n1958# x3.x2.GP1 2.33e-21
C675 x4.clknet_1_0__leaf_clk x4._12_ 0.075464f
C676 VDD a_23675_n4933# 0.721856f
C677 a_26159_n7409# a_26593_n7906# 0.00484f
C678 a_27194_n8171# a_28197_n9259# 2.14e-19
C679 x4._11_ a_27591_n8991# 0.028602f
C680 a_28470_n8715# x4._15_ 0.001174f
C681 x4._11_ x4._14_ 0.007676f
C682 VDD a_25600_n8741# 0.17068f
C683 x4.net9 a_26147_n9107# 3.24e-20
C684 x4._11_ a_25709_n7109# 4.59e-19
C685 x4._06_ x4._16_ 0.064563f
C686 VDD a_24287_n8893# 0.004797f
C687 x4.clknet_0_clk a_26094_n7261# 1.49e-19
C688 a_23670_n8741# x4.net6 6.4e-20
C689 mux_out counter7 4.51509f
C690 a_23675_n5233# a_23615_n5995# 4.35e-19
C691 x4._11_ a_23994_n9687# 1e-19
C692 a_25211_n9231# x4.net6 4.93e-21
C693 VDD a_28399_n7627# 0.206381f
C694 x4.net8 a_28895_n8715# 1.1e-19
C695 a_23229_n8709# a_23670_n8741# 0.127288f
C696 x4._17_ x4._18_ 0.181987f
C697 a_24149_n7805# x4.clknet_1_0__leaf_clk 4.17e-19
C698 a_28031_n8709# a_28579_n7627# 6.06e-21
C699 a_23927_n8715# a_23946_n9147# 3.73e-19
C700 a_24095_n8741# a_23778_n8893# 0.005602f
C701 a_26725_n8715# a_26191_n8709# 0.001632f
C702 x4.net9 a_26559_n9259# 0.006834f
C703 x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_3.A 0.17253f
C704 x4._21_ a_26357_n8709# 0.002388f
C705 x4._08_ a_26630_n8715# 1.22e-20
C706 a_28197_n9259# a_28579_n7627# 3.03e-21
C707 a_24371_n8991# a_25639_n9259# 3.71e-21
C708 a_23946_n9147# a_23693_n9259# 3.39e-19
C709 VDD a_26998_n8893# 0.256044f
C710 x4._21_ x4.net5 2.83e-22
C711 VDD a_26816_n8171# 1.76e-19
C712 m3_18862_n5953# counter7 6.07e-21
C713 a_25779_n7395# a_26094_n7261# 7.84e-20
C714 x4._04_ a_23927_n8715# 0.001211f
C715 a_23615_n8171# a_24595_n8741# 0.002539f
C716 a_27175_n9437# a_26979_n9829# 0.00119f
C717 x4._12_ a_24525_n5745# 0.001754f
C718 x3.x1.nSEL0 select0 0.324822f
C719 x4._17_ a_26191_n8709# 1.12e-20
C720 VDD a_23851_n9829# 0.377321f
C721 x4.net4 a_24625_n8715# 0.005199f
C722 x4.net4 a_23969_n8171# 0.011292f
C723 a_24222_n8059# a_24647_n7903# 1.28e-19
C724 a_23781_n8171# a_24479_n7805# 0.194203f
C725 a_28031_n9259# a_27807_n9829# 2.81e-20
C726 x4.net7 a_27755_n7261# 0.168744f
C727 VDD x1.sky130_fd_sc_hd__inv_2_4.A 0.636314f
C728 x4._06_ x4.net9 0.017291f
C729 a_26885_n10182# x4.net7 0.201574f
C730 x4.clknet_1_1__leaf_clk x4.net6 0.323735f
C731 a_25834_n7921# x4.clknet_0_clk 2.03e-19
C732 a_22837_n10182# x4.counter[0] 0.109791f
C733 x4._17_ x4._24_ 0.004444f
C734 a_28551_n9803# a_28470_n8893# 7.6e-20
C735 a_23505_n4363# a_23295_n4755# 3.08e-19
C736 a_24222_n8059# a_24605_n8171# 4.67e-20
C737 a_25297_n9465# x4._15_ 0.001523f
C738 a_24054_n7805# x4._11_ 0.054008f
C739 VDD a_23628_n8337# 4.21e-19
C740 x4.net9 a_28895_n8893# 0.020729f
C741 VDD a_27549_n9259# 2.75e-19
C742 a_18585_n1958# x3.x2.GN4 0.003699f
C743 a_25709_n7109# x4._17_ 7.15e-19
C744 x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__inv_2_12.A 0.001676f
C745 x3.x1.nSEL0 x3.x2.GP1 6.21e-20
C746 x4._16_ a_24316_n9803# 0.00427f
C747 a_24229_n4907# a_23682_n5329# 4.5e-20
C748 x4.clknet_1_0__leaf_clk a_23675_n5233# 0.683552f
C749 x4._11_ x4._20_ 0.174111f
C750 a_24229_n5073# x4.net2 1.01e-21
C751 a_25900_n8197# a_25875_n7395# 0.006438f
C752 a_25834_n7921# a_25779_n7395# 3.4e-19
C753 x4.net8 a_27175_n9437# 0.005557f
C754 a_26191_n8709# x4._23_ 1.94e-21
C755 a_24229_n4907# x4._00_ 0.139872f
C756 a_26357_n8709# x4.net7 0.456298f
C757 a_25875_n7395# x4._15_ 1.09e-20
C758 a_26357_n8709# a_26885_n10182# 7.09e-22
C759 a_28895_n8715# x4.net10 0.00375f
C760 a_25823_n8395# a_25729_n8715# 1.26e-19
C761 x1.sky130_fd_sc_hd__inv_2_4.A select1 4.96e-21
C762 x4.net1 x4.net2 0.722672f
C763 VDD a_24222_n8059# 0.177502f
C764 a_26159_n7409# x4._16_ 1.49e-19
C765 x4._23_ x4._24_ 0.206353f
C766 x4.net2 a_23339_n9259# 5.19e-20
C767 a_23670_n8741# a_23339_n9259# 0.001425f
C768 a_23229_n8709# x4._03_ 1.23e-19
C769 a_23063_n8709# a_23946_n9147# 0.001786f
C770 x4._11_ a_28003_n9437# 7.08e-19
C771 x4.net8 x4._09_ 2.1e-20
C772 x3.x2.GN2 a_17985_n1898# 0.002418f
C773 drv_out x3.x2.GN4 0.071598f
C774 a_23339_n9259# a_25211_n9231# 7.98e-21
C775 x4._03_ a_24203_n8893# 0.001345f
C776 a_23682_n4633# a_24229_n4907# 0.095025f
C777 x4.net8 a_26166_n7505# 4.93e-19
C778 VDD a_24329_n9259# 4.65e-19
C779 a_23675_n4933# a_24058_n4541# 0.002698f
C780 a_25729_n8715# x4._16_ 0.008193f
C781 a_27591_n8991# x4._23_ 1.37e-20
C782 x4._13_ x4.net2 0.197255f
C783 m2_17442_n2443# x3.x1.nSEL0 3.43e-19
C784 a_27055_n8715# a_26559_n9259# 0.004606f
C785 a_27223_n8741# a_26725_n9259# 0.002689f
C786 a_28385_n8715# a_28565_n8715# 0.001229f
C787 a_27423_n8893# x4.net7 0.040127f
C788 x4._04_ a_23063_n8709# 0.001469f
C789 VDD a_24075_n5995# 0.292813f
C790 x4.clknet_1_0__leaf_clk a_23927_n8715# 0.004501f
C791 a_27805_n10182# a_27591_n8991# 2.93e-21
C792 counter7 x4.net7 6.88e-20
C793 x4.clknet_1_0__leaf_clk a_23693_n9259# 0.003207f
C794 a_26191_n8709# a_26798_n8741# 0.136009f
C795 a_24647_n7903# x4._21_ 1.76e-19
C796 counter7 a_26885_n10182# 2.81e-20
C797 x3.x2.GP2 x3.x2.GP3 0.031766f
C798 VDD mux_out 14.7592f
C799 a_23615_n8171# a_23781_n8171# 0.966818f
C800 x4._15_ x4._25_ 0.003323f
C801 x4.net6 a_26117_n7627# 1.73e-19
C802 x4._22_ a_26559_n9259# 0.019806f
C803 VDD x4._05_ 0.240335f
C804 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_3.A 5.04e-19
C805 a_26593_n7906# a_26375_n8171# 0.004465f
C806 a_28197_n8709# x4.clknet_1_1__leaf_clk 0.026802f
C807 a_27181_n8337# x4._07_ 5.27e-19
C808 a_25762_n7921# a_25667_n8171# 0.002032f
C809 a_28638_n9147# x4.clknet_1_1__leaf_clk 2.7e-19
C810 a_23610_n4907# x4.net2 2.28e-19
C811 x4.net4 a_24095_n8741# 0.110738f
C812 x4.net2 x4.counter[1] 0.015257f
C813 a_23255_n4363# a_23337_n4363# 0.006406f
C814 a_27055_n8715# x4._06_ 9.38e-20
C815 x4.clknet_0_clk x4.net6 0.087511f
C816 a_25709_n7109# a_26798_n8741# 8.05e-21
C817 x4.net9 a_28031_n9259# 0.11266f
C818 x4._17_ x4._20_ 1.89e-19
C819 x3.x2.GN1 x3.x2.GN3 0.002857f
C820 a_28031_n8709# a_28470_n8715# 0.273138f
C821 a_28197_n8709# a_28638_n8741# 0.118966f
C822 a_18537_n1898# x3.x2.GP3 4.39e-19
C823 a_23225_n7109# a_23670_n8741# 3.17e-20
C824 counter7 x4.net5 6.88e-20
C825 a_26159_n7409# x4.net9 6.06e-20
C826 x4._11_ x4._17_ 0.113734f
C827 a_28638_n8741# a_28638_n9147# 0.012451f
C828 a_28470_n8715# a_28197_n9259# 1.54e-19
C829 a_28197_n8709# a_28470_n8893# 1.54e-19
C830 VDD a_26295_n7249# 0.191062f
C831 a_26630_n8715# x4._19_ 6.46e-21
C832 x4._06_ x4._22_ 0.004416f
C833 a_28638_n9147# a_28470_n8893# 0.239923f
C834 a_28197_n9259# a_29063_n8991# 0.034054f
C835 VDD x1.sky130_fd_sc_hd__inv_2_3.A 0.636314f
C836 a_24595_n9571# x4.net5 0.081136f
C837 a_25779_n7395# x4.net6 1.76e-19
C838 VDD x4._21_ 0.492491f
C839 x4.net2 a_23295_n4755# 0.092265f
C840 a_26998_n8893# a_27093_n8893# 0.007724f
C841 x4._16_ a_24125_n10182# 4.24e-19
C842 x4.net10 x4._09_ 0.081678f
C843 a_24625_n8715# x4.net6 0.007899f
C844 x3.x1.nSEL1 a_18409_n2290# 7.84e-19
C845 a_23969_n8171# x4.net6 5.63e-21
C846 x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_12.A 0.025028f
C847 x4.clknet_1_1__leaf_clk a_26713_n7249# 3.41e-20
C848 x4.counter[5] a_25965_n10182# 4.98e-19
C849 a_25729_n8395# a_25600_n8741# 0.010132f
C850 a_23597_n8715# a_23502_n8715# 0.007724f
C851 a_24011_n8715# a_23670_n8741# 9.73e-19
C852 a_23969_n8171# a_23229_n8709# 2.83e-19
C853 a_23339_n9259# x4._03_ 0.095111f
C854 a_26979_n9829# a_26998_n8893# 1.83e-19
C855 a_24479_n7805# x4._18_ 3.43e-19
C856 a_25834_n7921# a_26147_n9107# 2.49e-20
C857 x4._14_ a_25211_n9465# 9.06e-21
C858 a_23927_n8715# x4._15_ 7.5e-20
C859 x4.clknet_1_0__leaf_clk a_23063_n8709# 0.318658f
C860 x4._11_ x4._23_ 0.090724f
C861 x1.sky130_fd_sc_hd__inv_2_3.A select1 4.96e-21
C862 x4._08_ x4.net9 0.003243f
C863 x4._04_ a_24180_n8171# 2.91e-19
C864 x4._11_ a_27805_n10182# 2.18e-19
C865 x4._18_ a_25667_n8171# 0.002103f
C866 x4._16_ a_24595_n8741# 0.243866f
C867 x4.net11 x4._24_ 0.002712f
C868 x4.net6 a_28999_n7408# 1.17e-21
C869 x4.net8 a_25600_n8741# 2.76e-19
C870 a_26725_n9259# x4._15_ 2.57e-20
C871 a_28099_n9437# x4.net7 5.42e-19
C872 a_25359_n7627# x4.clknet_1_1__leaf_clk 1.19e-21
C873 a_18585_n1958# select0 0.279858f
C874 a_28565_n8715# x4._24_ 7.21e-19
C875 x4._12_ a_24031_n5085# 0.002771f
C876 VDD x4._01_ 0.468919f
C877 VDD a_27755_n7261# 0.455589f
C878 counter3 a_24125_n10182# 5.4e-19
C879 a_29063_n8741# a_29103_n9829# 1.35e-20
C880 VDD x4.net7 1.83862f
C881 x4._11_ a_26798_n8741# 7.26e-20
C882 x4._16_ a_27166_n9147# 8.82e-22
C883 VDD a_26885_n10182# 0.315151f
C884 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_2.A 0.159172f
C885 a_28895_n8893# a_29103_n9829# 0.003595f
C886 a_27194_n8171# x4.clknet_1_1__leaf_clk 1.80017f
C887 x4._16_ a_26375_n8171# 0.036674f
C888 x4.net8 a_26998_n8893# 0.001808f
C889 a_22962_n5131# x4.net1 0.001512f
C890 a_23295_n5219# x4.net2 0.004306f
C891 x4.net8 a_26816_n8171# 1.76e-19
C892 a_25834_n7921# x4._06_ 0.111795f
C893 x4.net1 a_23391_n4933# 0.017118f
C894 a_27223_n8741# a_27181_n8337# 7.84e-20
C895 x4._20_ a_26913_n9259# 5.09e-20
C896 x1.sky130_fd_sc_hd__inv_2_12.A select0 1.1e-22
C897 a_27139_n8715# x4.net7 0.001255f
C898 x4._22_ a_28031_n9259# 4.68e-20
C899 a_27194_n8171# a_28638_n8741# 0.006157f
C900 a_18585_n1958# x3.x2.GP1 2.87e-20
C901 a_19061_n2032# a_19235_n1926# 0.006584f
C902 x4._07_ a_26998_n8893# 0.008539f
C903 drv_out a_27251_n7408# 0.012863f
C904 VDD a_23811_n4907# 0.211499f
C905 a_26366_n7350# a_26593_n7906# 3.7e-19
C906 a_26159_n7409# x4._22_ 1.01e-19
C907 a_28895_n8715# x4._15_ 2.78e-19
C908 a_27194_n8171# a_28470_n8893# 6.58e-20
C909 x4._11_ a_26913_n9259# 0.016192f
C910 a_25709_n7109# a_25667_n8171# 1.78e-20
C911 x3.x2.GN2 x3.x2.GP2 2.14737f
C912 VDD a_26357_n8709# 0.300379f
C913 x4.clknet_1_1__leaf_clk a_28579_n7627# 3.65e-19
C914 a_28385_n9259# x4._15_ 0.005742f
C915 VDD x4.net5 0.923749f
C916 VDD x1.sky130_fd_sc_hd__inv_2_2.A 0.63819f
C917 x4.clknet_0_clk a_26713_n7249# 0.004448f
C918 a_23615_n8171# x4._18_ 7.56e-20
C919 x4._17_ x4._23_ 0.082072f
C920 a_23417_n8715# x4._16_ 4.26e-21
C921 x4.net4 a_24316_n9803# 0.003167f
C922 a_24095_n8741# x4.net6 6.37e-19
C923 a_23063_n8709# x4._15_ 8.17e-21
C924 x4.net3 a_23769_n5995# 8.45e-20
C925 a_23682_n5329# x4._10_ 6.77e-19
C926 x4._11_ a_25211_n9465# 0.002917f
C927 a_23882_n5174# a_23615_n5995# 0.0033f
C928 a_26147_n9107# x4.net6 0.173962f
C929 x4._16_ x4._19_ 0.001191f
C930 ring_out x3.x2.GP2 0.080385f
C931 a_23670_n8741# a_23502_n8715# 0.239923f
C932 a_23229_n8709# a_24095_n8741# 0.034054f
C933 x4._13_ a_23969_n8171# 5.97e-20
C934 a_24180_n8171# x4.clknet_1_0__leaf_clk 3.26e-19
C935 a_28031_n8709# x4._25_ 1.01e-19
C936 a_28638_n8741# a_28579_n7627# 2.48e-20
C937 x4.net3 a_24220_n9483# 9.94e-20
C938 a_27139_n8715# a_26357_n8709# 3.14e-19
C939 x4.net8 a_27549_n9259# 5.67e-20
C940 x4.net9 a_27166_n9147# 0.007121f
C941 x4._16_ x4._02_ 3.22e-20
C942 x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_13.A 0.001676f
C943 a_23225_n7109# x4.clknet_0_clk 0.317755f
C944 a_17985_n1898# x3.x2.GN3 5.17e-20
C945 x4._08_ a_27055_n8715# 7.33e-20
C946 x3.x2.GN2 a_18537_n1898# 3.11e-20
C947 a_23778_n8893# a_23873_n8893# 0.007724f
C948 a_23946_n9147# a_24287_n8893# 9.73e-19
C949 a_23505_n9259# a_23904_n9259# 0.001351f
C950 a_25211_n9231# a_25639_n9259# 0.00155f
C951 VDD a_27423_n8893# 0.1878f
C952 x4.net9 a_26375_n8171# 0.063508f
C953 drv_out x3.x2.GP1 0.125793f
C954 VDD a_17405_n2032# 0.211635f
C955 a_23610_n4907# a_23391_n4933# 0.006169f
C956 VDD counter7 2.34126f
C957 a_27377_n9437# a_26979_n9829# 0.005781f
C958 a_26559_n9259# x4.net6 0.083542f
C959 a_23781_n8171# x4._16_ 1.01e-19
C960 x4._08_ x4._22_ 1.19e-20
C961 x4.net9 a_29021_n9259# 6.87e-19
C962 x4._11_ x4.net11 2.31e-19
C963 x1.sky130_fd_sc_hd__inv_2_2.A select1 4.1e-20
C964 x4._17_ a_26798_n8741# 1.03e-20
C965 VDD a_24595_n9571# 0.201367f
C966 a_24222_n8059# x4.net8 1.22e-20
C967 ring_out a_18537_n1898# 2.99e-20
C968 x4.clknet_0_clk a_25359_n7627# 8e-19
C969 a_25211_n9231# a_25297_n9231# 0.006584f
C970 x4._14_ a_23505_n9259# 5.98e-19
C971 x4._09_ a_28457_n9803# 0.001692f
C972 a_27805_n10182# x4._23_ 2.99e-20
C973 a_27194_n8171# x4.clknet_0_clk 0.316676f
C974 a_23391_n5219# x4.net1 0.030538f
C975 a_29133_n9803# a_29063_n8991# 1.25e-19
C976 a_27175_n9437# x4._15_ 2.85e-21
C977 a_24647_n7903# a_24605_n8171# 7.84e-20
C978 a_23295_n4755# a_23391_n4933# 0.310858f
C979 a_24479_n7805# x4._11_ 0.043928f
C980 a_23851_n9829# a_23946_n9147# 1.66e-20
C981 a_23994_n9687# a_23505_n9259# 0.010312f
C982 a_17405_n2032# select1 0.02803f
C983 VDD a_24053_n8337# 0.002609f
C984 x4.net1 a_23255_n4363# 0.224922f
C985 a_25639_n9259# x4.clknet_1_1__leaf_clk 2.42e-19
C986 a_25359_n7627# a_25779_n7395# 0.017007f
C987 x4.net9 x4._19_ 4.58e-20
C988 x4._06_ x4.net6 0.037389f
C989 VDD a_28596_n9259# -4.73e-35
C990 x3.x2.GN1 x3.x2.GN4 0.001072f
C991 a_25667_n8171# x4._20_ 6.22e-20
C992 x4.clknet_1_0__leaf_clk a_23882_n5174# 0.037641f
C993 counter3 x4._02_ 0.001266f
C994 x4._11_ a_25667_n8171# 3.73e-19
C995 a_25834_n7921# a_26159_n7409# 0.001895f
C996 x4._09_ x4._15_ 0.030214f
C997 x4.net8 a_27377_n9437# 1.72e-20
C998 a_26630_n8715# a_26191_n8709# 0.260055f
C999 a_26166_n7505# x4._15_ 1.53e-20
C1000 x4.clknet_0_clk a_28579_n7627# 1.5e-20
C1001 x4._21_ a_25729_n8395# 2.03e-19
C1002 a_28031_n7261# x4.clknet_0_clk 6.75e-20
C1003 VDD a_24647_n7903# 0.386139f
C1004 a_27181_n8337# x4._15_ 0.00162f
C1005 x1.sky130_fd_sc_hd__inv_2_13.A select0 0.001551f
C1006 a_26366_n7350# x4._16_ 1.35e-21
C1007 a_26593_n7906# a_26191_n8709# 0.004179f
C1008 x4._11_ a_28205_n9437# 0.001561f
C1009 a_24095_n8741# a_23339_n9259# 0.00142f
C1010 a_23502_n8715# x4._03_ 0.001262f
C1011 a_23882_n4933# a_24229_n4907# 0.037333f
C1012 a_23675_n4933# x4.clknet_1_0__leaf_clk 0.308902f
C1013 x4.net8 a_26295_n7249# 0.00192f
C1014 x4.net4 a_24125_n10182# 0.202764f
C1015 VDD x1.sky130_fd_sc_hd__inv_2_8.Y 0.92605f
C1016 a_22837_n10182# x4.counter[1] 0.057818f
C1017 a_27055_n8715# a_27166_n9147# 0.001204f
C1018 a_27223_n8741# a_26998_n8893# 0.003655f
C1019 a_27093_n8893# x4.net7 5.23e-19
C1020 a_26630_n8715# a_25709_n7109# 5.07e-19
C1021 a_28197_n9259# a_26725_n9259# 0.002814f
C1022 x4.net8 x4._21_ 0.333812f
C1023 counter7 a_28725_n10182# 0.110188f
C1024 x4._04_ a_24222_n8059# 0.04931f
C1025 a_23615_n8171# a_24054_n7805# 0.269567f
C1026 x4._22_ a_27166_n9147# 0.001181f
C1027 x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_13.A 0.025028f
C1028 x4.net9 a_27271_n9437# 6.97e-19
C1029 a_26979_n9829# x4.net7 0.212284f
C1030 a_23946_n9147# a_24329_n9259# 4.67e-20
C1031 x4._22_ a_26375_n8171# 9.75e-19
C1032 a_25709_n7109# a_26593_n7906# 1.03e-20
C1033 a_28470_n8715# x4.clknet_1_1__leaf_clk 0.001015f
C1034 a_26885_n10182# a_26979_n9829# 3.27e-19
C1035 VDD a_28099_n9437# 0.001259f
C1036 a_23391_n5219# a_23295_n4755# 6.79e-19
C1037 a_23295_n5219# a_23391_n4933# 6.79e-19
C1038 x4._21_ x4._07_ 4.77e-20
C1039 x4._11_ a_23505_n9259# 0.03376f
C1040 a_29063_n8991# x4.clknet_1_1__leaf_clk 1.1e-19
C1041 x4.counter[4] a_25721_n9259# 4.37e-20
C1042 x4.net3 x4.net2 1.28152f
C1043 a_24479_n7805# x4._17_ 1.03e-20
C1044 m3_18866_n4909# counter3 2.1e-20
C1045 x4.net4 a_24595_n8741# 0.005124f
C1046 a_29321_n9483# x4._09_ 0.002954f
C1047 x4._00_ a_23337_n4363# 6.18e-19
C1048 a_23255_n4363# a_23295_n4755# 1.32e-19
C1049 a_23615_n8171# x4._11_ 0.205946f
C1050 x1.sky130_fd_sc_hd__inv_2_8.Y select1 0.008686f
C1051 a_28197_n8709# a_29063_n8741# 0.034054f
C1052 a_28579_n7627# a_28999_n7408# 0.017591f
C1053 a_28638_n8741# a_28470_n8715# 0.239923f
C1054 a_28031_n8709# a_28895_n8715# 0.032244f
C1055 a_26366_n7350# x4.net9 4.56e-19
C1056 x4._17_ a_25667_n8171# 0.060488f
C1057 x4.net11 x4._23_ 0.257634f
C1058 a_28895_n8715# a_28197_n9259# 1.3e-19
C1059 a_28669_n7261# a_28579_n7627# 0.004764f
C1060 a_28197_n8709# a_28895_n8893# 1.3e-19
C1061 a_28470_n8715# a_28470_n8893# 0.013839f
C1062 x4.counter[4] x4._15_ 9.07e-20
C1063 a_25823_n8395# x4._18_ 6.01e-19
C1064 x4._12_ x4.net2 0.10227f
C1065 a_28197_n9259# a_28385_n9259# 0.097994f
C1066 a_23927_n8715# a_24220_n9483# 3.78e-21
C1067 a_28638_n9147# a_28895_n8893# 0.036838f
C1068 a_28031_n9259# x4.net6 5.6e-22
C1069 a_23615_n5995# a_24075_n5995# 0.001479f
C1070 a_26979_n9829# x4.net5 1.18e-20
C1071 VDD a_27139_n8715# 0.004428f
C1072 a_26159_n7409# x4.net6 0.001597f
C1073 a_28895_n8715# a_28979_n8715# 0.008508f
C1074 a_28565_n8715# x4._23_ 8.32e-19
C1075 x4._22_ x4._19_ 7e-20
C1076 a_26381_n9259# a_26147_n9107# 0.005167f
C1077 select0 a_17579_n1926# 9.55e-19
C1078 VDD a_23421_n7921# 0.006535f
C1079 a_25729_n8715# x4.net6 0.044713f
C1080 x4.net8 x4.net7 1.22349f
C1081 x4._18_ x4._16_ 0.283975f
C1082 VDD select1 3.78574f
C1083 x3.x2.GN3 x3.x2.GP2 2.65608f
C1084 x4.clknet_1_0__leaf_clk a_23628_n8337# 0.001807f
C1085 x4.net8 a_26885_n10182# 3.76e-19
C1086 a_25900_n8197# a_25600_n8741# 8.74e-19
C1087 a_27807_n9829# a_27591_n8991# 0.001105f
C1088 a_25600_n8741# x4._15_ 0.229149f
C1089 x4._07_ x4.net7 0.047771f
C1090 a_26381_n9259# a_26559_n9259# 1.43e-19
C1091 a_26630_n8715# x4._11_ 2.99e-20
C1092 x4._07_ a_26885_n10182# 7.51e-19
C1093 x1.sky130_fd_sc_hd__inv_2_14.A select0 1.61e-19
C1094 x4._16_ a_26191_n8709# 1.57e-19
C1095 x4._14_ a_24769_n9465# 5.76e-19
C1096 x4.net4 a_23417_n8715# 1.97e-19
C1097 a_23295_n5219# a_23391_n5219# 0.310858f
C1098 a_24222_n8059# x4.clknet_1_0__leaf_clk 5.16e-19
C1099 x3.x2.GN3 a_18537_n1898# 0.001073f
C1100 x4._19_ a_26094_n7261# 1.38e-19
C1101 x4._15_ a_28399_n7627# 0.001697f
C1102 x3.x2.GN2 a_19235_n1926# 8.14e-21
C1103 x4._08_ x4.net6 5.42e-20
C1104 x4.counter[5] a_26798_n8741# 2.7e-21
C1105 x4.net8 a_26357_n8709# 0.031957f
C1106 a_26529_n7849# a_26725_n9259# 8.41e-19
C1107 a_27194_n8171# a_26559_n9259# 4.21e-21
C1108 x4._11_ a_26593_n7906# 0.004209f
C1109 a_25834_n7921# a_26375_n8171# 4.72e-19
C1110 a_28205_n9437# x4._23_ 1.08e-20
C1111 x4.net8 x4.net5 0.002187f
C1112 a_27124_n9259# x4.clknet_1_1__leaf_clk 4.82e-19
C1113 a_23615_n8171# x4._17_ 1.5e-21
C1114 x4.net4 x4._02_ 1.19e-19
C1115 a_25875_n7395# x4.clknet_1_1__leaf_clk 1.54e-20
C1116 x3.x2.GN1 select0 0.021168f
C1117 x4.net3 x4._03_ 0.019455f
C1118 x4._12_ a_23633_n5451# 1.13e-19
C1119 a_24229_n4907# x4._11_ 2.48e-19
C1120 x4.clknet_1_0__leaf_clk a_24075_n5995# 0.00537f
C1121 x4._07_ a_26357_n8709# 0.029939f
C1122 ring_out a_19235_n1926# 1.86e-19
C1123 a_24981_n8715# x4.clknet_1_1__leaf_clk 8.24e-20
C1124 VDD a_28725_n10182# 0.303091f
C1125 x4._22_ a_27271_n9437# 0.002353f
C1126 x4._16_ x4._14_ 0.202586f
C1127 x4.net4 a_23781_n8171# 0.34974f
C1128 a_23851_n9829# x4._15_ 3.5e-20
C1129 x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_14.A 0.001676f
C1130 a_25709_n7109# x4._16_ 4.51e-19
C1131 a_25297_n9465# x4._03_ 5.07e-20
C1132 a_28031_n8709# x4._09_ 1.11e-19
C1133 a_28197_n8709# a_28031_n9259# 2.64e-19
C1134 x4.net8 a_27423_n8893# 0.007067f
C1135 a_23675_n5233# x4.net2 3.07e-19
C1136 x4.net8 counter7 6.32e-19
C1137 x4._09_ a_28197_n9259# 0.413296f
C1138 a_28031_n9259# a_28638_n9147# 0.141453f
C1139 VDD a_19207_65# 0.006305f
C1140 x4._16_ a_23994_n9687# 0.146025f
C1141 x4.net2 a_23205_n10182# 0.016821f
C1142 a_26630_n8715# a_26725_n8715# 0.007724f
C1143 x4.net10 x4.net7 6.54e-19
C1144 x4._07_ a_27423_n8893# 5.62e-20
C1145 x3.x2.GN1 x3.x2.GP1 1.51569f
C1146 x4._09_ a_28979_n8715# 1.2e-19
C1147 VDD a_24058_n4541# 0.005789f
C1148 x4.net9 a_26191_n8709# 5.55e-19
C1149 x3.x1.nSEL0 a_17405_n2032# 0.081627f
C1150 x3.x1.nSEL1 x3.nselect2 0.047548f
C1151 a_23597_n8715# a_23063_n8709# 0.002698f
C1152 a_28743_n9483# x4._24_ 0.002926f
C1153 x4.clknet_0_clk a_27837_n7261# 5.18e-20
C1154 a_26630_n8715# x4._17_ 9.6e-21
C1155 a_24595_n8741# x4.net6 0.080758f
C1156 x4._11_ a_27807_n9829# 0.19543f
C1157 x4.net9 x4._24_ 0.165357f
C1158 x4._01_ a_23615_n5995# 3.94e-19
C1159 a_23811_n5073# x4._10_ 6.67e-19
C1160 a_23670_n8741# a_23927_n8715# 0.036838f
C1161 a_23781_n8171# a_25834_n7921# 1.23e-20
C1162 a_23670_n8741# a_23693_n9259# 6.87e-19
C1163 a_24595_n8741# a_24203_n8893# 0.006202f
C1164 x4.net9 a_27591_n8991# 0.115737f
C1165 x4._08_ a_28197_n8709# 0.415957f
C1166 a_23778_n8893# a_23904_n9259# 0.005525f
C1167 x4._17_ a_26593_n7906# 2.72e-19
C1168 a_23946_n9147# x4.net5 0.001073f
C1169 a_25639_n9259# a_26147_n9107# 0.017774f
C1170 x4._11_ a_24769_n9465# 8.14e-19
C1171 VDD a_27093_n8893# 0.003234f
C1172 a_25709_n7109# x4.net9 1.97e-19
C1173 a_26159_n7409# a_26713_n7249# 0.057611f
C1174 VDD a_18033_n1958# 0.192568f
C1175 x4.counter[6] a_27591_n8991# 4.54e-21
C1176 a_25875_n7395# a_26117_n7627# 0.008508f
C1177 m2_17442_n2443# x3.x2.GN1 0.06935f
C1178 a_28003_n9437# a_27807_n9829# 0.00119f
C1179 x4._04_ x4.net5 0.003846f
C1180 a_24054_n7805# x4._16_ 1.81e-20
C1181 a_25823_n8395# x4._11_ 5.64e-19
C1182 a_27166_n9147# x4.net6 6.78e-21
C1183 a_26375_n8171# x4.net6 0.00514f
C1184 VDD a_26979_n9829# 0.405792f
C1185 a_23682_n5329# a_24229_n5073# 0.099725f
C1186 a_23882_n5174# a_24031_n5085# 0.005525f
C1187 a_22962_n5131# x4._12_ 0.001776f
C1188 drv_out mux_out 4.52048f
C1189 a_24647_n7903# x4.net8 5.45e-19
C1190 x1.sky130_fd_sc_hd__inv_2_15.A select0 5.64e-20
C1191 x4.clknet_0_clk a_25875_n7395# 0.00222f
C1192 drv_out x4._05_ 0.0016f
C1193 a_25639_n9259# a_26559_n9259# 2.37e-21
C1194 x4._16_ x4._20_ 0.011071f
C1195 x4._14_ a_23778_n8893# 9.43e-20
C1196 a_27223_n8741# x4.net7 0.08513f
C1197 x4._12_ a_23391_n4933# 1.23e-19
C1198 a_24229_n5073# x4._00_ 0.001531f
C1199 x4.net10 counter7 5.8e-20
C1200 a_29319_n10347# x4._23_ 9.55e-20
C1201 x4._11_ x4._16_ 0.223435f
C1202 x4._05_ x4._15_ 9.02e-20
C1203 a_23682_n5329# x4.net1 0.00338f
C1204 a_27377_n9437# x4._15_ 5.62e-21
C1205 a_22885_n8715# counter3 1.26e-20
C1206 a_23994_n9687# a_23778_n8893# 0.003601f
C1207 a_18033_n1958# select1 0.254026f
C1208 VDD a_25729_n8395# 5.6e-19
C1209 x4.net1 x4._00_ 0.056053f
C1210 x4.net9 a_28979_n8893# 1.5e-19
C1211 a_25779_n7395# a_25875_n7395# 0.310858f
C1212 a_25359_n7627# a_26159_n7409# 2.3e-20
C1213 a_24125_n10182# a_23339_n9259# 8.97e-21
C1214 x4._04_ a_24595_n9571# 1.25e-20
C1215 x4.clknet_1_0__leaf_clk x4._01_ 0.05158f
C1216 a_23682_n4633# a_24229_n5073# 4.5e-20
C1217 a_27194_n8171# a_28031_n9259# 6.92e-20
C1218 a_23417_n8715# x4.net6 1.35e-20
C1219 x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_14.A 0.025028f
C1220 a_26529_n7849# a_26166_n7505# 6.47e-19
C1221 x4._19_ x4.net6 0.04173f
C1222 a_27055_n8715# a_26191_n8709# 0.030894f
C1223 a_27223_n8741# a_26357_n8709# 0.034054f
C1224 a_23417_n8715# a_23229_n8709# 0.097818f
C1225 a_26630_n8715# a_26798_n8741# 0.239923f
C1226 a_26295_n7249# x4._15_ 2.35e-21
C1227 a_23682_n4633# x4.net1 0.006588f
C1228 a_23675_n4933# a_23941_n3056# 6.9e-23
C1229 x4._02_ x4.net6 0.001309f
C1230 a_26725_n9259# x4.clknet_1_1__leaf_clk 0.486375f
C1231 a_26542_n7627# x4.clknet_0_clk 4.01e-19
C1232 a_25900_n8197# x4._21_ 0.114705f
C1233 a_25834_n7921# a_25762_n7921# 0.005941f
C1234 a_23969_n8171# a_24149_n7805# 0.001229f
C1235 VDD x4.net8 1.78891f
C1236 a_28596_n8337# x4._15_ 4.15e-19
C1237 x4.net2 a_23063_n8709# 3.28e-19
C1238 x4._21_ x4._15_ 0.054317f
C1239 a_23063_n8709# a_23670_n8741# 0.141453f
C1240 x4._02_ a_23229_n8709# 0.275992f
C1241 x4._22_ a_26191_n8709# 0.016414f
C1242 a_26593_n7906# a_26798_n8741# 1.06e-19
C1243 x3.x2.GN4 x3.x2.GP2 8.45e-19
C1244 x4.net7 a_25449_n7261# 5.91e-19
C1245 x4.net3 a_23391_n5219# 0.006429f
C1246 x4.net9 x4._20_ 1.35e-20
C1247 a_23781_n8171# x4.net6 0.004467f
C1248 x4._03_ a_23693_n9259# 0.13856f
C1249 a_28031_n9259# a_28579_n7627# 3.35e-21
C1250 a_23339_n9259# a_23873_n8893# 0.002698f
C1251 a_23811_n4907# x4.clknet_1_0__leaf_clk 0.050329f
C1252 m3_18866_n4909# x3.x2.GP3 9.67e-19
C1253 x4._11_ counter3 1.13e-19
C1254 x4.net3 a_22837_n10182# 0.006292f
C1255 a_25823_n8395# x4._17_ 3.09e-20
C1256 VDD x4._07_ 0.322336f
C1257 x4._11_ x4.net9 0.233741f
C1258 VDD x3.x1.nSEL0 0.5228f
C1259 a_23781_n8171# a_23229_n8709# 5.5e-20
C1260 a_27223_n8741# a_27423_n8893# 4.17e-19
C1261 a_26630_n8715# a_26913_n9259# 0.001307f
C1262 x4.net4 x4._18_ 3.06e-19
C1263 x4._01_ a_24525_n5745# 0.012244f
C1264 a_24222_n8059# a_24371_n8991# 8.5e-21
C1265 a_24054_n7805# a_23778_n8893# 9.19e-21
C1266 a_23781_n8171# a_24203_n8893# 0.001133f
C1267 x4.counter[6] x4._11_ 0.002692f
C1268 x4._22_ x4._24_ 0.01067f
C1269 x4.net8 a_27139_n8715# 9.28e-20
C1270 x4.clknet_1_0__leaf_clk x4.net5 6.12e-20
C1271 a_23391_n5219# x4._12_ 0.036321f
C1272 a_23615_n8171# a_24479_n7805# 0.030894f
C1273 x4._04_ a_24647_n7903# 0.003723f
C1274 x4._08_ a_27194_n8171# 0.011527f
C1275 a_27807_n9829# x4._23_ 0.130093f
C1276 x4._22_ a_27591_n8991# 3.11e-19
C1277 x3.x2.GN3 a_19235_n1926# 1.07e-20
C1278 a_24371_n8991# a_24329_n9259# 7.84e-20
C1279 a_18537_n1898# x3.x2.GN4 3.22e-19
C1280 x4._17_ x4._16_ 0.048058f
C1281 x3.x1.nSEL1 x3.x2.GN2 0.209956f
C1282 a_25709_n7109# x4._22_ 7.51e-19
C1283 a_28895_n8715# x4.clknet_1_1__leaf_clk 1.84e-19
C1284 a_27805_n10182# a_27807_n9829# 0.01226f
C1285 a_23675_n5233# a_23391_n4933# 9.64e-20
C1286 a_28638_n9147# a_29021_n9259# 4.67e-20
C1287 x4._12_ a_23255_n4363# 1.27e-21
C1288 x4._11_ a_23778_n8893# 0.00274f
C1289 a_28385_n9259# x4.clknet_1_1__leaf_clk 6.27e-19
C1290 enable_counter a_23675_n4933# 1.25e-19
C1291 x4.clknet_1_1__leaf_clk a_27251_n7408# 0.035969f
C1292 m3_18876_n6983# counter3 8.01e-20
C1293 a_29133_n9803# x4._09_ 0.07143f
C1294 x4._04_ a_24605_n8171# 6.79e-19
C1295 a_23615_n8171# a_25667_n8171# 9.88e-21
C1296 x4.net4 a_23904_n9259# 6.57e-19
C1297 x4._00_ a_23295_n4755# 0.001095f
C1298 drv_out a_27755_n7261# 1.34e-19
C1299 x3.x1.nSEL0 select1 0.137394f
C1300 drv_out x4.net7 6.87e-19
C1301 x1.sky130_fd_sc_hd__inv_2_16.A select0 9.57e-20
C1302 a_28638_n8741# a_28895_n8715# 0.036838f
C1303 a_28999_n7408# x4._25_ 0.227897f
C1304 a_26545_n8715# x4.net7 0.014734f
C1305 a_25900_n8197# x4.net7 0.003377f
C1306 x4._08_ a_28579_n7627# 0.001905f
C1307 a_28669_n7261# x4._25_ 8.17e-20
C1308 a_29063_n8741# a_29063_n8991# 0.026048f
C1309 x4._15_ a_27755_n7261# 0.142876f
C1310 x4.net7 x4._15_ 0.590844f
C1311 a_29319_n10347# x4.net11 0.250513f
C1312 a_25834_n7921# x4._18_ 5.77e-19
C1313 a_28470_n8893# a_28385_n9259# 0.037333f
C1314 a_29063_n8991# a_28895_n8893# 0.310858f
C1315 x4._10_ x4._11_ 0.033565f
C1316 a_23675_n4933# a_23505_n4363# 5.23e-20
C1317 VDD a_23946_n9147# 0.219675f
C1318 a_23682_n4633# a_23295_n4755# 0.034054f
C1319 VDD x4.net10 1.28398f
C1320 a_26366_n7350# x4.net6 6.81e-19
C1321 x4.net4 x4._14_ 0.209869f
C1322 a_23417_n8715# a_23339_n9259# 2.5e-19
C1323 x4._16_ x4._23_ 3.32e-22
C1324 VDD x4._04_ 0.27578f
C1325 a_28385_n8715# x4.net6 3.93e-20
C1326 a_25762_n7921# x4.net6 0.002624f
C1327 a_29103_n9829# x4._24_ 0.003347f
C1328 a_25875_n7395# a_26147_n9107# 5.98e-21
C1329 x4.clknet_0_clk a_26725_n9259# 3.43e-21
C1330 x4.clknet_1_0__leaf_clk a_24053_n8337# 4.11e-19
C1331 x1.sky130_fd_sc_hd__inv_2_5.A x1.sky130_fd_sc_hd__inv_2_15.A 0.001676f
C1332 x4.net8 a_28725_n10182# 7.5e-19
C1333 x4.net4 a_23994_n9687# 0.007901f
C1334 x4._02_ a_23339_n9259# 3.71e-19
C1335 x4._17_ x4.net9 7.02e-19
C1336 a_23063_n8709# x4._03_ 0.001727f
C1337 a_26545_n8715# a_26357_n8709# 0.095025f
C1338 a_25834_n7921# a_26191_n8709# 4.26e-19
C1339 a_25729_n8715# a_25639_n9259# 8.68e-19
C1340 x4._21_ a_24371_n8991# 1.79e-21
C1341 a_26357_n8709# x4._15_ 0.027322f
C1342 counter7 a_28457_n9803# 1.91e-19
C1343 x4._13_ x4._02_ 0.053355f
C1344 VDD a_23615_n5995# 0.266078f
C1345 x4.net5 x4._15_ 0.016962f
C1346 a_27507_n8893# a_26725_n9259# 3.14e-19
C1347 a_23781_n8171# a_23339_n9259# 1.21e-19
C1348 a_23615_n8171# a_23505_n9259# 3.23e-21
C1349 a_27055_n8715# x4._11_ 7.12e-21
C1350 x4._16_ a_26798_n8741# 0.001117f
C1351 a_23851_n9829# a_24220_n9483# 0.046138f
C1352 a_23295_n5219# a_23682_n5329# 0.034054f
C1353 a_23391_n5219# a_23675_n5233# 0.030894f
C1354 a_24647_n7903# x4.clknet_1_0__leaf_clk 1.77e-20
C1355 x4._13_ a_23781_n8171# 7.99e-20
C1356 x4._19_ a_26713_n7249# 0.014678f
C1357 x4._22_ x4._20_ 2.69e-20
C1358 drv_out counter7 2.39e-19
C1359 a_27194_n8171# a_27166_n9147# 2.72e-20
C1360 a_26529_n7849# a_26998_n8893# 5.18e-21
C1361 x4._11_ x4._22_ 0.420712f
C1362 a_26529_n7849# a_26816_n8171# 3.14e-19
C1363 a_25834_n7921# a_25709_n7109# 1.01e-19
C1364 VDD x1.sky130_fd_sc_hd__inv_2_11.A 0.639695f
C1365 a_28743_n9483# x4._23_ 2.44e-19
C1366 x4._09_ x4.clknet_1_1__leaf_clk 0.003413f
C1367 a_27423_n8893# x4._15_ 1.98e-20
C1368 a_22837_n10182# a_23205_n10182# 2.48e-19
C1369 a_26166_n7505# x4.clknet_1_1__leaf_clk 0.013843f
C1370 counter7 x4._15_ 0.003538f
C1371 a_23255_n4363# a_23505_n4043# 0.007234f
C1372 VDD a_23610_n5085# 3.44e-19
C1373 x4.net9 x4._23_ 0.065132f
C1374 x4.clknet_0_clk a_27251_n7408# 0.012442f
C1375 VDD a_27223_n8741# 0.406789f
C1376 x4.net9 a_27805_n10182# 7.77e-19
C1377 x4._16_ a_26913_n9259# 1.98e-21
C1378 VDD a_29645_n10182# 0.276039f
C1379 x4.net11 a_27807_n9829# 1.29e-21
C1380 x4._22_ a_28003_n9437# 0.001961f
C1381 x4.net4 a_24054_n7805# 0.034877f
C1382 a_24595_n9571# x4._15_ 1.84e-19
C1383 x4.counter[6] a_27805_n10182# 0.1107f
C1384 a_28470_n8715# a_28031_n9259# 1.73e-19
C1385 a_23882_n5174# x4.net2 3.35e-21
C1386 x4._09_ a_28470_n8893# 0.0221f
C1387 a_28031_n9259# a_29063_n8991# 0.048748f
C1388 a_25965_n10182# x4.net6 0.195979f
C1389 VDD a_26457_n7849# 0.001301f
C1390 m3_18866_n4909# x3.x2.GN2 0.099332f
C1391 a_23781_n8171# a_23225_n7109# 1.63e-19
C1392 x4._16_ a_25211_n9465# 0.039613f
C1393 x4._18_ x4.net6 0.081404f
C1394 a_25359_n7627# x4._19_ 0.082191f
C1395 select0 x3.x2.GP2 5.28e-19
C1396 x4.net4 x4._11_ 0.952686f
C1397 a_28197_n8709# a_28385_n8715# 0.097994f
C1398 x1.sky130_fd_sc_hd__inv_2_11.A select1 9.08e-20
C1399 x4.net10 a_28725_n10182# 2.65e-20
C1400 x4._07_ a_27093_n8893# 2.91e-19
C1401 x4.net8 a_26979_n9829# 0.1454f
C1402 VDD x4.clknet_1_0__leaf_clk 3.74806f
C1403 x1.sky130_fd_sc_hd__inv_2_17.A select0 9.57e-20
C1404 x4.net9 a_26798_n8741# 2.05e-20
C1405 a_27194_n8171# x4._19_ 6.04e-19
C1406 x3.x1.nSEL0 a_18033_n1958# 0.001174f
C1407 a_24625_n8715# a_23063_n8709# 2.77e-19
C1408 x4._11_ a_23697_n5995# 1.17e-19
C1409 a_23969_n8171# a_23063_n8709# 3.23e-19
C1410 a_24813_n8395# x4._16_ 3.98e-19
C1411 x4.net3 a_24316_n9803# 1.66e-19
C1412 a_27055_n8715# x4._17_ 8.73e-21
C1413 x4._07_ a_26979_n9829# 9.24e-19
C1414 a_26191_n8709# x4.net6 0.0618f
C1415 a_23675_n4933# x4.net2 4.59e-19
C1416 x3.x2.GN1 mux_out 0.430121f
C1417 x4._11_ a_29103_n9829# 2.01e-20
C1418 VDD a_25449_n7261# 0.002157f
C1419 a_25793_n9259# x4._20_ 0.001506f
C1420 select0 a_18537_n1898# 0.001558f
C1421 a_24095_n8741# a_23927_n8715# 0.310858f
C1422 a_24647_n7903# a_25900_n8197# 2.22e-20
C1423 x4._11_ a_25793_n9259# 0.001879f
C1424 x3.x2.GP1 x3.x2.GP2 0.043302f
C1425 x4.net9 a_26913_n9259# 1.61e-19
C1426 x4._08_ a_28470_n8715# 0.030723f
C1427 x4._17_ x4._22_ 1.76e-19
C1428 a_24371_n8991# x4.net5 0.13266f
C1429 a_23421_n7921# x4.clknet_1_0__leaf_clk 0.001585f
C1430 x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_15.A 0.025028f
C1431 x4.net6 x4._24_ 0.002355f
C1432 a_26366_n7350# a_26713_n7249# 0.037333f
C1433 VDD a_18585_n1958# 0.26222f
C1434 a_26295_n7249# a_26515_n7261# 4.62e-19
C1435 a_26166_n7505# a_26117_n7627# 4.04e-19
C1436 a_25834_n7921# x4._20_ 4.3e-20
C1437 a_28205_n9437# a_27807_n9829# 0.005781f
C1438 VDD a_24525_n5745# 0.006514f
C1439 a_27591_n8991# x4.net6 3.96e-21
C1440 a_24479_n7805# x4._16_ 0.003542f
C1441 a_25834_n7921# x4._11_ 0.043142f
C1442 a_25709_n7109# x4.net6 8.49e-19
C1443 VDD a_28457_n9803# 0.152186f
C1444 a_23811_n5073# a_24229_n5073# 3.39e-19
C1445 x4.clknet_0_clk a_26166_n7505# 0.025079f
C1446 x4._14_ a_23229_n8709# 4.89e-20
C1447 a_26147_n9107# a_26725_n9259# 0.00145f
C1448 x3.x2.GN4 a_19235_n1926# 0.001562f
C1449 x4._14_ a_24203_n8893# 0.002114f
C1450 VDD a_25721_n9259# 2.86e-19
C1451 x3.x1.nSEL1 x3.x2.GN3 0.012418f
C1452 a_26529_n7849# x4._05_ 3.16e-19
C1453 x4._16_ a_25667_n8171# 0.061172f
C1454 a_28031_n8709# x4.net7 8.61e-20
C1455 a_28197_n9259# x4.net7 0.001362f
C1456 a_23811_n5073# x4.net1 0.001727f
C1457 VDD x1.sky130_fd_sc_hd__inv_2_12.A 0.637448f
C1458 x4.net8 x4._07_ 0.001136f
C1459 a_28099_n9437# x4._15_ 0.00403f
C1460 VDD drv_out 16.4224f
C1461 x4.net4 x4._17_ 9.08e-20
C1462 a_25600_n8741# x4.clknet_1_1__leaf_clk 0.048773f
C1463 a_24595_n9571# a_24371_n8991# 0.001036f
C1464 a_18585_n1958# select1 0.127717f
C1465 VDD a_26545_n8715# 0.084103f
C1466 x4._22_ x4._23_ 0.511385f
C1467 VDD a_25900_n8197# 0.084816f
C1468 a_26630_n8715# a_26593_n7906# 1.41e-19
C1469 x4.net9 x4.net11 0.055197f
C1470 a_25875_n7395# a_26159_n7409# 0.030894f
C1471 a_25779_n7395# a_26166_n7505# 0.034054f
C1472 a_26559_n9259# a_26725_n9259# 0.966391f
C1473 x4._22_ a_27805_n10182# 2.78e-19
C1474 VDD x4._15_ 1.72333f
C1475 a_25729_n8715# a_25875_n7395# 4.21e-21
C1476 a_26529_n7849# a_26295_n7249# 1.61e-19
C1477 x4.clknet_1_1__leaf_clk a_28399_n7627# 7.87e-19
C1478 a_28197_n8709# a_26191_n8709# 3.42e-21
C1479 a_23628_n8337# a_23670_n8741# 4.62e-19
C1480 a_27055_n8715# a_26798_n8741# 0.036838f
C1481 a_23417_n8715# a_23502_n8715# 0.037333f
C1482 a_28031_n8709# a_26357_n8709# 1.33e-19
C1483 a_23882_n4933# x4.net1 0.002893f
C1484 a_26998_n8893# x4.clknet_1_1__leaf_clk 0.042872f
C1485 a_27194_n8171# a_28385_n8715# 9.53e-19
C1486 a_26529_n7849# x4._21_ 0.001146f
C1487 x1.sky130_fd_sc_hd__inv_2_12.A select1 0.001652f
C1488 x4.counter[5] x4.counter[6] 0.070133f
C1489 a_23063_n8709# a_24095_n8741# 0.048748f
C1490 x4._02_ a_23502_n8715# 8.22e-19
C1491 x1.sky130_fd_sc_hd__inv_2_17.Y select0 9.57e-20
C1492 drv_out select1 1.17e-19
C1493 x4._22_ a_26798_n8741# 0.01767f
C1494 a_28197_n8709# x4._24_ 0.035946f
C1495 x4._11_ a_28551_n9803# 0.039972f
C1496 x4.net3 a_23682_n5329# 0.005586f
C1497 x4.net7 a_26515_n7261# 0.002551f
C1498 a_24054_n7805# x4.net6 3.12e-19
C1499 a_28638_n9147# x4._24_ 0.014122f
C1500 x4._16_ a_23505_n9259# 2.51e-21
C1501 m3_18876_n6983# x3.x2.GP3 0.006132f
C1502 x4.net3 a_24125_n10182# 0.001252f
C1503 a_25834_n7921# x4._17_ 0.076419f
C1504 x4._18_ a_26713_n7249# 2.19e-20
C1505 a_23781_n8171# a_23502_n8715# 0.001124f
C1506 a_26542_n7627# a_26159_n7409# 0.001632f
C1507 a_23811_n5073# a_23225_n7109# 1.29e-20
C1508 a_28197_n9259# a_27423_n8893# 2.56e-19
C1509 a_28385_n9259# a_26559_n9259# 4.76e-21
C1510 a_24054_n7805# a_24203_n8893# 1.06e-19
C1511 a_23615_n8171# x4._16_ 6.86e-20
C1512 x4._20_ x4.net6 0.00624f
C1513 x4.net8 x4.net10 1.02e-19
C1514 counter7 a_28197_n9259# 5.88e-20
C1515 x4._11_ x4.net6 2.01574f
C1516 x4._04_ x4.net8 7.52e-21
C1517 a_23682_n5329# x4._12_ 0.206007f
C1518 x4._22_ a_26913_n9259# 0.012798f
C1519 a_29103_n9829# x4._23_ 0.220841f
C1520 x4.clknet_0_clk a_25179_n7627# 2.32e-20
C1521 x4.net2 a_24075_n5995# 3.45e-20
C1522 a_17405_n2032# a_17579_n1926# 0.006584f
C1523 x4._11_ a_23229_n8709# 0.008371f
C1524 VDD a_29321_n9483# 0.003335f
C1525 x4._14_ a_23339_n9259# 0.008544f
C1526 x1.sky130_fd_sc_hd__inv_2_4.A x1.sky130_fd_sc_hd__inv_2_16.A 0.001676f
C1527 a_28725_n10182# a_28457_n9803# 1.23e-19
C1528 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_13.A 3.14e-21
C1529 a_29063_n8991# a_29021_n9259# 7.84e-20
C1530 x4._12_ x4._00_ 4.17e-19
C1531 x4._11_ a_24203_n8893# 0.045224f
C1532 enable_counter a_23811_n4907# 2.79e-20
C1533 a_26309_n9259# x4.net7 1.98e-19
C1534 x4._13_ x4._14_ 0.074354f
C1535 a_23851_n9829# x4._03_ 0.112166f
C1536 a_23994_n9687# a_23339_n9259# 0.00127f
C1537 x4._18_ a_25359_n7627# 0.190808f
C1538 a_29063_n8741# a_28895_n8715# 0.310858f
C1539 x4.clknet_0_clk a_25600_n8741# 8.98e-21
C1540 a_26529_n7849# x4.net7 6.37e-20
C1541 x4._08_ x4._25_ 0.208467f
C1542 x4.net10 a_28647_n9483# 8.38e-19
C1543 a_23682_n4633# x4._12_ 0.003541f
C1544 a_28895_n8715# a_28895_n8893# 0.01464f
C1545 x1.sky130_fd_sc_hd__inv_2_14.A a_17405_n2032# 6.58e-22
C1546 a_28638_n9147# a_28979_n8893# 9.73e-19
C1547 a_28725_n10182# x4._15_ 0.006207f
C1548 a_24125_n10182# x4.counter[2] 0.1107f
C1549 m3_18866_n4909# x3.x2.GN3 0.001446f
C1550 VDD x1.sky130_fd_sc_hd__inv_2_13.A 0.637284f
C1551 a_25709_n7109# a_26713_n7249# 8.9e-19
C1552 a_24220_n9483# x4.net5 0.075434f
C1553 a_23675_n4933# a_23391_n4933# 0.032244f
C1554 VDD a_24371_n8991# 0.391294f
C1555 x4.clknet_0_clk a_28399_n7627# 2.96e-20
C1556 x4._14_ x4.counter[1] 1.03e-21
C1557 a_26630_n8715# x4._16_ 0.00213f
C1558 x4._22_ x4.net11 1.96e-19
C1559 a_25779_n7395# a_25600_n8741# 8.51e-20
C1560 a_17405_n2032# x3.x2.GN1 0.12869f
C1561 a_26725_n8715# x4.net6 0.001259f
C1562 x4.clknet_0_clk a_26998_n8893# 4.63e-19
C1563 a_26166_n7505# a_26147_n9107# 2.42e-19
C1564 x4.net8 a_27223_n8741# 0.084103f
C1565 x4.net4 a_25211_n9465# 0.083888f
C1566 a_24981_n8715# a_24595_n8741# 0.006406f
C1567 a_26756_n8337# a_26798_n8741# 4.62e-19
C1568 a_26529_n7849# a_26357_n8709# 1.08e-19
C1569 a_27925_n7261# a_27755_n7261# 0.001675f
C1570 a_26593_n7906# x4._16_ 0.060109f
C1571 a_27925_n7261# x4.net7 0.00717f
C1572 a_23505_n9259# a_23778_n8893# 0.081834f
C1573 x4._05_ x4.clknet_1_1__leaf_clk 0.143201f
C1574 a_24229_n5073# x4._11_ 0.001319f
C1575 a_27223_n8741# x4._07_ 0.008579f
C1576 a_28031_n9259# a_26725_n9259# 3.23e-19
C1577 a_23615_n8171# a_23778_n8893# 8.98e-19
C1578 a_28197_n8709# x4._11_ 2.03e-20
C1579 x4._17_ x4.net6 0.277113f
C1580 a_27124_n9259# a_27166_n9147# 4.62e-19
C1581 a_24054_n7805# a_23339_n9259# 5.5e-20
C1582 select0 a_19235_n1926# 1.4e-19
C1583 a_26159_n7409# a_26725_n9259# 4.79e-20
C1584 x1.sky130_fd_sc_hd__inv_2_13.A select1 1.79e-19
C1585 a_27194_n8171# x4._24_ 0.025563f
C1586 x4._11_ a_28638_n9147# 8.51e-19
C1587 a_24595_n9571# a_24220_n9483# 4e-20
C1588 x4.net4 a_24813_n8395# 5.3e-19
C1589 a_23675_n5233# a_23682_n5329# 0.969092f
C1590 x4.net3 a_23417_n8715# 0.003111f
C1591 a_23295_n5219# a_23811_n5073# 1.28e-19
C1592 x4._13_ a_24054_n7805# 5.02e-20
C1593 x1.sky130_fd_sc_hd__inv_2_12.A a_18033_n1958# 2.34e-20
C1594 x4.net1 x4._11_ 0.002334f
C1595 a_23339_n9259# x4._20_ 1.9e-21
C1596 x4._03_ a_24329_n9259# 9.96e-20
C1597 a_27194_n8171# a_27591_n8991# 0.001883f
C1598 a_23675_n5233# x4._00_ 8.76e-20
C1599 x4._11_ a_23339_n9259# 0.005486f
C1600 a_28551_n9803# x4._23_ 0.038842f
C1601 x4.net3 x4._02_ 0.031079f
C1602 a_26295_n7249# x4.clknet_1_1__leaf_clk 1.17e-20
C1603 a_23205_n10182# a_24125_n10182# 1.37e-20
C1604 a_23505_n4043# x4._00_ 0.002065f
C1605 VDD a_24031_n5085# 0.002269f
C1606 x4._13_ x4._11_ 0.217373f
C1607 a_26630_n8715# x4.net9 6.38e-21
C1608 VDD a_28031_n8709# 0.714632f
C1609 x4.net9 a_29319_n10347# 0.003439f
C1610 VDD a_28197_n9259# 0.31984f
C1611 x4.net4 a_24479_n7805# 0.002624f
C1612 x4.net11 a_29103_n9829# 0.088145f
C1613 x4._22_ a_28205_n9437# 2.76e-20
C1614 x4._24_ a_28579_n7627# 0.197975f
C1615 x4._21_ x4.clknet_1_1__leaf_clk 0.038033f
C1616 a_26166_n7505# x4._06_ 1.63e-21
C1617 a_26979_n9829# x4._15_ 1.2e-20
C1618 a_23682_n4633# a_23675_n5233# 3.36e-19
C1619 a_28895_n8715# a_28031_n9259# 1.29e-19
C1620 a_29063_n8741# x4._09_ 5.87e-19
C1621 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_14.A 7.08e-21
C1622 a_23675_n4933# a_23391_n5219# 9.64e-20
C1623 x4.net6 x4._23_ 0.023006f
C1624 x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_16.A 0.025028f
C1625 VDD a_23941_n3056# 0.305606f
C1626 x4._01_ x4.net2 9.85e-20
C1627 x4.net9 a_26593_n7906# 0.122363f
C1628 a_28031_n9259# a_28385_n9259# 0.062224f
C1629 x4._09_ a_28895_n8893# 0.024482f
C1630 VDD a_17579_n1926# 9.25e-19
C1631 a_23675_n4933# a_23255_n4363# 0.001828f
C1632 VDD a_28979_n8715# 0.00533f
C1633 a_25875_n7395# x4._19_ 0.046625f
C1634 a_26159_n7409# a_27251_n7408# 5.23e-20
C1635 x4._11_ a_26713_n7249# 7.39e-21
C1636 a_28470_n8715# a_28385_n8715# 0.037333f
C1637 a_28638_n8741# a_28596_n8337# 4.62e-19
C1638 x4.net8 a_28457_n9803# 4.33e-20
C1639 x4.net10 a_29645_n10182# 0.219068f
C1640 a_25729_n8395# x4._15_ 0.005043f
C1641 x3.x1.nSEL0 a_18585_n1958# 1.21e-20
C1642 x4._11_ a_23225_n7109# 0.055744f
C1643 x4.net8 a_25721_n9259# 4.38e-20
C1644 VDD x1.sky130_fd_sc_hd__inv_2_14.A 0.637855f
C1645 a_25823_n8395# x4._16_ 3.31e-19
C1646 a_26798_n8741# x4.net6 0.012704f
C1647 a_23811_n4907# x4.net2 3.46e-19
C1648 VDD a_26515_n7261# 0.002269f
C1649 x4.clknet_1_0__leaf_clk a_23946_n9147# 0.001507f
C1650 a_24095_n8741# a_25600_n8741# 1e-20
C1651 x4.net8 a_26545_n8715# 0.005878f
C1652 x4.clknet_0_clk x4._05_ 0.067252f
C1653 x4.net8 a_25900_n8197# 0.028641f
C1654 a_24222_n8059# a_23969_n8171# 3.39e-19
C1655 x4.net2 x4.net5 7.09e-21
C1656 x4._11_ a_26381_n9259# 0.001398f
C1657 x4.counter[9] x4._23_ 7.62e-19
C1658 VDD enable_counter 0.254269f
C1659 x4.net8 x4._15_ 0.048599f
C1660 x4._08_ a_28895_n8715# 0.013878f
C1661 a_25211_n9231# x4.net5 4.5e-19
C1662 x4._11_ a_25359_n7627# 0.001495f
C1663 a_23693_n9259# a_23873_n8893# 0.001229f
C1664 x4.counter[9] a_27805_n10182# 2.37e-20
C1665 x4._04_ x4.clknet_1_0__leaf_clk 0.005301f
C1666 x4._19_ x4._25_ 9.05e-21
C1667 a_26295_n7249# a_26117_n7627# 9.73e-19
C1668 VDD x3.x2.GN1 1.47002f
C1669 x4.clknet_1_1__leaf_clk a_27755_n7261# 0.001522f
C1670 a_28647_n9483# a_28457_n9803# 0.011458f
C1671 x4.clknet_1_1__leaf_clk x4.net7 0.397702f
C1672 VDD a_23769_n5995# 3.14e-19
C1673 a_25834_n7921# a_25667_n8171# 0.046138f
C1674 a_26885_n10182# x4.clknet_1_1__leaf_clk 4.13e-21
C1675 a_24011_n8715# x4._11_ 7.61e-19
C1676 a_26913_n9259# x4.net6 0.00565f
C1677 a_27194_n8171# x4._11_ 0.049204f
C1678 mux_out x3.x2.GP2 0.349381f
C1679 x4.net9 a_27807_n9829# 9.8e-19
C1680 x4._07_ x4._15_ 0.022092f
C1681 a_25779_n7395# x4._05_ 1.85e-19
C1682 x4._21_ a_26117_n7627# 1.26e-19
C1683 x4.net4 a_23505_n9259# 0.019846f
C1684 VDD a_24220_n9483# 0.007674f
C1685 x4._01_ a_23633_n5451# 2.39e-19
C1686 x4.clknet_1_0__leaf_clk a_23615_n5995# 0.024338f
C1687 x1.sky130_fd_sc_hd__inv_2_14.A select1 1.03e-20
C1688 x4.net2 counter7 6.88e-20
C1689 x4.clknet_0_clk a_26295_n7249# 0.003343f
C1690 a_28197_n8709# x4._23_ 0.031087f
C1691 x4.net4 a_23615_n8171# 0.071607f
C1692 VDD a_26309_n9259# 4.84e-19
C1693 VDD a_23505_n4363# 0.262851f
C1694 a_25211_n9465# x4.net6 1.4e-20
C1695 a_28638_n9147# x4._23_ 0.005759f
C1696 a_28470_n8893# x4.net7 4.39e-19
C1697 m3_18862_n5953# x3.x2.GP2 0.005314f
C1698 x4._21_ x4.clknet_0_clk 4.86e-19
C1699 x4._17_ a_26713_n7249# 0.016586f
C1700 a_28647_n9483# x4._15_ 0.004129f
C1701 a_28031_n9259# x4._09_ 0.098799f
C1702 a_24095_n8741# a_23851_n9829# 2.52e-20
C1703 a_26357_n8709# x4.clknet_1_1__leaf_clk 0.079788f
C1704 x4.net10 a_28457_n9803# 0.27342f
C1705 x3.x2.GN1 select1 0.312198f
C1706 VDD a_23597_n8715# 0.003619f
C1707 a_26630_n8715# x4._22_ 0.006172f
C1708 VDD a_26529_n7849# 0.2552f
C1709 a_25779_n7395# a_26295_n7249# 1.28e-19
C1710 a_26159_n7409# a_26166_n7505# 0.961627f
C1711 a_28031_n7261# x4._11_ 0.005861f
C1712 a_26559_n9259# a_26998_n8893# 0.273138f
C1713 a_26725_n9259# a_27166_n9147# 0.110715f
C1714 x4.clknet_1_0__leaf_clk a_23610_n5085# 0.001172f
C1715 a_24813_n8395# x4.net6 0.001315f
C1716 x4._06_ a_25600_n8741# 0.002127f
C1717 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_15.A 1.11e-20
C1718 counter3 x4._16_ 1.05e-19
C1719 x1.sky130_fd_sc_hd__inv_2_3.A x1.sky130_fd_sc_hd__inv_2_17.A 0.001676f
C1720 x4._21_ a_25779_n7395# 0.001295f
C1721 x4.net9 x4._16_ 0.243936f
C1722 a_26593_n7906# x4._22_ 0.155189f
C1723 a_24053_n8337# a_23670_n8741# 4.67e-20
C1724 m3_18866_n4909# x3.x2.GN4 7.17e-19
C1725 a_23633_n4541# x4.net1 8.57e-19
C1726 a_27423_n8893# x4.clknet_1_1__leaf_clk 0.044904f
C1727 x4.net10 x4._15_ 0.289356f
C1728 x4._02_ a_23927_n8715# 3.18e-19
C1729 a_23063_n8709# a_24595_n8741# 1.05e-19
C1730 x4._04_ a_25900_n8197# 8.65e-21
C1731 a_23615_n8171# a_25834_n7921# 1.89e-21
C1732 x4._17_ a_25359_n7627# 0.043588f
C1733 VDD a_27925_n7261# 0.002069f
C1734 a_28470_n8715# x4._24_ 0.010979f
C1735 x4.net7 a_26117_n7627# 6.13e-20
C1736 x1.sky130_fd_sc_hd__inv_2_11.A a_18585_n1958# 9.97e-21
C1737 x4.net3 a_23811_n5073# 2.06e-19
C1738 a_24479_n7805# x4.net6 0.021756f
C1739 x4._04_ x4._15_ 3.75e-19
C1740 x4.counter[5] x4.net6 0.080069f
C1741 a_29063_n8991# x4._24_ 0.009415f
C1742 x4._03_ x4.net5 3.86e-19
C1743 x4._06_ a_26816_n8171# 6.53e-20
C1744 x4._16_ a_23778_n8893# 2.79e-19
C1745 x4._08_ x4._09_ 0.013938f
C1746 a_27194_n8171# x4._17_ 0.002308f
C1747 a_24222_n8059# a_24095_n8741# 0.002135f
C1748 a_23781_n8171# a_23927_n8715# 3.42e-19
C1749 VDD x1.sky130_fd_sc_hd__inv_2_15.A 0.637064f
C1750 a_26542_n7627# a_26366_n7350# 0.007724f
C1751 a_24479_n7805# a_24203_n8893# 2.6e-20
C1752 x4.clknet_0_clk a_27755_n7261# 1.5e-19
C1753 x4.clknet_0_clk x4.net7 0.043959f
C1754 a_25667_n8171# x4.net6 4.02e-19
C1755 x3.x1.nSEL1 select0 0.168464f
C1756 a_23811_n5073# x4._12_ 0.039032f
C1757 x4.counter[9] x4.net11 0.066386f
C1758 a_25639_n9259# x4._20_ 0.237238f
C1759 x4._11_ a_23502_n8715# 0.003174f
C1760 a_17857_n2290# x3.x2.GN2 0.106178f
C1761 x1.sky130_fd_sc_hd__inv_2_12.A x1.sky130_fd_sc_hd__inv_2_11.A 0.173286f
C1762 a_29319_n10347# a_29103_n9829# 1.29e-21
C1763 x1.sky130_fd_sc_hd__inv_2_13.A x3.x1.nSEL0 1.14e-19
C1764 VDD a_29133_n9803# 0.283149f
C1765 a_23811_n4907# a_24031_n4907# 4.62e-19
C1766 x4._11_ a_25639_n9259# 0.222369f
C1767 a_27507_n8893# x4.net7 0.002598f
C1768 x4._17_ a_28579_n7627# 8.24e-19
C1769 a_25779_n7395# x4.net7 0.114197f
C1770 x4.counter[6] x4.net9 3.69e-19
C1771 x4._22_ a_27807_n9829# 0.191159f
C1772 a_28031_n7261# x4._17_ 3.01e-19
C1773 a_24595_n9571# x4._03_ 1.19e-19
C1774 drv_out a_27223_n8741# 1.4e-22
C1775 x4._18_ a_25875_n7395# 2.33e-19
C1776 a_25179_n7627# a_26159_n7409# 6.46e-21
C1777 x1.sky130_fd_sc_hd__inv_2_15.A select1 7.73e-20
C1778 a_25729_n8715# x4.counter[4] 4.47e-20
C1779 a_26630_n8715# a_26756_n8337# 0.005525f
C1780 x4.clknet_0_clk a_26357_n8709# 5.94e-19
C1781 a_27194_n8171# x4._23_ 0.042503f
C1782 x3.x1.nSEL1 x3.x2.GP1 1.21e-19
C1783 x4.net10 a_29321_n9483# 0.002502f
C1784 a_23882_n4933# x4._12_ 5.69e-20
C1785 x4._11_ a_25297_n9231# 0.003027f
C1786 a_27223_n8741# x4._15_ 0.031321f
C1787 VDD x4.net2 2.41286f
C1788 a_24981_n8715# x4._18_ 2.06e-20
C1789 VDD a_23670_n8741# 0.200136f
C1790 a_28470_n8893# a_28596_n9259# 0.005525f
C1791 a_28385_n9259# a_28565_n8893# 0.001229f
C1792 a_27251_n7408# x4._19_ 0.214472f
C1793 a_23417_n8715# a_23063_n8709# 0.062224f
C1794 VDD a_17985_n1898# 2.96e-19
C1795 VDD a_25211_n9231# 0.254188f
C1796 m3_18876_n6983# x3.x2.GN3 0.016026f
C1797 a_23811_n4907# a_23391_n4933# 0.036838f
C1798 x4.net3 x4._14_ 0.471315f
C1799 a_25875_n7395# a_26191_n8709# 1.16e-21
C1800 a_18033_n1958# x3.x2.GN1 1.46e-19
C1801 a_23063_n8709# x4._02_ 0.184941f
C1802 x4.net8 a_28031_n8709# 0.001229f
C1803 x4._23_ a_28579_n7627# 0.007723f
C1804 x4.net7 a_28999_n7408# 2.85e-19
C1805 x4.net3 a_23994_n9687# 8.22e-19
C1806 a_23229_n8709# a_23505_n9259# 6.25e-19
C1807 x4.net8 a_28197_n9259# 1.04e-19
C1808 a_25729_n8715# a_25600_n8741# 0.062574f
C1809 a_23615_n8171# x4.net6 0.006287f
C1810 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_16.A 1.99e-20
C1811 x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_17.A 0.025028f
C1812 x4._22_ x4._16_ 0.135659f
C1813 a_28669_n7261# x4.net7 1.83e-19
C1814 a_23946_n9147# a_24371_n8991# 1.28e-19
C1815 a_23505_n9259# a_24203_n8893# 0.195152f
C1816 x4._21_ a_26147_n9107# 0.011629f
C1817 m2_17442_n2443# x3.x1.nSEL1 0.00815f
C1818 a_23781_n8171# a_23063_n8709# 9.16e-19
C1819 a_23615_n8171# a_23229_n8709# 1.36e-19
C1820 a_24316_n9803# a_23851_n9829# 0.005941f
C1821 x4._04_ a_24371_n8991# 7.11e-19
C1822 x4.net8 a_28979_n8715# 2.29e-20
C1823 a_28099_n9437# x4.clknet_1_1__leaf_clk 3.29e-19
C1824 a_27507_n8893# a_27423_n8893# 0.008508f
C1825 a_23615_n8171# a_24203_n8893# 0.001131f
C1826 a_28470_n8715# x4._11_ 6.96e-20
C1827 a_26159_n7409# a_26998_n8893# 7.91e-22
C1828 x4._11_ a_29063_n8991# 5.38e-21
C1829 a_25709_n7109# a_25875_n7395# 0.017149f
C1830 a_23675_n5233# a_23811_n5073# 0.136009f
C1831 a_23391_n5219# x4._01_ 8.93e-19
C1832 a_23682_n5329# a_23882_n5174# 0.080195f
C1833 x3.x2.GP2 counter7 1.13e-20
C1834 VDD x4.clknet_1_1__leaf_clk 3.34801f
C1835 x4._17_ a_25639_n9259# 1e-20
C1836 x4._21_ a_26559_n9259# 5.62e-21
C1837 x4._09_ a_29021_n9259# 0.001794f
C1838 a_29489_n9803# x4._23_ 0.009249f
C1839 VDD x1.sky130_fd_sc_hd__inv_2_16.A 0.636224f
C1840 a_24125_n10182# a_25229_n10182# 9e-21
C1841 a_27055_n8715# x4.net9 0.002503f
C1842 x4.net4 x4._16_ 0.442589f
C1843 VDD a_23633_n5451# 0.004522f
C1844 counter3 x4.counter[0] 0.117902f
C1845 VDD a_28638_n8741# 0.182123f
C1846 a_24625_n8715# a_24595_n9571# 6.77e-20
C1847 a_27139_n8715# x4.clknet_1_1__leaf_clk 0.001538f
C1848 x4._24_ x4._25_ 0.095329f
C1849 x4._22_ a_28743_n9483# 3.67e-19
C1850 VDD a_28470_n8893# 0.248502f
C1851 a_26295_n7249# x4._06_ 4.29e-19
C1852 a_28457_n9803# x4._15_ 0.087822f
C1853 a_23675_n4933# a_23682_n5329# 3.36e-19
C1854 x1.sky130_fd_sc_hd__inv_2_13.A x1.sky130_fd_sc_hd__inv_2_11.A 5.04e-19
C1855 a_23682_n4633# a_23882_n5174# 1.26e-19
C1856 x4.counter[2] a_23994_n9687# 6.46e-19
C1857 a_23882_n4933# a_23675_n5233# 6.88e-20
C1858 a_26630_n8715# x4.net6 0.019975f
C1859 x4.net9 x4._22_ 0.369389f
C1860 a_25721_n9259# x4._15_ 1.25e-19
C1861 VDD x4._03_ 0.393273f
C1862 x4._21_ x4._06_ 0.224771f
C1863 a_23675_n4933# x4._00_ 0.118744f
C1864 a_24647_n7903# x4.clknet_0_clk 3.43e-19
C1865 x4.counter[6] x4._22_ 9.35e-22
C1866 x4._11_ a_27837_n7261# 2.28e-19
C1867 a_26166_n7505# x4._19_ 0.457296f
C1868 a_28031_n8709# x4.net10 4.73e-19
C1869 a_26147_n9107# x4.net7 0.084753f
C1870 x4.net3 x4._11_ 0.005186f
C1871 a_26593_n7906# x4.net6 0.027058f
C1872 drv_out x4._15_ 0.005511f
C1873 x4.net10 a_28197_n9259# 0.003321f
C1874 x1.sky130_fd_sc_hd__inv_2_16.A select1 1.2e-19
C1875 a_18409_n2290# x3.x2.GP3 0.00144f
C1876 x4._16_ a_25793_n9259# 5.12e-19
C1877 a_26545_n8715# x4._15_ 0.019231f
C1878 x3.nselect2 a_18409_n2290# 1.29e-19
C1879 x3.x1.nSEL0 x3.x2.GN1 0.004375f
C1880 a_25900_n8197# x4._15_ 6.77e-20
C1881 x4._11_ a_25297_n9465# 6.46e-19
C1882 x4.net8 a_26309_n9259# 0.002158f
C1883 a_23339_n9259# a_23505_n9259# 0.970278f
C1884 m3_18866_n4909# x3.x2.GP1 5.81e-19
C1885 x4.net10 a_28979_n8715# 3.67e-19
C1886 a_23682_n4633# a_23675_n4933# 0.966391f
C1887 a_25834_n7921# x4._16_ 0.029136f
C1888 a_26559_n9259# x4.net7 0.003956f
C1889 x4._12_ x4._11_ 0.214271f
C1890 a_26885_n10182# a_26559_n9259# 1.63e-21
C1891 x4.net4 counter3 8.11e-19
C1892 a_23615_n8171# a_23339_n9259# 2.82e-20
C1893 VDD a_26117_n7627# 0.004852f
C1894 x4.clknet_1_0__leaf_clk a_24371_n8991# 1.1e-19
C1895 a_24222_n8059# a_24563_n7805# 9.73e-19
C1896 x4.net8 a_26529_n7849# 0.003186f
C1897 a_24054_n7805# a_24149_n7805# 0.007724f
C1898 counter7 a_22837_n10182# 2.81e-20
C1899 a_25875_n7395# x4._20_ 1.76e-19
C1900 VDD a_24031_n4907# 0.003202f
C1901 a_24095_n8741# x4.net5 6.71e-21
C1902 x4._11_ a_27124_n9259# 0.002651f
C1903 x4._13_ a_23615_n8171# 0.002226f
C1904 x4._11_ a_25875_n7395# 1.82e-19
C1905 x4.counter[9] a_29319_n10347# 0.109832f
C1906 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_17.A 5.48e-19
C1907 x1.sky130_fd_sc_hd__inv_2_2.A x1.sky130_fd_sc_hd__inv_2_17.Y 0.001676f
C1908 a_24125_n10182# a_23851_n9829# 4.71e-19
C1909 VDD x4.clknet_0_clk 2.53166f
C1910 a_26529_n7849# x4._07_ 0.096566f
C1911 a_24981_n8715# x4._11_ 0.00137f
C1912 a_24149_n7805# x4._11_ 0.00121f
C1913 x4.net9 a_29103_n9829# 0.001158f
C1914 a_26159_n7409# x4._05_ 0.196756f
C1915 x4.net4 a_23778_n8893# 0.004091f
C1916 VDD a_22962_n5131# 4.93e-19
C1917 a_26357_n8709# a_26559_n9259# 0.003672f
C1918 a_26191_n8709# a_26725_n9259# 0.003047f
C1919 x4._06_ x4.net7 0.141876f
C1920 x4._14_ a_23927_n8715# 2.97e-21
C1921 a_28470_n8715# x4._23_ 0.012578f
C1922 a_17857_n2290# x3.x2.GN3 6.68e-19
C1923 a_27223_n8741# a_28031_n8709# 4.62e-19
C1924 VDD a_27507_n8893# 0.004788f
C1925 VDD a_23391_n4933# 0.19379f
C1926 a_27807_n9829# x4.net6 0.009771f
C1927 a_29063_n8991# x4._23_ 2.3e-19
C1928 VDD a_25779_n7395# 0.376761f
C1929 a_28895_n8893# x4.net7 1.49e-19
C1930 VDD x3.x2.GP2 1.81711f
C1931 a_28725_n10182# a_28470_n8893# 6.36e-19
C1932 a_29489_n9803# x4.net11 0.004987f
C1933 VDD x1.sky130_fd_sc_hd__inv_2_17.A 0.636188f
C1934 a_23615_n8171# a_23225_n7109# 5.49e-20
C1935 VDD a_24625_n8715# 0.261491f
C1936 a_25179_n7627# x4._19_ 0.001413f
C1937 x4._11_ x4._25_ 2.54e-20
C1938 a_27055_n8715# x4._22_ 1.1e-21
C1939 VDD a_23969_n8171# 0.093135f
C1940 a_26166_n7505# a_26366_n7350# 0.074815f
C1941 a_26159_n7409# a_26295_n7249# 0.136009f
C1942 a_27166_n9147# a_26998_n8893# 0.239923f
C1943 a_26559_n9259# a_27423_n8893# 0.032244f
C1944 a_26725_n9259# a_27591_n8991# 0.034054f
C1945 x4.counter[8] x4._23_ 9.18e-19
C1946 x4._18_ a_23063_n8709# 3.08e-21
C1947 x4.clknet_1_0__leaf_clk a_24031_n5085# 4.64e-19
C1948 x4._06_ a_26357_n8709# 0.183131f
C1949 x4._21_ a_26159_n7409# 8.19e-20
C1950 x1.sky130_fd_sc_hd__inv_2_13.A x1.sky130_fd_sc_hd__inv_2_12.A 0.173286f
C1951 a_24053_n8337# a_24095_n8741# 7.84e-20
C1952 x4._10_ a_23697_n5995# 4.63e-20
C1953 a_23615_n5995# a_23769_n5995# 0.004009f
C1954 VDD a_18537_n1898# 0.001127f
C1955 m3_18876_n6983# x3.x2.GN4 0.084813f
C1956 a_24229_n4907# x4.net1 5.53e-20
C1957 a_25600_n8741# x4._19_ 8.51e-20
C1958 a_27093_n8893# x4.clknet_1_1__leaf_clk 0.001835f
C1959 a_23682_n5329# a_24075_n5995# 0.011211f
C1960 a_23675_n5233# x4._11_ 9.54e-19
C1961 select1 x3.x2.GP2 1.37e-19
C1962 a_24371_n8991# x4._15_ 2.99e-20
C1963 x4._16_ x4.net6 0.291584f
C1964 VDD a_28999_n7408# 0.28996f
C1965 x4._17_ a_25875_n7395# 0.036473f
C1966 x1.sky130_fd_sc_hd__inv_2_17.A select1 1.2e-19
C1967 a_28895_n8715# x4._24_ 0.013075f
C1968 VDD a_28669_n7261# 6.35e-19
C1969 x4._00_ a_24075_n5995# 5.19e-20
C1970 x4._16_ a_23229_n8709# 8.97e-20
C1971 x3.x2.GP3 counter3 4.0653f
C1972 a_28385_n9259# x4._24_ 3.3e-19
C1973 x4._16_ a_24203_n8893# 6.21e-20
C1974 a_26979_n9829# x4.clknet_1_1__leaf_clk 1.84e-19
C1975 a_27251_n7408# x4._24_ 1.86e-20
C1976 a_24054_n7805# a_23927_n8715# 0.002298f
C1977 a_27549_n9259# a_27166_n9147# 4.67e-20
C1978 a_28743_n9483# a_28551_n9803# 6.96e-20
C1979 a_25709_n7109# a_27251_n7408# 1.59e-19
C1980 x4._08_ a_28596_n8337# 0.001882f
C1981 VDD a_23391_n5219# 0.181976f
C1982 a_23682_n4633# a_24075_n5995# 6.42e-21
C1983 x4._14_ a_23063_n8709# 0.001276f
C1984 x4.net9 a_28551_n9803# 0.003753f
C1985 x4._11_ a_23927_n8715# 0.017838f
C1986 a_18409_n2290# x3.x2.GN2 1.63e-19
C1987 VDD a_22837_n10182# 0.25802f
C1988 x4._07_ a_25211_n9231# 2.73e-21
C1989 x3.x1.nSEL0 a_17985_n1898# 2.51e-19
C1990 VDD a_23255_n4363# 0.260172f
C1991 a_28197_n9259# a_28457_n9803# 0.008374f
C1992 x1.sky130_fd_sc_hd__inv_2_8.Y x1.sky130_fd_sc_hd__inv_2_17.Y 0.174714f
C1993 x4._11_ a_23693_n9259# 4.78e-19
C1994 a_28031_n9259# x4.net7 0.007864f
C1995 x4._17_ x4._25_ 1.89e-19
C1996 a_26159_n7409# a_27755_n7261# 2.69e-21
C1997 a_26159_n7409# x4.net7 0.035144f
C1998 x4._22_ a_29103_n9829# 4.31e-19
C1999 a_26542_n7627# x4._17_ 0.002153f
C2000 x4.clknet_1_0__leaf_clk a_23769_n5995# 3.8e-19
C2001 counter3 x4.net6 1.1e-21
C2002 x4.net9 x4.net6 0.566537f
C2003 x4._18_ a_26166_n7505# 1.59e-19
C2004 ring_out a_18409_n2290# 5.47e-20
C2005 x4._20_ a_26725_n9259# 0.003428f
C2006 a_25729_n8715# x4.net7 0.006434f
C2007 x4.net10 a_29133_n9803# 0.001384f
C2008 x4._11_ a_26725_n9259# 0.042209f
C2009 a_28031_n8709# x4._15_ 0.069151f
C2010 x4.net8 x4.clknet_1_1__leaf_clk 0.073766f
C2011 VDD a_24095_n8741# 0.421579f
C2012 a_29063_n8991# x4.net11 0.092457f
C2013 a_28197_n9259# x4._15_ 0.036316f
C2014 VDD a_26147_n9107# 0.226919f
C2015 a_22885_n8715# a_23063_n8709# 5.87e-19
C2016 x4.clknet_1_0__leaf_clk a_23505_n4363# 2.59e-19
C2017 VDD x1.sky130_fd_sc_hd__inv_2_17.Y 0.638508f
C2018 a_24647_n7903# x4._06_ 1.81e-20
C2019 a_28470_n8715# a_28565_n8715# 0.007724f
C2020 a_26159_n7409# a_26357_n8709# 3.93e-19
C2021 a_26166_n7505# a_26191_n8709# 1.6e-20
C2022 x4._07_ x4.clknet_1_1__leaf_clk 0.44529f
C2023 a_18585_n1958# x3.x2.GN1 3.78e-20
C2024 x4.net8 a_28638_n8741# 8.61e-20
C2025 x4.clknet_1_0__leaf_clk a_23597_n8715# 0.001355f
C2026 x4.counter[8] x4.net11 0.024563f
C2027 x4._23_ x4._25_ 0.0063f
C2028 a_23229_n8709# a_23778_n8893# 0.002f
C2029 a_23502_n8715# a_23505_n9259# 0.004962f
C2030 x4._09_ x4._24_ 0.151845f
C2031 x1.sky130_fd_sc_hd__inv_2_14.A x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C2032 x4._08_ x4.net7 1.97e-19
C2033 VDD a_26559_n9259# 0.727748f
C2034 x4._16_ a_23339_n9259# 1.96e-20
C2035 x4._04_ x4.net2 4.09e-22
C2036 a_23615_n8171# a_23502_n8715# 0.002054f
C2037 x4._04_ a_23670_n8741# 8.38e-20
C2038 a_25297_n9465# a_25211_n9465# 0.006584f
C2039 x4.counter[9] x4.net9 5.19e-19
C2040 x4._09_ a_27591_n8991# 0.001669f
C2041 a_28031_n9259# a_27423_n8893# 3.54e-19
C2042 counter7 a_28031_n9259# 2.09e-20
C2043 x4._11_ a_28385_n9259# 2.79e-20
C2044 x4._11_ a_27251_n7408# 0.004334f
C2045 a_26295_n7249# a_26375_n8171# 1.71e-20
C2046 x1.sky130_fd_sc_hd__inv_2_17.Y select1 2.29e-19
C2047 a_25709_n7109# a_26166_n7505# 0.016444f
C2048 drv_out enable_counter 0.391919f
C2049 a_23882_n5174# a_23811_n5073# 0.239923f
C2050 a_23682_n5329# x4._01_ 0.239739f
C2051 a_23781_n8171# a_24222_n8059# 0.111047f
C2052 x4.net2 a_23615_n5995# 0.165774f
C2053 x4._11_ a_23063_n8709# 0.00462f
C2054 drv_out x3.x2.GN1 3.11e-19
C2055 x4._01_ x4._00_ 0.014628f
C2056 x4._21_ a_26375_n8171# 0.053333f
C2057 a_25965_n10182# x4.counter[4] 0.110403f
C2058 x4._08_ a_26357_n8709# 8.29e-20
C2059 x4._05_ x4._19_ 0.284135f
C2060 VDD x4._06_ 0.276236f
C2061 a_25229_n10182# a_25965_n10182# 2.31e-20
C2062 a_28197_n8709# x4.net9 0.001054f
C2063 VDD a_29063_n8741# 0.48745f
C2064 x4.net9 a_28638_n9147# 0.022365f
C2065 a_27194_n8171# a_27807_n9829# 4.57e-20
C2066 a_25179_n7627# x4._18_ 0.09549f
C2067 x4.net10 x4.clknet_1_1__leaf_clk 6.99e-20
C2068 x4._17_ a_26725_n9259# 6.74e-21
C2069 x4._22_ a_28551_n9803# 0.063386f
C2070 VDD a_28895_n8893# 0.215619f
C2071 a_24220_n9483# x4._15_ 8.81e-20
C2072 a_23882_n4933# a_23882_n5174# 0.013851f
C2073 a_23682_n4633# x4._01_ 8.68e-20
C2074 a_23675_n4933# a_23811_n5073# 5.28e-20
C2075 a_27055_n8715# x4.net6 8.63e-19
C2076 x4._04_ x4.clknet_1_1__leaf_clk 1.67e-21
C2077 x3.x2.GN2 counter3 0.004367f
C2078 x4._09_ a_28979_n8893# 6.12e-19
C2079 x4.net8 x4.clknet_0_clk 8.45e-19
C2080 a_23811_n4907# x4._00_ 0.005564f
C2081 a_26295_n7249# x4._19_ 0.040707f
C2082 x4._13_ counter3 0.003357f
C2083 a_28638_n8741# x4.net10 2.56e-19
C2084 x4._22_ x4.net6 0.641715f
C2085 x4._18_ a_25600_n8741# 0.079699f
C2086 x4.net10 a_28470_n8893# 5.45e-19
C2087 x3.nselect2 a_19061_n2032# 9.77e-20
C2088 a_26529_n7849# x4._15_ 2.91e-20
C2089 x4._21_ x4._19_ 7.87e-20
C2090 a_25359_n7627# x4._16_ 1.86e-20
C2091 x4.clknet_0_clk x4._07_ 0.114561f
C2092 x4._03_ a_23946_n9147# 0.006259f
C2093 a_23339_n9259# a_23778_n8893# 0.273138f
C2094 x4.net8 a_25779_n7395# 1.16e-19
C2095 VDD a_19235_n1926# 7.45e-19
C2096 a_23675_n4933# a_23882_n4933# 0.273138f
C2097 a_23682_n4633# a_23811_n4907# 0.110715f
C2098 a_27194_n8171# x4._16_ 0.001016f
C2099 x4.clknet_1_0__leaf_clk x4.net2 0.026712f
C2100 a_27166_n9147# x4.net7 0.005145f
C2101 x4.clknet_1_0__leaf_clk a_23670_n8741# 0.01796f
C2102 a_26375_n8171# x4.net7 2.13e-20
C2103 x4._17_ a_27251_n7408# 0.019971f
C2104 a_25600_n8741# a_26191_n8709# 0.044245f
C2105 a_23781_n8171# x4._21_ 2.75e-21
C2106 counter3 x4.counter[1] 0.099026f
C2107 a_24054_n7805# a_24180_n8171# 0.005525f
C2108 counter7 a_24125_n10182# 2.81e-20
C2109 x4._11_ x4._09_ 0.004259f
C2110 a_24595_n8741# x4.net5 0.001034f
C2111 a_25875_n7395# a_25667_n8171# 9.42e-20
C2112 x4._11_ a_26166_n7505# 3.7e-19
C2113 x4.net1 x4._10_ 0.033245f
C2114 x4.net6 a_26094_n7261# 1.91e-20
C2115 x1.sky130_fd_sc_hd__inv_2_14.A x1.sky130_fd_sc_hd__inv_2_13.A 0.173286f
C2116 x4.net4 x4.net6 0.008308f
C2117 a_27223_n8741# x4.clknet_1_1__leaf_clk 0.005058f
C2118 VDD a_24316_n9803# 0.012117f
C2119 a_24180_n8171# x4._11_ 0.003523f
C2120 x4.net4 a_23229_n8709# 0.002039f
C2121 a_26366_n7350# x4._05_ 3.36e-19
C2122 x4.net4 a_24203_n8893# 0.022715f
C2123 m3_18866_n4909# m3_18862_n5953# 0.003764f
C2124 select1 a_19235_n1926# 8.84e-19
C2125 x4.net3 a_23505_n9259# 0.00115f
C2126 a_26357_n8709# a_27166_n9147# 6.74e-19
C2127 a_26191_n8709# a_26998_n8893# 4.58e-19
C2128 a_26798_n8741# a_26725_n9259# 0.001607f
C2129 a_25709_n7109# a_25600_n8741# 4.81e-21
C2130 a_27055_n8715# a_28197_n8709# 8.68e-20
C2131 a_18409_n2290# x3.x2.GN3 0.104151f
C2132 a_28399_n7627# x4._24_ 0.095435f
C2133 VDD a_28031_n9259# 0.667506f
C2134 a_23615_n8171# x4.net3 1.48e-19
C2135 a_29103_n9829# x4.net6 4.97e-21
C2136 a_28385_n9259# x4._23_ 0.012973f
C2137 VDD a_26159_n7409# 0.438492f
C2138 a_28031_n8709# a_28197_n9259# 2.64e-19
C2139 a_28565_n8893# x4.net7 1.13e-19
C2140 a_27251_n7408# x4._23_ 1.03e-19
C2141 a_22879_n5451# x4.net1 0.060735f
C2142 x4._19_ x4.net7 0.552257f
C2143 a_29319_n10347# a_29063_n8991# 3.35e-20
C2144 a_24595_n8741# a_24595_n9571# 8.07e-19
C2145 a_27194_n8171# x4.net9 0.111158f
C2146 a_24220_n9483# a_24371_n8991# 0.001062f
C2147 VDD a_25729_n8715# 0.206364f
C2148 a_28197_n8709# x4._22_ 4.96e-21
C2149 VDD a_24563_n7805# 0.004177f
C2150 a_26366_n7350# a_26295_n7249# 0.239923f
C2151 a_26559_n9259# a_27093_n8893# 0.002698f
C2152 a_26725_n9259# a_26913_n9259# 0.095025f
C2153 a_27166_n9147# a_27423_n8893# 0.036838f
C2154 x4._22_ a_28638_n9147# 8.71e-19
C2155 x4.clknet_1_0__leaf_clk a_23633_n5451# 0.002574f
C2156 a_26756_n8337# x4.net6 0.001426f
C2157 a_25834_n7921# x4.net6 0.074355f
C2158 x3.x1.nSEL1 a_17405_n2032# 0.193944f
C2159 x4.counter[8] a_29319_n10347# 0.006251f
C2160 x4._21_ a_26366_n7350# 0.0043f
C2161 x4._13_ x4.counter[0] 3.39e-20
C2162 a_24222_n8059# x4._18_ 1.41e-19
C2163 a_26979_n9829# a_26559_n9259# 0.009169f
C2164 a_26357_n8709# x4._19_ 4.93e-21
C2165 x4._14_ a_23851_n9829# 0.134293f
C2166 x4.net9 a_28579_n7627# 7.48e-22
C2167 a_25211_n9231# x4._15_ 0.22097f
C2168 x4.clknet_1_0__leaf_clk x4._03_ 0.00668f
C2169 x4._11_ x4.counter[4] 6.77e-20
C2170 x4._04_ a_24625_n8715# 0.072162f
C2171 x4._04_ a_23969_n8171# 0.126198f
C2172 a_23615_n8171# a_24149_n7805# 0.002698f
C2173 x4._17_ a_26166_n7505# 0.050404f
C2174 VDD x4._08_ 0.467036f
C2175 x4._16_ a_23502_n8715# 1.68e-20
C2176 a_23851_n9829# a_23994_n9687# 0.221119f
C2177 x4._11_ a_25179_n7627# 0.001422f
C2178 x4._16_ a_25639_n9259# 0.105405f
C2179 a_24647_n7903# a_24595_n8741# 0.004132f
C2180 x4.counter[0] x4.counter[1] 0.079742f
C2181 x4.net8 a_26147_n9107# 0.236033f
C2182 a_27549_n9259# a_27591_n8991# 7.84e-20
C2183 a_23781_n8171# x4.net5 3.57e-21
C2184 x4._22_ a_26713_n7249# 0.001069f
C2185 a_27271_n9437# x4.net7 0.006602f
C2186 enable_counter a_23941_n3056# 0.231636f
C2187 a_27223_n8741# x4.clknet_0_clk 0.01296f
C2188 x4._18_ x4._05_ 1.11e-19
C2189 a_17857_n2290# select0 0.246189f
C2190 x4.net4 a_23339_n9259# 0.008383f
C2191 VDD a_23682_n5329# 0.309635f
C2192 a_25600_n8741# x4._20_ 3.36e-20
C2193 a_23675_n4933# x4._11_ 8.58e-21
C2194 drv_out x4.clknet_1_1__leaf_clk 0.008913f
C2195 x4.net9 a_29489_n9803# 3.29e-19
C2196 x4.net1 a_23697_n5995# 0.00162f
C2197 a_19061_n2032# x3.x2.GN2 7.58e-21
C2198 x4._16_ a_25297_n9231# 5.76e-19
C2199 x3.x2.GN1 a_17579_n1926# 0.001144f
C2200 x4._11_ a_25600_n8741# 0.058411f
C2201 a_26545_n8715# x4.clknet_1_1__leaf_clk 0.017223f
C2202 VDD a_24125_n10182# 0.317416f
C2203 a_28470_n8893# a_28457_n9803# 2.47e-19
C2204 x4._07_ a_26147_n9107# 1.81e-19
C2205 x4.net4 x4._13_ 0.050083f
C2206 VDD x4._00_ 0.655201f
C2207 x4.clknet_0_clk a_26457_n7849# 2.68e-20
C2208 x4.clknet_1_0__leaf_clk a_24031_n4907# 0.002297f
C2209 x4._11_ a_24287_n8893# 0.002515f
C2210 x1.sky130_fd_sc_hd__inv_2_15.A x1.sky130_fd_sc_hd__inv_2_13.A 5.04e-19
C2211 x4._09_ x4._23_ 0.130147f
C2212 x4.clknet_1_1__leaf_clk x4._15_ 0.471647f
C2213 x4.net8 a_26559_n9259# 0.009204f
C2214 a_28725_n10182# a_28031_n9259# 4.75e-20
C2215 a_28551_n9803# x4.net6 7.2e-20
C2216 a_26366_n7350# x4.net7 0.026259f
C2217 x4.clknet_1_0__leaf_clk x4.clknet_0_clk 0.004956f
C2218 x4.net1 a_23337_n4363# 0.010028f
C2219 ring_out a_19061_n2032# 0.001281f
C2220 x4._18_ a_26295_n7249# 7.52e-20
C2221 x4._20_ a_26998_n8893# 9.2e-20
C2222 a_27194_n8171# a_27055_n8715# 5.73e-19
C2223 a_17857_n2290# x3.x2.GP1 9.92e-19
C2224 x4._07_ a_26559_n9259# 0.112051f
C2225 VDD a_23682_n4633# 0.335402f
C2226 x4._11_ a_26998_n8893# 0.026293f
C2227 a_28638_n8741# x4._15_ 4.57e-19
C2228 VDD a_24595_n8741# 0.252112f
C2229 x3.x2.GN3 counter3 3.89796f
C2230 x4._21_ x4._18_ 0.005609f
C2231 x4.net4 x4.counter[1] 3.68e-19
C2232 a_28470_n8893# x4._15_ 0.001788f
C2233 x4._05_ x4._24_ 2.08e-20
C2234 VDD a_23873_n8893# 0.005794f
C2235 x4.clknet_1_0__leaf_clk a_23391_n4933# 0.038899f
C2236 a_27194_n8171# x4._22_ 8.12e-19
C2237 x4.clknet_0_clk a_25449_n7261# 9.48e-20
C2238 x4.net8 x4._06_ 0.209874f
C2239 a_23229_n8709# x4.net6 1.26e-19
C2240 x4.net4 a_23225_n7109# 4.87e-19
C2241 ring_out enable_ring 0.549705f
C2242 a_26366_n7350# a_26357_n8709# 8.21e-21
C2243 x4._11_ a_23851_n9829# 7.66e-19
C2244 a_26295_n7249# a_26191_n8709# 5.48e-20
C2245 a_25709_n7109# x4._05_ 0.005813f
C2246 x4.net8 a_29063_n8741# 4.93e-20
C2247 a_23969_n8171# x4.clknet_1_0__leaf_clk 0.003123f
C2248 x4._17_ a_25179_n7627# 0.250762f
C2249 a_23255_n4363# a_23615_n5995# 2.44e-21
C2250 a_23927_n8715# a_23505_n9259# 0.003824f
C2251 a_23502_n8715# a_23778_n8893# 4.47e-19
C2252 a_24095_n8741# a_23946_n9147# 0.001344f
C2253 a_27181_n8337# a_26798_n8741# 4.67e-20
C2254 x4._21_ a_26191_n8709# 0.016583f
C2255 a_23505_n9259# a_23693_n9259# 0.097994f
C2256 a_24371_n8991# a_25211_n9231# 7.43e-20
C2257 x4._06_ x4._07_ 5.11e-20
C2258 VDD a_27166_n9147# 0.183641f
C2259 VDD x3.x1.nSEL1 0.646724f
C2260 VDD a_26375_n8171# 0.011033f
C2261 a_23615_n8171# a_23927_n8715# 0.001393f
C2262 x4._04_ a_24095_n8741# 0.008333f
C2263 a_23628_n8337# x4._11_ 4.01e-19
C2264 a_28596_n8337# x4._24_ 9.29e-19
C2265 x4._11_ a_27549_n9259# 2.44e-19
C2266 x4._17_ a_25600_n8741# 1.33e-19
C2267 VDD a_29021_n9259# 4.71e-19
C2268 a_25709_n7109# a_26295_n7249# 0.013455f
C2269 a_23295_n5219# a_22879_n5451# 5.03e-19
C2270 a_18585_n1958# x3.x2.GP2 3.2e-20
C2271 a_24222_n8059# a_24054_n7805# 0.239923f
C2272 a_23391_n5219# a_23610_n5085# 0.006169f
C2273 a_23811_n5073# x4._01_ 0.00226f
C2274 a_23781_n8171# a_24647_n7903# 0.034054f
C2275 x3.x2.GN2 x3.x2.GP3 0.004296f
C2276 drv_out x4.clknet_0_clk 0.00889f
C2277 x4._21_ a_25709_n7109# 0.001038f
C2278 a_25900_n8197# x4.clknet_0_clk 7.65e-20
C2279 a_25965_n10182# a_26885_n10182# 1.37e-20
C2280 a_28551_n9803# a_28638_n9147# 5.71e-20
C2281 x4._17_ a_28399_n7627# 0.056144f
C2282 x4._18_ x4.net7 0.004371f
C2283 a_24222_n8059# x4._11_ 0.032361f
C2284 x4.net3 x4._16_ 6.72e-19
C2285 x4.clknet_0_clk x4._15_ 4.05e-19
C2286 VDD a_23417_n8715# 0.075425f
C2287 x3.x1.nSEL1 select1 0.272823f
C2288 ring_out x3.x2.GP3 0.080819f
C2289 x4.net9 a_29063_n8991# 0.001937f
C2290 ring_out x3.nselect2 0.006614f
C2291 VDD a_28565_n8893# 0.002923f
C2292 a_18409_n2290# x3.x2.GN4 6.84e-19
C2293 VDD x4._19_ 0.197759f
C2294 x4._16_ a_25297_n9465# 8.82e-20
C2295 x4._11_ a_24329_n9259# 5.7e-19
C2296 x4.clknet_1_0__leaf_clk a_23391_n5219# 0.044938f
C2297 a_23811_n4907# a_23811_n5073# 0.013661f
C2298 a_28197_n8709# x4.net6 1.27e-19
C2299 drv_out x3.x2.GP2 4.09557f
C2300 VDD x4._02_ 0.325572f
C2301 x1.sky130_fd_sc_hd__inv_2_15.A x1.sky130_fd_sc_hd__inv_2_14.A 0.173286f
C2302 x4._09_ x4.net11 0.071633f
C2303 a_25900_n8197# a_25779_n7395# 0.002561f
C2304 a_24075_n5995# x4._11_ 0.201886f
C2305 a_24058_n4541# x4._00_ 8.32e-19
C2306 x4.clknet_1_0__leaf_clk a_23255_n4363# 3.24e-19
C2307 a_26191_n8709# x4.net7 0.088061f
C2308 a_25779_n7395# x4._15_ 1.78e-19
C2309 x4.counter[8] x4.net9 2.39e-19
C2310 a_26191_n8709# a_26885_n10182# 1.7e-21
C2311 a_25729_n8395# a_25729_n8715# 6.96e-20
C2312 a_28895_n8715# a_29021_n8337# 0.006169f
C2313 a_29063_n8741# x4.net10 0.084593f
C2314 a_25965_n10182# x4.net5 0.001724f
C2315 VDD a_23781_n8171# 0.304738f
C2316 x4.net10 a_28895_n8893# 0.003817f
C2317 x4._11_ x4._05_ 0.023537f
C2318 a_25875_n7395# x4._16_ 1.29e-20
C2319 x1.sky130_fd_sc_hd__inv_2_15.A x3.x2.GN1 2.09e-20
C2320 a_27755_n7261# x4._24_ 4.18e-19
C2321 x4._23_ a_28399_n7627# 0.213625f
C2322 a_23063_n8709# a_23505_n9259# 2.24e-19
C2323 a_23229_n8709# a_23339_n9259# 0.010101f
C2324 x4.net7 x4._24_ 2.68e-19
C2325 x4.net8 a_28031_n9259# 3.27e-19
C2326 x4._13_ x4.net6 2.81e-21
C2327 a_23339_n9259# a_24203_n8893# 0.032244f
C2328 x4._03_ a_24371_n8991# 3.08e-19
C2329 a_23882_n4933# a_23811_n4907# 0.239923f
C2330 x4.net8 a_26159_n7409# 0.001356f
C2331 a_24981_n8715# x4._16_ 0.010038f
C2332 a_26630_n8715# a_26725_n9259# 8.92e-19
C2333 a_27223_n8741# a_26559_n9259# 0.002274f
C2334 a_23615_n8171# a_23063_n8709# 0.002682f
C2335 x4._13_ a_23229_n8709# 1.58e-19
C2336 a_27591_n8991# x4.net7 0.064911f
C2337 x4.clknet_1_0__leaf_clk a_24095_n8741# 0.002373f
C2338 x1.sky130_fd_sc_hd__nand2_2_0.B enable_ring 0.108977f
C2339 a_25709_n7109# x4.net7 0.002812f
C2340 x4.net8 a_25729_n8715# 2.79e-20
C2341 x4.net3 counter3 6.21e-20
C2342 a_26191_n8709# a_26357_n8709# 0.961627f
C2343 x4._16_ x4.counter[2] 3.86e-19
C2344 counter7 a_25965_n10182# 2.81e-20
C2345 a_26159_n7409# x4._07_ 5.99e-19
C2346 a_23904_n9259# x4.net5 3e-19
C2347 x4._11_ a_26295_n7249# 5.19e-20
C2348 x4._15_ a_28999_n7408# 8.98e-20
C2349 x4.net6 a_26713_n7249# 9.51e-20
C2350 x4._21_ x4._20_ 0.296715f
C2351 a_29489_n9803# a_29103_n9829# 0.006406f
C2352 a_28031_n8709# x4.clknet_1_1__leaf_clk 0.285659f
C2353 a_28197_n9259# x4.clknet_1_1__leaf_clk 0.031849f
C2354 x4._21_ x4._11_ 0.059807f
C2355 a_24222_n8059# x4._17_ 2.52e-22
C2356 x4.net4 a_23502_n8715# 4.27e-19
C2357 x4.net3 a_23778_n8893# 3.32e-20
C2358 m3_18862_n5953# m3_18876_n6983# 0.003741f
C2359 a_27223_n8741# x4._06_ 1.75e-19
C2360 a_25709_n7109# a_26357_n8709# 4.98e-20
C2361 x4.net9 a_27124_n9259# 3.93e-19
C2362 a_28031_n8709# a_28638_n8741# 0.141453f
C2363 a_19061_n2032# x3.x2.GN3 1.07e-20
C2364 x4._14_ x4.net5 0.258421f
C2365 x3.x2.GN1 a_17985_n1898# 1.22e-20
C2366 x4._08_ x4.net8 2.38e-19
C2367 a_23225_n7109# a_23229_n8709# 1.82e-21
C2368 a_28197_n8709# a_28638_n9147# 2.96e-21
C2369 a_28638_n8741# a_28197_n9259# 2.96e-21
C2370 a_28031_n8709# a_28470_n8893# 1.73e-19
C2371 VDD a_26366_n7350# 0.266088f
C2372 a_28979_n8893# x4.net7 3.05e-20
C2373 a_24229_n5073# x4.net1 6.38e-20
C2374 a_28197_n9259# a_28470_n8893# 0.078545f
C2375 a_26381_n9259# x4.net6 7.29e-19
C2376 a_23994_n9687# x4.net5 3.95e-20
C2377 VDD a_28385_n8715# 0.078044f
C2378 VDD a_25762_n7921# 0.011634f
C2379 a_25359_n7627# x4.net6 1.5e-19
C2380 x4.net2 a_23505_n4363# 0.008042f
C2381 x4._08_ x4._07_ 9.41e-21
C2382 a_28638_n8741# a_28979_n8715# 9.73e-19
C2383 a_27591_n8991# a_27423_n8893# 0.310858f
C2384 x4._17_ x4._05_ 0.0576f
C2385 x4.net3 x4._10_ 0.003052f
C2386 a_26998_n8893# a_26913_n9259# 0.037333f
C2387 counter3 x4.counter[2] 0.16993f
C2388 a_25793_n9259# a_25639_n9259# 0.004009f
C2389 x1.sky130_fd_sc_hd__nand2_2_0.B x3.nselect2 2.88e-20
C2390 a_29021_n8337# x4._09_ 1.66e-19
C2391 x4.net10 a_28031_n9259# 0.001924f
C2392 x3.x1.nSEL1 a_18033_n1958# 0.041068f
C2393 a_27194_n8171# x4.net6 0.047825f
C2394 x4.counter[5] x4.counter[4] 0.068962f
C2395 x3.x2.GN4 counter3 0.237196f
C2396 a_24011_n8715# a_23229_n8709# 6.32e-19
C2397 x1.sky130_fd_sc_hd__inv_2_16.A x1.sky130_fd_sc_hd__inv_2_14.A 5.04e-19
C2398 a_24625_n8715# a_24371_n8991# 0.001352f
C2399 a_24647_n7903# x4._18_ 0.001543f
C2400 a_26979_n9829# a_27166_n9147# 3.07e-19
C2401 a_25834_n7921# a_25639_n9259# 5.65e-20
C2402 x4._14_ a_24595_n9571# 0.112679f
C2403 a_24095_n8741# x4._15_ 1.37e-19
C2404 x4._20_ x4.net7 0.035834f
C2405 x4._12_ x4._10_ 0.002721f
C2406 x4._01_ x4._11_ 0.20957f
C2407 a_26147_n9107# x4._15_ 2.8e-19
C2408 x4._11_ a_27755_n7261# 0.087773f
C2409 x4.counter[2] a_23778_n8893# 1.99e-20
C2410 x4._13_ a_23339_n9259# 6.65e-20
C2411 x4._11_ x4.net7 0.966176f
C2412 x4._17_ a_26295_n7249# 0.016441f
C2413 x4.net3 a_22879_n5451# 0.042192f
C2414 ring_out x3.x2.GN2 0.23158f
C2415 x4._16_ a_23927_n8715# 1.35e-19
C2416 a_28596_n9259# x4._24_ 6.57e-19
C2417 x4.net6 a_28579_n7627# 7.38e-20
C2418 x4._21_ x4._17_ 0.019243f
C2419 x4._05_ x4._23_ 9.36e-20
C2420 a_24054_n7805# x4.net5 1.47e-19
C2421 a_23610_n4907# x4.net1 2.14e-19
C2422 a_26559_n9259# x4._15_ 4.49e-20
C2423 a_28003_n9437# x4.net7 6.49e-19
C2424 x1.sky130_fd_sc_hd__inv_2_9.A enable_ring 6.29e-19
C2425 a_18409_n2290# select0 0.086353f
C2426 x4._12_ a_22879_n5451# 0.090947f
C2427 x4._08_ x4.net10 0.001321f
C2428 VDD a_23811_n5073# 0.211083f
C2429 counter3 a_23205_n10182# 4.27e-20
C2430 x4.net1 a_23225_n7109# 0.001584f
C2431 x4.net5 x4._20_ 8.42e-21
C2432 x3.x2.GN3 x3.x2.GP3 2.86851f
C2433 x4._16_ a_26725_n9259# 4.88e-21
C2434 x4._11_ a_26357_n8709# 8.46e-20
C2435 x3.nselect2 x3.x2.GN3 7.39e-21
C2436 VDD a_25965_n10182# 0.287214f
C2437 a_28895_n8893# a_28457_n9803# 2.58e-19
C2438 a_29063_n8991# a_29103_n9829# 0.005283f
C2439 a_26529_n7849# x4.clknet_1_1__leaf_clk 7.2e-19
C2440 x4._11_ x4.net5 0.388184f
C2441 VDD x4._18_ 0.686881f
C2442 x4.net8 a_27166_n9147# 0.00264f
C2443 a_26630_n8715# a_26166_n7505# 9.47e-20
C2444 x4.net8 a_26375_n8171# 0.009814f
C2445 a_26545_n8715# x4._06_ 0.114717f
C2446 a_25900_n8197# x4._06_ 0.004838f
C2447 a_26798_n8741# x4._05_ 8.7e-19
C2448 a_24220_n9483# x4._03_ 9.33e-19
C2449 x4.net1 a_23295_n4755# 0.045364f
C2450 a_28596_n8337# x4._23_ 9.59e-19
C2451 x4._06_ x4._15_ 0.139237f
C2452 x4.counter[8] a_29103_n9829# 0.001844f
C2453 x4._20_ a_27423_n8893# 1.2e-20
C2454 a_27194_n8171# a_28197_n8709# 0.008007f
C2455 x4._22_ a_27124_n9259# 6.82e-19
C2456 x4._07_ a_27166_n9147# 0.004454f
C2457 a_18409_n2290# x3.x2.GP1 1.21e-20
C2458 VDD a_23882_n4933# 0.286747f
C2459 a_29063_n8741# x4._15_ 1.61e-19
C2460 a_27194_n8171# a_28638_n9147# 7.13e-20
C2461 x4._11_ a_27423_n8893# 0.045045f
C2462 a_26166_n7505# a_26593_n7906# 0.003687f
C2463 x3.x1.nSEL0 x3.x1.nSEL1 0.352716f
C2464 x4.net4 x4.net3 0.0313f
C2465 VDD a_26191_n8709# 0.421866f
C2466 x4._11_ counter7 2.85e-19
C2467 VDD a_23904_n9259# 0.003212f
C2468 x4.clknet_0_clk a_26515_n7261# 4.62e-19
C2469 x4._17_ a_27755_n7261# 0.139841f
C2470 a_23502_n8715# x4.net6 6.57e-20
C2471 x4._17_ x4.net7 0.072785f
C2472 x4.net3 a_23697_n5995# 1.25e-19
C2473 a_23682_n5329# a_23615_n5995# 1.58e-19
C2474 a_23675_n5233# x4._10_ 0.011255f
C2475 x4._11_ a_24595_n9571# 0.159397f
C2476 a_25639_n9259# x4.net6 0.005791f
C2477 VDD x4._24_ 0.6956f
C2478 a_23229_n8709# a_23502_n8715# 0.078737f
C2479 x1.sky130_fd_sc_hd__inv_2_9.A x3.nselect2 5.69e-21
C2480 a_28031_n8709# a_28999_n7408# 7.7e-20
C2481 a_28197_n8709# a_28579_n7627# 6.98e-21
C2482 a_24095_n8741# a_24371_n8991# 0.007214f
C2483 a_23927_n8715# a_23778_n8893# 0.001152f
C2484 x4._16_ a_23063_n8709# 0.001516f
C2485 x4.net9 a_26725_n9259# 0.017191f
C2486 x4.net8 x4._19_ 2.14e-19
C2487 x4._08_ a_27223_n8741# 9.54e-19
C2488 a_28638_n9147# a_28579_n7627# 1.02e-20
C2489 a_23505_n9259# a_24287_n8893# 3.14e-19
C2490 a_23778_n8893# a_23693_n9259# 0.037333f
C2491 VDD a_27591_n8991# 0.400861f
C2492 x1.sky130_fd_sc_hd__inv_2_16.A x1.sky130_fd_sc_hd__inv_2_15.A 0.173286f
C2493 VDD x4._14_ 0.685574f
C2494 a_25875_n7395# a_26094_n7261# 0.006169f
C2495 VDD a_25709_n7109# 1.29479f
C2496 m3_18876_n6983# counter7 0.117708f
C2497 a_23610_n4907# a_23295_n4755# 7.84e-20
C2498 x4._04_ a_24595_n8741# 0.171873f
C2499 a_27271_n9437# a_26979_n9829# 0.001675f
C2500 enable_counter a_23391_n4933# 2.06e-20
C2501 a_24053_n8337# x4._11_ 6.78e-19
C2502 x4._11_ a_28596_n9259# 4.03e-21
C2503 VDD a_23994_n9687# 0.108977f
C2504 x4._17_ a_26357_n8709# 1.22e-20
C2505 x3.x2.GN1 x3.x2.GP2 0.005192f
C2506 x4.net4 a_24981_n8715# 6.79e-19
C2507 a_24222_n8059# a_24479_n7805# 0.036838f
C2508 a_23781_n8171# x4.net8 0.001542f
C2509 a_27755_n7261# x4._23_ 0.026998f
C2510 x4.net7 x4._23_ 0.074369f
C2511 a_28031_n9259# a_28457_n9803# 9.12e-19
C2512 x4._09_ a_27807_n9829# 1.89e-19
C2513 x4.net4 x4.counter[2] 0.006188f
C2514 a_27805_n10182# x4.net7 4.41e-19
C2515 a_26529_n7849# x4.clknet_0_clk 0.034583f
C2516 a_23295_n5219# x4.net1 0.081622f
C2517 a_26885_n10182# a_27805_n10182# 1.37e-20
C2518 a_23505_n4363# a_23391_n4933# 1.96e-19
C2519 a_28895_n8715# x4.net9 2.45e-19
C2520 a_24647_n7903# x4._11_ 0.052724f
C2521 a_23851_n9829# a_23505_n9259# 0.010515f
C2522 x1.sky130_fd_sc_hd__inv_2_7.Y enable_ring 3.49e-19
C2523 VDD a_22885_n8715# 0.006911f
C2524 x1.sky130_fd_sc_hd__nand2_2_0.B ring_out 0.083309f
C2525 x4.net9 a_28385_n9259# 0.016338f
C2526 a_25211_n9231# x4.clknet_1_1__leaf_clk 2.67e-20
C2527 x4.net9 a_27251_n7408# 3.61e-20
C2528 VDD a_28979_n8893# 0.005629f
C2529 a_19061_n2032# x3.x2.GN4 0.134079f
C2530 x4.clknet_1_0__leaf_clk a_23682_n5329# 0.083453f
C2531 drv_out a_26159_n7409# 4.16e-19
C2532 a_26545_n8715# a_26159_n7409# 6.17e-21
C2533 x4._11_ a_24605_n8171# 8.02e-19
C2534 a_25834_n7921# a_25875_n7395# 0.001715f
C2535 a_28031_n9259# x4._15_ 0.02569f
C2536 x4.net8 a_27271_n9437# 0.001229f
C2537 x4.clknet_1_0__leaf_clk x4._00_ 0.144154f
C2538 a_26798_n8741# x4.net7 0.040813f
C2539 a_26159_n7409# x4._15_ 3.85e-20
C2540 a_25900_n8197# a_25729_n8715# 1.06e-19
C2541 a_27925_n7261# x4.clknet_0_clk 9.17e-20
C2542 VDD a_24054_n7805# 0.255338f
C2543 a_25729_n8715# x4._15_ 0.046541f
C2544 x4._04_ a_23417_n8715# 3.27e-21
C2545 a_26166_n7505# x4._16_ 6.29e-20
C2546 x4._11_ a_28099_n9437# 0.006396f
C2547 x4.net2 x4._03_ 5.34e-20
C2548 a_23502_n8715# a_23339_n9259# 4.57e-19
C2549 a_23063_n8709# a_23778_n8893# 0.001041f
C2550 a_23670_n8741# x4._03_ 0.009555f
C2551 x3.x2.GP1 counter3 5.62e-21
C2552 x3.x2.GN2 x3.x2.GN3 0.067463f
C2553 a_28725_n10182# x4._24_ 0.00116f
C2554 a_23339_n9259# a_25639_n9259# 1.62e-21
C2555 x4._03_ a_25211_n9231# 2.2e-20
C2556 VDD x4._20_ 0.175404f
C2557 a_23682_n4633# x4.clknet_1_0__leaf_clk 0.470509f
C2558 a_23675_n4933# a_24229_n4907# 0.062224f
C2559 a_23882_n4933# a_24058_n4541# 0.007724f
C2560 a_23811_n4907# a_23633_n4541# 9.73e-19
C2561 x4.net8 a_26366_n7350# 5.83e-19
C2562 x4.net4 a_23205_n10182# 7.77e-19
C2563 a_24180_n8171# x4._16_ 2.63e-21
C2564 a_27423_n8893# x4._23_ 0.001187f
C2565 a_27223_n8741# a_27166_n9147# 6.84e-19
C2566 a_27055_n8715# a_26725_n9259# 1.5e-19
C2567 x4._04_ x4._02_ 1.6e-19
C2568 x4.clknet_1_0__leaf_clk a_24595_n8741# 1.95e-19
C2569 a_26913_n9259# x4.net7 4.68e-19
C2570 VDD x4._11_ 5.18499f
C2571 counter7 x4._23_ 0.004833f
C2572 a_26885_n10182# a_26913_n9259# 7.39e-20
C2573 a_27805_n10182# a_27423_n8893# 3.85e-20
C2574 a_28197_n9259# a_26559_n9259# 8.05e-21
C2575 x4.clknet_1_0__leaf_clk a_23873_n8893# 5.04e-19
C2576 x4.net8 a_28385_n8715# 1.28e-19
C2577 a_26357_n8709# a_26798_n8741# 0.110715f
C2578 counter7 a_27805_n10182# 8.66e-19
C2579 a_24479_n7805# x4._21_ 8.88e-21
C2580 x4.net8 a_25762_n7921# 0.001644f
C2581 a_27194_n8171# a_28579_n7627# 0.006666f
C2582 ring_out x3.x2.GN3 0.080584f
C2583 x4._04_ a_23781_n8171# 0.215918f
C2584 a_23615_n8171# a_24222_n8059# 0.136461f
C2585 x4._22_ a_26725_n9259# 0.02378f
C2586 a_25211_n9465# x4.net7 2.04e-20
C2587 x4.net9 a_27175_n9437# 0.001755f
C2588 a_26593_n7906# a_26816_n8171# 3.74e-19
C2589 a_26457_n7849# a_26375_n8171# 2.78e-19
C2590 x4._08_ x4._15_ 0.030258f
C2591 a_28638_n8741# x4.clknet_1_1__leaf_clk 5.16e-19
C2592 VDD a_28003_n9437# 0.001618f
C2593 x1.sky130_fd_sc_hd__inv_2_17.A x1.sky130_fd_sc_hd__inv_2_15.A 5.04e-19
C2594 a_23295_n5219# a_23295_n4755# 0.025128f
C2595 x4._21_ a_25667_n8171# 0.002821f
C2596 a_28470_n8893# x4.clknet_1_1__leaf_clk 3.02e-19
C2597 a_24647_n7903# x4._17_ 1.35e-20
C2598 a_24031_n4907# x4.net2 1.37e-19
C2599 x4.net3 a_23229_n8709# 0.007798f
C2600 x4.net4 a_23927_n8715# 0.006897f
C2601 a_23255_n4363# a_23505_n4363# 0.025037f
C2602 x4.net4 a_23693_n9259# 4.45e-19
C2603 x4.net3 a_24203_n8893# 1.53e-21
C2604 a_28031_n8709# x4._06_ 4.19e-21
C2605 a_24229_n5073# a_24058_n5451# 0.001229f
C2606 a_23421_n7921# x4._11_ 0.002118f
C2607 x4.counter[9] x4.counter[8] 0.299988f
C2608 x4.net9 x4._09_ 0.571636f
C2609 a_23225_n7109# a_23502_n8715# 7.35e-19
C2610 a_28031_n8709# a_29063_n8741# 0.048748f
C2611 a_28197_n8709# a_28470_n8715# 0.078545f
C2612 x3.x2.GN4 x3.x2.GP3 3.4436f
C2613 x3.nselect2 x3.x2.GN4 1.53e-20
C2614 a_26166_n7505# x4.net9 1.52e-20
C2615 a_28596_n9259# x4._23_ 6.82e-19
C2616 a_28031_n8709# a_28895_n8893# 1.29e-19
C2617 a_28638_n8741# a_28470_n8893# 3.15e-19
C2618 a_28470_n8715# a_28638_n9147# 3.15e-19
C2619 x4.net11 x4.net7 2.47e-20
C2620 a_22962_n5131# x4.net2 0.010623f
C2621 a_25729_n8395# x4._18_ 9.76e-19
C2622 a_28638_n9147# a_29063_n8991# 1.28e-19
C2623 a_28197_n9259# a_28895_n8893# 0.194892f
C2624 a_27181_n8337# x4.net9 3.81e-19
C2625 a_25211_n9465# x4.net5 0.201023f
C2626 a_25875_n7395# x4.net6 8.38e-19
C2627 VDD a_26725_n8715# 0.004219f
C2628 x4.net2 a_23391_n4933# 0.019416f
C2629 x1.sky130_fd_sc_hd__inv_2_7.A enable_ring 1.67e-19
C2630 x1.sky130_fd_sc_hd__inv_2_9.A ring_out 0.025177f
C2631 x4._16_ a_25229_n10182# 3.59e-21
C2632 a_26309_n9259# a_26147_n9107# 0.004009f
C2633 a_24981_n8715# x4.net6 7.79e-20
C2634 a_17405_n2032# a_17857_n2290# 0.002207f
C2635 x3.x1.nSEL1 a_18585_n1958# 1.59e-19
C2636 x4.clknet_1_0__leaf_clk a_23417_n8715# 0.03291f
C2637 x4.counter[5] x4.net7 0.002945f
C2638 x4.counter[5] a_26885_n10182# 0.1107f
C2639 a_25823_n8395# a_25600_n8741# 0.011458f
C2640 VDD x4._17_ 2.38225f
C2641 x4.net8 x4._18_ 0.01511f
C2642 a_28385_n8715# x4.net10 6.3e-20
C2643 a_24595_n8741# x4._15_ 8.84e-19
C2644 x4.clknet_1_0__leaf_clk x4._02_ 0.254839f
C2645 x4.clknet_0_clk x4.clknet_1_1__leaf_clk 0.335671f
C2646 x4.net3 a_24229_n5073# 4.27e-20
C2647 x4._16_ a_25600_n8741# 0.01721f
C2648 a_24595_n9571# a_25211_n9465# 0.013543f
C2649 x4._19_ a_25449_n7261# 8.17e-20
C2650 x4.net6 x4._25_ 2.22e-20
C2651 a_23781_n8171# x4.clknet_1_0__leaf_clk 0.020113f
C2652 x1.sky130_fd_sc_hd__inv_2_12.A x3.x1.nSEL1 1.23e-19
C2653 a_26529_n7849# a_26559_n9259# 5.07e-21
C2654 a_26630_n8715# x4._05_ 6.05e-21
C2655 x4.net8 a_26191_n8709# 0.036074f
C2656 a_24479_n7805# x4.net5 4.89e-20
C2657 x4.net3 x4.net1 0.313425f
C2658 a_27507_n8893# x4.clknet_1_1__leaf_clk 1.62e-19
C2659 a_27166_n9147# x4._15_ 4.59e-21
C2660 a_28205_n9437# x4.net7 6.33e-20
C2661 x4.net4 a_23063_n8709# 0.007432f
C2662 counter7 x4.net11 1.31e-19
C2663 a_25779_n7395# x4.clknet_1_1__leaf_clk 1.77e-20
C2664 a_19061_n2032# select0 0.220366f
C2665 x4.net3 a_23339_n9259# 0.005671f
C2666 counter3 x4.counter[4] 0.07836f
C2667 x4._12_ a_24229_n5073# 0.023132f
C2668 a_24229_n4907# a_24075_n5995# 9.03e-20
C2669 VDD x4._23_ 1.70159f
C2670 a_28895_n8715# a_29103_n9829# 9.49e-21
C2671 counter3 a_25229_n10182# 0.110188f
C2672 x4._07_ a_26191_n8709# 0.022853f
C2673 a_26593_n7906# x4._05_ 2.43e-19
C2674 x4.net8 x4._24_ 1.23e-20
C2675 x4._16_ a_26998_n8893# 7.37e-22
C2676 a_24625_n8715# x4.clknet_1_1__leaf_clk 7.11e-20
C2677 VDD a_27805_n10182# 0.309637f
C2678 x4._22_ a_27175_n9437# 0.002279f
C2679 x4._16_ a_26816_n8171# 3.12e-19
C2680 x4._13_ x4.net3 0.031667f
C2681 a_28031_n8709# a_28031_n9259# 0.037572f
C2682 x4.net8 a_27591_n8991# 0.020836f
C2683 x4._12_ x4.net1 0.312817f
C2684 x1.sky130_fd_sc_hd__inv_2_17.A x1.sky130_fd_sc_hd__inv_2_16.A 0.173286f
C2685 a_23391_n5219# x4.net2 0.00144f
C2686 x4.counter[5] counter7 0.007023f
C2687 a_28031_n9259# a_28197_n9259# 0.970499f
C2688 x4.net8 a_25709_n7109# 0.001938f
C2689 a_26529_n7849# x4._06_ 0.003245f
C2690 x4._16_ a_23851_n9829# 0.184103f
C2691 x4.net2 a_22837_n10182# 0.223155f
C2692 x4.net2 a_23255_n4363# 0.107098f
C2693 a_27055_n8715# a_27181_n8337# 0.006169f
C2694 a_27194_n8171# a_28470_n8715# 0.01166f
C2695 x4._22_ x4._09_ 0.009594f
C2696 x4._07_ a_27591_n8991# 3.3e-20
C2697 drv_out x4._19_ 0.013619f
C2698 a_24479_n7805# a_24595_n9571# 3.06e-22
C2699 VDD a_23633_n4541# 0.005315f
C2700 a_26166_n7505# x4._22_ 8.56e-19
C2701 VDD a_26798_n8741# 0.185172f
C2702 x4.net3 x4.counter[1] 0.103986f
C2703 x4._19_ x4._15_ 6.2e-22
C2704 a_28647_n9483# x4._24_ 9.33e-19
C2705 x4.clknet_0_clk a_26117_n7627# 2.01e-19
C2706 x4._21_ a_26593_n7906# 1.69e-19
C2707 x4._04_ x4._18_ 0.003255f
C2708 a_23927_n8715# x4.net6 5.09e-19
C2709 x4.net3 a_23225_n7109# 0.011213f
C2710 x4._11_ a_26979_n9829# 2.67e-19
C2711 a_23882_n5174# x4._10_ 2.11e-19
C2712 x1.sky130_fd_sc_hd__inv_2_6.A enable_ring 5.64e-20
C2713 a_23229_n8709# a_23927_n8715# 0.196846f
C2714 a_23670_n8741# a_24095_n8741# 1.28e-19
C2715 x1.sky130_fd_sc_hd__inv_2_9.A x1.sky130_fd_sc_hd__nand2_2_0.B 0.163894f
C2716 a_23781_n8171# a_25900_n8197# 8.39e-21
C2717 a_28197_n8709# x4._25_ 1.11e-19
C2718 a_23927_n8715# a_24203_n8893# 5.06e-19
C2719 a_24595_n8741# a_24371_n8991# 0.002391f
C2720 a_27139_n8715# a_26798_n8741# 9.73e-19
C2721 x4.net9 a_26998_n8893# 0.003585f
C2722 x4._08_ a_28031_n8709# 0.097891f
C2723 x3.x2.GN2 x3.x2.GN4 8.82e-19
C2724 a_23505_n9259# x4.net5 8.3e-19
C2725 a_23946_n9147# a_23904_n9259# 4.62e-19
C2726 VDD a_26913_n9259# 0.079731f
C2727 VDD a_17857_n2290# 0.161536f
C2728 x4._08_ a_28197_n9259# 0.001269f
C2729 x4.net3 a_23295_n4755# 9.98e-20
C2730 a_24316_n9803# a_24220_n9483# 0.002032f
C2731 x4._12_ a_23225_n7109# 4.42e-19
C2732 a_23615_n8171# x4.net5 1.51e-20
C2733 a_24222_n8059# x4._16_ 1.01e-19
C2734 a_26725_n9259# x4.net6 0.045685f
C2735 select0 x3.x2.GP3 2.82e-19
C2736 x4.net10 x4._24_ 0.13484f
C2737 x3.nselect2 select0 1.88e-19
C2738 x4._08_ a_28979_n8715# 2.34e-19
C2739 VDD a_25211_n9465# 0.2419f
C2740 a_23391_n5219# a_23633_n5451# 0.008508f
C2741 a_23675_n5233# a_24229_n5073# 0.057611f
C2742 a_23811_n5073# a_23610_n5085# 4.67e-20
C2743 a_23682_n5329# a_24031_n5085# 2.36e-19
C2744 a_24054_n7805# x4.net8 4.11e-20
C2745 a_24647_n7903# a_24479_n7805# 0.310858f
C2746 ring_out x3.x2.GN4 0.080391f
C2747 x4.clknet_0_clk a_25779_n7395# 0.002548f
C2748 x4._14_ a_23946_n9147# 1.1e-19
C2749 x1.sky130_fd_sc_hd__inv_2_13.A x3.x1.nSEL1 2.53e-21
C2750 x4._09_ a_29103_n9829# 0.17213f
C2751 a_26630_n8715# x4.net7 0.034093f
C2752 x4._12_ a_23295_n4755# 6.08e-20
C2753 a_28725_n10182# x4._23_ 7.52e-20
C2754 x4.counter[1] x4.counter[2] 0.070133f
C2755 a_26630_n8715# a_26885_n10182# 3e-19
C2756 a_23675_n5233# x4.net1 0.002755f
C2757 x4.net8 x4._20_ 0.027217f
C2758 a_27805_n10182# a_28725_n10182# 1.37e-20
C2759 a_29133_n9803# a_28895_n8893# 3.93e-20
C2760 a_24647_n7903# a_25667_n8171# 3.28e-20
C2761 a_27271_n9437# x4._15_ 3.42e-21
C2762 x4._04_ x4._14_ 4.63e-22
C2763 a_24479_n7805# a_24605_n8171# 0.006169f
C2764 m3_18866_n4909# drv_out 0.132758f
C2765 x4.net8 x4._11_ 0.418201f
C2766 a_23851_n9829# a_23778_n8893# 3.53e-19
C2767 a_23994_n9687# a_23946_n9147# 5.83e-19
C2768 VDD a_24813_n8395# 0.001324f
C2769 a_17857_n2290# select1 0.03417f
C2770 a_23941_n3056# x4._00_ 4.57e-22
C2771 x4.net1 a_23505_n4043# 0.003019f
C2772 a_26593_n7906# x4.net7 1.85e-20
C2773 a_26147_n9107# x4.clknet_1_1__leaf_clk 0.050301f
C2774 x4.net9 a_27549_n9259# 0.001933f
C2775 x4._16_ x4._05_ 0.001611f
C2776 VDD x4.net11 0.794015f
C2777 x3.x2.GP1 x3.x2.GP3 0.001226f
C2778 x4._07_ x4._20_ 1.72e-19
C2779 a_26542_n7627# a_26713_n7249# 0.001229f
C2780 x4.clknet_1_0__leaf_clk a_23811_n5073# 0.024273f
C2781 x4.counter[8] a_29489_n9803# 1.28e-20
C2782 x4._11_ x4._07_ 0.161717f
C2783 a_26529_n7849# a_26159_n7409# 0.007926f
C2784 a_25834_n7921# a_26166_n7505# 0.002652f
C2785 a_27251_n7408# x4.net6 0.019537f
C2786 x1.sky130_fd_sc_hd__inv_2_17.Y x1.sky130_fd_sc_hd__inv_2_16.A 5.04e-19
C2787 a_26630_n8715# a_26357_n8709# 0.074815f
C2788 a_27223_n8741# a_26191_n8709# 0.048748f
C2789 a_26366_n7350# x4._15_ 1.61e-21
C2790 VDD a_28565_n8715# 0.002923f
C2791 a_23682_n4633# a_23941_n3056# 4.65e-23
C2792 a_23063_n8709# x4.net6 1.88e-19
C2793 x4._21_ a_25823_n8395# 4.25e-19
C2794 a_26559_n9259# x4.clknet_1_1__leaf_clk 0.319108f
C2795 x4.counter[5] VDD 0.450193f
C2796 x4.net10 a_28979_n8893# 3.08e-19
C2797 VDD a_24479_n7805# 0.169689f
C2798 a_28385_n8715# x4._15_ 0.007874f
C2799 a_23063_n8709# a_23229_n8709# 0.968904f
C2800 a_26295_n7249# x4._16_ 2.16e-20
C2801 a_26593_n7906# a_26357_n8709# 0.003413f
C2802 a_23927_n8715# a_23339_n9259# 0.002525f
C2803 x4.net3 a_23295_n5219# 0.115857f
C2804 a_23339_n9259# a_23693_n9259# 0.062224f
C2805 a_23882_n4933# x4.clknet_1_0__leaf_clk 0.040993f
C2806 a_23811_n4907# a_24229_n4907# 3.39e-19
C2807 x4.net4 a_25229_n10182# 0.003224f
C2808 x4._21_ x4._16_ 0.249175f
C2809 VDD a_25667_n8171# 0.004487f
C2810 a_23205_n10182# x4.counter[1] 0.1107f
C2811 a_27055_n8715# a_26998_n8893# 7.26e-19
C2812 enable_counter x4._00_ 2.67e-19
C2813 a_23675_n5233# a_23225_n7109# 6.92e-20
C2814 a_23781_n8171# a_24371_n8991# 8.13e-20
C2815 x4.net8 a_26725_n8715# 4.84e-19
C2816 counter7 a_29319_n10347# 3.7e-19
C2817 mux_out counter3 4.52136f
C2818 x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__nand2_2_0.B 5.04e-19
C2819 x4._06_ x4.clknet_1_1__leaf_clk 0.005269f
C2820 x4.net9 x4._05_ 1.93e-19
C2821 a_23295_n5219# x4._12_ 0.027335f
C2822 a_23615_n8171# a_24647_n7903# 0.048608f
C2823 x4._04_ a_24054_n7805# 0.01404f
C2824 a_26979_n9829# x4._23_ 2.79e-19
C2825 x4._22_ a_26998_n8893# 0.002895f
C2826 x4.net9 a_27377_n9437# 6.77e-19
C2827 a_27807_n9829# x4.net7 0.023542f
C2828 x4._22_ a_26816_n8171# 0.006962f
C2829 x3.x1.nSEL1 a_17579_n1926# 0.00175f
C2830 VDD a_28205_n9437# 1.16e-19
C2831 a_29063_n8741# x4.clknet_1_1__leaf_clk 9.45e-20
C2832 a_23391_n5219# a_23391_n4933# 0.015931f
C2833 x4._11_ a_23946_n9147# 0.004479f
C2834 a_28895_n8893# x4.clknet_1_1__leaf_clk 2.2e-19
C2835 x4.net10 x4._11_ 0.36244f
C2836 x4.net8 x4._17_ 0.172731f
C2837 enable_counter a_23682_n4633# 4.56e-21
C2838 x4.counter[4] a_25793_n9259# 4.17e-20
C2839 x4.net4 a_25600_n8741# 1.34e-19
C2840 m3_18862_n5953# counter3 0.119717f
C2841 x4.net3 a_23502_n8715# 8.21e-19
C2842 a_28551_n9803# x4._09_ 2.04e-21
C2843 a_23255_n4363# a_23391_n4933# 7.31e-19
C2844 x4.net4 a_24287_n8893# 8.77e-19
C2845 x4._00_ a_23505_n4363# 0.07841f
C2846 x4.clknet_1_0__leaf_clk x4._14_ 0.088295f
C2847 x4._04_ x4._11_ 0.257603f
C2848 a_28638_n8741# a_29063_n8741# 1.28e-19
C2849 a_28197_n8709# a_28895_n8715# 0.194892f
C2850 a_28579_n7627# x4._25_ 0.082413f
C2851 a_26295_n7249# x4.net9 0.004659f
C2852 x4._17_ x4._07_ 3.97e-20
C2853 a_28197_n8709# a_28385_n9259# 1.41e-20
C2854 a_28725_n10182# x4.net11 3.2e-20
C2855 a_25900_n8197# x4._18_ 7.58e-19
C2856 a_28638_n9147# a_28385_n9259# 3.39e-19
C2857 x4._09_ x4.net6 1.5e-20
C2858 x4._10_ a_24075_n5995# 0.423817f
C2859 a_23615_n5995# x4._11_ 0.005192f
C2860 x4._21_ x4.net9 0.170283f
C2861 VDD a_23505_n9259# 0.342267f
C2862 a_23682_n4633# a_23505_n4363# 0.001655f
C2863 VDD a_29021_n8337# 7.83e-19
C2864 a_26166_n7505# x4.net6 0.001918f
C2865 x4._18_ x4._15_ 0.045245f
C2866 a_26913_n9259# a_27093_n8893# 0.001229f
C2867 x4._16_ x4.net7 5.07e-19
C2868 x4._22_ a_27549_n9259# 7.63e-20
C2869 select0 x3.x2.GN2 0.114345f
C2870 VDD a_23615_n8171# 0.6434f
C2871 x3.x1.nSEL1 x3.x2.GN1 0.034862f
C2872 x4.net8 x4._23_ 0.011201f
C2873 a_28457_n9803# x4._24_ 0.085832f
C2874 a_17857_n2290# a_18033_n1958# 0.185422f
C2875 x4.clknet_0_clk a_26559_n9259# 1.17e-21
C2876 a_24769_n9465# x4.net5 0.002311f
C2877 x4.clknet_1_0__leaf_clk a_22885_n8715# 1.21e-20
C2878 x4.net8 a_27805_n10182# 0.2272f
C2879 x4.net4 a_23851_n9829# 0.021386f
C2880 a_23063_n8709# a_23339_n9259# 0.001876f
C2881 a_26545_n8715# a_26191_n8709# 0.057611f
C2882 a_24625_n8715# a_24095_n8741# 2.84e-19
C2883 a_24011_n8715# a_23927_n8715# 0.008508f
C2884 a_27807_n9829# a_27423_n8893# 0.009905f
C2885 x1.sky130_fd_sc_hd__inv_2_17.Y x1.sky130_fd_sc_hd__inv_2_17.A 0.173286f
C2886 a_26191_n8709# x4._15_ 0.034785f
C2887 x4._13_ a_23063_n8709# 3.88e-19
C2888 ring_out select0 3.69e-19
C2889 a_27223_n8741# x4._11_ 1.18e-19
C2890 x4._16_ a_26357_n8709# 9.89e-20
C2891 x4.net4 a_23628_n8337# 1.81e-19
C2892 a_23295_n5219# a_23675_n5233# 0.048748f
C2893 a_23421_n7921# a_23615_n8171# 5.05e-19
C2894 a_24054_n7805# x4.clknet_1_0__leaf_clk 0.002436f
C2895 x4._15_ x4._24_ 0.032103f
C2896 x3.x2.GN2 x3.x2.GP1 2.56189f
C2897 x4._16_ x4.net5 0.096932f
C2898 x4._19_ a_26515_n7261# 2.79e-19
C2899 x3.x2.GN3 x3.x2.GN4 0.071282f
C2900 x4.clknet_0_clk x4._06_ 2.8e-19
C2901 x4.net8 a_26798_n8741# 0.001066f
C2902 drv_out a_25709_n7109# 0.318051f
C2903 a_27194_n8171# a_26725_n9259# 1.98e-20
C2904 x4._11_ a_26457_n7849# 4.38e-19
C2905 a_23391_n5219# a_23255_n4363# 6.59e-20
C2906 a_26545_n8715# a_25709_n7109# 2.19e-20
C2907 a_26529_n7849# a_26375_n8171# 0.049785f
C2908 a_25900_n8197# a_25709_n7109# 3.15e-19
C2909 a_28647_n9483# x4._23_ 4.18e-19
C2910 a_28031_n9259# x4.clknet_1_1__leaf_clk 0.306202f
C2911 a_27591_n8991# x4._15_ 7.77e-19
C2912 x4._04_ x4._17_ 6.62e-21
C2913 a_24769_n9465# a_24595_n9571# 0.006584f
C2914 x4._14_ x4._15_ 1.65e-19
C2915 a_25709_n7109# x4._15_ 2.08e-20
C2916 a_26159_n7409# x4.clknet_1_1__leaf_clk 0.228247f
C2917 x4.clknet_1_0__leaf_clk x4._11_ 0.317456f
C2918 x4.net9 x4.net7 0.742565f
C2919 x4._07_ a_26798_n8741# 0.011124f
C2920 ring_out x3.x2.GP1 4.09516f
C2921 x1.sky130_fd_sc_hd__inv_2_7.Y x1.sky130_fd_sc_hd__inv_2_9.A 0.17253f
C2922 VDD a_26630_n8715# 0.255475f
C2923 x4._22_ x4._05_ 0.001519f
C2924 VDD a_29319_n10347# 0.293517f
C2925 a_25729_n8715# x4.clknet_1_1__leaf_clk 0.001857f
C2926 x4.counter[6] x4.net7 1.8e-19
C2927 x4._22_ a_27377_n9437# 0.002069f
C2928 x4.net4 a_24222_n8059# 0.034264f
C2929 a_23994_n9687# x4._15_ 4.86e-20
C2930 x4.counter[6] a_26885_n10182# 4.98e-19
C2931 a_28638_n8741# a_28031_n9259# 1.99e-20
C2932 x4.counter[4] x4.net6 0.003133f
C2933 a_23682_n5329# x4.net2 8.79e-19
C2934 x4._09_ a_28638_n9147# 0.039926f
C2935 a_28031_n9259# a_28470_n8893# 0.273138f
C2936 a_25229_n10182# x4.net6 3.58e-19
C2937 VDD a_26593_n7906# 0.129866f
C2938 x4.net4 a_24329_n9259# 0.00133f
C2939 x4._16_ a_24595_n9571# 0.01632f
C2940 x4._11_ a_25449_n7261# 1.46e-19
C2941 x4.net2 x4._00_ 0.002662f
C2942 x4.net10 x4._23_ 0.188811f
C2943 a_28031_n8709# a_28385_n8715# 0.062224f
C2944 a_23417_n8715# a_23597_n8715# 0.001229f
C2945 x4._07_ a_26913_n9259# 0.128255f
C2946 VDD a_24229_n4907# 0.080219f
C2947 a_28385_n8715# a_28197_n9259# 1.41e-20
C2948 x4.net8 a_25211_n9465# 9.57e-20
C2949 x4.net9 a_26357_n8709# 0.002182f
C2950 a_27194_n8171# a_28385_n9259# 1.26e-19
C2951 a_26529_n7849# x4._19_ 1.87e-20
C2952 x3.x1.nSEL0 a_17857_n2290# 0.03096f
C2953 counter3 x4.net5 0.082815f
C2954 x4._11_ a_24525_n5745# 0.002858f
C2955 x4._08_ x4.clknet_1_1__leaf_clk 0.00277f
C2956 a_29321_n9483# x4._24_ 5.3e-19
C2957 x4._21_ x4._22_ 2.96e-19
C2958 a_25600_n8741# x4.net6 0.050235f
C2959 a_27223_n8741# x4._17_ 4.35e-22
C2960 a_23682_n4633# x4.net2 4.89e-19
C2961 x4._11_ a_28457_n9803# 0.054652f
C2962 x4._01_ x4._10_ 0.002197f
C2963 x4._13_ a_24180_n8171# 2.65e-20
C2964 x4._11_ a_25721_n9259# 0.002312f
C2965 x4.net3 x4._12_ 0.271994f
C2966 x4.net9 a_27423_n8893# 0.031858f
C2967 x4._08_ a_28638_n8741# 0.047112f
C2968 x4._17_ a_26457_n7849# 4.44e-20
C2969 a_24203_n8893# a_24287_n8893# 0.008508f
C2970 a_23778_n8893# x4.net5 4.4e-19
C2971 counter3 counter7 3.44556f
C2972 counter7 x4.net9 0.006102f
C2973 x4.net6 a_28399_n7627# 2.84e-19
C2974 VDD a_18409_n2290# 0.179803f
C2975 m3_18866_n4909# x3.x2.GN1 6.03e-20
C2976 a_26295_n7249# a_26094_n7261# 4.67e-20
C2977 a_26366_n7350# a_26515_n7261# 0.005525f
C2978 x4.counter[6] a_27423_n8893# 2e-19
C2979 a_26166_n7505# a_26713_n7249# 0.095025f
C2980 a_28099_n9437# a_27807_n9829# 0.001675f
C2981 drv_out x4._11_ 1.2e-19
C2982 x4.counter[6] counter7 0.087745f
C2983 a_24647_n7903# x4._16_ 0.001048f
C2984 a_26998_n8893# x4.net6 6.05e-21
C2985 a_25900_n8197# x4._11_ 0.002559f
C2986 x4._20_ x4._15_ 0.093509f
C2987 x4.clknet_1_0__leaf_clk x4._17_ 3.38e-20
C2988 x4.net8 a_28565_n8715# 7.49e-20
C2989 counter3 a_24595_n9571# 8.56e-20
C2990 a_26816_n8171# x4.net6 0.001357f
C2991 x4._11_ x4._15_ 1.40124f
C2992 VDD a_27807_n9829# 0.419035f
C2993 a_23675_n5233# a_24058_n5451# 0.001632f
C2994 a_23682_n5329# a_23633_n5451# 4.04e-19
C2995 a_23882_n5174# a_24229_n5073# 0.037333f
C2996 a_23811_n5073# a_24031_n5085# 4.62e-19
C2997 a_24479_n7805# x4.net8 3.5e-19
C2998 x4.clknet_0_clk a_26159_n7409# 0.043419f
C2999 a_26147_n9107# a_26559_n9259# 0.020429f
C3000 x4._14_ a_24371_n8991# 1.14e-20
C3001 x3.x1.nSEL1 a_17985_n1898# 9.57e-19
C3002 x4._16_ a_24605_n8171# 4.87e-20
C3003 a_27055_n8715# x4.net7 0.054488f
C3004 x4.net3 x4.counter[2] 7.38e-19
C3005 VDD a_24769_n9465# 3.83e-21
C3006 a_23882_n5174# x4.net1 1.33e-19
C3007 x4._17_ a_25449_n7261# 7.93e-19
C3008 x4.net8 a_25667_n8171# 0.057781f
C3009 x4.counter[5] x4._07_ 1.62e-19
C3010 a_28003_n9437# x4._15_ 0.006963f
C3011 a_24595_n8741# x4.clknet_1_1__leaf_clk 1.5e-19
C3012 VDD a_25823_n8395# 2.25e-21
C3013 a_18409_n2290# select1 0.261734f
C3014 x4.net9 a_28596_n9259# 0.002793f
C3015 x4._22_ x4.net7 0.179589f
C3016 a_25779_n7395# a_26159_n7409# 0.048635f
C3017 x4._22_ a_26885_n10182# 8.8e-19
C3018 x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_9.A 5.04e-19
C3019 a_27194_n8171# x4._09_ 3.55e-20
C3020 a_25729_n8715# a_25779_n7395# 2.76e-21
C3021 x4._06_ a_26147_n9107# 2.49e-19
C3022 a_23628_n8337# a_23229_n8709# 8.12e-19
C3023 a_27055_n8715# a_26357_n8709# 0.192206f
C3024 a_27223_n8741# a_26798_n8741# 1.28e-19
C3025 a_28031_n8709# a_26191_n8709# 0.002059f
C3026 a_23417_n8715# a_23670_n8741# 3.39e-19
C3027 VDD x4._16_ 2.17996f
C3028 a_23882_n4933# a_23941_n3056# 2.02e-20
C3029 a_26545_n8715# a_26725_n8715# 0.001229f
C3030 a_23675_n4933# x4.net1 0.003904f
C3031 mux_out x3.x2.GP3 0.357364f
C3032 a_27166_n9147# x4.clknet_1_1__leaf_clk 0.046669f
C3033 a_25834_n7921# x4._21_ 0.128337f
C3034 a_26375_n8171# x4.clknet_1_1__leaf_clk 3.57e-20
C3035 x4.net10 x4.net11 0.310558f
C3036 select0 x3.x2.GN3 0.254198f
C3037 x4.net2 x4._02_ 0.035742f
C3038 x4._04_ a_24813_n8395# 0.002919f
C3039 a_23063_n8709# a_23502_n8715# 0.273138f
C3040 x4._02_ a_23670_n8741# 4.65e-19
C3041 x4._22_ a_26357_n8709# 0.015364f
C3042 a_28031_n8709# x4._24_ 0.031818f
C3043 x4.net7 a_26094_n7261# 0.001683f
C3044 x4.net3 a_23675_n5233# 0.008811f
C3045 a_24222_n8059# x4.net6 3.85e-19
C3046 x4._22_ x4.net5 4.26e-20
C3047 a_28197_n9259# x4._24_ 0.03707f
C3048 drv_out x4._17_ 1.68e-19
C3049 x4._09_ a_28579_n7627# 2.51e-21
C3050 a_24058_n4541# a_24229_n4907# 0.001229f
C3051 a_23633_n4541# x4.clknet_1_0__leaf_clk 7.44e-19
C3052 m3_18862_n5953# x3.x2.GP3 0.002824f
C3053 x4.net3 a_23205_n10182# 0.233128f
C3054 a_27055_n8715# a_27423_n8893# 3.78e-19
C3055 x4.net10 a_28565_n8715# 8.52e-20
C3056 a_25900_n8197# x4._17_ 0.062168f
C3057 a_23882_n5174# a_23225_n7109# 2.84e-19
C3058 a_28197_n9259# a_27591_n8991# 8.52e-19
C3059 a_24054_n7805# a_24371_n8991# 2.18e-19
C3060 x4._17_ x4._15_ 0.083602f
C3061 counter7 x4.counter[0] 0.003899f
C3062 a_28979_n8715# x4._24_ 8.56e-19
C3063 a_23615_n8171# x4.net8 9.67e-20
C3064 x4._04_ a_24479_n7805# 0.006456f
C3065 a_23675_n5233# x4._12_ 0.062549f
C3066 x4._22_ a_27423_n8893# 6.29e-19
C3067 a_28457_n9803# x4._23_ 0.04546f
C3068 a_24203_n8893# a_24329_n9259# 0.006169f
C3069 x3.x2.GN3 x3.x2.GP1 0.001426f
C3070 counter7 x4._22_ 1.31e-20
C3071 VDD a_28743_n9483# 4.51e-19
C3072 a_23682_n5329# a_23391_n4933# 1.53e-19
C3073 x4._11_ a_24371_n8991# 0.065594f
C3074 enable_counter a_23882_n4933# 1.46e-21
C3075 x4._05_ x4.net6 0.03493f
C3076 x4.clknet_1_1__leaf_clk x4._19_ 0.060342f
C3077 VDD counter3 2.4239f
C3078 VDD x4.net9 0.964697f
C3079 a_29489_n9803# x4._09_ 2.25e-19
C3080 x4.net3 a_23693_n9259# 7.76e-19
C3081 x4._00_ a_23391_n4933# 0.001635f
C3082 x4.net4 x4.net5 0.483177f
C3083 x4.counter[6] VDD 0.462317f
C3084 a_23851_n9829# a_23339_n9259# 2.64e-19
C3085 a_25179_n7627# a_25359_n7627# 0.185422f
C3086 x4.clknet_0_clk a_24595_n8741# 4.87e-21
C3087 a_26756_n8337# x4.net7 2.79e-19
C3088 a_25834_n7921# x4.net7 3.79e-19
C3089 x4._08_ a_28999_n7408# 0.109717f
C3090 a_28895_n8715# a_29063_n8991# 7.04e-19
C3091 a_29063_n8741# a_28895_n8893# 7.04e-19
C3092 x4._15_ x4._23_ 0.683594f
C3093 a_29645_n10182# x4.net11 0.003661f
C3094 a_28470_n8893# a_28565_n8893# 0.007724f
C3095 a_28197_n9259# a_28979_n8893# 6.32e-19
C3096 a_23205_n10182# x4.counter[2] 4.98e-19
C3097 VDD a_23778_n8893# 0.286549f
C3098 a_23682_n4633# a_23391_n4933# 0.194892f
C3099 a_23675_n4933# a_23295_n4755# 0.048748f
C3100 a_26295_n7249# x4.net6 0.001158f
C3101 x4.net4 counter7 6.88e-20
C3102 a_25359_n7627# a_25600_n8741# 6.83e-19
C3103 a_25793_n9259# x4.net5 1.04e-20
C3104 x1.sky130_fd_sc_hd__inv_2_7.A x1.sky130_fd_sc_hd__inv_2_7.Y 0.17253f
C3105 a_18033_n1958# a_18409_n2290# 3.02e-19
C3106 x4._21_ x4.net6 0.083542f
C3107 x4.clknet_0_clk a_27166_n9147# 8.09e-19
C3108 a_26159_n7409# a_26147_n9107# 8.37e-20
C3109 x4.net8 a_26630_n8715# 0.003635f
C3110 x4.clknet_1_0__leaf_clk a_24813_n8395# 1.8e-20
C3111 x4.net4 a_24595_n9571# 0.130038f
C3112 a_25729_n8715# a_24095_n8741# 2.67e-21
C3113 a_26545_n8715# a_26798_n8741# 3.39e-19
C3114 a_24625_n8715# a_24595_n8741# 0.025037f
C3115 a_26529_n7849# a_26191_n8709# 0.001396f
C3116 a_23505_n9259# a_23946_n9147# 0.127288f
C3117 x4._14_ a_24220_n9483# 0.122283f
C3118 a_26798_n8741# x4._15_ 0.03519f
C3119 VDD x4._10_ 0.249351f
C3120 a_24229_n5073# a_24075_n5995# 6.31e-19
C3121 x4.net8 a_26593_n7906# 0.003744f
C3122 a_26630_n8715# x4._07_ 0.002926f
C3123 a_23781_n8171# x4._03_ 3.92e-19
C3124 a_28031_n9259# a_26559_n9259# 0.003146f
C3125 a_27507_n8893# a_27166_n9147# 9.73e-19
C3126 a_28031_n8709# x4._11_ 3.54e-20
C3127 a_26159_n7409# a_26559_n9259# 2.6e-21
C3128 a_27194_n8171# a_28399_n7627# 0.010673f
C3129 x4._11_ a_28197_n9259# 7.13e-19
C3130 a_23994_n9687# a_24220_n9483# 0.005961f
C3131 x4.net4 a_24053_n8337# 3.33e-19
C3132 a_23391_n5219# a_23682_n5329# 0.192341f
C3133 a_23615_n8171# x4._04_ 0.09532f
C3134 a_24479_n7805# x4.clknet_1_0__leaf_clk 6.75e-21
C3135 x4._19_ a_26117_n7627# 1.83e-19
C3136 x4.net1 a_24075_n5995# 4.64e-19
C3137 a_26593_n7906# x4._07_ 0.001092f
C3138 a_29321_n9483# x4._23_ 3.52e-19
C3139 a_26529_n7849# a_25709_n7109# 6.61e-19
C3140 a_26913_n9259# x4._15_ 7.24e-21
C3141 x4.net3 a_23063_n8709# 0.023332f
C3142 a_26366_n7350# x4.clknet_1_1__leaf_clk 4.65e-20
C3143 a_23255_n4363# x4._00_ 0.167554f
C3144 VDD a_22879_n5451# 0.229121f
C3145 x4.clknet_0_clk x4._19_ 0.038005f
C3146 mux_out x3.x2.GN2 0.42933f
C3147 VDD a_27055_n8715# 0.182006f
C3148 x4.net9 a_28725_n10182# 0.202772f
C3149 VDD x4.counter[0] 0.524238f
C3150 a_28385_n8715# x4.clknet_1_1__leaf_clk 3.58e-19
C3151 x4.net11 a_28457_n9803# 2.78e-19
C3152 a_28399_n7627# a_28579_n7627# 0.185422f
C3153 x4.net4 a_24647_n7903# 7.5e-19
C3154 x4._22_ a_28099_n9437# 6.12e-20
C3155 a_26159_n7409# x4._06_ 0.002324f
C3156 x3.x1.nSEL1 a_18537_n1898# 4.08e-19
C3157 a_25211_n9465# x4._15_ 0.110742f
C3158 x4.net6 a_27755_n7261# 0.157729f
C3159 a_23682_n4633# a_23391_n5219# 1.53e-19
C3160 x4.net6 x4.net7 0.905861f
C3161 a_23811_n5073# x4.net2 8.2e-21
C3162 x4._09_ a_29063_n8991# 0.010518f
C3163 a_28031_n9259# a_28895_n8893# 0.032244f
C3164 a_26885_n10182# x4.net6 0.013611f
C3165 m3_18862_n5953# x3.x2.GN2 0.016745f
C3166 VDD x4._22_ 0.56354f
C3167 a_25729_n8715# x4._06_ 2.02e-19
C3168 a_23682_n4633# a_23255_n4363# 0.00324f
C3169 ring_out mux_out 4.51997f
C3170 a_25779_n7395# x4._19_ 0.065395f
C3171 x4.counter[4] a_25639_n9259# 2.6e-19
C3172 a_28638_n8741# a_28385_n8715# 3.39e-19
C3173 a_27055_n8715# a_27139_n8715# 0.008508f
C3174 x4.net8 a_27807_n9829# 0.004343f
C3175 x4.net10 a_29319_n10347# 1.3e-21
C3176 a_24054_n7805# a_24220_n9483# 4.44e-21
C3177 x3.x2.GP3 counter7 0.165274f
C3178 a_24813_n8395# x4._15_ 1.54e-19
C3179 x3.x1.nSEL0 a_18409_n2290# 1.91e-20
C3180 x4._18_ a_25211_n9231# 1.7e-19
C3181 x4._05_ a_26713_n7249# 0.114695f
C3182 x4.net11 x4._15_ 1.7e-19
C3183 a_24981_n8715# a_23063_n8709# 4.04e-20
C3184 x4._11_ a_23769_n5995# 2.12e-19
C3185 a_25729_n8395# x4._16_ 0.001343f
C3186 a_26357_n8709# x4.net6 0.048602f
C3187 a_23882_n4933# x4.net2 1.88e-19
C3188 x4._11_ a_24220_n9483# 9.44e-19
C3189 x4.net5 x4.net6 0.003368f
C3190 x4.clknet_1_0__leaf_clk a_23505_n9259# 0.021572f
C3191 VDD a_26094_n7261# 7.65e-20
C3192 select0 x3.x2.GN4 0.218716f
C3193 a_24095_n8741# a_24595_n8741# 0.016344f
C3194 a_24647_n7903# a_25834_n7921# 1.25e-19
C3195 a_23781_n8171# a_23969_n8171# 0.095025f
C3196 VDD x4.net4 1.18326f
C3197 a_25600_n8741# a_25639_n9259# 2.2e-19
C3198 x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_7.Y 5.04e-19
C3199 x4._11_ a_26309_n9259# 0.001677f
C3200 x4._08_ a_29063_n8741# 0.004928f
C3201 a_24203_n8893# x4.net5 0.019334f
C3202 a_23615_n8171# x4.clknet_1_0__leaf_clk 0.245743f
C3203 a_27251_n7408# x4._25_ 6.03e-21
C3204 x4._08_ a_28895_n8893# 3.02e-19
C3205 VDD a_19061_n2032# 0.217593f
C3206 a_26295_n7249# a_26713_n7249# 3.39e-19
C3207 VDD a_23697_n5995# 2.01e-19
C3208 a_25900_n8197# a_25667_n8171# 0.005961f
C3209 a_23597_n8715# x4._11_ 3.45e-19
C3210 a_27423_n8893# x4.net6 4.38e-19
C3211 x4.net8 x4._16_ 0.193029f
C3212 a_26529_n7849# x4._11_ 0.042839f
C3213 x4.net9 a_26979_n9829# 0.125008f
C3214 a_25667_n8171# x4._15_ 9.44e-19
C3215 counter7 x4.net6 6.88e-20
C3216 x4._18_ x4.clknet_1_1__leaf_clk 3.06e-19
C3217 a_25359_n7627# x4._05_ 4.91e-20
C3218 VDD a_29103_n9829# 0.230416f
C3219 a_23811_n5073# a_23633_n5451# 9.73e-19
C3220 a_23882_n5174# a_24058_n5451# 0.007724f
C3221 x4._01_ a_24229_n5073# 0.121379f
C3222 x4.net2 x4._14_ 0.45134f
C3223 x4._14_ a_23670_n8741# 8.48e-21
C3224 x4.clknet_0_clk a_26366_n7350# 0.004436f
C3225 x3.x2.GN4 x3.x2.GP1 8.08e-19
C3226 a_28031_n8709# x4._23_ 0.029216f
C3227 x1.sky130_fd_sc_hd__inv_2_13.A a_17857_n2290# 2.51e-19
C3228 VDD a_23337_n4363# 0.008578f
C3229 a_28197_n8709# x4.net7 2.99e-20
C3230 a_27194_n8171# x4._05_ 0.003024f
C3231 VDD enable_ring 0.618517f
C3232 VDD a_25793_n9259# 3.08e-19
C3233 x4._16_ x4._07_ 0.003808f
C3234 a_24595_n9571# x4.net6 5.34e-20
C3235 a_28197_n9259# x4._23_ 0.031117f
C3236 m3_18866_n4909# x3.x2.GP2 0.004119f
C3237 a_28638_n9147# x4.net7 1.23e-19
C3238 x4._01_ x4.net1 1.96e-19
C3239 a_29319_n10347# a_29645_n10182# 0.024477f
C3240 a_29321_n9483# x4.net11 0.001149f
C3241 a_28205_n9437# x4._15_ 0.002119f
C3242 a_26191_n8709# x4.clknet_1_1__leaf_clk 0.670964f
C3243 a_24595_n9571# a_24203_n8893# 0.001309f
C3244 x4.net10 a_27807_n9829# 0.158335f
C3245 VDD a_26756_n8337# 0.001185f
C3246 a_19061_n2032# select1 0.125445f
C3247 VDD a_25834_n7921# 0.316019f
C3248 a_25875_n7395# a_26166_n7505# 0.192261f
C3249 a_27925_n7261# x4._11_ 0.001703f
C3250 a_26559_n9259# a_27166_n9147# 0.141453f
C3251 x4._22_ a_28725_n10182# 1.85e-19
C3252 x4._06_ a_24595_n8741# 1.6e-20
C3253 x4._05_ a_28579_n7627# 4.21e-20
C3254 x4.clknet_1_1__leaf_clk x4._24_ 0.041474f
C3255 x4.net2 a_22885_n8715# 0.002977f
C3256 a_23628_n8337# a_23502_n8715# 0.005525f
C3257 a_28197_n8709# a_26357_n8709# 0.001861f
C3258 x4.counter[9] counter7 2.14e-19
C3259 a_23811_n4907# x4.net1 0.002441f
C3260 x4.net8 x4.net9 0.748324f
C3261 a_27591_n8991# x4.clknet_1_1__leaf_clk 0.084941f
C3262 a_27194_n8171# x4._21_ 3.33e-20
C3263 a_25709_n7109# x4.clknet_1_1__leaf_clk 0.002451f
C3264 a_26147_n9107# x4._19_ 4.85e-22
C3265 a_29021_n8337# x4._15_ 6.51e-20
C3266 x4.counter[6] x4.net8 0.079257f
C3267 x4._02_ a_24095_n8741# 1.8e-19
C3268 a_23063_n8709# a_23927_n8715# 0.032244f
C3269 a_23615_n8171# a_25900_n8197# 1.55e-21
C3270 a_28638_n8741# x4._24_ 0.015657f
C3271 x1.sky130_fd_sc_hd__inv_2_11.A a_18409_n2290# 2.51e-19
C3272 x4.net3 a_23882_n5174# 3.02e-19
C3273 x4.net7 a_26713_n7249# 0.019182f
C3274 a_24647_n7903# x4.net6 0.129987f
C3275 a_28470_n8893# x4._24_ 0.010089f
C3276 x4._03_ a_23904_n9259# 0.001074f
C3277 a_23339_n9259# x4.net5 8.46e-19
C3278 a_24229_n4907# x4.clknet_1_0__leaf_clk 0.012004f
C3279 x4._06_ a_26375_n8171# 0.046896f
C3280 x4._16_ a_23946_n9147# 0.005579f
C3281 x4.net9 x4._07_ 0.03749f
C3282 VDD x3.x2.GP3 1.79155f
C3283 x4._08_ a_28031_n9259# 1.13e-19
C3284 VDD x3.nselect2 1.23654f
C3285 a_26529_n7849# x4._17_ 7.49e-19
C3286 a_23781_n8171# a_24095_n8741# 0.003783f
C3287 x4._01_ a_23225_n7109# 3.77e-19
C3288 x4._04_ x4._16_ 0.025302f
C3289 counter7 a_28638_n9147# 1.4e-19
C3290 a_24605_n8171# x4.net6 5.88e-19
C3291 a_23882_n5174# x4._12_ 0.032034f
C3292 x1.sky130_fd_sc_hd__inv_2_6.A x1.sky130_fd_sc_hd__inv_2_7.A 0.17253f
C3293 x4.clknet_0_clk x4._18_ 0.002702f
C3294 a_27055_n8715# a_26979_n9829# 3.32e-21
C3295 x4.net2 x4._11_ 0.001125f
C3296 a_25211_n9231# x4._20_ 3.41e-19
C3297 a_17405_n2032# x3.x2.GN2 0.039612f
C3298 x4._11_ a_23670_n8741# 0.005658f
C3299 VDD a_28551_n9803# 0.191262f
C3300 x4._14_ x4._03_ 0.071143f
C3301 a_28895_n8893# a_29021_n9259# 0.006169f
C3302 a_23811_n4907# a_23610_n4907# 4.67e-20
C3303 a_23882_n4933# a_24031_n4907# 0.005525f
C3304 x4._11_ a_25211_n9231# 0.163973f
C3305 a_26357_n8709# a_26713_n7249# 1.11e-20
C3306 a_25359_n7627# x4.net7 0.002934f
C3307 x4._22_ a_26979_n9829# 0.106132f
C3308 select1 x3.x2.GP3 0.003259f
C3309 a_23994_n9687# x4._03_ 0.005187f
C3310 mux_out x3.x2.GN3 0.429944f
C3311 x3.nselect2 select1 0.001177f
C3312 x4._18_ a_25779_n7395# 0.006776f
C3313 a_26630_n8715# a_26545_n8715# 0.037333f
C3314 x4._06_ x4._19_ 7.42e-21
C3315 x4.clknet_0_clk a_26191_n8709# 0.009291f
C3316 a_27194_n8171# a_27755_n7261# 0.010774f
C3317 a_27194_n8171# x4.net7 0.037674f
C3318 VDD x4.net6 3.11824f
C3319 a_19207_65# enable_ring 0.040112f
C3320 x4.net10 a_28743_n9483# 0.002966f
C3321 a_23675_n4933# x4._12_ 2.52e-19
C3322 a_26630_n8715# x4._15_ 0.026278f
C3323 a_24625_n8715# x4._18_ 4.57e-20
C3324 VDD a_23229_n8709# 0.341027f
C3325 a_28197_n9259# x4.net11 2.58e-19
C3326 a_28638_n9147# a_28596_n9259# 4.62e-19
C3327 x4.net10 x4.net9 0.022804f
C3328 m3_18862_n5953# x3.x2.GN3 0.087318f
C3329 VDD a_24203_n8893# 0.183311f
C3330 a_23811_n4907# a_23295_n4755# 1.28e-19
C3331 a_26545_n8715# a_26593_n7906# 1.39e-19
C3332 counter7 x4.counter[1] 0.003115f
C3333 mux_out VSS 13.574714f
C3334 enable_counter VSS 2.79528f
C3335 select1 VSS 7.705475f
C3336 select0 VSS 7.106359f
C3337 enable_ring VSS 1.66173f
C3338 VDD VSS 0.459367p
C3339 m3_18876_n6983# VSS 0.075151f $ **FLOATING
C3340 m3_18862_n5953# VSS 0.073094f $ **FLOATING
C3341 m3_18866_n4909# VSS 0.148749f $ **FLOATING
C3342 m2_17442_n2443# VSS 0.070212f $ **FLOATING
C3343 x4.counter[8] VSS 0.58641f
C3344 x4.counter[9] VSS 0.871549f
C3345 x4.counter[6] VSS 0.660698f
C3346 x4.counter[5] VSS 0.63746f
C3347 x4.counter[4] VSS 0.792045f
C3348 x4.counter[2] VSS 0.607552f
C3349 x4.counter[1] VSS 0.592623f
C3350 x4.counter[0] VSS 0.939839f
C3351 a_29645_n10182# VSS 0.269609f
C3352 a_29319_n10347# VSS 0.257101f
C3353 a_28725_n10182# VSS 0.296141f
C3354 a_27805_n10182# VSS 0.269288f
C3355 a_26885_n10182# VSS 0.278393f
C3356 a_25965_n10182# VSS 0.327843f
C3357 a_25229_n10182# VSS 0.269041f
C3358 a_24125_n10182# VSS 0.276333f
C3359 a_23205_n10182# VSS 0.316834f
C3360 a_22837_n10182# VSS 0.25238f
C3361 a_29489_n9803# VSS 8.84e-19
C3362 a_29133_n9803# VSS 0.004608f
C3363 a_28551_n9803# VSS 0.01879f
C3364 a_29321_n9483# VSS 0.005268f
C3365 a_28743_n9483# VSS 0.00969f
C3366 a_28647_n9483# VSS 0.006323f
C3367 a_28205_n9437# VSS 0.001553f
C3368 a_28099_n9437# VSS 0.003693f
C3369 a_28003_n9437# VSS 0.003656f
C3370 a_27377_n9437# VSS 0.003203f
C3371 a_27271_n9437# VSS 0.005457f
C3372 a_27175_n9437# VSS 0.005167f
C3373 a_24316_n9803# VSS 0.001114f
C3374 a_25297_n9465# VSS 0.004685f
C3375 a_24769_n9465# VSS 0.007506f
C3376 a_24220_n9483# VSS 0.183329f
C3377 a_29103_n9829# VSS 0.363777f
C3378 a_28457_n9803# VSS 0.343017f
C3379 a_27807_n9829# VSS 0.260798f
C3380 a_26979_n9829# VSS 0.294745f
C3381 a_25211_n9465# VSS 0.255389f
C3382 a_24595_n9571# VSS 0.284107f
C3383 a_23994_n9687# VSS 0.207092f
C3384 a_23851_n9829# VSS 0.20644f
C3385 a_29021_n9259# VSS 0.004786f
C3386 x4.net11 VSS 0.755509f
C3387 a_28596_n9259# VSS 0.009087f
C3388 a_28979_n8893# VSS 3.75e-19
C3389 a_27549_n9259# VSS 0.004164f
C3390 a_28565_n8893# VSS 0.002645f
C3391 a_28385_n9259# VSS 0.063765f
C3392 a_28895_n8893# VSS 0.268634f
C3393 a_29063_n8991# VSS 0.376509f
C3394 a_28470_n8893# VSS 0.227724f
C3395 a_28638_n9147# VSS 0.257495f
C3396 a_28197_n9259# VSS 0.334487f
C3397 x4._09_ VSS 0.540883f
C3398 a_28031_n9259# VSS 0.496464f
C3399 a_27124_n9259# VSS 0.008691f
C3400 a_27507_n8893# VSS 2.5e-19
C3401 a_26381_n9259# VSS 7.68e-19
C3402 a_26309_n9259# VSS 0.002515f
C3403 a_25793_n9259# VSS 0.002664f
C3404 a_25721_n9259# VSS 7.95e-19
C3405 a_27093_n8893# VSS 7.5e-19
C3406 a_26913_n9259# VSS 0.062716f
C3407 a_27423_n8893# VSS 0.275541f
C3408 a_27591_n8991# VSS 0.356576f
C3409 a_26998_n8893# VSS 0.218254f
C3410 a_27166_n9147# VSS 0.278138f
C3411 a_26725_n9259# VSS 0.323857f
C3412 a_26559_n9259# VSS 0.485385f
C3413 a_25297_n9231# VSS 0.004685f
C3414 x4._20_ VSS 0.296302f
C3415 a_24329_n9259# VSS 0.004794f
C3416 x4.net5 VSS 1.52232f
C3417 a_23904_n9259# VSS 0.007478f
C3418 a_24287_n8893# VSS 3.28e-19
C3419 a_23693_n9259# VSS 0.069011f
C3420 a_26147_n9107# VSS 0.233023f
C3421 a_25639_n9259# VSS 0.25233f
C3422 a_25211_n9231# VSS 0.250617f
C3423 a_24203_n8893# VSS 0.29125f
C3424 a_24371_n8991# VSS 0.405228f
C3425 a_23778_n8893# VSS 0.210325f
C3426 a_23946_n9147# VSS 0.255348f
C3427 a_23505_n9259# VSS 0.417108f
C3428 x4._03_ VSS 0.578555f
C3429 a_23339_n9259# VSS 0.557931f
C3430 a_28979_n8715# VSS 0.001033f
C3431 a_28565_n8715# VSS 0.002645f
C3432 x4.net10 VSS 1.52118f
C3433 a_29021_n8337# VSS 0.005282f
C3434 a_27139_n8715# VSS 0.002002f
C3435 a_28596_n8337# VSS 0.010952f
C3436 a_28385_n8715# VSS 0.070151f
C3437 a_27181_n8337# VSS 0.005844f
C3438 a_25729_n8715# VSS 0.014804f
C3439 a_24981_n8715# VSS 0.001519f
C3440 a_24625_n8715# VSS 0.026188f
C3441 a_24011_n8715# VSS 4.07e-19
C3442 a_23597_n8715# VSS 6.93e-19
C3443 a_26756_n8337# VSS 0.006941f
C3444 a_26545_n8715# VSS 0.060618f
C3445 a_25823_n8395# VSS 0.006538f
C3446 a_25729_n8395# VSS 0.008165f
C3447 a_24813_n8395# VSS 0.007253f
C3448 a_24053_n8337# VSS 0.004473f
C3449 a_22885_n8715# VSS 4.64e-19
C3450 a_23628_n8337# VSS 0.008558f
C3451 a_23417_n8715# VSS 0.080622f
C3452 a_28895_n8715# VSS 0.275172f
C3453 a_29063_n8741# VSS 0.371259f
C3454 a_28470_n8715# VSS 0.237292f
C3455 a_28638_n8741# VSS 0.266551f
C3456 a_28197_n8709# VSS 0.344626f
C3457 a_28031_n8709# VSS 0.532322f
C3458 a_27055_n8715# VSS 0.288597f
C3459 a_27223_n8741# VSS 0.391747f
C3460 a_26630_n8715# VSS 0.200127f
C3461 a_26798_n8741# VSS 0.247676f
C3462 a_26357_n8709# VSS 0.312142f
C3463 a_26191_n8709# VSS 0.480598f
C3464 a_25600_n8741# VSS 0.352433f
C3465 a_24595_n8741# VSS 0.430766f
C3466 a_23927_n8715# VSS 0.280567f
C3467 a_24095_n8741# VSS 0.367396f
C3468 a_23502_n8715# VSS 0.214988f
C3469 a_23670_n8741# VSS 0.263107f
C3470 a_23229_n8709# VSS 0.41156f
C3471 x4._02_ VSS 0.384112f
C3472 a_23063_n8709# VSS 0.551857f
C3473 x4._14_ VSS 1.2474f
C3474 a_26816_n8171# VSS 0.004249f
C3475 a_26375_n8171# VSS 0.154917f
C3476 x4._07_ VSS 0.467795f
C3477 a_25667_n8171# VSS 0.204157f
C3478 a_24605_n8171# VSS 0.00681f
C3479 x4._16_ VSS 2.102403f
C3480 x4._22_ VSS 1.56987f
C3481 a_26457_n7849# VSS 8.25e-20
C3482 a_26593_n7906# VSS 0.189132f
C3483 x4.net9 VSS 1.97499f
C3484 x4._06_ VSS 0.355082f
C3485 x4._21_ VSS 0.491639f
C3486 a_25762_n7921# VSS 9.9e-19
C3487 a_24180_n8171# VSS 0.007439f
C3488 a_24563_n7805# VSS 0.002478f
C3489 a_24149_n7805# VSS 5.31e-19
C3490 a_23969_n8171# VSS 0.062654f
C3491 a_27194_n8171# VSS 2.07482f
C3492 a_26529_n7849# VSS 0.166512f
C3493 a_25834_n7921# VSS 0.208373f
C3494 a_25900_n8197# VSS 0.228425f
C3495 x4.net8 VSS 1.78641f
C3496 a_24479_n7805# VSS 0.331871f
C3497 a_24647_n7903# VSS 0.427232f
C3498 a_24054_n7805# VSS 0.220057f
C3499 a_24222_n8059# VSS 0.267836f
C3500 a_23781_n8171# VSS 0.384412f
C3501 x4._04_ VSS 0.647447f
C3502 a_23615_n8171# VSS 0.561386f
C3503 a_23421_n7921# VSS 0.005123f
C3504 x4._13_ VSS 1.13412f
C3505 x4.net4 VSS 1.31635f
C3506 x4._08_ VSS 0.727548f
C3507 a_28669_n7261# VSS 0.00819f
C3508 a_28031_n7261# VSS 0.003851f
C3509 a_27925_n7261# VSS 0.003674f
C3510 a_27837_n7261# VSS 0.001688f
C3511 a_26117_n7627# VSS 7.93e-19
C3512 a_26713_n7249# VSS 0.060853f
C3513 a_26515_n7261# VSS 0.006624f
C3514 a_26094_n7261# VSS 0.005539f
C3515 a_25449_n7261# VSS 0.005238f
C3516 x4._25_ VSS 0.366822f
C3517 a_28999_n7408# VSS 0.272105f
C3518 a_28579_n7627# VSS 0.262291f
C3519 x4._24_ VSS 0.696921f
C3520 a_28399_n7627# VSS 0.271218f
C3521 x4._23_ VSS 0.973323f
C3522 a_27755_n7261# VSS 0.264312f
C3523 x4._15_ VSS 3.54853f
C3524 x4.net7 VSS 2.72071f
C3525 x4.net6 VSS 3.218643f
C3526 x4._19_ VSS 0.32708f
C3527 a_27251_n7408# VSS 0.252712f
C3528 x4.clknet_1_1__leaf_clk VSS 3.414301f
C3529 x4._05_ VSS 0.318608f
C3530 a_26295_n7249# VSS 0.241882f
C3531 a_26366_n7350# VSS 0.198121f
C3532 a_26166_n7505# VSS 0.303545f
C3533 a_26159_n7409# VSS 0.46613f
C3534 a_25875_n7395# VSS 0.281525f
C3535 a_25779_n7395# VSS 0.378965f
C3536 a_25359_n7627# VSS 0.234926f
C3537 x4._18_ VSS 0.468402f
C3538 a_25179_n7627# VSS 0.254342f
C3539 x4._17_ VSS 0.622186f
C3540 counter7 VSS 17.74957f
C3541 a_25709_n7109# VSS 2.29287f
C3542 x4.clknet_0_clk VSS 4.193551f
C3543 a_23225_n7109# VSS 2.29289f
C3544 a_23769_n5995# VSS 0.002457f
C3545 a_23697_n5995# VSS 0.001303f
C3546 a_24525_n5745# VSS 0.005104f
C3547 counter3 VSS 14.305035f
C3548 x4._11_ VSS 5.669386f
C3549 a_24075_n5995# VSS 0.298451f
C3550 x4._10_ VSS 0.339714f
C3551 a_23615_n5995# VSS 0.252154f
C3552 a_23633_n5451# VSS 6.89e-19
C3553 a_24229_n5073# VSS 0.064411f
C3554 a_24031_n5085# VSS 0.006624f
C3555 a_22879_n5451# VSS 0.017559f
C3556 a_23610_n5085# VSS 0.004183f
C3557 x4._12_ VSS 1.2616f
C3558 a_22962_n5131# VSS 0.004429f
C3559 x4._01_ VSS 0.405148f
C3560 a_23811_n5073# VSS 0.238144f
C3561 a_23882_n5174# VSS 0.195482f
C3562 a_23682_n5329# VSS 0.31379f
C3563 a_23675_n5233# VSS 0.552106f
C3564 a_23391_n5219# VSS 0.279727f
C3565 a_23295_n5219# VSS 0.390267f
C3566 x4.net3 VSS 2.298238f
C3567 a_24031_n4907# VSS 0.007478f
C3568 a_23610_n4907# VSS 0.004654f
C3569 x4.clknet_1_0__leaf_clk VSS 4.010709f
C3570 a_24229_n4907# VSS 0.069779f
C3571 a_23633_n4541# VSS 6.84e-19
C3572 a_23811_n4907# VSS 0.264386f
C3573 a_23882_n4933# VSS 0.210923f
C3574 a_23675_n4933# VSS 0.580201f
C3575 a_23682_n4633# VSS 0.340144f
C3576 a_23391_n4933# VSS 0.287469f
C3577 a_23295_n4755# VSS 0.412387f
C3578 a_23505_n4363# VSS 0.013142f
C3579 a_23337_n4363# VSS 0.006974f
C3580 x4._00_ VSS 0.757573f
C3581 a_23505_n4043# VSS 0.006222f
C3582 a_23255_n4363# VSS 0.393994f
C3583 x4.net2 VSS 3.500251f
C3584 x4.net1 VSS 1.81106f
C3585 a_23941_n3056# VSS 0.293097f
C3586 x3.x2.GP3 VSS 1.64575f
C3587 x3.x2.GP2 VSS 5.54164f
C3588 x3.x2.GP1 VSS 4.63625f
C3589 a_19235_n1926# VSS 0.006782f
C3590 x3.x2.GN4 VSS 3.79271f
C3591 a_18537_n1898# VSS 0.007327f
C3592 x3.x2.GN3 VSS 3.64172f
C3593 a_17985_n1898# VSS 0.004704f
C3594 x3.x2.GN2 VSS 3.91967f
C3595 a_17579_n1926# VSS 0.006793f
C3596 x3.x2.GN1 VSS 4.84443f
C3597 a_19061_n2032# VSS 0.3167f
C3598 a_18585_n1958# VSS 0.251626f
C3599 a_18409_n2290# VSS 0.236732f
C3600 a_18033_n1958# VSS 0.236633f
C3601 a_17857_n2290# VSS 0.222621f
C3602 a_17405_n2032# VSS 0.270062f
C3603 x3.nselect2 VSS 0.455447f
C3604 x3.x1.nSEL1 VSS 0.740163f
C3605 x3.x1.nSEL0 VSS 0.685116f
C3606 x1.sky130_fd_sc_hd__inv_2_11.A VSS 0.505562f
C3607 x1.sky130_fd_sc_hd__inv_2_12.A VSS 0.498424f
C3608 x1.sky130_fd_sc_hd__inv_2_13.A VSS 0.498285f
C3609 x1.sky130_fd_sc_hd__inv_2_14.A VSS 0.499488f
C3610 x1.sky130_fd_sc_hd__inv_2_15.A VSS 0.500758f
C3611 x1.sky130_fd_sc_hd__inv_2_16.A VSS 0.50136f
C3612 x1.sky130_fd_sc_hd__inv_2_17.A VSS 0.501617f
C3613 x1.sky130_fd_sc_hd__inv_2_17.Y VSS 0.52312f
C3614 drv_out VSS 29.368395f
C3615 a_19207_65# VSS 0.332619f
C3616 ring_out VSS 16.291151f
C3617 x1.sky130_fd_sc_hd__nand2_2_0.B VSS 0.632983f
C3618 x1.sky130_fd_sc_hd__inv_2_9.A VSS 0.508122f
C3619 x1.sky130_fd_sc_hd__inv_2_7.Y VSS 0.498331f
C3620 x1.sky130_fd_sc_hd__inv_2_7.A VSS 0.498331f
C3621 x1.sky130_fd_sc_hd__inv_2_6.A VSS 0.498339f
C3622 x1.sky130_fd_sc_hd__inv_2_5.A VSS 0.498632f
C3623 x1.sky130_fd_sc_hd__inv_2_4.A VSS 0.498682f
C3624 x1.sky130_fd_sc_hd__inv_2_3.A VSS 0.498707f
C3625 x1.sky130_fd_sc_hd__inv_2_2.A VSS 0.507755f
C3626 x1.sky130_fd_sc_hd__inv_2_8.Y VSS 0.971227f
C3627 x3.x2.GP1.t3 VSS 0.012908f
C3628 x3.x2.GP1.t2 VSS 0.012908f
C3629 x3.x2.GP1.n0 VSS 0.028358f
C3630 x3.x2.GP1.n1 VSS 0.018329f
C3631 x3.x2.GP1.t5 VSS 0.653268f
C3632 x3.x2.GP1.t4 VSS 0.671486f
C3633 x3.x2.GP1.n2 VSS 2.37213f
C3634 x3.x2.GP1.t1 VSS 0.019859f
C3635 x3.x2.GP1.t0 VSS 0.019859f
C3636 x3.x2.GP1.n3 VSS 0.04092f
C3637 x3.x2.GP1.n4 VSS 0.100085f
C3638 x3.x2.GP1.n5 VSS 0.021877f
C3639 x4._16_.t1 VSS 0.046376f
C3640 x4._16_.n0 VSS 0.026397f
C3641 x4._16_.t2 VSS 0.021164f
C3642 x4._16_.t6 VSS 0.017507f
C3643 x4._16_.n1 VSS 0.047954f
C3644 x4._16_.n2 VSS 0.154756f
C3645 x4._16_.t7 VSS 0.020065f
C3646 x4._16_.t9 VSS 0.031953f
C3647 x4._16_.n3 VSS 0.045672f
C3648 x4._16_.n4 VSS 0.0375f
C3649 x4._16_.t4 VSS 0.020065f
C3650 x4._16_.t5 VSS 0.031953f
C3651 x4._16_.n5 VSS 0.058943f
C3652 x4._16_.n6 VSS 0.063595f
C3653 x4._16_.n7 VSS 0.426096f
C3654 x4._16_.t8 VSS 0.012893f
C3655 x4._16_.t3 VSS 0.013824f
C3656 x4._16_.n8 VSS 0.03796f
C3657 x4._16_.n9 VSS 0.022428f
C3658 x4._16_.n10 VSS 0.327394f
C3659 x4._16_.n11 VSS 0.020414f
C3660 x4._16_.t0 VSS 0.119992f
C3661 x4._16_.n12 VSS 0.021583f
C3662 x4._16_.n13 VSS 0.021194f
C3663 counter3.t2 VSS 0.033645f
C3664 counter3.n0 VSS 0.005854f
C3665 counter3.t3 VSS 0.023271f
C3666 counter3.n1 VSS 0.028526f
C3667 counter3.n2 VSS 0.0367f
C3668 counter3.n3 VSS 0.369569f
C3669 counter3.t0 VSS 0.736319f
C3670 counter3.t1 VSS 0.520878f
C3671 counter3.n4 VSS 4.03837f
C3672 counter3.t5 VSS 0.40872f
C3673 counter3.t4 VSS 0.757526f
C3674 counter3.n5 VSS 4.27416f
C3675 counter3.n6 VSS 0.668836f
C3676 x3.x2.GP2.t2 VSS 0.016198f
C3677 x3.x2.GP2.t3 VSS 0.016198f
C3678 x3.x2.GP2.n0 VSS 0.035585f
C3679 x3.x2.GP2.n1 VSS 0.023f
C3680 x3.x2.GP2.t5 VSS 0.819754f
C3681 x3.x2.GP2.t4 VSS 0.842614f
C3682 x3.x2.GP2.n2 VSS 2.98946f
C3683 x3.x2.GP2.t1 VSS 0.02492f
C3684 x3.x2.GP2.t0 VSS 0.02492f
C3685 x3.x2.GP2.n3 VSS 0.051391f
C3686 x3.x2.GP2.n4 VSS 0.120168f
C3687 x3.x2.GP2.n5 VSS 0.027176f
C3688 counter7.t0 VSS 0.030185f
C3689 counter7.n0 VSS 0.005252f
C3690 counter7.t1 VSS 0.020878f
C3691 counter7.n1 VSS 0.025593f
C3692 counter7.n2 VSS 0.0377f
C3693 counter7.n3 VSS 0.369403f
C3694 counter7.t5 VSS 0.660605f
C3695 counter7.t4 VSS 0.467316f
C3696 counter7.n4 VSS 3.62311f
C3697 counter7.t3 VSS 0.366915f
C3698 counter7.t2 VSS 0.672936f
C3699 counter7.n5 VSS 3.76478f
C3700 counter7.n6 VSS 0.600061f
C3701 x4.net3.t0 VSS 0.067779f
C3702 x4.net3.t6 VSS 0.019614f
C3703 x4.net3.t3 VSS 0.031428f
C3704 x4.net3.n0 VSS 0.061838f
C3705 x4.net3.n1 VSS 0.008618f
C3706 x4.net3.n2 VSS 0.005246f
C3707 x4.net3.t4 VSS 0.029572f
C3708 x4.net3.t5 VSS 0.018443f
C3709 x4.net3.n3 VSS 0.059457f
C3710 x4.net3.n4 VSS 0.019056f
C3711 x4.net3.t2 VSS 0.030361f
C3712 x4.net3.t7 VSS 0.055573f
C3713 x4.net3.n5 VSS 0.744487f
C3714 x4.net3.n6 VSS 0.124162f
C3715 x4.net3.n7 VSS 0.092279f
C3716 x4.net3.t1 VSS 0.037792f
C3717 x4.net3.n8 VSS 0.040884f
C3718 select0.t9 VSS 0.029056f
C3719 select0.t5 VSS 0.017122f
C3720 select0.t7 VSS 0.029056f
C3721 select0.t4 VSS 0.017122f
C3722 select0.n0 VSS 0.048752f
C3723 select0.n1 VSS 0.072053f
C3724 select0.n2 VSS 0.022642f
C3725 select0.t6 VSS 0.014311f
C3726 select0.t3 VSS 0.020786f
C3727 select0.n3 VSS 0.049512f
C3728 select0.n4 VSS 0.027499f
C3729 select0.t0 VSS 0.016946f
C3730 select0.t1 VSS 0.024957f
C3731 select0.n5 VSS 0.058963f
C3732 select0.n6 VSS 0.012245f
C3733 select0.n7 VSS 0.004774f
C3734 select0.n8 VSS 0.436077f
C3735 select0.t8 VSS 0.028355f
C3736 select0.t2 VSS 0.013445f
C3737 select0.n9 VSS 0.101818f
C3738 select0.n10 VSS 0.019731f
C3739 select0.n11 VSS 0.500298f
C3740 select0.n12 VSS 0.325096f
C3741 x4.net6.t13 VSS 0.023291f
C3742 x4.net6.t12 VSS 0.034395f
C3743 x4.net6.n0 VSS 0.095831f
C3744 x4.net6.t2 VSS 0.040459f
C3745 x4.net6.t5 VSS 0.025233f
C3746 x4.net6.n1 VSS 0.081347f
C3747 x4.net6.n2 VSS 0.124436f
C3748 x4.net6.t3 VSS 0.023291f
C3749 x4.net6.t8 VSS 0.034395f
C3750 x4.net6.n3 VSS 0.095831f
C3751 x4.net6.n4 VSS 0.41789f
C3752 x4.net6.t14 VSS 0.021456f
C3753 x4.net6.t15 VSS 0.017754f
C3754 x4.net6.n5 VSS 0.093771f
C3755 x4.net6.n6 VSS 0.080526f
C3756 x4.net6.n7 VSS 0.286209f
C3757 x4.net6.t4 VSS 0.027524f
C3758 x4.net6.t7 VSS 0.043832f
C3759 x4.net6.n8 VSS 0.059723f
C3760 x4.net6.n9 VSS 0.146037f
C3761 x4.net6.n10 VSS 0.772479f
C3762 x4.net6.n11 VSS 0.732404f
C3763 x4.net6.t6 VSS 0.023842f
C3764 x4.net6.t10 VSS 0.040459f
C3765 x4.net6.n12 VSS 0.051672f
C3766 x4.net6.t9 VSS 0.023842f
C3767 x4.net6.t11 VSS 0.040459f
C3768 x4.net6.n13 VSS 0.057394f
C3769 x4.net6.n14 VSS 0.027196f
C3770 x4.net6.n15 VSS 0.1061f
C3771 x4.net6.n16 VSS 0.491563f
C3772 x4.net6.t0 VSS 0.092732f
C3773 x4.net6.n17 VSS 0.127274f
C3774 x4.net6.t1 VSS 0.050895f
C3775 x4.net6.n18 VSS 0.064268f
C3776 select1.t2 VSS 0.033091f
C3777 select1.t9 VSS 0.0195f
C3778 select1.t4 VSS 0.033091f
C3779 select1.t1 VSS 0.0195f
C3780 select1.n0 VSS 0.055522f
C3781 select1.n1 VSS 0.082032f
C3782 select1.n2 VSS 0.050049f
C3783 select1.t8 VSS 0.032292f
C3784 select1.t0 VSS 0.015312f
C3785 select1.n3 VSS 0.115956f
C3786 select1.n4 VSS 0.022483f
C3787 select1.n5 VSS 0.019193f
C3788 select1.t7 VSS 0.016031f
C3789 select1.t3 VSS 0.023329f
C3790 select1.n6 VSS 0.067792f
C3791 select1.n7 VSS 0.015616f
C3792 select1.n8 VSS 0.111838f
C3793 select1.n9 VSS 0.405177f
C3794 select1.t5 VSS 0.0193f
C3795 select1.t6 VSS 0.028423f
C3796 select1.n10 VSS 0.067151f
C3797 select1.n11 VSS 0.008745f
C3798 select1.n12 VSS 0.098822f
C3799 select1.n13 VSS 0.467651f
C3800 select1.n14 VSS 0.610841f
C3801 x4.net2.t6 VSS 0.015381f
C3802 x4.net2.t10 VSS 0.026101f
C3803 x4.net2.n0 VSS 0.037026f
C3804 x4.net2.t4 VSS 0.015381f
C3805 x4.net2.t9 VSS 0.026101f
C3806 x4.net2.n1 VSS 0.033335f
C3807 x4.net2.n2 VSS 0.017289f
C3808 x4.net2.n3 VSS 0.0837f
C3809 x4.net2.t5 VSS 0.026101f
C3810 x4.net2.t7 VSS 0.016278f
C3811 x4.net2.n4 VSS 0.052479f
C3812 x4.net2.n5 VSS 0.259642f
C3813 x4.net2.t2 VSS 0.013842f
C3814 x4.net2.t3 VSS 0.011454f
C3815 x4.net2.n6 VSS 0.060494f
C3816 x4.net2.n7 VSS 0.03533f
C3817 x4.net2.n8 VSS 0.650991f
C3818 x4.net2.t8 VSS 0.017756f
C3819 x4.net2.t11 VSS 0.028277f
C3820 x4.net2.n9 VSS 0.038818f
C3821 x4.net2.n10 VSS 0.03575f
C3822 x4.net2.n11 VSS 0.11929f
C3823 x4.net2.n12 VSS 0.278364f
C3824 x4.net2.n13 VSS 0.037886f
C3825 x4.net2.t0 VSS 0.08709f
C3826 x4.net2.n14 VSS 0.10636f
C3827 x4.net2.t1 VSS 0.032833f
C3828 x4.clknet_0_clk.t31 VSS 0.004717f
C3829 x4.clknet_0_clk.t18 VSS 0.004717f
C3830 x4.clknet_0_clk.n0 VSS 0.016749f
C3831 x4.clknet_0_clk.t23 VSS 0.004717f
C3832 x4.clknet_0_clk.t17 VSS 0.004717f
C3833 x4.clknet_0_clk.n1 VSS 0.010767f
C3834 x4.clknet_0_clk.n2 VSS 0.068037f
C3835 x4.clknet_0_clk.t22 VSS 0.004717f
C3836 x4.clknet_0_clk.t28 VSS 0.004717f
C3837 x4.clknet_0_clk.n3 VSS 0.010767f
C3838 x4.clknet_0_clk.n4 VSS 0.040895f
C3839 x4.clknet_0_clk.t20 VSS 0.004717f
C3840 x4.clknet_0_clk.t26 VSS 0.004717f
C3841 x4.clknet_0_clk.n5 VSS 0.010774f
C3842 x4.clknet_0_clk.n6 VSS 0.042184f
C3843 x4.clknet_0_clk.t19 VSS 0.004717f
C3844 x4.clknet_0_clk.t25 VSS 0.004717f
C3845 x4.clknet_0_clk.n7 VSS 0.010767f
C3846 x4.clknet_0_clk.n8 VSS 0.040895f
C3847 x4.clknet_0_clk.t16 VSS 0.004717f
C3848 x4.clknet_0_clk.t24 VSS 0.004717f
C3849 x4.clknet_0_clk.n9 VSS 0.009573f
C3850 x4.clknet_0_clk.t45 VSS 0.015823f
C3851 x4.clknet_0_clk.t47 VSS 0.0074f
C3852 x4.clknet_0_clk.t38 VSS 0.015823f
C3853 x4.clknet_0_clk.t39 VSS 0.0074f
C3854 x4.clknet_0_clk.t42 VSS 0.015823f
C3855 x4.clknet_0_clk.t44 VSS 0.0074f
C3856 x4.clknet_0_clk.t36 VSS 0.015823f
C3857 x4.clknet_0_clk.t37 VSS 0.0074f
C3858 x4.clknet_0_clk.n10 VSS 0.036121f
C3859 x4.clknet_0_clk.n11 VSS 0.047576f
C3860 x4.clknet_0_clk.n12 VSS 0.047576f
C3861 x4.clknet_0_clk.n13 VSS 0.057784f
C3862 x4.clknet_0_clk.n14 VSS 0.075138f
C3863 x4.clknet_0_clk.t32 VSS 0.015823f
C3864 x4.clknet_0_clk.t33 VSS 0.0074f
C3865 x4.clknet_0_clk.t40 VSS 0.015823f
C3866 x4.clknet_0_clk.t41 VSS 0.0074f
C3867 x4.clknet_0_clk.t34 VSS 0.015823f
C3868 x4.clknet_0_clk.t35 VSS 0.0074f
C3869 x4.clknet_0_clk.t43 VSS 0.015823f
C3870 x4.clknet_0_clk.t46 VSS 0.0074f
C3871 x4.clknet_0_clk.n15 VSS 0.036121f
C3872 x4.clknet_0_clk.n16 VSS 0.047576f
C3873 x4.clknet_0_clk.n17 VSS 0.047576f
C3874 x4.clknet_0_clk.n18 VSS 0.057941f
C3875 x4.clknet_0_clk.n19 VSS 0.038186f
C3876 x4.clknet_0_clk.n20 VSS 0.145873f
C3877 x4.clknet_0_clk.n21 VSS 0.015919f
C3878 x4.clknet_0_clk.n22 VSS 0.026375f
C3879 x4.clknet_0_clk.t30 VSS 0.004717f
C3880 x4.clknet_0_clk.t21 VSS 0.004717f
C3881 x4.clknet_0_clk.n23 VSS 0.010767f
C3882 x4.clknet_0_clk.n24 VSS 0.035304f
C3883 x4.clknet_0_clk.t12 VSS 0.01123f
C3884 x4.clknet_0_clk.t14 VSS 0.01123f
C3885 x4.clknet_0_clk.n25 VSS 0.023364f
C3886 x4.clknet_0_clk.t0 VSS 0.01123f
C3887 x4.clknet_0_clk.t3 VSS 0.01123f
C3888 x4.clknet_0_clk.n26 VSS 0.028528f
C3889 x4.clknet_0_clk.t8 VSS 0.01123f
C3890 x4.clknet_0_clk.t2 VSS 0.01123f
C3891 x4.clknet_0_clk.n27 VSS 0.023672f
C3892 x4.clknet_0_clk.n28 VSS 0.107879f
C3893 x4.clknet_0_clk.t7 VSS 0.01123f
C3894 x4.clknet_0_clk.t13 VSS 0.01123f
C3895 x4.clknet_0_clk.n29 VSS 0.023672f
C3896 x4.clknet_0_clk.n30 VSS 0.062143f
C3897 x4.clknet_0_clk.t5 VSS 0.01123f
C3898 x4.clknet_0_clk.t11 VSS 0.01123f
C3899 x4.clknet_0_clk.n31 VSS 0.023672f
C3900 x4.clknet_0_clk.n32 VSS 0.061854f
C3901 x4.clknet_0_clk.t4 VSS 0.01123f
C3902 x4.clknet_0_clk.t10 VSS 0.01123f
C3903 x4.clknet_0_clk.n33 VSS 0.023672f
C3904 x4.clknet_0_clk.n34 VSS 0.061854f
C3905 x4.clknet_0_clk.t1 VSS 0.01123f
C3906 x4.clknet_0_clk.t9 VSS 0.01123f
C3907 x4.clknet_0_clk.n35 VSS 0.023672f
C3908 x4.clknet_0_clk.n36 VSS 0.062143f
C3909 x4.clknet_0_clk.t15 VSS 0.01123f
C3910 x4.clknet_0_clk.t6 VSS 0.01123f
C3911 x4.clknet_0_clk.n37 VSS 0.023672f
C3912 x4.clknet_0_clk.n38 VSS 0.053374f
C3913 x4.clknet_0_clk.n39 VSS 0.073498f
C3914 x4.clknet_0_clk.n40 VSS 0.034156f
C3915 x4.clknet_0_clk.t27 VSS 0.004717f
C3916 x4.clknet_0_clk.t29 VSS 0.004717f
C3917 x4.clknet_0_clk.n41 VSS 0.010394f
C3918 x4.clknet_1_1__leaf_clk.t18 VSS 0.005541f
C3919 x4.clknet_1_1__leaf_clk.t20 VSS 0.005541f
C3920 x4.clknet_1_1__leaf_clk.n0 VSS 0.019676f
C3921 x4.clknet_1_1__leaf_clk.t21 VSS 0.005541f
C3922 x4.clknet_1_1__leaf_clk.t28 VSS 0.005541f
C3923 x4.clknet_1_1__leaf_clk.n1 VSS 0.01265f
C3924 x4.clknet_1_1__leaf_clk.n2 VSS 0.07993f
C3925 x4.clknet_1_1__leaf_clk.t23 VSS 0.005541f
C3926 x4.clknet_1_1__leaf_clk.t30 VSS 0.005541f
C3927 x4.clknet_1_1__leaf_clk.n3 VSS 0.01265f
C3928 x4.clknet_1_1__leaf_clk.n4 VSS 0.048044f
C3929 x4.clknet_1_1__leaf_clk.t26 VSS 0.005541f
C3930 x4.clknet_1_1__leaf_clk.t16 VSS 0.005541f
C3931 x4.clknet_1_1__leaf_clk.n5 VSS 0.012657f
C3932 x4.clknet_1_1__leaf_clk.n6 VSS 0.049559f
C3933 x4.clknet_1_1__leaf_clk.t27 VSS 0.005541f
C3934 x4.clknet_1_1__leaf_clk.t17 VSS 0.005541f
C3935 x4.clknet_1_1__leaf_clk.n7 VSS 0.01265f
C3936 x4.clknet_1_1__leaf_clk.n8 VSS 0.048044f
C3937 x4.clknet_1_1__leaf_clk.t29 VSS 0.005541f
C3938 x4.clknet_1_1__leaf_clk.t19 VSS 0.005541f
C3939 x4.clknet_1_1__leaf_clk.n9 VSS 0.011247f
C3940 x4.clknet_1_1__leaf_clk.t33 VSS 0.013817f
C3941 x4.clknet_1_1__leaf_clk.t32 VSS 0.020651f
C3942 x4.clknet_1_1__leaf_clk.n10 VSS 0.038168f
C3943 x4.clknet_1_1__leaf_clk.t36 VSS 0.020651f
C3944 x4.clknet_1_1__leaf_clk.t35 VSS 0.013817f
C3945 x4.clknet_1_1__leaf_clk.n11 VSS 0.037785f
C3946 x4.clknet_1_1__leaf_clk.n12 VSS 0.039947f
C3947 x4.clknet_1_1__leaf_clk.t37 VSS 0.013817f
C3948 x4.clknet_1_1__leaf_clk.t34 VSS 0.020651f
C3949 x4.clknet_1_1__leaf_clk.n13 VSS 0.038168f
C3950 x4.clknet_1_1__leaf_clk.n14 VSS 0.30833f
C3951 x4.clknet_1_1__leaf_clk.t40 VSS 0.020651f
C3952 x4.clknet_1_1__leaf_clk.t39 VSS 0.013817f
C3953 x4.clknet_1_1__leaf_clk.n15 VSS 0.037785f
C3954 x4.clknet_1_1__leaf_clk.n16 VSS 0.030886f
C3955 x4.clknet_1_1__leaf_clk.n17 VSS 0.118422f
C3956 x4.clknet_1_1__leaf_clk.t41 VSS 0.013817f
C3957 x4.clknet_1_1__leaf_clk.t38 VSS 0.020651f
C3958 x4.clknet_1_1__leaf_clk.n18 VSS 0.037832f
C3959 x4.clknet_1_1__leaf_clk.n19 VSS 0.022005f
C3960 x4.clknet_1_1__leaf_clk.n20 VSS 0.128874f
C3961 x4.clknet_1_1__leaf_clk.n21 VSS 0.280206f
C3962 x4.clknet_1_1__leaf_clk.n22 VSS 0.023331f
C3963 x4.clknet_1_1__leaf_clk.n23 VSS 0.030986f
C3964 x4.clknet_1_1__leaf_clk.t31 VSS 0.005541f
C3965 x4.clknet_1_1__leaf_clk.t22 VSS 0.005541f
C3966 x4.clknet_1_1__leaf_clk.n24 VSS 0.01265f
C3967 x4.clknet_1_1__leaf_clk.n25 VSS 0.041476f
C3968 x4.clknet_1_1__leaf_clk.t8 VSS 0.013193f
C3969 x4.clknet_1_1__leaf_clk.t9 VSS 0.013193f
C3970 x4.clknet_1_1__leaf_clk.n26 VSS 0.027449f
C3971 x4.clknet_1_1__leaf_clk.t2 VSS 0.013193f
C3972 x4.clknet_1_1__leaf_clk.t4 VSS 0.013193f
C3973 x4.clknet_1_1__leaf_clk.n27 VSS 0.033515f
C3974 x4.clknet_1_1__leaf_clk.t5 VSS 0.013193f
C3975 x4.clknet_1_1__leaf_clk.t12 VSS 0.013193f
C3976 x4.clknet_1_1__leaf_clk.n28 VSS 0.02781f
C3977 x4.clknet_1_1__leaf_clk.n29 VSS 0.126738f
C3978 x4.clknet_1_1__leaf_clk.t7 VSS 0.013193f
C3979 x4.clknet_1_1__leaf_clk.t14 VSS 0.013193f
C3980 x4.clknet_1_1__leaf_clk.n30 VSS 0.02781f
C3981 x4.clknet_1_1__leaf_clk.n31 VSS 0.073006f
C3982 x4.clknet_1_1__leaf_clk.t10 VSS 0.013193f
C3983 x4.clknet_1_1__leaf_clk.t0 VSS 0.013193f
C3984 x4.clknet_1_1__leaf_clk.n32 VSS 0.02781f
C3985 x4.clknet_1_1__leaf_clk.n33 VSS 0.072667f
C3986 x4.clknet_1_1__leaf_clk.t11 VSS 0.013193f
C3987 x4.clknet_1_1__leaf_clk.t1 VSS 0.013193f
C3988 x4.clknet_1_1__leaf_clk.n34 VSS 0.02781f
C3989 x4.clknet_1_1__leaf_clk.n35 VSS 0.072667f
C3990 x4.clknet_1_1__leaf_clk.t13 VSS 0.013193f
C3991 x4.clknet_1_1__leaf_clk.t3 VSS 0.013193f
C3992 x4.clknet_1_1__leaf_clk.n36 VSS 0.02781f
C3993 x4.clknet_1_1__leaf_clk.n37 VSS 0.073006f
C3994 x4.clknet_1_1__leaf_clk.t15 VSS 0.013193f
C3995 x4.clknet_1_1__leaf_clk.t6 VSS 0.013193f
C3996 x4.clknet_1_1__leaf_clk.n38 VSS 0.02781f
C3997 x4.clknet_1_1__leaf_clk.n39 VSS 0.062704f
C3998 x4.clknet_1_1__leaf_clk.n40 VSS 0.086346f
C3999 x4.clknet_1_1__leaf_clk.n41 VSS 0.040127f
C4000 x4.clknet_1_1__leaf_clk.t24 VSS 0.005541f
C4001 x4.clknet_1_1__leaf_clk.t25 VSS 0.005541f
C4002 x4.clknet_1_1__leaf_clk.n42 VSS 0.012211f
C4003 mux_out.t15 VSS 0.469199f
C4004 mux_out.n0 VSS 0.583543f
C4005 mux_out.t2 VSS 0.363309f
C4006 mux_out.t14 VSS 0.482119f
C4007 mux_out.n1 VSS 2.43292f
C4008 mux_out.n2 VSS 0.823196f
C4009 mux_out.t3 VSS 0.35616f
C4010 mux_out.n3 VSS 0.53181f
C4011 mux_out.n4 VSS 0.741524f
C4012 mux_out.t0 VSS 0.469199f
C4013 mux_out.n5 VSS 0.583543f
C4014 mux_out.t6 VSS 0.363309f
C4015 mux_out.t1 VSS 0.482119f
C4016 mux_out.n6 VSS 2.43292f
C4017 mux_out.n7 VSS 0.823196f
C4018 mux_out.t7 VSS 0.35616f
C4019 mux_out.n8 VSS 0.53181f
C4020 mux_out.n9 VSS 0.72062f
C4021 mux_out.n10 VSS 0.393629f
C4022 mux_out.t12 VSS 0.469199f
C4023 mux_out.n11 VSS 0.583543f
C4024 mux_out.t10 VSS 0.363309f
C4025 mux_out.t13 VSS 0.482119f
C4026 mux_out.n12 VSS 2.43292f
C4027 mux_out.n13 VSS 0.823196f
C4028 mux_out.t11 VSS 0.35616f
C4029 mux_out.n14 VSS 0.53181f
C4030 mux_out.n15 VSS 0.721457f
C4031 mux_out.n16 VSS 0.390909f
C4032 mux_out.n17 VSS 1.16541f
C4033 mux_out.t4 VSS 0.469199f
C4034 mux_out.n18 VSS 0.583543f
C4035 mux_out.t9 VSS 0.363309f
C4036 mux_out.t5 VSS 0.482119f
C4037 mux_out.n19 VSS 2.43292f
C4038 mux_out.n20 VSS 0.823196f
C4039 mux_out.t8 VSS 0.35616f
C4040 mux_out.n21 VSS 0.53181f
C4041 mux_out.n22 VSS 0.727887f
C4042 mux_out.n23 VSS 0.384347f
C4043 mux_out.n24 VSS 0.557092f
C4044 drv_out.t2 VSS 0.591341f
C4045 drv_out.t3 VSS 0.418319f
C4046 drv_out.n0 VSS 3.24323f
C4047 drv_out.t0 VSS 0.328444f
C4048 drv_out.t1 VSS 0.602379f
C4049 drv_out.n1 VSS 3.37005f
C4050 drv_out.n2 VSS 0.537145f
C4051 drv_out.n3 VSS 0.110148f
C4052 drv_out.t24 VSS 0.015262f
C4053 drv_out.t25 VSS 0.007138f
C4054 drv_out.t20 VSS 0.015262f
C4055 drv_out.t21 VSS 0.007138f
C4056 drv_out.t26 VSS 0.015262f
C4057 drv_out.t27 VSS 0.007138f
C4058 drv_out.t22 VSS 0.015262f
C4059 drv_out.t23 VSS 0.007138f
C4060 drv_out.n4 VSS 0.034841f
C4061 drv_out.n5 VSS 0.04589f
C4062 drv_out.n6 VSS 0.04589f
C4063 drv_out.n7 VSS 0.055736f
C4064 drv_out.n8 VSS 0.015444f
C4065 drv_out.n9 VSS 0.346765f
C4066 drv_out.n10 VSS 0.764086f
C4067 drv_out.n11 VSS 5.53733f
C4068 drv_out.t4 VSS 0.1149f
C4069 drv_out.t6 VSS 0.1149f
C4070 drv_out.n12 VSS 0.273611f
C4071 drv_out.t8 VSS 0.1149f
C4072 drv_out.t7 VSS 0.1149f
C4073 drv_out.n13 VSS 0.273611f
C4074 drv_out.t10 VSS 0.1149f
C4075 drv_out.t9 VSS 0.1149f
C4076 drv_out.n14 VSS 0.273611f
C4077 drv_out.t11 VSS 0.1149f
C4078 drv_out.t5 VSS 0.1149f
C4079 drv_out.n15 VSS 0.273611f
C4080 drv_out.n16 VSS 4.32f
C4081 drv_out.t17 VSS 0.0383f
C4082 drv_out.t18 VSS 0.0383f
C4083 drv_out.n17 VSS 0.093269f
C4084 drv_out.t12 VSS 0.0383f
C4085 drv_out.t19 VSS 0.0383f
C4086 drv_out.n18 VSS 0.093269f
C4087 drv_out.t15 VSS 0.0383f
C4088 drv_out.t14 VSS 0.0383f
C4089 drv_out.n19 VSS 0.093269f
C4090 drv_out.t16 VSS 0.0383f
C4091 drv_out.t13 VSS 0.0383f
C4092 drv_out.n20 VSS 0.093269f
C4093 drv_out.n21 VSS 1.9949f
C4094 drv_out.n22 VSS 2.14485f
C4095 x4._11_.t0 VSS 0.02558f
C4096 x4._11_.t1 VSS 0.02558f
C4097 x4._11_.n0 VSS 0.053419f
C4098 x4._11_.t7 VSS 0.042601f
C4099 x4._11_.t11 VSS 0.026392f
C4100 x4._11_.n1 VSS 0.086305f
C4101 x4._11_.n2 VSS 0.024278f
C4102 x4._11_.t8 VSS 0.027069f
C4103 x4._11_.t10 VSS 0.043108f
C4104 x4._11_.n3 VSS 0.058737f
C4105 x4._11_.n4 VSS 0.032841f
C4106 x4._11_.t14 VSS 0.023619f
C4107 x4._11_.t17 VSS 0.034667f
C4108 x4._11_.n5 VSS 0.06984f
C4109 x4._11_.n6 VSS 0.034707f
C4110 x4._11_.n7 VSS 0.494881f
C4111 x4._11_.t6 VSS 0.027069f
C4112 x4._11_.t9 VSS 0.043108f
C4113 x4._11_.n8 VSS 0.058739f
C4114 x4._11_.n9 VSS 0.133927f
C4115 x4._11_.n10 VSS 0.765831f
C4116 x4._11_.t15 VSS 0.021102f
C4117 x4._11_.t16 VSS 0.017461f
C4118 x4._11_.n11 VSS 0.092223f
C4119 x4._11_.n12 VSS 0.043963f
C4120 x4._11_.n13 VSS 0.150035f
C4121 x4._11_.t20 VSS 0.028052f
C4122 x4._11_.t18 VSS 0.019277f
C4123 x4._11_.n14 VSS 0.081517f
C4124 x4._11_.n15 VSS 0.011369f
C4125 x4._11_.n16 VSS 0.03744f
C4126 x4._11_.n17 VSS 0.156255f
C4127 x4._11_.t13 VSS 0.019598f
C4128 x4._11_.t19 VSS 0.028465f
C4129 x4._11_.n18 VSS 0.067767f
C4130 x4._11_.n19 VSS 0.143997f
C4131 x4._11_.n20 VSS 0.492685f
C4132 x4._11_.t21 VSS 0.042359f
C4133 x4._11_.t4 VSS 0.026451f
C4134 x4._11_.n21 VSS 0.080165f
C4135 x4._11_.n22 VSS 0.023455f
C4136 x4._11_.n23 VSS 0.356691f
C4137 x4._11_.t12 VSS 0.023619f
C4138 x4._11_.t5 VSS 0.034667f
C4139 x4._11_.n24 VSS 0.06984f
C4140 x4._11_.n25 VSS 0.014495f
C4141 x4._11_.n26 VSS 0.490885f
C4142 x4._11_.n27 VSS 1.19049f
C4143 x4._11_.n28 VSS 0.353781f
C4144 x4._11_.n29 VSS 0.021904f
C4145 x4._11_.t2 VSS 0.010743f
C4146 x4._11_.t3 VSS 0.010743f
C4147 x4._11_.n30 VSS 0.02648f
C4148 x3.x2.x4.GP VSS 2.5438f
C4149 x3.x1.gpo3 VSS 1.19037f
C4150 x3.x2.GP4.t2 VSS 0.012213f
C4151 x3.x2.GP4.t3 VSS 0.012213f
C4152 x3.x2.GP4.n0 VSS 0.026831f
C4153 x3.x1.x14.Y VSS 0.075955f
C4154 x3.x2.GP4.n1 VSS 0.010383f
C4155 x3.x2.GP4.t5 VSS 0.618091f
C4156 x3.x2.GP4.t4 VSS 0.635327f
C4157 x3.x2.GP4.n2 VSS 2.25863f
C4158 x3.x2.GP4.n3 VSS 0.047772f
C4159 x3.x2.GP4.t1 VSS 0.01879f
C4160 x3.x2.GP4.t0 VSS 0.01879f
C4161 x3.x2.GP4.n4 VSS 0.043205f
C4162 x3.x2.GP4.n5 VSS 0.087626f
C4163 a_21119_n968.t9 VSS 0.136375f
C4164 a_21119_n968.t7 VSS 0.13635f
C4165 a_21119_n968.n0 VSS 0.157675f
C4166 a_21119_n968.t6 VSS 0.13635f
C4167 a_21119_n968.n1 VSS 0.086028f
C4168 a_21119_n968.t14 VSS 0.13635f
C4169 a_21119_n968.n2 VSS 0.160734f
C4170 a_21119_n968.t2 VSS 0.049796f
C4171 a_21119_n968.t15 VSS 0.049764f
C4172 a_21119_n968.n3 VSS 0.09498f
C4173 a_21119_n968.t3 VSS 0.049764f
C4174 a_21119_n968.n4 VSS 0.055718f
C4175 a_21119_n968.t16 VSS 0.049764f
C4176 a_21119_n968.n5 VSS 0.086134f
C4177 a_21119_n968.t1 VSS 0.098833f
C4178 a_21119_n968.n6 VSS 0.831842f
C4179 a_21119_n968.t17 VSS 0.049771f
C4180 a_21119_n968.t10 VSS 0.13635f
C4181 a_21119_n968.n7 VSS 0.503671f
C4182 a_21119_n968.t11 VSS 0.049764f
C4183 a_21119_n968.n8 VSS 0.212248f
C4184 a_21119_n968.t8 VSS 0.13635f
C4185 a_21119_n968.n9 VSS 0.242932f
C4186 a_21119_n968.t4 VSS 0.049764f
C4187 a_21119_n968.n10 VSS 0.212248f
C4188 a_21119_n968.t13 VSS 0.13635f
C4189 a_21119_n968.n11 VSS 0.242932f
C4190 a_21119_n968.t5 VSS 0.049764f
C4191 a_21119_n968.n12 VSS 0.212248f
C4192 a_21119_n968.t12 VSS 0.13635f
C4193 a_21119_n968.n13 VSS 0.494157f
C4194 a_21119_n968.n14 VSS 1.47337f
C4195 a_21119_n968.n15 VSS 2.33573f
C4196 a_21119_n968.t0 VSS 0.309542f
C4197 ring_out.t10 VSS 0.143976f
C4198 ring_out.t12 VSS 0.066482f
C4199 ring_out.n0 VSS 1.43742f
C4200 ring_out.t3 VSS 0.011895f
C4201 ring_out.t2 VSS 0.011895f
C4202 ring_out.n1 VSS 0.036116f
C4203 ring_out.t0 VSS 0.011895f
C4204 ring_out.t4 VSS 0.011895f
C4205 ring_out.n2 VSS 0.026441f
C4206 ring_out.n3 VSS 0.119642f
C4207 ring_out.t1 VSS 0.007732f
C4208 ring_out.t5 VSS 0.007732f
C4209 ring_out.n4 VSS 0.017154f
C4210 ring_out.n5 VSS 0.032249f
C4211 ring_out.n6 VSS 0.009203f
C4212 ring_out.t13 VSS 0.010903f
C4213 ring_out.t14 VSS 0.018503f
C4214 ring_out.t15 VSS 0.010903f
C4215 ring_out.t11 VSS 0.018503f
C4216 ring_out.n7 VSS 0.031045f
C4217 ring_out.n8 VSS 0.04596f
C4218 ring_out.n9 VSS 0.181049f
C4219 ring_out.n10 VSS 0.421446f
C4220 ring_out.t6 VSS 0.673389f
C4221 ring_out.t7 VSS 0.47636f
C4222 ring_out.n11 VSS 3.69323f
C4223 ring_out.t8 VSS 0.374016f
C4224 ring_out.t9 VSS 0.685959f
C4225 ring_out.n12 VSS 3.83764f
C4226 ring_out.n13 VSS 0.611674f
C4227 x4.clknet_1_0__leaf_clk.t36 VSS 0.022262f
C4228 x4.clknet_1_0__leaf_clk.t34 VSS 0.014894f
C4229 x4.clknet_1_0__leaf_clk.n0 VSS 0.04068f
C4230 x4.clknet_1_0__leaf_clk.n1 VSS 0.107083f
C4231 x4.clknet_1_0__leaf_clk.t40 VSS 0.014894f
C4232 x4.clknet_1_0__leaf_clk.t38 VSS 0.022262f
C4233 x4.clknet_1_0__leaf_clk.n2 VSS 0.041145f
C4234 x4.clknet_1_0__leaf_clk.n3 VSS 0.437523f
C4235 x4.clknet_1_0__leaf_clk.t10 VSS 0.014222f
C4236 x4.clknet_1_0__leaf_clk.t0 VSS 0.014222f
C4237 x4.clknet_1_0__leaf_clk.n4 VSS 0.029978f
C4238 x4.clknet_1_0__leaf_clk.t4 VSS 0.014222f
C4239 x4.clknet_1_0__leaf_clk.t9 VSS 0.014222f
C4240 x4.clknet_1_0__leaf_clk.n5 VSS 0.029589f
C4241 x4.clknet_1_0__leaf_clk.t23 VSS 0.005973f
C4242 x4.clknet_1_0__leaf_clk.t29 VSS 0.005973f
C4243 x4.clknet_1_0__leaf_clk.n6 VSS 0.021211f
C4244 x4.clknet_1_0__leaf_clk.t21 VSS 0.005973f
C4245 x4.clknet_1_0__leaf_clk.t27 VSS 0.005973f
C4246 x4.clknet_1_0__leaf_clk.n7 VSS 0.013636f
C4247 x4.clknet_1_0__leaf_clk.n8 VSS 0.086164f
C4248 x4.clknet_1_0__leaf_clk.t19 VSS 0.005973f
C4249 x4.clknet_1_0__leaf_clk.t24 VSS 0.005973f
C4250 x4.clknet_1_0__leaf_clk.n9 VSS 0.013636f
C4251 x4.clknet_1_0__leaf_clk.n10 VSS 0.051791f
C4252 x4.clknet_1_0__leaf_clk.t31 VSS 0.005973f
C4253 x4.clknet_1_0__leaf_clk.t18 VSS 0.005973f
C4254 x4.clknet_1_0__leaf_clk.n11 VSS 0.013644f
C4255 x4.clknet_1_0__leaf_clk.n12 VSS 0.053424f
C4256 x4.clknet_1_0__leaf_clk.t30 VSS 0.005973f
C4257 x4.clknet_1_0__leaf_clk.t22 VSS 0.005973f
C4258 x4.clknet_1_0__leaf_clk.n13 VSS 0.013636f
C4259 x4.clknet_1_0__leaf_clk.n14 VSS 0.051791f
C4260 x4.clknet_1_0__leaf_clk.t28 VSS 0.005973f
C4261 x4.clknet_1_0__leaf_clk.t17 VSS 0.005973f
C4262 x4.clknet_1_0__leaf_clk.n15 VSS 0.013636f
C4263 x4.clknet_1_0__leaf_clk.n16 VSS 0.05205f
C4264 x4.clknet_1_0__leaf_clk.t26 VSS 0.005973f
C4265 x4.clknet_1_0__leaf_clk.t16 VSS 0.005973f
C4266 x4.clknet_1_0__leaf_clk.n17 VSS 0.013636f
C4267 x4.clknet_1_0__leaf_clk.n18 VSS 0.04471f
C4268 x4.clknet_1_0__leaf_clk.t20 VSS 0.005973f
C4269 x4.clknet_1_0__leaf_clk.t25 VSS 0.005973f
C4270 x4.clknet_1_0__leaf_clk.n19 VSS 0.013163f
C4271 x4.clknet_1_0__leaf_clk.n20 VSS 0.043256f
C4272 x4.clknet_1_0__leaf_clk.n21 VSS 0.09308f
C4273 x4.clknet_1_0__leaf_clk.n22 VSS 0.067594f
C4274 x4.clknet_1_0__leaf_clk.t14 VSS 0.014222f
C4275 x4.clknet_1_0__leaf_clk.t6 VSS 0.014222f
C4276 x4.clknet_1_0__leaf_clk.n23 VSS 0.029978f
C4277 x4.clknet_1_0__leaf_clk.t7 VSS 0.014222f
C4278 x4.clknet_1_0__leaf_clk.t13 VSS 0.014222f
C4279 x4.clknet_1_0__leaf_clk.n24 VSS 0.036128f
C4280 x4.clknet_1_0__leaf_clk.t5 VSS 0.014222f
C4281 x4.clknet_1_0__leaf_clk.t11 VSS 0.014222f
C4282 x4.clknet_1_0__leaf_clk.n25 VSS 0.029978f
C4283 x4.clknet_1_0__leaf_clk.n26 VSS 0.136621f
C4284 x4.clknet_1_0__leaf_clk.t3 VSS 0.014222f
C4285 x4.clknet_1_0__leaf_clk.t8 VSS 0.014222f
C4286 x4.clknet_1_0__leaf_clk.n27 VSS 0.029978f
C4287 x4.clknet_1_0__leaf_clk.n28 VSS 0.0787f
C4288 x4.clknet_1_0__leaf_clk.t15 VSS 0.014222f
C4289 x4.clknet_1_0__leaf_clk.t2 VSS 0.014222f
C4290 x4.clknet_1_0__leaf_clk.n29 VSS 0.029978f
C4291 x4.clknet_1_0__leaf_clk.n30 VSS 0.078334f
C4292 x4.clknet_1_0__leaf_clk.n31 VSS 0.078334f
C4293 x4.clknet_1_0__leaf_clk.n32 VSS 0.04742f
C4294 x4.clknet_1_0__leaf_clk.t12 VSS 0.014222f
C4295 x4.clknet_1_0__leaf_clk.t1 VSS 0.014222f
C4296 x4.clknet_1_0__leaf_clk.n33 VSS 0.028445f
C4297 x4.clknet_1_0__leaf_clk.n34 VSS 0.022411f
C4298 x4.clknet_1_0__leaf_clk.n35 VSS 0.171468f
C4299 x4.clknet_1_0__leaf_clk.t41 VSS 0.014894f
C4300 x4.clknet_1_0__leaf_clk.t39 VSS 0.022262f
C4301 x4.clknet_1_0__leaf_clk.n36 VSS 0.040782f
C4302 x4.clknet_1_0__leaf_clk.n37 VSS 0.024896f
C4303 x4.clknet_1_0__leaf_clk.t33 VSS 0.022262f
C4304 x4.clknet_1_0__leaf_clk.t32 VSS 0.014894f
C4305 x4.clknet_1_0__leaf_clk.n38 VSS 0.040732f
C4306 x4.clknet_1_0__leaf_clk.n39 VSS 0.086433f
C4307 x4.clknet_1_0__leaf_clk.n40 VSS 0.225449f
C4308 x4.clknet_1_0__leaf_clk.t35 VSS 0.022262f
C4309 x4.clknet_1_0__leaf_clk.t37 VSS 0.014894f
C4310 x4.clknet_1_0__leaf_clk.n41 VSS 0.04068f
C4311 x4.clknet_1_0__leaf_clk.n42 VSS 0.027948f
C4312 x4.clknet_1_0__leaf_clk.n43 VSS 0.145937f
.ends

