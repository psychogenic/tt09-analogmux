magic
tech sky130A
magscale 1 2
timestamp 1729136545
<< pwell >>
rect 3936 -650 3986 -522
rect 7518 -550 7576 -506
rect 5742 -664 5890 -584
rect 5756 -828 5876 -664
<< locali >>
rect 8002 -318 8070 36
rect 7868 -320 8070 -318
rect 3522 -390 8070 -320
rect 7868 -412 8070 -390
rect 3800 -650 3970 -428
rect 7868 -526 7878 -412
rect 8050 -578 8070 -412
rect 3860 -792 3970 -650
rect 3860 -812 7700 -792
rect 3702 -880 7700 -812
<< viali >>
rect 7878 -580 8050 -412
rect 3702 -812 3860 -650
<< metal1 >>
rect 3508 34 7950 88
rect 3508 -404 3582 34
rect 3714 -92 3724 -20
rect 5498 -92 5508 -20
rect 3724 -112 5498 -92
rect 5692 -126 5782 34
rect 5990 -76 6000 -4
rect 7774 -76 7784 -4
rect 5996 -106 7770 -76
rect 5662 -192 5808 -126
rect 7896 -194 7950 34
rect 3780 -298 5362 -206
rect 6032 -292 7614 -200
rect 3436 -604 3636 -404
rect 3682 -512 3882 -404
rect 4264 -480 4524 -298
rect 5050 -356 5310 -298
rect 6102 -356 6362 -292
rect 5050 -438 6362 -356
rect 5050 -480 5310 -438
rect 6102 -478 6362 -438
rect 6970 -478 7230 -292
rect 7460 -400 7576 -292
rect 7460 -478 7826 -400
rect 3682 -590 3986 -512
rect 4126 -572 5708 -480
rect 5938 -494 7826 -478
rect 5938 -550 7576 -494
rect 5938 -570 7520 -550
rect 3682 -604 4078 -590
rect 3434 -660 3634 -632
rect 3434 -802 3460 -660
rect 3600 -802 3634 -660
rect 3434 -832 3634 -802
rect 3684 -650 3884 -632
rect 3936 -650 4078 -604
rect 3684 -812 3702 -650
rect 3860 -812 3884 -650
rect 3684 -832 3884 -812
rect 4016 -792 4072 -650
rect 5742 -664 5890 -584
rect 4152 -684 5636 -666
rect 4142 -760 4152 -684
rect 5636 -760 5646 -684
rect 5756 -792 5876 -664
rect 5986 -688 7470 -668
rect 5984 -764 5994 -688
rect 7478 -764 7488 -688
rect 7560 -792 7620 -586
rect 7720 -642 7826 -494
rect 7866 -412 8066 -398
rect 7866 -580 7878 -412
rect 8050 -580 8066 -412
rect 7866 -598 8066 -580
rect 4016 -864 7622 -792
rect 7720 -842 7972 -642
<< via1 >>
rect 3724 -92 5498 -20
rect 6000 -76 7774 -4
rect 3460 -802 3600 -660
rect 4152 -760 5636 -684
rect 5994 -764 7478 -688
<< metal2 >>
rect 3356 71 7073 137
rect 3356 -654 3422 71
rect 4096 -10 4998 71
rect 6168 6 7070 71
rect 6000 -4 7774 6
rect 3724 -20 5498 -10
rect 6000 -86 7774 -76
rect 3724 -102 5498 -92
rect 3460 -654 3600 -650
rect 3356 -660 3600 -654
rect 3356 -772 3460 -660
rect 3358 -776 3460 -772
rect 4152 -684 5636 -674
rect 4152 -770 5636 -760
rect 5994 -688 7478 -678
rect 3460 -820 3600 -802
rect 4348 -820 5504 -770
rect 5994 -774 7478 -764
rect 6096 -820 7252 -774
rect 3460 -886 7396 -820
rect 3460 -888 3600 -886
rect 3460 -890 3570 -888
use sky130_fd_pr__nfet_01v8_lvt_PEJ72P  XM1 std
timestamp 1725636896
transform 0 -1 5819 1 0 -621
box -231 -1919 231 1919
use sky130_fd_pr__pfet_01v8_lvt_4QFMR3  XM3 std
timestamp 1725636896
transform 0 -1 5735 1 0 -157
box -231 -2337 231 2337
<< labels >>
flabel metal1 3434 -832 3634 -632 0 FreeSans 256 0 0 0 A
port 0 nsew
flabel metal1 3682 -604 3882 -404 0 FreeSans 256 0 0 0 GN
port 1 nsew
flabel metal1 3436 -604 3636 -404 0 FreeSans 256 0 0 0 GP
port 2 nsew
flabel metal1 7772 -842 7972 -642 0 FreeSans 256 0 0 0 Z
port 3 nsew
flabel metal1 7866 -598 8066 -398 0 FreeSans 256 0 0 0 VDD
port 4 nsew
flabel metal1 3684 -832 3884 -632 0 FreeSans 256 0 0 0 VSS
port 5 nsew
<< end >>
