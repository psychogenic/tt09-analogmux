** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sch
.subckt muxtest VSS VDD SELECT0 SELECT1 VRES RSEL0 RSEL1 RSEL2 OUT LADDEROUT
*.PININFO VSS:I VDD:I SELECT0:I SELECT1:I VRES:I RSEL0:I RSEL1:I RSEL2:I OUT:O LADDEROUT:O
x1 VDD VSS RSEL0 RSEL1 A1 A5 A6 A2 A7 A3 RSEL2 VRES A4 LADDEROUT mux8onehot
x2 SELECT0 SELECT1 VDD LADDEROUT VRES A5 A1 OUT OUT OUT OUT net1 VDD VSS mux4onehot_b
XR1 A7 VRES VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR2 A6 A7 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR3 A5 A6 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR4 A4 A5 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR5 A3 A4 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR6 A2 A3 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR7 A1 A2 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR8 VSS A1 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
.ends

* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sch
.subckt mux8onehot VDD VSS select0 select1 A1 A5 A6 A2 A7 A3 select2 A8 A4 Z
*.PININFO select0:I select1:I select2:I VDD:I VSS:I Z:B A1:B A2:B A3:B A4:B A5:B A6:B A7:B A8:B
x4 OUT_HIGH select2 nSEL2 Z VDD VSS passgate
x5 OUT_LOW nSEL2 select2 Z VDD VSS passgate
x2 A1 gno0 gpo0 OUT_LOW A2 gno1 gpo1 OUT_LOW A3 gno2 gpo2 OUT_LOW A4 gno3 gpo3 OUT_LOW VDD VSS passgatex4
x1 select0 select1 select2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nSEL2 VDD VSS passgatesCtrlManual
x3 A5 gno0 gpo0 OUT_HIGH A6 gno1 gpo1 OUT_HIGH A7 gno2 gpo2 OUT_HIGH A8 gno3 gpo3 OUT_HIGH VDD VSS passgatex4
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sch
.subckt mux4onehot_b select0 select1 select2 A1 A2 A3 A4 Z1 Z2 Z3 Z4 nselect2 VDD VSS
*.PININFO select0:I select1:I select2:I A1:B A2:B A3:B A4:B Z1:B Z2:B Z3:B Z4:B nselect2:O VDD:I VSS:I
x2 A1 gno0 gpo0 Z1 A2 gno1 gpo1 Z2 A3 gno2 gpo2 Z3 A4 gno3 gpo3 Z4 VDD VSS passgatex4
x1 select0 select1 select2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nselect2 VDD VSS passgatesCtrlManual
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym # of pins=6
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sch
.subckt passgate A GN GP Z VCCBPIN VSSBPIN
*.PININFO GN:I VCCBPIN:I VSSBPIN:I GP:I A:B Z:B
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 m=2
XM3 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=2
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym # of pins=18
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sch
.subckt passgatex4 A1 GN1 GP1 Z1 A2 GN2 GP2 Z2 A3 GN3 GP3 Z3 A4 GN4 GP4 Z4 VDD VSS
*.PININFO VDD:I VSS:I GP1:I GN1:I A1:B Z1:B GP2:I GN2:I A2:B Z2:B GP3:I GN3:I A3:B Z3:B GP4:I GN4:I A4:B Z4:B
x1 Z1 A1 GP1 GN1 VSS VDD passgate
x2 Z2 A2 GP2 GN2 VSS VDD passgate
x3 Z3 A3 GP3 GN3 VSS VDD passgate
x4 Z4 A4 GP4 GN4 VSS VDD passgate
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sch
.subckt passgatesCtrlManual SEL0 SEL1 SEL2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nSEL2 VPWR VGND
*.PININFO SEL0:I SEL1:I SEL2:I gno0:O gpo0:O gno1:O gpo1:O gno2:O gpo2:O gno3:O gpo3:O nSEL2:O VPWR:I VGND:I
x1 SEL0 VGND VGND VPWR VPWR nSEL0 sky130_fd_sc_hd__inv_2
x2 SEL1 VGND VGND VPWR VPWR nSEL1 sky130_fd_sc_hd__inv_2
x7 nSEL0 nSEL1 VGND VGND VPWR VPWR gno0 sky130_fd_sc_hd__and2_1
x10 SEL1 SEL0 VGND VGND VPWR VPWR gno3 sky130_fd_sc_hd__and2_1
x11 gno0 VGND VGND VPWR VPWR gpo0 sky130_fd_sc_hd__inv_2
x12 gno1 VGND VGND VPWR VPWR gpo1 sky130_fd_sc_hd__inv_2
x13 gno2 VGND VGND VPWR VPWR gpo2 sky130_fd_sc_hd__inv_2
x14 gno3 VGND VGND VPWR VPWR gpo3 sky130_fd_sc_hd__inv_2
x15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x8 SEL1 SEL0 VGND VGND VPWR VPWR gno1 sky130_fd_sc_hd__and2b_1
x9 SEL0 SEL1 VGND VGND VPWR VPWR gno2 sky130_fd_sc_hd__and2b_1
x18 SEL2 VGND VGND VPWR VPWR nSEL2 sky130_fd_sc_hd__inv_2
x19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

.end
