* NGSPICE file created from passgate_parax.ext - technology: sky130A

.subckt passgate_parax Z A GP VSSBPIN VCCBPIN
X0 Z.t1 a_4022_n656# A.t0 VSSBPIN.t1 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X1 A.t2 GP.t0 Z.t2 VCCBPIN.t1 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X2 Z.t0 a_4022_n656# A.t1 VSSBPIN.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X3 A.t3 GP.t1 Z.t3 VCCBPIN.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
R0 A.n0 A.t3 26.3998
R1 A.n0 A.t2 23.5483
R2 A.n1 A.t0 12.7127
R3 A.n1 A.t1 10.8578
R4 A.n2 A.n0 3.06895
R5 A.n2 A.n1 1.84731
R6 A A.n2 1.18948
R7 Z.n1 Z.t2 23.6581
R8 Z.n0 Z.t3 23.3739
R9 Z.n1 Z.t0 10.7528
R10 Z.n3 Z.t1 10.6417
R11 Z.n2 Z.n1 1.30064
R12 Z Z.n4 0.958687
R13 Z.n2 Z.n0 0.726502
R14 Z.n3 Z.n2 0.512491
R15 Z.n4 Z.n3 0.359663
R16 Z.n4 Z.n0 0.216071
R17 VSSBPIN.n6 VSSBPIN.n4 11744.7
R18 VSSBPIN.n8 VSSBPIN.n4 11744.7
R19 VSSBPIN.n8 VSSBPIN.n3 11744.7
R20 VSSBPIN.n6 VSSBPIN.n3 11744.7
R21 VSSBPIN.t1 VSSBPIN.n3 8583.05
R22 VSSBPIN.t0 VSSBPIN.n4 8583.05
R23 VSSBPIN.n7 VSSBPIN.t1 7967.33
R24 VSSBPIN.n7 VSSBPIN.t0 7967.33
R25 VSSBPIN.n5 VSSBPIN.n2 763.09
R26 VSSBPIN.n5 VSSBPIN.n0 732.236
R27 VSSBPIN.n9 VSSBPIN.n2 304.553
R28 VSSBPIN.n10 VSSBPIN.n9 266.349
R29 VSSBPIN.n3 VSSBPIN.n2 195
R30 VSSBPIN.n4 VSSBPIN.n1 195
R31 VSSBPIN.n10 VSSBPIN.n1 54.2123
R32 VSSBPIN.n1 VSSBPIN.n0 30.8711
R33 VSSBPIN.n6 VSSBPIN.n5 11.0382
R34 VSSBPIN.n7 VSSBPIN.n6 11.0382
R35 VSSBPIN.n9 VSSBPIN.n8 11.0382
R36 VSSBPIN.n8 VSSBPIN.n7 11.0382
R37 VSSBPIN.n11 VSSBPIN.n0 10.4476
R38 VSSBPIN VSSBPIN.n11 7.23036
R39 VSSBPIN.n11 VSSBPIN.n10 3.78485
R40 GP.n0 GP.t1 450.938
R41 GP.n0 GP.t0 445.666
R42 GP GP.n0 3.23793
R43 VCCBPIN.n8 VCCBPIN.n2 8629.41
R44 VCCBPIN.n8 VCCBPIN.n3 8629.41
R45 VCCBPIN.n6 VCCBPIN.n2 8629.41
R46 VCCBPIN.n6 VCCBPIN.n3 8629.41
R47 VCCBPIN.n8 VCCBPIN.t0 2459.29
R48 VCCBPIN.t1 VCCBPIN.n6 2459.29
R49 VCCBPIN.t0 VCCBPIN.n7 2298.92
R50 VCCBPIN.n7 VCCBPIN.t1 2298.92
R51 VCCBPIN.n5 VCCBPIN.n4 920.471
R52 VCCBPIN.n4 VCCBPIN.n0 914.447
R53 VCCBPIN.n5 VCCBPIN.n1 480.764
R54 VCCBPIN.n10 VCCBPIN.n1 379.2
R55 VCCBPIN.n11 VCCBPIN.n0 105.788
R56 VCCBPIN.n10 VCCBPIN.n9 63.3551
R57 VCCBPIN.n6 VCCBPIN.n5 61.6672
R58 VCCBPIN.n9 VCCBPIN.n8 61.6672
R59 VCCBPIN VCCBPIN.n11 7.60782
R60 VCCBPIN.n9 VCCBPIN.n0 6.02403
R61 VCCBPIN.n11 VCCBPIN.n10 5.18145
R62 VCCBPIN.n3 VCCBPIN.n1 2.84665
R63 VCCBPIN.n7 VCCBPIN.n3 2.84665
R64 VCCBPIN.n4 VCCBPIN.n2 2.84665
R65 VCCBPIN.n7 VCCBPIN.n2 2.84665
C0 Z a_4022_n656# 0.415547f
C1 VCCBPIN a_4022_n656# 0.06934f
C2 GP A 3.81669f
C3 Z GP 0.278468f
C4 VCCBPIN GP 1.13434f
C5 a_4022_n656# GP 0.092899f
C6 Z A 4.51796f
C7 VCCBPIN A 1.49242f
C8 Z VCCBPIN 2.3841f
C9 a_4022_n656# A 3.41074f
C10 Z VSSBPIN 2.587317f
C11 GP VSSBPIN 2.214785f
C12 A VSSBPIN 4.20282f
C13 VCCBPIN VSSBPIN 9.990746f
C14 a_4022_n656# VSSBPIN 2.75176f
C15 VCCBPIN.n0 VSSBPIN 0.041049f
C16 VCCBPIN.n1 VSSBPIN 0.13325f
C17 VCCBPIN.n2 VSSBPIN 0.064566f
C18 VCCBPIN.n3 VSSBPIN 0.064566f
C19 VCCBPIN.n4 VSSBPIN 0.064356f
C20 VCCBPIN.n5 VSSBPIN 0.089219f
C21 VCCBPIN.n6 VSSBPIN 0.287635f
C22 VCCBPIN.t1 VSSBPIN 0.415127f
C23 VCCBPIN.n7 VSSBPIN 0.400805f
C24 VCCBPIN.t0 VSSBPIN 0.415127f
C25 VCCBPIN.n8 VSSBPIN 0.287635f
C26 VCCBPIN.n9 VSSBPIN 0.002528f
C27 VCCBPIN.n10 VSSBPIN 0.070642f
C28 VCCBPIN.n11 VSSBPIN 0.021449f
C29 GP.t0 VSSBPIN 0.508073f
C30 GP.t1 VSSBPIN 0.522241f
C31 GP.n0 VSSBPIN 1.91856f
C32 Z.t3 VSSBPIN 0.452527f
C33 Z.n0 VSSBPIN 0.562808f
C34 Z.t2 VSSBPIN 0.464987f
C35 Z.t0 VSSBPIN 0.350399f
C36 Z.n1 VSSBPIN 2.34646f
C37 Z.n2 VSSBPIN 0.793945f
C38 Z.t1 VSSBPIN 0.343504f
C39 Z.n3 VSSBPIN 0.512912f
C40 Z.n4 VSSBPIN 0.705679f
C41 A.t3 VSSBPIN 0.768569f
C42 A.t2 VSSBPIN 0.543692f
C43 A.n0 VSSBPIN 4.21525f
C44 A.t0 VSSBPIN 0.742571f
C45 A.t1 VSSBPIN 0.426296f
C46 A.n1 VSSBPIN 4.13493f
C47 A.n2 VSSBPIN 0.675541f
.ends

