* NGSPICE file created from tt_um_patdeegan_anamux_parax.ext - technology: sky130A

.subckt tt_um_patdeegan_anamux_parax clk ena rst_n ua[4] ua[5] ua[6] ua[7] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ ui_in[5] ua[0] ua[3] ui_in[1] ua[1] ui_in[4] ui_in[2] ui_in[6] ui_in[0] ua[2] ui_in[3]
+ VDPWR VSS
X0 a_21007_3867# ringtest_0.x4.net2.t2 VSS.t701 VSS.t700 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VSS.t445 VDPWR.t1166 VSS.t444 VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2 VSS.t447 VDPWR.t1167 VSS.t446 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3 a_24527_5340# a_24361_5340# VSS.t663 VSS.t662 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 ua[2].t15 muxtest_0.x2.x2.GP1.t4 ua[3].t9 VDPWR.t535 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X5 ringtest_0.x4.clknet_0_clk.t31 a_23879_6940# VSS.t1105 VSS.t1104 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_24135_3867# ringtest_0.x4.net6.t2 VDPWR.t250 VDPWR.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7 VSS.t656 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t31 VSS.t655 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VDPWR.t351 ui_in[1].t0 muxtest_0.x1.x1.nSEL1 VDPWR.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 a_22399_8976# a_21852_8720# a_22052_8875# VDPWR.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X10 muxtest_0.x1.x3.GP1.t1 muxtest_0.x1.x3.GN1 VDPWR.t345 VDPWR.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_27491_4566# ringtest_0.x4._23_ ringtest_0.x4._09_ VSS.t1114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X12 VSS.t607 a_27065_5156# a_27233_5058# VSS.t606 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VDPWR.t771 ringtest_0.x4._05_ a_24883_6800# VDPWR.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X14 VDPWR.t698 a_16579_11759# ringtest_0.x3.x2.GN3 VDPWR.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X15 VDPWR.t1159 VSS.t1127 VDPWR.t1158 VDPWR.t1157 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X16 a_25309_5334# a_24527_5340# a_25225_5334# VDPWR.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_12019_24012# muxtest_0.x2.x1.nSEL1 VSS.t309 VSS.t308 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X18 a_26913_4566# ringtest_0.x4._15_ a_26817_4566# VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X19 VSS.t1022 ringtest_0.x4._21_ a_24545_5878# VSS.t1021 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 muxtest_0.x1.x3.GP4.t1 muxtest_0.x1.x3.GN4 VDPWR.t775 VDPWR.t774 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR.t784 VDPWR.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 VDPWR.t34 ringtest_0.x4._15_ a_25925_6788# VDPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_24004_6128# ringtest_0.x4._17_ a_23932_6128# VDPWR.t821 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X24 VSS.t450 VDPWR.t1168 VSS.t449 VSS.t448 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X25 a_23467_4818# ringtest_0.x4._11_.t4 a_23381_4818# VSS.t908 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X26 a_19114_31955# a_19290_32287# a_19242_32347# VSS.t988 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 VSS.t452 VDPWR.t1169 VSS.t451 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X28 ringtest_0.x4.clknet_1_1__leaf_clk.t30 a_25364_5878# VSS.t654 VSS.t653 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 VDPWR.t1161 a_21375_3867# ringtest_0.x4.counter[1] VDPWR.t1160 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X30 VDPWR.t750 ringtest_0.x4.net5 a_22486_4246# VDPWR.t749 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X31 muxtest_0.x1.x1.nSEL0 ui_in[0].t0 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X32 VDPWR.t239 a_19842_32287# a_19666_31955# VDPWR.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X33 muxtest_0.R3R4.t7 muxtest_0.x2.x2.GN3 ua[2].t9 VSS.t684 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X34 VDPWR.t1156 VSS.t1128 VDPWR.t1155 VDPWR.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X35 a_12473_23980# ui_in[4].t0 VDPWR.t417 VDPWR.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X36 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP3 muxtest_0.R1R2.t3 VDPWR.t714 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X37 a_16579_11759# a_16755_12091# a_16707_12151# VSS.t904 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X38 VDPWR.t36 a_13501_23906# muxtest_0.x2.x2.GN4 VDPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X39 VDPWR.t716 a_19289_13081.t2 ringtest_0.drv_out.t8 VDPWR.t715 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X40 VSS.t3 a_21465_9294# ringtest_0.x4.net2.t0 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X41 ringtest_0.x4.clknet_0_clk.t15 a_23879_6940# VDPWR.t818 VDPWR.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X42 VDPWR.t680 a_22021_4220# ringtest_0.x4._03_ VDPWR.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
X43 VSS.t1031 ringtest_0.x4.net5 a_23467_4584# VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X44 muxtest_0.x2.nselect2 VDPWR.t708 VDPWR.t710 VDPWR.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X45 a_16707_12151# ui_in[4].t1 VSS.t665 VSS.t664 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X46 VSS.t455 VDPWR.t1170 VSS.t454 VSS.t453 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X47 VDPWR.t1153 VSS.t1129 VDPWR.t1152 VDPWR.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X48 ringtest_0.x4._15_ a_23381_4584# VSS.t1047 VSS.t496 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X49 a_23899_5334# ringtest_0.x4._15_ VDPWR.t32 VDPWR.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X50 VDPWR.t366 a_27065_5156# a_27233_5058# VDPWR.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X51 muxtest_0.x1.x3.GP3 muxtest_0.x1.x3.GN3 VDPWR.t759 VDPWR.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X52 VSS.t458 VDPWR.t1171 VSS.t457 VSS.t456 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X53 VSS.t711 ringtest_0.x4.net3.t2 ringtest_0.x4._12_ VSS.t710 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X54 VSS.t1046 a_25975_3867# ringtest_0.x4.counter[6] VSS.t1045 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X55 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk.t32 VDPWR.t538 VDPWR.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X56 muxtest_0.x1.x5.A ui_in[2].t0 ua[3].t10 VDPWR.t362 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X57 ua[1].t5 ringtest_0.x3.x2.GP4.t4 ringtest_0.counter7.t5 VDPWR.t363 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X58 a_22392_5990# a_22224_6244# VDPWR.t70 VDPWR.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X59 ringtest_0.x4.clknet_1_0__leaf_clk.t15 a_21395_6940# VDPWR.t318 VDPWR.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X60 VSS.t825 ringtest_0.x4._22_ a_26913_4566# VSS.t824 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X61 a_26640_5334# a_26367_5340# a_26555_5334# VDPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X62 ringtest_0.x4.clknet_1_1__leaf_clk.t15 a_25364_5878# VDPWR.t409 VDPWR.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X63 VDPWR.t1151 VSS.t1130 VDPWR.t1150 VDPWR.t1149 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X64 VSS.t461 VDPWR.t1172 VSS.t460 VSS.t459 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X65 a_21785_8054# ringtest_0.x4.net3.t3 VDPWR.t455 VDPWR.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X66 ringtest_0.x4._17_ a_25925_6788# VSS.t1049 VSS.t1048 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X67 VSS.t583 a_19114_31955# muxtest_0.x1.x3.GN2 VSS.t582 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VDPWR.t138 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X69 VDPWR.t707 VDPWR.t705 ringtest_0.x3.nselect2 VDPWR.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X70 VDPWR.t816 a_23879_6940# ringtest_0.x4.clknet_0_clk.t14 VDPWR.t815 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X71 VSS.t910 ringtest_0.x4.net4 ringtest_0.x4._13_ VSS.t909 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 a_24317_4942# ringtest_0.x4.net6.t3 a_24551_4790# VSS.t442 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X73 VSS.t790 ringtest_0.x4.clknet_0_clk.t32 a_25364_5878# VSS.t789 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X74 VSS.t396 a_22111_10993# ringtest_0.x4.net1 VSS.t395 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X75 VSS.t464 VDPWR.t1173 VSS.t463 VSS.t462 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X76 VDPWR.t353 a_27815_3867# ringtest_0.x4.counter[8] VDPWR.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X77 ringtest_0.x4._00_ a_21425_9686# a_21675_9686# VDPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X78 VDPWR.t1148 VSS.t1131 VDPWR.t1147 VDPWR.t1007 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X79 VDPWR.t1146 VSS.t1132 VDPWR.t1145 VDPWR.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X80 VDPWR.t215 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X81 VDPWR.t282 ringtest_0.x4._00_ a_22399_9142# VDPWR.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X82 VSS.t1103 a_23879_6940# ringtest_0.x4.clknet_0_clk.t30 VSS.t1102 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X83 a_21675_4790# a_21509_4790# VSS.t747 VSS.t746 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X84 VSS.t299 ui_in[0].t1 a_19842_32287# VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X85 VSS.t467 VDPWR.t1174 VSS.t466 VSS.t465 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X86 VDPWR.t316 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t14 VDPWR.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X87 VSS.t73 a_23399_3867# ringtest_0.counter3.t1 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X88 VDPWR.t119 a_18662_32213# muxtest_0.x1.x3.GN1 VDPWR.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X89 VDPWR.t445 ringtest_0.x4.net2.t3 a_21507_9686# VDPWR.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 VDPWR.t1143 VSS.t1133 VDPWR.t1142 VDPWR.t1141 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X91 a_27659_4246# ringtest_0.x4.net11 VDPWR.t377 VDPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X92 a_22390_4566# ringtest_0.x4.net5 VSS.t1030 VSS.t1029 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X93 ringtest_0.x3.x1.nSEL1 ui_in[4].t2 VSS.t667 VSS.t666 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X94 ringtest_0.x4.clknet_1_0__leaf_clk.t31 a_21395_6940# VSS.t557 VSS.t556 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X95 a_22649_6244# a_21785_5878# a_22392_5990# VDPWR.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X96 muxtest_0.x1.x3.GP2.t1 muxtest_0.x1.x3.GN2 VDPWR.t134 VDPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X97 ua[3].t11 ui_in[2].t1 muxtest_0.x1.x4.A VSS.t604 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X98 muxtest_0.R5R6.t5 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A VSS.t1042 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X99 VSS.t431 a_24329_6640# a_24336_6544# VSS.t430 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X100 a_27303_4246# a_27273_4220# ringtest_0.x4._09_ VDPWR.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X101 VDPWR.t1140 VSS.t1134 VDPWR.t1139 VDPWR.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X102 ringtest_0.x4.clknet_1_0__leaf_clk.t13 a_21395_6940# VDPWR.t314 VDPWR.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X103 VSS.t699 ringtest_0.x4.net2.t4 a_21425_9686# VSS.t698 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X104 a_19666_31955# a_19842_32287# a_19794_32347# VSS.t432 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X105 muxtest_0.R3R4.t5 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A VSS.t591 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X106 VDPWR.t357 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X107 a_21845_8816# ringtest_0.x4.clknet_1_0__leaf_clk.t32 VDPWR.t87 VDPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X108 VSS.t555 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t30 VSS.t554 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X109 a_21672_5334# a_21399_5340# a_21587_5334# VDPWR.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X110 ringtest_0.x4.clknet_1_1__leaf_clk.t14 a_25364_5878# VDPWR.t407 VDPWR.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X111 VDPWR.t1137 VSS.t1135 VDPWR.t1136 VDPWR.t1135 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X112 a_18662_32213# muxtest_0.x1.x1.nSEL0 a_18836_32319# VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X113 a_16203_12091# ui_in[4].t3 VDPWR.t419 VDPWR.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X114 a_19794_32347# ui_in[1].t1 VSS.t688 VSS.t687 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X115 VDPWR.t1134 VSS.t1136 VDPWR.t1133 VDPWR.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X116 VDPWR.t93 a_22817_6146# a_22733_6244# VDPWR.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X117 VDPWR.t144 a_17231_12017# ringtest_0.x3.x2.GN4 VDPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X118 VDPWR.t814 a_23879_6940# ringtest_0.x4.clknet_0_clk.t13 VDPWR.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X119 VSS.t652 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t29 VSS.t651 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X120 ringtest_0.x3.nselect2 VDPWR.t702 VDPWR.t704 VDPWR.t703 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X121 a_25925_6788# ringtest_0.x4.net6.t4 VDPWR.t726 VDPWR.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X122 a_25975_3867# ringtest_0.x4.net8 VDPWR.t84 VDPWR.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X123 ringtest_0.x4.net10 a_27233_5308# VDPWR.t125 VDPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X124 a_11845_23906# muxtest_0.x2.x1.nSEL1 VDPWR.t117 VDPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X125 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VSS.t757 VSS.t756 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X126 VDPWR.t551 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X127 a_21939_8054# ringtest_0.x4.net3.t4 a_21867_8054# VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X128 a_26721_4246# ringtest_0.x4.net10 a_26627_4246# VDPWR.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X129 a_22116_4902# a_21948_5156# VSS.t292 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X130 VDPWR.t312 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t12 VDPWR.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X131 a_25149_4220# ringtest_0.x4.net7 VDPWR.t671 VDPWR.t670 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X132 VDPWR.t546 a_21840_5308# a_21767_5334# VDPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X133 VSS.t470 VDPWR.t1175 VSS.t469 VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X134 VSS.t473 VDPWR.t1176 VSS.t472 VSS.t471 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X135 VDPWR.t585 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR.t584 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X136 VDPWR.t1131 VSS.t1137 VDPWR.t1130 VDPWR.t1129 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X137 a_24627_6200# ringtest_0.x4._21_ VDPWR.t734 VDPWR.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X138 VSS.t130 ringtest_0.x4._16_.t2 a_24986_5878# VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.06615 ps=0.735 w=0.42 l=0.15
X139 VSS.t476 VDPWR.t1177 VSS.t475 VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X140 VDPWR.t14 a_22245_8054# ringtest_0.x4._11_.t1 VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X141 a_25977_4220# ringtest_0.x4._11_.t5 VDPWR.t487 VDPWR.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X142 VSS.t479 VDPWR.t1178 VSS.t478 VSS.t477 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X143 a_26367_4790# a_26201_4790# VSS.t436 VSS.t435 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X144 VDPWR.t1128 VSS.t1138 VDPWR.t1127 VDPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X145 a_25677_5156# a_24895_4790# a_25593_5156# VDPWR.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 VDPWR.t820 ringtest_0.x4._17_ a_23349_6422# VDPWR.t819 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 VDPWR.t30 ringtest_0.x4._15_ a_25977_4220# VDPWR.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X148 VDPWR.t1126 VSS.t1139 VDPWR.t1125 VDPWR.t903 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X149 VDPWR.t534 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2.t1 VDPWR.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X150 VDPWR.t570 a_24070_5852# a_24004_6128# VDPWR.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X151 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP2.t4 muxtest_0.R6R7.t3 VDPWR.t49 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X152 ua[0].t4 muxtest_0.x2.x2.GN2 ua[2].t11 VSS.t767 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X153 VSS.t848 a_25977_4220# ringtest_0.x4._23_ VSS.t847 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X154 VDPWR.t1124 VSS.t1140 VDPWR.t1123 VDPWR.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X155 VDPWR.t1121 VSS.t1141 VDPWR.t1120 VDPWR.t1119 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X156 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VSS.t334 VSS.t333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X157 VDPWR.t324 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X158 a_21425_9686# ringtest_0.x4.net1 VSS.t403 VSS.t402 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X159 VSS.t109 a_24317_4942# ringtest_0.x4._20_ VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X160 muxtest_0.x1.x1.nSEL1 ui_in[1].t2 VDPWR.t433 VDPWR.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X161 a_21465_8830# a_21561_8830# VSS.t376 VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X162 ringtest_0.x4.clknet_0_clk.t29 a_23879_6940# VSS.t1101 VSS.t1100 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X163 a_22295_3867# ringtest_0.x4.net4 VDPWR.t640 VDPWR.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X164 muxtest_0.R7R8.t9 muxtest_0.R6R7.t5 VSS.t419 sky130_fd_pr__res_high_po_1p41 l=1.75
X165 VDPWR.t1118 VSS.t1142 VDPWR.t1117 VDPWR.t1116 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X166 a_26808_4902# a_26640_5156# VDPWR.t271 VDPWR.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X167 VSS.t482 VDPWR.t1179 VSS.t481 VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X168 ringtest_0.x4.clknet_1_1__leaf_clk.t13 a_25364_5878# VDPWR.t405 VDPWR.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X169 VSS.t384 a_26808_5308# a_26766_5712# VSS.t383 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X170 a_25351_5712# a_24361_5340# a_25225_5334# VSS.t661 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X171 VSS.t553 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t29 VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X172 VSS.t485 VDPWR.t1180 VSS.t484 VSS.t483 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X173 muxtest_0.R7R8.t4 muxtest_0.x2.x2.GN4 ua[2].t7 VSS.t425 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X174 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VSS.t407 VSS.t406 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X175 VSS.t488 VDPWR.t1181 VSS.t487 VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X176 a_21007_3867# ringtest_0.x4.net2.t5 VDPWR.t443 VDPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X177 ringtest_0.x4.net4 a_22265_5308# VDPWR.t196 VDPWR.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X178 VDPWR.t616 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X179 VSS.t1004 a_19289_13081.t3 ringtest_0.drv_out.t16 VSS.t1003 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X180 a_22373_5156# a_21509_4790# a_22116_4902# VDPWR.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X181 VDPWR.t1115 VSS.t1143 VDPWR.t1114 VDPWR.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X182 a_26895_3867# ringtest_0.x4.net9 VSS.t364 VSS.t363 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X183 a_27191_4790# a_26201_4790# a_27065_5156# VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X184 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR.t219 VDPWR.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X185 VDPWR.t1113 VSS.t1144 VDPWR.t1112 VDPWR.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X186 VSS.t491 VDPWR.t1182 VSS.t490 VSS.t489 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X187 a_22116_4902# a_21948_5156# VDPWR.t98 VDPWR.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X188 VSS.t124 ringtest_0.x4.net8 a_23837_5878# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X189 VDPWR.t310 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t11 VDPWR.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X190 a_16755_12091# ui_in[3].t0 VDPWR.t648 VDPWR.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X191 VDPWR.t403 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t12 VDPWR.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X192 VDPWR.t778 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 VDPWR.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X193 ringtest_0.x4.clknet_1_0__leaf_clk.t28 a_21395_6940# VSS.t551 VSS.t550 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X194 VSS.t22 VDPWR.t1183 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X195 VSS.t503 a_21007_3867# ringtest_0.x4.counter[0] VSS.t502 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X196 a_22181_5334# a_21399_5340# a_22097_5334# VDPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X197 a_20318_32213# ui_in[1].t3 a_20492_32319# VSS.t689 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X198 VSS.t521 ringtest_0.x4._00_ a_22399_9142# VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X199 a_22224_6244# a_21951_5878# a_22139_5878# VDPWR.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X200 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VSS.t761 VSS.t756 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X201 VSS.t840 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1.t3 VSS.t839 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X202 VDPWR.t748 ringtest_0.x4.net5 a_23381_4584# VDPWR.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X203 a_26555_5334# ringtest_0.x4._08_ VSS.t350 VSS.t349 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X204 ua[2].t3 muxtest_0.x2.x2.GP3 muxtest_0.R3R4.t1 VDPWR.t76 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X205 a_16027_11759# ui_in[3].t1 VDPWR.t458 VDPWR.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X206 VDPWR.t115 a_22541_5058# a_22457_5156# VDPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X207 ringtest_0.x4.clknet_1_1__leaf_clk.t28 a_25364_5878# VSS.t650 VSS.t649 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X208 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VSS.t599 VSS.t566 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X209 ringtest_0.x4._19_ a_23529_6422# VSS.t392 VSS.t391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X210 a_26569_6422# ringtest_0.x4._23_ VSS.t1113 VSS.t1112 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X211 a_24895_4790# a_24729_4790# VDPWR.t560 VDPWR.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X212 VDPWR.t530 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 ringtest_0.ring_out.t3 ringtest_0.x3.x2.GN1 ua[1].t13 VSS.t838 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X214 ringtest_0.drv_out.t15 a_19289_13081.t4 VSS.t1006 VSS.t1005 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X215 a_23899_5334# ringtest_0.x4.net6.t5 VDPWR.t728 VDPWR.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X216 VDPWR.t1111 VSS.t1145 VDPWR.t1110 VDPWR.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X217 a_24045_6654# a_24336_6544# a_24287_6422# VDPWR.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X218 a_24800_5334# a_24527_5340# a_24715_5334# VDPWR.t829 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X219 muxtest_0.R7R8.t6 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A VSS.t590 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X220 muxtest_0.x2.x2.GP3 muxtest_0.x2.x2.GN3 VSS.t683 VSS.t682 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X221 VSS.t25 VDPWR.t1184 VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X222 a_25925_6788# ringtest_0.x4._11_.t6 VDPWR.t489 VDPWR.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X223 ringtest_0.x4.net10 a_27233_5308# VSS.t317 VSS.t316 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X224 VSS.t771 a_21840_5308# a_21798_5712# VSS.t770 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X225 VSS.t716 ui_in[3].t2 muxtest_0.x2.x1.nSEL0 VSS.t715 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X226 VDPWR.t1108 VSS.t1146 VDPWR.t1107 VDPWR.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X227 VDPWR.t72 a_22392_5990# a_22319_6244# VDPWR.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X228 VSS.t28 VDPWR.t1185 VSS.t27 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X229 VSS.t707 a_15575_12017# ringtest_0.x3.x2.GN1 VSS.t706 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X230 a_22201_9142# a_21981_9142# VSS.t1034 VSS.t961 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X231 ringtest_0.counter7.t1 ringtest_0.x3.x2.GN4 ua[1].t2 VSS.t346 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X232 VDPWR.t669 ringtest_0.x4.net7 a_25925_6788# VDPWR.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X233 VDPWR.t761 a_25975_3867# ringtest_0.x4.counter[6] VDPWR.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X234 VSS.t737 ringtest_0.x4.clknet_0_clk.t33 a_25364_5878# VSS.t736 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X235 VDPWR.t1106 VSS.t1147 VDPWR.t1105 VDPWR.t1104 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X236 VSS.t739 ringtest_0.x4.clknet_0_clk.t34 a_21395_6940# VSS.t738 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X237 a_19114_31955# ui_in[0].t2 VDPWR.t108 VDPWR.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X238 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VSS.t1051 VSS.t333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X239 VDPWR.t1103 VSS.t1148 VDPWR.t1102 VDPWR.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X240 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR.t614 VDPWR.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X241 VDPWR.t591 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2.t1 VDPWR.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X242 VDPWR.t89 ringtest_0.x4.clknet_1_0__leaf_clk.t33 a_21509_4790# VDPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X243 VDPWR.t1100 VSS.t1149 VDPWR.t1099 VDPWR.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X244 a_21803_9508# a_21465_9294# VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X245 a_22052_9116# a_21852_9416# a_22201_9142# VSS.t617 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X246 VSS.t31 VDPWR.t1186 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X247 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VSS.t778 VSS.t406 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X248 ringtest_0.x4._12_ ringtest_0.x4.net2.t6 a_21132_8918# VSS.t697 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X249 a_22052_8875# a_21852_8720# a_22201_8964# VSS.t617 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X250 a_27065_5156# a_26201_4790# a_26808_4902# VDPWR.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X251 ringtest_0.x4.clknet_1_0__leaf_clk.t27 a_21395_6940# VSS.t549 VSS.t548 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X252 a_21587_5334# ringtest_0.x4._02_ VSS.t814 VSS.t813 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X253 VSS.t301 ui_in[0].t3 muxtest_0.x1.x1.nSEL0 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X254 VSS.t34 VDPWR.t1187 VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X255 VDPWR.t1 a_21465_9294# ringtest_0.x4.net2.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X256 ringtest_0.x4._25_ a_26749_6422# VDPWR.t7 VDPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X257 VDPWR.t22 a_23399_3867# ringtest_0.counter3.t0 VDPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X258 VDPWR.t401 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t11 VDPWR.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X259 muxtest_0.x2.x2.GP2.t3 muxtest_0.x2.x2.GN2 VSS.t766 VSS.t765 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X260 ringtest_0.x3.x2.GP1.t2 ringtest_0.x3.x2.GN1 VSS.t837 VSS.t836 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X261 VSS.t37 VDPWR.t1188 VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X262 VDPWR.t1098 VSS.t1150 VDPWR.t1097 VDPWR.t988 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X263 a_26817_4566# ringtest_0.x4._11_.t7 a_26627_4246# VSS.t729 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X264 a_22649_6244# a_21951_5878# a_22392_5990# VSS.t751 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X265 VDPWR.t757 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 VDPWR.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X266 VDPWR.t1096 VSS.t1151 VDPWR.t1095 VDPWR.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X267 VSS.t759 a_21845_9116# a_21852_9416# VSS.t523 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X268 a_21591_6128# ringtest_0.x4._11_.t8 ringtest_0.x4._13_ VDPWR.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X269 VDPWR.t28 ringtest_0.x4._15_ a_23381_4818# VDPWR.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X270 a_21981_9142# a_21845_9116# a_21561_9116# VDPWR.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X271 VDPWR.t1094 VSS.t1152 VDPWR.t1093 VDPWR.t1092 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X272 VSS.t648 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t27 VSS.t647 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X273 VSS.t589 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1.t3 VSS.t588 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X274 muxtest_0.R6R7.t1 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A VSS.t330 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X275 VDPWR.t1091 VSS.t1153 VDPWR.t1090 VDPWR.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X276 ringtest_0.x4.clknet_0_clk.t28 a_23879_6940# VSS.t1099 VSS.t1098 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X277 VDPWR.t828 a_27233_5058# a_27149_5156# VDPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X278 VDPWR.t1088 VSS.t1154 VDPWR.t1087 VDPWR.t1086 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X279 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VSS.t567 VSS.t566 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X280 VDPWR.t1085 VSS.t1155 VDPWR.t1084 VDPWR.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X281 ringtest_0.x4.clknet_1_1__leaf_clk.t10 a_25364_5878# VDPWR.t399 VDPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X282 a_26839_6788# a_26569_6422# a_26749_6422# VSS.t758 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X283 VSS.t40 VDPWR.t1189 VSS.t39 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X284 VSS.t547 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t26 VSS.t546 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X285 VSS.t43 VDPWR.t1190 VSS.t42 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X286 ringtest_0.x4.net8 a_25393_5308# VDPWR.t190 VDPWR.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X287 VSS.t1061 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP4.t3 VSS.t1060 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X288 a_24479_4790# ringtest_0.x4.net8 VSS.t122 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X289 ringtest_0.x4.net9 a_25761_5058# VSS.t579 VSS.t578 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X290 a_27191_5712# a_26201_5340# a_27065_5334# VSS.t573 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X291 VSS.t1111 ringtest_0.x4._23_ a_27273_4220# VSS.t1110 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X292 a_25593_5156# a_24895_4790# a_25336_4902# VSS.t336 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X293 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR.t583 VDPWR.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X294 VSS.t624 ringtest_0.x4.net11 a_27489_3702# VSS.t623 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X295 ringtest_0.drv_out.t14 a_19289_13081.t5 VSS.t1008 VSS.t1007 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X296 ringtest_0.x3.x2.GP3 ringtest_0.x3.x2.GN3 VSS.t1067 VSS.t1066 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X297 VSS.t46 VDPWR.t1191 VSS.t45 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X298 ringtest_0.counter3.t5 ringtest_0.x3.x2.GN3 ua[1].t15 VSS.t1065 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X299 ringtest_0.x4.clknet_0_clk.t12 a_23879_6940# VDPWR.t812 VDPWR.t811 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X300 a_24699_6200# ringtest_0.x4.net9 a_24627_6200# VDPWR.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0441 ps=0.63 w=0.42 l=0.15
X301 VSS.t49 VDPWR.t1192 VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X302 VDPWR.t1082 VSS.t1156 VDPWR.t1081 VDPWR.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X303 VSS.t51 VDPWR.t1193 muxtest_0.x2.nselect2 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X304 ringtest_0.x4.clknet_1_0__leaf_clk.t25 a_21395_6940# VSS.t545 VSS.t544 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X305 a_24264_6788# a_23949_6654# VSS.t417 VSS.t416 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X306 VSS.t501 a_24135_3867# ringtest_0.x4.counter[4] VSS.t500 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X307 VSS.t54 VDPWR.t1194 VSS.t53 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X308 VDPWR.t540 ringtest_0.x4.clknet_1_1__leaf_clk.t33 a_26201_4790# VDPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X309 a_21465_8830# a_21561_8830# VDPWR.t182 VDPWR.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X310 a_19666_31955# ui_in[1].t4 VDPWR.t435 VDPWR.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X311 VDPWR.t132 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2.t0 VDPWR.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X312 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP2.t5 muxtest_0.R6R7.t2 VDPWR.t246 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X313 ua[0].t8 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A VSS.t1059 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X314 ringtest_0.x4.net5 a_22541_5058# VSS.t307 VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X315 VSS.t681 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 VSS.t680 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X316 VDPWR.t198 a_16027_11759# ringtest_0.x3.x2.GN2 VDPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X317 VDPWR.t397 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t9 VDPWR.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X318 VSS.t57 VDPWR.t1195 VSS.t56 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X319 a_21395_6940# ringtest_0.x4.clknet_0_clk.t35 VSS.t741 VSS.t740 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X320 a_23949_6654# a_24045_6654# VDPWR.t604 VDPWR.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X321 VDPWR.t542 ringtest_0.x4.clknet_1_1__leaf_clk.t34 a_24361_5340# VDPWR.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X322 VDPWR.t696 a_23770_5308# ringtest_0.x4._18_ VDPWR.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X323 VSS.t992 a_22765_4478# ringtest_0.x4._14_ VSS.t991 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X324 VDPWR.t171 ringtest_0.ring_out.t10 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X325 VSS.t990 ringtest_0.x4._10_ a_22245_8054# VSS.t989 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X326 a_21675_10006# ringtest_0.x4.net2.t7 VSS.t696 VSS.t695 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X327 VSS.t609 a_22052_8875# a_21981_8976# VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X328 ringtest_0.x4.net9 a_25761_5058# VDPWR.t337 VDPWR.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X329 VDPWR.t1080 VSS.t1157 VDPWR.t1079 VDPWR.t1078 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X330 VSS.t726 a_19289_13081.t6 ringtest_0.drv_out.t13 VSS.t725 sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X331 VSS.t427 a_24968_5308# a_24926_5712# VSS.t426 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X332 VSS.t691 ui_in[1].t5 muxtest_0.x1.x1.nSEL1 VSS.t690 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X333 muxtest_0.x1.x3.GP1.t2 muxtest_0.x1.x3.GN1 VSS.t587 VSS.t586 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X334 a_16027_11759# a_16203_12091# a_16155_12151# VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X335 ringtest_0.x4.clknet_0_clk.t27 a_23879_6940# VSS.t1097 VSS.t1096 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X336 VDPWR.t211 ringtest_0.x4.net1 a_21049_8598# VDPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X337 VDPWR.t1077 VSS.t1158 VDPWR.t1076 VDPWR.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X338 VSS.t60 VDPWR.t1196 VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X339 VSS.t850 a_20318_32213# muxtest_0.x1.x3.GN4 VSS.t849 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X340 muxtest_0.x2.x1.nSEL0 ui_in[3].t3 VDPWR.t460 VDPWR.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X341 a_16155_12151# ui_in[3].t4 VSS.t718 VSS.t717 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X342 a_26269_4612# ringtest_0.x4._15_ a_26173_4612# VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X343 VDPWR.t1074 VSS.t1159 VDPWR.t1073 VDPWR.t1072 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X344 VDPWR.t1071 VSS.t1160 VDPWR.t1070 VDPWR.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X345 VSS.t543 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t24 VSS.t542 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X346 a_25149_4220# ringtest_0.x4.net9 VDPWR.t164 VDPWR.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X347 a_22223_5712# a_21233_5340# a_22097_5334# VSS.t1126 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X348 muxtest_0.x1.x3.GP4.t2 muxtest_0.x1.x3.GN4 VSS.t1058 VSS.t1057 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X349 VSS.t62 VDPWR.t1197 VSS.t61 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X350 VSS.t65 VDPWR.t1198 VSS.t64 VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X351 ringtest_0.x4.net5 a_22541_5058# VDPWR.t113 VDPWR.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X352 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR.t322 VDPWR.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X353 VSS.t68 VDPWR.t1199 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X354 VSS.t735 ringtest_0.x4._11_.t9 ringtest_0.x4._01_ VSS.t734 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X355 a_22765_5308# ringtest_0.x4._16_.t3 a_23151_5334# VDPWR.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X356 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP1.t4 muxtest_0.R7R8.t8 VDPWR.t659 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X357 a_25977_4220# ringtest_0.x4._22_ VDPWR.t597 VDPWR.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X358 a_25083_4790# ringtest_0.x4._07_ VDPWR.t544 VDPWR.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X359 VSS.t71 VDPWR.t1200 VSS.t70 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X360 VDPWR.t1068 VSS.t1161 VDPWR.t1067 VDPWR.t1066 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X361 a_22983_5654# ringtest_0.x4._16_.t4 ringtest_0.x4._04_ VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X362 VSS.t244 VDPWR.t1201 VSS.t243 VSS.t242 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X363 VDPWR.t462 ui_in[3].t5 ringtest_0.x3.x1.nSEL0 VDPWR.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X364 a_23879_6940# ringtest_0.drv_out.t20 VDPWR.t63 VDPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X365 a_22164_4362# ringtest_0.x4._16_.t5 VSS.t1010 VSS.t1009 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X366 a_25168_5156# a_24729_4790# a_25083_4790# VSS.t782 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X367 VDPWR.t1065 VSS.t1162 VDPWR.t1064 VDPWR.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X368 VSS.t115 a_22392_5990# a_22350_5878# VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X369 VDPWR.t150 ringtest_0.x4._20_ a_23809_4790# VDPWR.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X370 muxtest_0.x2.nselect2 VDPWR.t1202 VSS.t246 VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X371 a_21780_8964# a_21465_8830# VSS.t378 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X372 ringtest_0.x4._11_.t3 a_22245_8054# VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X373 a_26895_3867# ringtest_0.x4.net9 VDPWR.t162 VDPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X374 a_24715_5334# ringtest_0.x4._06_ VSS.t808 VSS.t807 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X375 VSS.t248 VDPWR.t1203 VSS.t247 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X376 VDPWR.t502 ringtest_0.x4._11_.t10 a_23899_5334# VDPWR.t501 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X377 VDPWR.t395 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t8 VDPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X378 VDPWR.t269 a_25421_6641# ringtest_0.x4._05_ VDPWR.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X379 muxtest_0.x1.x3.GP3 muxtest_0.x1.x3.GN3 VSS.t1041 VSS.t1040 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X380 muxtest_0.x1.x4.A muxtest_0.x1.x5.GN ua[3].t5 VDPWR.t547 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X381 ua[2].t14 muxtest_0.x2.x2.GP1.t5 ua[3].t8 VDPWR.t536 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X382 ua[0].t3 muxtest_0.x2.x2.GN2 ua[2].t10 VSS.t764 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X383 a_25294_4790# a_24895_4790# a_25168_5156# VSS.t335 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X384 a_21863_4790# ringtest_0.x4._03_ VDPWR.t682 VDPWR.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X385 VDPWR.t1062 VSS.t1163 VDPWR.t1061 VDPWR.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X386 VDPWR.t261 a_21007_3867# ringtest_0.x4.counter[0] VDPWR.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X387 VSS.t251 VDPWR.t1204 VSS.t250 VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X388 a_21948_5156# a_21509_4790# a_21863_4790# VSS.t745 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X389 VSS.t254 VDPWR.t1205 VSS.t253 VSS.t252 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X390 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.ring_out.t11 VDPWR.t173 VDPWR.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X391 VSS.t622 ringtest_0.x4.net11 a_27491_4566# VSS.t621 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X392 ringtest_0.x4.net11 a_27233_5058# VSS.t1118 VSS.t1117 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X393 ringtest_0.x4._21_ a_23809_4790# VDPWR.t158 VDPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X394 VSS.t332 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VSS.t331 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X395 VSS.t256 VDPWR.t1206 ringtest_0.x3.nselect2 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X396 VDPWR.t676 ringtest_0.x4._01_ a_22399_8976# VDPWR.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X397 VDPWR.t810 a_23879_6940# ringtest_0.x4.clknet_0_clk.t11 VDPWR.t809 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X398 a_25149_4220# ringtest_0.x4.net6.t6 a_25547_4612# VSS.t1015 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X399 ringtest_0.x4.net8 a_25393_5308# VSS.t382 VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X400 VSS.t9 a_21425_9686# ringtest_0.x4._00_ VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X401 VSS.t581 a_25336_4902# a_25294_4790# VSS.t580 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X402 VDPWR.t808 a_23879_6940# ringtest_0.x4.clknet_0_clk.t10 VDPWR.t807 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X403 ua[2].t0 muxtest_0.x2.x2.GP4.t4 muxtest_0.R7R8.t0 VDPWR.t4 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X404 a_22139_5878# ringtest_0.x4._04_ VSS.t806 VSS.t805 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X405 ringtest_0.x3.x2.GP2.t0 ringtest_0.x3.x2.GN2 VDPWR.t589 VDPWR.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X406 ringtest_0.x4.clknet_0_clk.t26 a_23879_6940# VSS.t1095 VSS.t1094 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X407 a_25977_4220# ringtest_0.x4.net10 a_26375_4612# VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X408 VSS.t259 VDPWR.t1207 VSS.t258 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X409 VSS.t508 a_25421_6641# ringtest_0.x4._05_ VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X410 VDPWR.t678 ringtest_0.x4._24_ a_26749_6422# VDPWR.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X411 VSS.t107 ringtest_0.x4.clknet_1_0__leaf_clk.t34 a_21785_5878# VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X412 VSS.t405 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VSS.t404 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 VDPWR.t481 a_19289_13081.t7 ringtest_0.drv_out.t7 VDPWR.t480 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X414 a_22021_4220# a_22164_4362# VDPWR.t280 VDPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X415 VDPWR.t217 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X416 VSS.t262 VDPWR.t1208 VSS.t261 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X417 VDPWR.t504 ringtest_0.x4._11_.t11 a_23809_4790# VDPWR.t503 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X418 ua[3].t6 muxtest_0.x2.x2.GN1 ua[2].t13 VSS.t968 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X419 VDPWR.t1060 VSS.t1164 VDPWR.t1059 VDPWR.t1058 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X420 a_19242_32347# ui_in[0].t4 VSS.t303 VSS.t302 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X421 muxtest_0.x1.x3.GP2.t3 muxtest_0.x1.x3.GN2 VSS.t329 VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X422 ringtest_0.x4.clknet_1_0__leaf_clk.t23 a_21395_6940# VSS.t541 VSS.t540 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X423 VSS.t982 ringtest_0.x4._24_ a_26839_6788# VSS.t981 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X424 VDPWR.t59 ringtest_0.x4.clknet_1_0__leaf_clk.t35 a_21785_5878# VDPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X425 VSS.t728 a_19289_13081.t8 ringtest_0.drv_out.t12 VSS.t727 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X426 VDPWR.t1057 VSS.t1165 VDPWR.t1056 VDPWR.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X427 ringtest_0.x4.net11 a_27233_5058# VDPWR.t827 VDPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X428 muxtest_0.x2.x1.nSEL1 ui_in[4].t4 VDPWR.t421 VDPWR.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X429 a_15575_12017# ringtest_0.x3.x1.nSEL0 a_15749_12123# VSS.t987 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X430 a_25083_4790# ringtest_0.x4._07_ VSS.t769 VSS.t768 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X431 VDPWR.t568 a_19666_31955# muxtest_0.x1.x3.GN3 VDPWR.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X432 VSS.t996 ringtest_0.x4._14_ ringtest_0.x4._02_ VSS.t995 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 muxtest_0.R1R2.t1 ua[0].t2 VSS.t519 sky130_fd_pr__res_high_po_1p41 l=1.75
X434 VSS.t265 VDPWR.t1209 VSS.t264 VSS.t263 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X435 VSS.t1093 a_23879_6940# ringtest_0.x4.clknet_0_clk.t25 VSS.t1092 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X436 VSS.t795 ringtest_0.x4.clknet_1_1__leaf_clk.t35 a_24729_4790# VSS.t794 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X437 a_26808_5308# a_26640_5334# VSS.t714 VSS.t713 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X438 VDPWR.t393 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t7 VDPWR.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X439 VDPWR.t1054 VSS.t1166 VDPWR.t1053 VDPWR.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X440 VDPWR.t1052 VSS.t1167 VDPWR.t1051 VDPWR.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X441 VSS.t268 VDPWR.t1210 VSS.t267 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X442 VSS.t271 VDPWR.t1211 VSS.t270 VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X443 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP4.t4 muxtest_0.R4R5.t2 VDPWR.t464 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X444 VDPWR.t638 ringtest_0.x4.net4 a_21591_6128# VDPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X445 a_21055_5334# ringtest_0.x4._13_ VDPWR.t642 VDPWR.t641 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X446 VDPWR.t516 a_11845_23906# muxtest_0.x2.x2.GN1 VDPWR.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X447 VSS.t598 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VSS.t564 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X448 VDPWR.t1050 VSS.t1168 VDPWR.t1049 VDPWR.t1048 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X449 a_21395_6940# ringtest_0.x4.clknet_0_clk.t36 VSS.t743 VSS.t742 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X450 VDPWR.t82 ringtest_0.x4.net8 a_25149_4220# VDPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X451 ringtest_0.drv_out.t6 a_19289_13081.t9 VDPWR.t483 VDPWR.t482 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X452 VDPWR.t361 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X453 VDPWR.t1047 VSS.t1169 VDPWR.t1046 VDPWR.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X454 a_25168_5156# a_24895_4790# a_25083_4790# VDPWR.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X455 VDPWR.t571 ringtest_0.x4.clknet_1_1__leaf_clk.t36 a_26201_5340# VDPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X456 VDPWR.t730 ringtest_0.x4.net6.t7 a_22795_5334# VDPWR.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X457 a_25364_5878# ringtest_0.x4.clknet_0_clk.t37 VDPWR.t740 VDPWR.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X458 a_21863_4790# ringtest_0.x4._03_ VSS.t986 VSS.t985 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X459 ringtest_0.x3.nselect2 VDPWR.t1212 VSS.t273 VSS.t272 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X460 a_23949_6654# a_24045_6654# VSS.t831 VSS.t830 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X461 a_23529_6422# a_23349_6422# VDPWR.t96 VDPWR.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X462 a_25055_3867# ringtest_0.x4.net7 VSS.t975 VSS.t974 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X463 a_26555_4790# ringtest_0.x4._09_ VDPWR.t257 VDPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X464 a_22795_5334# a_22765_5308# ringtest_0.x4._04_ VDPWR.t674 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X465 VDPWR.t231 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP4.t1 VDPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X466 VSS.t276 VDPWR.t1213 VSS.t275 VSS.t274 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X467 VDPWR.t472 ringtest_0.drv_out.t21 a_23879_6940# VDPWR.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X468 ringtest_0.x4._24_ a_26627_4246# VSS.t709 VSS.t708 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X469 a_26640_5156# a_26201_4790# a_26555_4790# VSS.t433 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X470 a_21675_9686# ringtest_0.x4.net2.t8 VDPWR.t441 VDPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X471 VDPWR.t372 a_22052_9116# a_21981_9142# VDPWR.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X472 VDPWR.t620 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X473 VSS.t1050 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VSS.t331 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X474 VDPWR.t1044 VSS.t1170 VDPWR.t1043 VDPWR.t1042 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X475 a_27303_4246# ringtest_0.x4._23_ VDPWR.t826 VDPWR.t825 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X476 a_21948_5156# a_21675_4790# a_21863_4790# VDPWR.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X477 a_13675_24012# ui_in[3].t6 VSS.t674 VSS.t673 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X478 VSS.t279 VDPWR.t1214 VSS.t278 VSS.t277 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X479 VSS.t282 VDPWR.t1215 VSS.t281 VSS.t280 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X480 VSS.t285 VDPWR.t1216 VSS.t284 VSS.t283 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X481 a_26766_4790# a_26367_4790# a_26640_5156# VSS.t438 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X482 VSS.t812 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VSS.t811 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X483 VDPWR.t1041 VSS.t1171 VDPWR.t1040 VDPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X484 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk.t37 VSS.t797 VSS.t796 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X485 VDPWR.t752 ui_in[2].t2 muxtest_0.x1.x5.GN VDPWR.t751 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X486 a_26721_4246# ringtest_0.x4._15_ VDPWR.t26 VDPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X487 VSS.t569 a_22295_3867# ringtest_0.x4.counter[2] VSS.t568 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X488 VSS.t799 ringtest_0.x4.clknet_1_1__leaf_clk.t38 a_24361_5340# VSS.t798 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X489 VSS.t777 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VSS.t404 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X490 VSS.t1053 ringtest_0.x4._05_ a_24883_6800# VSS.t1052 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X491 VDPWR.t339 a_25336_4902# a_25263_5156# VDPWR.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X492 a_20318_32213# ui_in[0].t5 VDPWR.t110 VDPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X493 VSS.t1002 a_16579_11759# ringtest_0.x3.x2.GN3 VSS.t1001 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X494 ringtest_0.counter7.t0 ringtest_0.x3.x2.GN4 ua[1].t1 VSS.t345 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X495 VDPWR.t1039 VSS.t1172 VDPWR.t1038 VDPWR.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X496 a_23879_6940# ringtest_0.drv_out.t22 VDPWR.t474 VDPWR.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X497 a_26808_5308# a_26640_5334# VDPWR.t456 VDPWR.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X498 ringtest_0.x4.clknet_1_1__leaf_clk.t26 a_25364_5878# VSS.t646 VSS.t645 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X499 a_26095_6788# ringtest_0.x4.net7 a_26007_6788# VSS.t973 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X500 ringtest_0.x4._07_ a_24699_6200# VDPWR.t601 VDPWR.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14575 ps=1.335 w=1 l=0.15
X501 a_21840_5308# a_21672_5334# VSS.t515 VSS.t514 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X502 a_15749_12123# ringtest_0.x3.x1.nSEL1 VSS.t91 VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X503 VSS.t288 VDPWR.t1217 VSS.t287 VSS.t286 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X504 VSS.t80 ringtest_0.x4._15_ a_26201_6788# VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X505 VDPWR.t376 ringtest_0.x4.net11 a_27489_3702# VDPWR.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X506 VSS.t512 a_26808_4902# a_26766_4790# VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X507 VDPWR.t1037 VSS.t1173 VDPWR.t1036 VDPWR.t1035 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X508 a_25263_5156# a_24729_4790# a_25168_5156# VDPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X509 VSS.t763 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2.t2 VSS.t762 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X510 ua[2].t1 muxtest_0.x2.x2.GP4.t5 muxtest_0.R7R8.t1 VDPWR.t5 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X511 VSS.t1091 a_23879_6940# ringtest_0.x4.clknet_0_clk.t24 VSS.t1090 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X512 VSS.t290 VDPWR.t1218 VSS.t289 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X513 a_21375_3867# ringtest_0.x4.net3.t5 VSS.t724 VSS.t723 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X514 VDPWR.t520 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X515 VSS.t196 VDPWR.t1219 VSS.t195 VSS.t194 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X516 ringtest_0.x4._15_ a_23381_4584# VDPWR.t763 VDPWR.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X517 VDPWR.t259 a_24135_3867# ringtest_0.x4.counter[4] VDPWR.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X518 VDPWR.t61 ringtest_0.x4.clknet_1_0__leaf_clk.t36 a_21233_5340# VDPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X519 muxtest_0.x1.x1.nSEL1 ui_in[1].t6 VSS.t693 VSS.t692 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X520 ringtest_0.ring_out.t2 ringtest_0.x3.x2.GN1 ua[1].t12 VSS.t835 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X521 ringtest_0.x4._10_ a_21785_8054# VDPWR.t74 VDPWR.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X522 ua[1].t8 ringtest_0.x3.x2.GP3 ringtest_0.counter3.t3 VDPWR.t557 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X523 a_22164_4362# ringtest_0.x4._16_.t6 VDPWR.t718 VDPWR.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X524 a_23467_4584# ringtest_0.x4.net4 a_23381_4584# VSS.t908 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X525 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP2.t6 muxtest_0.R2R3.t5 VDPWR.t247 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X526 VSS.t1026 ringtest_0.x4.clknet_0_clk.t38 a_21395_6940# VSS.t1025 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X527 VDPWR.t1034 VSS.t1174 VDPWR.t1033 VDPWR.t1032 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X528 VSS.t565 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VSS.t564 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X529 a_24685_6788# a_24465_6800# VSS.t703 VSS.t702 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X530 VDPWR.t1031 VSS.t1175 VDPWR.t1030 VDPWR.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X531 VDPWR.t650 ui_in[6].t0 ringtest_0.ring_out.t6 VDPWR.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X532 VSS.t199 VDPWR.t1220 VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X533 VSS.t202 VDPWR.t1221 VSS.t201 VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X534 VSS.t539 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t22 VSS.t538 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X535 VDPWR.t595 ringtest_0.x4._22_ a_26721_4246# VDPWR.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X536 VSS.t348 ringtest_0.x4._20_ a_23963_4790# VSS.t347 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X537 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP1.t5 muxtest_0.R7R8.t7 VDPWR.t660 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X538 a_22695_8304# ringtest_0.x4._12_ ringtest_0.x4._01_ VDPWR.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X539 ringtest_0.x4._17_ a_25925_6788# VDPWR.t765 VDPWR.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X540 muxtest_0.x2.x2.GP4.t0 muxtest_0.x2.x2.GN4 VDPWR.t229 VDPWR.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X541 ringtest_0.x4.clknet_0_clk.t23 a_23879_6940# VSS.t1089 VSS.t1088 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X542 a_26555_4790# ringtest_0.x4._09_ VSS.t499 VSS.t498 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X543 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VSS.t411 VSS.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X544 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR.t618 VDPWR.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X545 ringtest_0.x4.clknet_1_1__leaf_clk.t6 a_25364_5878# VDPWR.t391 VDPWR.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X546 VDPWR.t439 ringtest_0.x4.net2.t9 a_21785_8054# VDPWR.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X547 a_27169_6641# ringtest_0.x4._25_ VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X548 a_24317_4942# ringtest_0.x4.net8 VDPWR.t80 VDPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X549 ringtest_0.x4._16_.t1 a_23381_4818# VSS.t497 VSS.t496 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X550 ringtest_0.drv_out.t5 a_19289_13081.t10 VDPWR.t485 VDPWR.t484 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X551 muxtest_0.R5R6.t4 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A VSS.t1039 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X552 muxtest_0.R4R5.t0 muxtest_0.R3R4.t2 VSS.t138 sky130_fd_pr__res_high_po_1p41 l=1.75
X553 VSS.t1064 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 VSS.t1063 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X554 a_21845_8816# ringtest_0.x4.clknet_1_0__leaf_clk.t37 VSS.t439 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X555 a_27815_3867# ringtest_0.x4.net10 VSS.t321 VSS.t320 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X556 a_21561_9116# a_21845_9116# a_21780_9142# VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X557 a_21840_5308# a_21672_5334# VDPWR.t276 VDPWR.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X558 muxtest_0.x1.x5.GN ui_in[2].t3 VDPWR.t754 VDPWR.t753 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X559 VSS.t1024 a_12297_23648# muxtest_0.x2.x2.GN2 VSS.t1023 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X560 VDPWR.t684 ringtest_0.x3.x1.nSEL0 a_15575_12017# VDPWR.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X561 ringtest_0.x4.clknet_1_0__leaf_clk.t21 a_21395_6940# VSS.t537 VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X562 VSS.t977 a_25149_4220# ringtest_0.x4._22_ VSS.t976 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X563 VDPWR.t148 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP4.t1 VDPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X564 VDPWR.t1028 VSS.t1176 VDPWR.t1027 VDPWR.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X565 a_21561_8830# a_21845_8816# a_21780_8964# VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X566 VDPWR.t1026 VSS.t1177 VDPWR.t1025 VDPWR.t1024 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X567 VSS.t204 VDPWR.t1222 VSS.t203 VSS.t194 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X568 VDPWR.t1023 VSS.t1178 VDPWR.t1022 VDPWR.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X569 VSS.t1071 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VSS.t811 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X570 VSS.t311 a_18662_32213# muxtest_0.x1.x3.GN1 VSS.t310 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X571 VDPWR.t658 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1.t1 VDPWR.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X572 VDPWR.t1020 VSS.t1179 VDPWR.t1019 VDPWR.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X573 VSS.t207 VDPWR.t1223 VSS.t206 VSS.t205 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X574 VDPWR.t227 a_13025_23980# a_12849_23648# VDPWR.t226 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X575 a_21507_9686# ringtest_0.x4.net1 a_21425_9686# VDPWR.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X576 VDPWR.t1017 VSS.t1180 VDPWR.t1016 VDPWR.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X577 VSS.t210 VDPWR.t1224 VSS.t209 VSS.t208 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X578 a_24045_6654# a_24329_6640# a_24264_6788# VSS.t429 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X579 VSS.t994 ringtest_0.x4._14_ a_22390_4566# VSS.t993 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X580 a_25719_4790# a_24729_4790# a_25593_5156# VSS.t781 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X581 a_17405_12123# ui_in[3].t7 VSS.t676 VSS.t675 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X582 VDPWR.t1014 VSS.t1181 VDPWR.t1013 VDPWR.t864 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X583 ringtest_0.counter3.t4 ringtest_0.x3.x2.GN3 ua[1].t14 VSS.t1062 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X584 a_27169_6641# ringtest_0.x4._25_ VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X585 ringtest_0.drv_out.t11 a_19289_13081.t11 VSS.t93 VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X586 ringtest_0.x3.x1.nSEL0 ui_in[3].t8 VDPWR.t425 VDPWR.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X587 VSS.t212 VDPWR.t1225 VSS.t211 VSS.t200 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X588 VDPWR.t806 a_23879_6940# ringtest_0.x4.clknet_0_clk.t9 VDPWR.t805 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X589 VSS.t214 VDPWR.t1226 VSS.t213 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X590 ringtest_0.x4._00_ ringtest_0.x4.net1 a_21675_10006# VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X591 VDPWR.t720 ringtest_0.x4._16_.t7 a_24763_6143# VDPWR.t719 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.129 ps=1.18 w=0.42 l=0.15
X592 VSS.t217 VDPWR.t1227 VSS.t216 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X593 a_21803_8598# a_21465_8830# VDPWR.t186 VDPWR.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X594 a_22457_5156# a_21675_4790# a_22373_5156# VDPWR.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X595 a_18836_32319# muxtest_0.x1.x1.nSEL1 VSS.t593 VSS.t592 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X596 VSS.t220 VDPWR.t1228 VSS.t219 VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X597 VDPWR.t1012 VSS.t1182 VDPWR.t1011 VDPWR.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X598 a_25364_5878# ringtest_0.x4.clknet_0_clk.t39 VDPWR.t742 VDPWR.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X599 VDPWR.t44 a_19289_13081.t12 ringtest_0.drv_out.t4 VDPWR.t43 sky130_fd_pr__pfet_01v8 ad=2.79 pd=18.62 as=1.485 ps=9.33 w=9 l=0.15
X600 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP3 muxtest_0.R5R6.t2 VDPWR.t713 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X601 muxtest_0.R4R5.t5 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A VSS.t1056 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X602 ringtest_0.x4.net6.t1 a_22817_6146# VSS.t137 VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X603 a_24986_5878# ringtest_0.x4._22_ a_24763_6143# VSS.t823 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.1092 ps=1.36 w=0.42 l=0.15
X604 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP4.t5 muxtest_0.R4R5.t1 VDPWR.t465 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X605 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk.t38 VDPWR.t245 VDPWR.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X606 a_24287_6422# a_23949_6654# VDPWR.t225 VDPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X607 VDPWR.t272 a_26808_4902# a_26735_5156# VDPWR.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X608 a_26640_5334# a_26201_5340# a_26555_5334# VSS.t572 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X609 VSS.t820 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2.t3 VSS.t819 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X610 VDPWR.t476 ringtest_0.drv_out.t23 a_23879_6940# VDPWR.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X611 a_23837_5878# ringtest_0.x4._17_ VSS.t1109 VSS.t1108 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X612 ringtest_0.ring_out.t7 ui_in[6].t1 VDPWR.t652 VDPWR.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X613 VDPWR.t286 a_21845_8816# a_21852_8720# VDPWR.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X614 ringtest_0.x4.net4 a_22265_5308# VSS.t388 VSS.t387 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X615 VSS.t678 ui_in[3].t9 a_13025_23980# VSS.t677 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X616 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP4.t6 ua[0].t1 VDPWR.t466 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X617 VDPWR.t1009 VSS.t1183 VDPWR.t1008 VDPWR.t1007 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X618 VDPWR.t1006 VSS.t1184 VDPWR.t1005 VDPWR.t1004 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X619 a_13501_23906# ui_in[3].t10 VDPWR.t427 VDPWR.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X620 VSS.t222 VDPWR.t1229 VSS.t221 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X621 a_26735_5156# a_26201_4790# a_26640_5156# VDPWR.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X622 VSS.t225 VDPWR.t1230 VSS.t224 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X623 VDPWR.t1003 VSS.t1185 VDPWR.t1002 VDPWR.t1001 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X624 VSS.t340 a_17231_12017# ringtest_0.x3.x2.GN4 VSS.t339 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X625 ringtest_0.x4.clknet_0_clk.t22 a_23879_6940# VSS.t1087 VSS.t1086 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X626 VSS.t228 VDPWR.t1231 VSS.t227 VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X627 a_26766_5712# a_26367_5340# a_26640_5334# VSS.t358 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X628 VDPWR.t1000 VSS.t1186 VDPWR.t999 VDPWR.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X629 a_21981_8976# a_21845_8816# a_21561_8830# VDPWR.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X630 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VSS.t776 VSS.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X631 a_26007_6788# ringtest_0.x4.net6.t8 a_25925_6788# VSS.t1016 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X632 VDPWR.t998 VSS.t1187 VDPWR.t997 VDPWR.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X633 VDPWR.t732 ringtest_0.x4._21_ a_24070_5852# VDPWR.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.1176 ps=1.4 w=0.42 l=0.15
X634 VSS.t577 a_25761_5058# a_25719_4790# VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X635 VDPWR.t106 a_12473_23980# a_12297_23648# VDPWR.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X636 a_15575_12017# ringtest_0.x3.x1.nSEL1 VDPWR.t42 VDPWR.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X637 ringtest_0.x4.clknet_0_clk.t8 a_23879_6940# VDPWR.t804 VDPWR.t803 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X638 VSS.t230 VDPWR.t1232 VSS.t229 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X639 a_24465_6800# a_24329_6640# a_24045_6654# VDPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X640 VSS.t953 ringtest_0.x4.clknet_1_1__leaf_clk.t39 a_26201_5340# VSS.t952 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X641 VDPWR.t389 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t5 VDPWR.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X642 VDPWR.t996 VSS.t1188 VDPWR.t995 VDPWR.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X643 ringtest_0.x4._06_ a_24004_6128# VSS.t659 VSS.t658 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X644 VDPWR.t993 VSS.t1189 VDPWR.t992 VDPWR.t991 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X645 ringtest_0.x4.net6.t0 a_22817_6146# VDPWR.t91 VDPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X646 VSS.t1038 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 VSS.t1037 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X647 VSS.t232 VDPWR.t1233 VSS.t231 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X648 ringtest_0.x4.clknet_1_0__leaf_clk.t20 a_21395_6940# VSS.t535 VSS.t534 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X649 ringtest_0.x4.clknet_1_1__leaf_clk.t25 a_25364_5878# VSS.t644 VSS.t643 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X650 muxtest_0.x2.x2.GP1.t0 muxtest_0.x2.x2.GN1 VDPWR.t656 VDPWR.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X651 VSS.t1085 a_23879_6940# ringtest_0.x4.clknet_0_clk.t21 VSS.t1084 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X652 VDPWR.t180 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X653 muxtest_0.R1R2.t5 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A VSS.t1036 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X654 VSS.t235 VDPWR.t1234 VSS.t234 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X655 a_27065_5334# a_26201_5340# a_26808_5308# VDPWR.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X656 VSS.t1014 a_12849_23648# muxtest_0.x2.x2.GN3 VSS.t1013 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X657 VDPWR.t622 a_25977_4220# ringtest_0.x4._23_ VDPWR.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X658 VDPWR.t38 muxtest_0.x1.x1.nSEL0 a_18662_32213# VDPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X659 a_23349_6422# ringtest_0.x4._17_ VSS.t1107 VSS.t1106 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X660 ringtest_0.x4.clknet_1_1__leaf_clk.t4 a_25364_5878# VDPWR.t387 VDPWR.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X661 a_21675_4790# a_21509_4790# VDPWR.t509 VDPWR.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X662 a_21672_5334# a_21233_5340# a_21587_5334# VSS.t1125 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X663 a_22765_4478# ringtest_0.x4.net4 a_22939_4584# VSS.t907 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X664 VSS.t669 ui_in[4].t5 a_12473_23980# VSS.t668 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X665 VSS.t533 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t19 VSS.t532 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X666 VDPWR.t990 VSS.t1190 VDPWR.t989 VDPWR.t988 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X667 a_25441_4612# ringtest_0.x4.net8 a_25345_4612# VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X668 a_27149_5156# a_26367_4790# a_27065_5156# VDPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X669 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VSS.t810 VSS.t809 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X670 VSS.t377 a_21465_8830# ringtest_0.x4.net3.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X671 muxtest_0.R2R3.t2 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A VSS.t327 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X672 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR.t359 VDPWR.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X673 a_22224_6244# a_21785_5878# a_22139_5878# VSS.t786 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X674 a_25055_3867# ringtest_0.x4.net7 VDPWR.t667 VDPWR.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X675 VSS.t380 a_25393_5308# a_25351_5712# VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X676 a_21798_5712# a_21399_5340# a_21672_5334# VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X677 muxtest_0.R7R8.t5 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A VSS.t585 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X678 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP2.t7 muxtest_0.R2R3.t4 VDPWR.t248 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X679 VDPWR.t987 VSS.t1191 VDPWR.t986 VDPWR.t985 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X680 VDPWR.t365 a_24763_6143# a_24699_6200# VDPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.0672 ps=0.74 w=0.42 l=0.15
X681 VDPWR.t780 a_24536_6699# a_24465_6800# VDPWR.t779 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X682 VDPWR.t123 a_27233_5308# a_27149_5334# VDPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X683 VSS.t238 VDPWR.t1235 VSS.t237 VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X684 VSS.t326 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2.t2 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X685 VDPWR.t46 a_19289_13081.t13 ringtest_0.drv_out.t3 VDPWR.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X686 a_22350_5878# a_21951_5878# a_22224_6244# VSS.t750 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X687 VSS.t972 ringtest_0.x4.net7 a_23770_5308# VSS.t971 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X688 VSS.t441 ringtest_0.x4.clknet_1_0__leaf_clk.t39 a_21233_5340# VSS.t440 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X689 ringtest_0.x4.clknet_1_0__leaf_clk.t18 a_21395_6940# VSS.t531 VSS.t530 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X690 VDPWR.t423 ui_in[4].t6 muxtest_0.x2.x1.nSEL1 VDPWR.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X691 a_19289_13081.t0 ringtest_0.ring_out.t12 VSS.t370 VSS.t369 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X692 VDPWR.t984 VSS.t1192 VDPWR.t983 VDPWR.t982 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X693 VDPWR.t744 ringtest_0.x4.clknet_0_clk.t40 a_25364_5878# VDPWR.t743 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X694 ringtest_0.x4.counter[9] a_27489_3702# VSS.t368 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X695 ringtest_0.x4.clknet_1_1__leaf_clk.t24 a_25364_5878# VSS.t642 VSS.t641 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X696 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR.t528 VDPWR.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X697 a_17231_12017# ui_in[3].t11 VDPWR.t55 VDPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X698 VDPWR.t981 VSS.t1193 VDPWR.t980 VDPWR.t979 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X699 VSS.t241 VDPWR.t1236 VSS.t240 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X700 VDPWR.t330 a_22295_3867# ringtest_0.x4.counter[2] VDPWR.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X701 VDPWR.t978 VSS.t1194 VDPWR.t977 VDPWR.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X702 a_22765_5308# ringtest_0.x4.net6.t9 VSS.t1018 VSS.t1017 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X703 ua[3].t3 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A VSS.t774 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X704 VSS.t1083 a_23879_6940# ringtest_0.x4.clknet_0_clk.t20 VSS.t1082 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X705 ua[2].t4 muxtest_0.x2.x2.GP2.t4 ua[0].t6 VDPWR.t94 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X706 a_22097_5334# a_21233_5340# a_21840_5308# VDPWR.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X707 muxtest_0.R3R4.t6 muxtest_0.x2.x2.GN3 ua[2].t8 VSS.t679 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X708 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR.t178 VDPWR.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X709 VSS.t142 VDPWR.t1237 VSS.t141 VSS.t140 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X710 VDPWR.t802 a_23879_6940# ringtest_0.x4.clknet_0_clk.t7 VDPWR.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X711 ringtest_0.x4._19_ a_23529_6422# VDPWR.t200 VDPWR.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X712 a_23381_4584# ringtest_0.x4.net4 VDPWR.t636 VDPWR.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X713 VSS.t338 a_25593_5156# a_25761_5058# VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X714 a_22139_5878# ringtest_0.x4._04_ VDPWR.t579 VDPWR.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X715 muxtest_0.x2.x1.nSEL0 ui_in[3].t12 VSS.t101 VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X716 VSS.t145 VDPWR.t1238 VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X717 a_21375_3867# ringtest_0.x4.net3.t6 VDPWR.t478 VDPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X718 a_24317_4942# ringtest_0.x4.net6.t10 VDPWR.t575 VDPWR.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X719 VDPWR.t40 a_16203_12091# a_16027_11759# VDPWR.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X720 VDPWR.t506 ringtest_0.x4._11_.t12 a_22695_8304# VDPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X721 ringtest_0.x4.clknet_1_0__leaf_clk.t10 a_21395_6940# VDPWR.t308 VDPWR.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X722 VSS.t148 VDPWR.t1239 VSS.t147 VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X723 VSS.t366 a_26895_3867# ringtest_0.counter7.t3 VSS.t365 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X724 ua[1].t7 ringtest_0.x3.x2.GP3 ringtest_0.counter3.t2 VDPWR.t556 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X725 VSS.t151 VDPWR.t1240 VSS.t150 VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X726 VSS.t529 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t17 VSS.t528 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X727 ua[2].t2 muxtest_0.x2.x2.GP3 muxtest_0.R3R4.t0 VDPWR.t75 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X728 VDPWR.t975 VSS.t1195 VDPWR.t974 VDPWR.t973 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X729 VDPWR.t972 VSS.t1196 VDPWR.t971 VDPWR.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X730 VSS.t154 VDPWR.t1241 VSS.t153 VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X731 a_26367_4790# a_26201_4790# VDPWR.t241 VDPWR.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X732 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR.t769 VDPWR.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X733 a_24545_5878# ringtest_0.x4.net9 VSS.t362 VSS.t361 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X734 muxtest_0.R6R7.t0 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A VSS.t324 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X735 muxtest_0.x1.x5.A muxtest_0.x1.x3.GP3 muxtest_0.R5R6.t1 VDPWR.t712 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X736 a_24968_5308# a_24800_5334# VSS.t801 VSS.t800 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X737 VDPWR.t194 a_22265_5308# a_22181_5334# VDPWR.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X738 a_13501_23906# ui_in[4].t7 a_13675_24012# VSS.t670 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X739 VSS.t103 ui_in[3].t13 ringtest_0.x3.x1.nSEL0 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X740 VDPWR.t223 a_23949_6654# ringtest_0.x4.net7 VDPWR.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X741 VSS.t157 VDPWR.t1242 VSS.t156 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X742 VDPWR.t969 VSS.t1197 VDPWR.t968 VDPWR.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X743 VSS.t78 ringtest_0.x4._15_ a_23467_4818# VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X744 VDPWR.t306 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t9 VDPWR.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X745 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VSS.t1070 VSS.t809 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X746 VSS.t672 ui_in[4].t8 a_16203_12091# VSS.t671 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X747 VDPWR.t966 VSS.t1198 VDPWR.t965 VDPWR.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X748 VSS.t160 VDPWR.t1243 VSS.t159 VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X749 VDPWR.t102 ui_in[1].t7 a_20318_32213# VDPWR.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X750 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP4.t7 ua[0].t0 VDPWR.t467 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X751 a_24004_6128# a_24070_5852# a_23837_5878# VSS.t793 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X752 VDPWR.t142 a_25593_5156# a_25761_5058# VDPWR.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X753 a_22373_5156# a_21675_4790# a_22116_4902# VSS.t749 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X754 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR.t555 VDPWR.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X755 a_21465_9294# a_21561_9116# VSS.t834 VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X756 VDPWR.t385 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t3 VDPWR.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X757 ua[3].t2 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A VSS.t774 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X758 a_23932_6128# ringtest_0.x4.net8 VDPWR.t78 VDPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X759 a_23399_3867# ringtest_0.x4.net5 VSS.t1028 VSS.t1027 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X760 a_27815_3867# ringtest_0.x4.net10 VDPWR.t129 VDPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X761 ringtest_0.x4.clknet_1_1__leaf_clk.t23 a_25364_5878# VSS.t640 VSS.t639 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X762 VSS.t84 a_13501_23906# muxtest_0.x2.x2.GN4 VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X763 VDPWR.t368 a_22052_8875# a_21981_8976# VDPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X764 VDPWR.t963 VSS.t1199 VDPWR.t962 VDPWR.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X765 ringtest_0.x3.x2.GP4.t0 ringtest_0.x3.x2.GN4 VDPWR.t146 VDPWR.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X766 VDPWR.t154 ringtest_0.x4._11_.t13 a_26721_4246# VDPWR.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X767 a_23899_5654# ringtest_0.x4._15_ VSS.t76 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X768 ringtest_0.x3.x2.GP2.t2 ringtest_0.x3.x2.GN2 VSS.t818 VSS.t817 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X769 VDPWR.t341 a_19114_31955# muxtest_0.x1.x3.GN2 VDPWR.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X770 VDPWR.t254 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.ring_out.t1 VDPWR.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X771 VDPWR.t263 ui_in[4].t9 ringtest_0.x3.x1.nSEL1 VDPWR.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X772 VDPWR.t960 VSS.t1200 VDPWR.t959 VDPWR.t958 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X773 a_24800_5334# a_24361_5340# a_24715_5334# VSS.t660 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X774 VSS.t163 VDPWR.t1244 VSS.t162 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X775 VSS.t527 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t16 VSS.t526 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X776 a_23381_4818# ringtest_0.x4._11_.t14 VDPWR.t156 VDPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X777 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR.t328 VDPWR.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X778 a_21561_9116# a_21852_9416# a_21803_9508# VDPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X779 VSS.t409 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VSS.t408 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X780 VSS.t638 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t22 VSS.t637 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X781 a_24968_5308# a_24800_5334# VDPWR.t573 VDPWR.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X782 a_24926_5712# a_24527_5340# a_24800_5334# VSS.t1120 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X783 VDPWR.t957 VSS.t1201 VDPWR.t956 VDPWR.t955 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X784 VSS.t11 a_22245_8054# ringtest_0.x4._11_.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X785 a_21132_8918# ringtest_0.x4.net1 VSS.t400 VSS.t399 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X786 ringtest_0.x4._09_ a_27273_4220# VSS.t686 VSS.t685 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X787 a_24551_4790# ringtest_0.x4.net7 a_24479_4790# VSS.t970 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X788 VSS.t166 VDPWR.t1245 VSS.t165 VSS.t164 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X789 muxtest_0.x2.x1.nSEL1 ui_in[4].t10 VSS.t505 VSS.t504 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X790 ua[0].t7 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A VSS.t1055 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X791 VDPWR.t632 a_16755_12091# a_16579_11759# VDPWR.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X792 a_27273_4220# ringtest_0.x4._23_ a_27659_4246# VDPWR.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X793 VDPWR.t66 a_24317_4942# ringtest_0.x4._20_ VDPWR.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X794 VSS.t315 a_27233_5308# a_27191_5712# VSS.t314 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X795 ua[2].t5 muxtest_0.x2.x2.GP2.t5 ua[0].t5 VDPWR.t111 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X796 VSS.t169 VDPWR.t1246 VSS.t168 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X797 ringtest_0.x4.clknet_0_clk.t6 a_23879_6940# VDPWR.t800 VDPWR.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X798 a_22733_6244# a_21951_5878# a_22649_6244# VDPWR.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X799 VDPWR.t954 VSS.t1202 VDPWR.t953 VDPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X800 VDPWR.t952 VSS.t1203 VDPWR.t951 VDPWR.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X801 a_27273_4220# ringtest_0.x4.net11 VSS.t620 VSS.t619 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X802 VDPWR.t786 a_25225_5334# a_25393_5308# VDPWR.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X803 a_25225_5334# a_24527_5340# a_24968_5308# VSS.t1119 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X804 a_22111_10993# ui_in[5].t0 VDPWR.t68 VDPWR.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X805 VDPWR.t304 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t8 VDPWR.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X806 VDPWR.t949 VSS.t1204 VDPWR.t948 VDPWR.t947 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X807 VDPWR.t208 ringtest_0.x4.net1 a_21785_8054# VDPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X808 a_27065_5156# a_26367_4790# a_26808_4902# VSS.t437 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X809 VSS.t601 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X810 a_17231_12017# ui_in[4].t11 a_17405_12123# VSS.t506 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X811 ringtest_0.x4._12_ ringtest_0.x4.net3.t7 a_21049_8598# VDPWR.t479 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X812 a_25225_5334# a_24361_5340# a_24968_5308# VDPWR.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X813 VDPWR.t946 VSS.t1205 VDPWR.t945 VDPWR.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X814 VDPWR.t943 VSS.t1206 VDPWR.t942 VDPWR.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X815 VDPWR.t184 a_21465_8830# ringtest_0.x4.net3.t0 VDPWR.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X816 VSS.t172 VDPWR.t1247 VSS.t171 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X817 muxtest_0.R5R6.t3 muxtest_0.R4R5.t3 VSS.t419 sky130_fd_pr__res_high_po_1p41 l=1.75
X818 ringtest_0.drv_out.t2 a_19289_13081.t14 VDPWR.t48 VDPWR.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=2.79 ps=18.62 w=9 l=0.15
X819 VDPWR.t690 a_22765_4478# ringtest_0.x4._14_ VDPWR.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X820 VSS.t390 a_16027_11759# ringtest_0.x3.x2.GN2 VSS.t389 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X821 VSS.t105 ui_in[3].t14 a_16755_12091# VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X822 VSS.t175 VDPWR.t1248 VSS.t174 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X823 VSS.t424 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP4.t3 VSS.t423 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X824 VDPWR.t634 ringtest_0.x4.net4 a_22765_4478# VDPWR.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X825 a_22074_4790# a_21675_4790# a_21948_5156# VSS.t748 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X826 a_21780_9142# a_21465_9294# VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X827 a_24763_6143# ringtest_0.x4._22_ VDPWR.t593 VDPWR.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.20925 ps=1.345 w=0.42 l=0.15
X828 VSS.t178 VDPWR.t1249 VSS.t177 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X829 ringtest_0.x4.clknet_1_0__leaf_clk.t7 a_21395_6940# VDPWR.t302 VDPWR.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X830 ringtest_0.ring_out.t0 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR.t252 VDPWR.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X831 VSS.t846 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VSS.t843 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X832 a_23809_4790# ringtest_0.x4._15_ VDPWR.t24 VDPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X833 VDPWR.t940 VSS.t1207 VDPWR.t939 VDPWR.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X834 VSS.t181 VDPWR.t1250 VSS.t180 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X835 VSS.t87 muxtest_0.R7R8.t2 VSS.t86 sky130_fd_pr__res_high_po_1p41 l=1.75
X836 VSS.t184 VDPWR.t1251 VSS.t183 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X837 VDPWR.t938 VSS.t1208 VDPWR.t937 VDPWR.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X838 a_22052_9116# a_21845_9116# a_22228_9508# VDPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X839 a_22939_4584# ringtest_0.x4._11_.t15 VSS.t352 VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X840 VSS.t294 a_22116_4902# a_22074_4790# VSS.t293 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X841 ringtest_0.x4.clknet_1_1__leaf_clk.t2 a_25364_5878# VDPWR.t383 VDPWR.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X842 VDPWR.t265 ui_in[4].t12 a_13501_23906# VDPWR.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X843 a_22228_9508# a_21981_9142# VDPWR.t756 VDPWR.t755 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X844 VSS.t1033 ui_in[2].t4 muxtest_0.x1.x5.GN VSS.t1032 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X845 VDPWR.t188 a_25393_5308# a_25309_5334# VDPWR.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X846 a_24895_4790# a_24729_4790# VSS.t780 VSS.t779 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X847 VSS.t386 a_22265_5308# a_22223_5712# VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X848 VSS.t636 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t21 VSS.t635 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X849 VSS.t187 VDPWR.t1252 VSS.t186 VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X850 VDPWR.t236 a_24329_6640# a_24336_6544# VDPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X851 VSS.t190 VDPWR.t1253 VSS.t189 VSS.t188 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X852 muxtest_0.R7R8.t3 muxtest_0.x2.x2.GN4 ua[2].t6 VSS.t422 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X853 a_26555_5334# ringtest_0.x4._08_ VDPWR.t152 VDPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X854 a_19290_32287# ui_in[1].t8 VDPWR.t104 VDPWR.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X855 muxtest_0.R6R7.t4 muxtest_0.R5R6.t0 VSS.t138 sky130_fd_pr__res_high_po_1p41 l=1.75
X856 VSS.t775 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VSS.t408 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X857 VDPWR.t935 VSS.t1209 VDPWR.t934 VDPWR.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X858 a_26627_4246# ringtest_0.x4.net10 VSS.t319 VSS.t318 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X859 VSS.t193 VDPWR.t1254 VSS.t192 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X860 a_22775_5878# a_21785_5878# a_22649_6244# VSS.t785 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X861 VSS.t855 VDPWR.t1255 VSS.t854 VSS.t853 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X862 a_22795_5334# ringtest_0.x4._16_.t8 VDPWR.t722 VDPWR.t721 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X863 ringtest_0.x4._13_ ringtest_0.x4._11_.t16 VSS.t354 VSS.t353 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X864 VSS.t755 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VSS.t754 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X865 VSS.t415 a_23949_6654# ringtest_0.x4.net7 VSS.t414 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X866 VDPWR.t496 ringtest_0.x4.clknet_0_clk.t41 a_25364_5878# VDPWR.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X867 a_26367_5340# a_26201_5340# VDPWR.t331 VDPWR.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X868 VDPWR.t498 ringtest_0.x4.clknet_0_clk.t42 a_21395_6940# VDPWR.t497 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X869 ringtest_0.drv_out.t10 a_19289_13081.t15 VSS.t95 VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X870 ua[1].t11 ringtest_0.x3.x2.GP1.t4 ringtest_0.ring_out.t5 VDPWR.t602 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X871 VSS.t998 ringtest_0.x4._18_ a_23619_6788# VSS.t997 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X872 VSS.t857 VDPWR.t1256 VSS.t856 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X873 a_12849_23648# ui_in[4].t13 VDPWR.t267 VDPWR.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X874 ringtest_0.x4.clknet_1_1__leaf_clk.t20 a_25364_5878# VSS.t634 VSS.t633 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X875 VDPWR.t932 VSS.t1210 VDPWR.t931 VDPWR.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X876 a_26640_5156# a_26367_4790# a_26555_4790# VDPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X877 muxtest_0.R3R4.t4 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A VSS.t584 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X878 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP1.t6 muxtest_0.R3R4.t9 VDPWR.t661 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X879 VSS.t860 VDPWR.t1257 VSS.t859 VSS.t858 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X880 VSS.t863 VDPWR.t1258 VSS.t862 VSS.t861 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X881 VDPWR.t929 VSS.t1211 VDPWR.t928 VDPWR.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X882 a_22399_9142# a_21852_9416# a_22052_9116# VDPWR.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X883 VDPWR.t206 ringtest_0.x4.net1 a_21675_9686# VDPWR.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X884 ringtest_0.x4.counter[9] a_27489_3702# VDPWR.t169 VDPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X885 VSS.t126 ringtest_0.x4.clknet_1_0__leaf_clk.t40 a_21509_4790# VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X886 a_22392_5990# a_22224_6244# VSS.t113 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X887 muxtest_0.x1.x1.nSEL0 ui_in[0].t6 VDPWR.t626 VDPWR.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X888 a_17377_14114# ui_in[6].t2 ringtest_0.ring_out.t8 VSS.t959 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X889 ua[1].t0 ringtest_0.x3.x2.GP2.t4 ringtest_0.drv_out.t0 VDPWR.t64 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X890 VDPWR.t374 ringtest_0.x4.net11 a_27303_4246# VDPWR.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X891 muxtest_0.x2.x2.GP4.t2 muxtest_0.x2.x2.GN4 VSS.t421 VSS.t420 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X892 muxtest_0.R2R3.t0 muxtest_0.R1R2.t0 VSS.t88 sky130_fd_pr__res_high_po_1p41 l=1.75
X893 VSS.t563 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X894 ringtest_0.x4.clknet_1_0__leaf_clk.t6 a_21395_6940# VDPWR.t300 VDPWR.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X895 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VSS.t845 VSS.t841 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X896 ringtest_0.x4.clknet_0_clk.t19 a_23879_6940# VSS.t1081 VSS.t1080 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X897 VDPWR.t665 ringtest_0.x4.net7 a_24317_4942# VDPWR.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X898 VSS.t135 a_22817_6146# a_22775_5878# VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X899 VSS.t866 VDPWR.t1259 VSS.t865 VSS.t864 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X900 VDPWR.t167 a_26895_3867# ringtest_0.counter7.t2 VDPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X901 VSS.t844 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VSS.t843 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X902 VDPWR.t926 VSS.t1212 VDPWR.t925 VDPWR.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X903 VDPWR.t688 ringtest_0.x4._10_ a_22245_8054# VDPWR.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X904 VSS.t1073 a_25225_5334# a_25393_5308# VSS.t1072 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X905 a_21587_5334# ringtest_0.x4._02_ VDPWR.t587 VDPWR.t586 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X906 muxtest_0.x1.x5.GN ui_in[2].t5 VSS.t603 VSS.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X907 a_25336_4902# a_25168_5156# VSS.t595 VSS.t594 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X908 VSS.t632 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t19 VSS.t631 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X909 VSS.t344 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP4.t3 VSS.t343 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X910 VDPWR.t381 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t1 VDPWR.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X911 VSS.t869 VDPWR.t1260 VSS.t868 VSS.t867 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X912 ringtest_0.x4.clknet_0_clk.t5 a_23879_6940# VDPWR.t798 VDPWR.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X913 VSS.t967 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1.t3 VSS.t966 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X914 ringtest_0.drv_out.t19 ringtest_0.x3.x2.GN2 ua[1].t10 VSS.t816 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X915 VSS.t398 ringtest_0.x4.net1 a_21939_8054# VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X916 a_21399_5340# a_21233_5340# VDPWR.t1164 VDPWR.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X917 muxtest_0.x1.x5.A ui_in[2].t6 ua[3].t0 VDPWR.t362 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X918 a_19289_13081.t1 ringtest_0.ring_out.t13 VDPWR.t175 VDPWR.t174 sky130_fd_pr__pfet_01v8 ad=2.61 pd=18.58 as=2.61 ps=18.58 w=9 l=0.15
X919 VDPWR.t923 VSS.t1213 VDPWR.t922 VDPWR.t921 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X920 a_12297_23648# ui_in[3].t15 VDPWR.t57 VDPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X921 a_25345_4612# ringtest_0.x4.net9 VSS.t360 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X922 VSS.t872 VDPWR.t1261 VSS.t871 VSS.t870 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X923 VSS.t875 VDPWR.t1262 VSS.t874 VSS.t873 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X924 VDPWR.t298 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t5 VDPWR.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X925 VSS.t878 VDPWR.t1263 VSS.t877 VSS.t876 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X926 ringtest_0.x3.x1.nSEL0 ui_in[3].t16 VSS.t97 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X927 a_25547_4612# ringtest_0.x4.net7 a_25441_4612# VSS.t969 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X928 VDPWR.t100 a_22116_4902# a_22043_5156# VDPWR.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X929 VDPWR.t16 ui_in[4].t14 a_17231_12017# VDPWR.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X930 VDPWR.t823 ringtest_0.x4._23_ a_26569_6422# VDPWR.t822 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X931 VDPWR.t333 a_27065_5334# a_27233_5308# VDPWR.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X932 a_27065_5334# a_26367_5340# a_26808_5308# VSS.t357 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X933 ringtest_0.x4._02_ ringtest_0.x4._14_ a_21055_5334# VDPWR.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X934 VDPWR.t920 VSS.t1214 VDPWR.t919 VDPWR.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X935 a_26173_4612# ringtest_0.x4._22_ VSS.t822 VSS.t821 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X936 VSS.t792 a_19666_31955# muxtest_0.x1.x3.GN3 VSS.t791 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X937 ringtest_0.x3.x1.nSEL1 ui_in[4].t15 VDPWR.t18 VDPWR.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X938 a_26375_4612# ringtest_0.x4._11_.t17 a_26269_4612# VSS.t956 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X939 VSS.t881 VDPWR.t1264 VSS.t880 VSS.t879 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X940 VSS.t884 VDPWR.t1265 VSS.t883 VSS.t882 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X941 a_22043_5156# a_21509_4790# a_21948_5156# VDPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X942 VSS.t760 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VSS.t754 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X943 a_26749_6422# a_26569_6422# VDPWR.t522 VDPWR.t521 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X944 a_23770_5308# ringtest_0.x4.net6.t11 a_23993_5654# VSS.t802 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X945 VSS.t618 a_22052_9116# a_21981_9142# VSS.t608 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X946 a_23399_3867# ringtest_0.x4.net5 VDPWR.t746 VDPWR.t745 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X947 VSS.t886 VDPWR.t1266 VSS.t885 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X948 ringtest_0.ring_out.t9 ui_in[6].t3 a_17377_14114# VSS.t960 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X949 VDPWR.t451 a_15575_12017# ringtest_0.x3.x2.GN1 VDPWR.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X950 ringtest_0.x4._11_.t0 a_22245_8054# VDPWR.t12 VDPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X951 ringtest_0.x4._02_ ringtest_0.x4._13_ VSS.t912 VSS.t911 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X952 ringtest_0.x4.clknet_1_0__leaf_clk.t4 a_21395_6940# VDPWR.t296 VDPWR.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X953 muxtest_0.x1.x4.A muxtest_0.x1.x5.GN ua[3].t4 VDPWR.t547 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X954 VSS.t984 a_22021_4220# ringtest_0.x4._03_ VSS.t983 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X955 VSS.t955 ringtest_0.x4.clknet_1_1__leaf_clk.t40 a_26201_4790# VSS.t954 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X956 VDPWR.t917 VSS.t1215 VDPWR.t916 VDPWR.t915 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X957 VDPWR.t914 VSS.t1216 VDPWR.t913 VDPWR.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X958 VDPWR.t911 VSS.t1217 VDPWR.t910 VDPWR.t909 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X959 a_23879_6940# ringtest_0.drv_out.t24 VSS.t722 VSS.t721 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X960 ringtest_0.x4._24_ a_26627_4246# VDPWR.t453 VDPWR.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X961 a_25593_5156# a_24729_4790# a_25336_4902# VDPWR.t558 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X962 a_22111_10993# ui_in[5].t1 VSS.t111 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X963 a_21395_6940# ringtest_0.x4.clknet_0_clk.t43 VDPWR.t500 VDPWR.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X964 VDPWR.t767 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X965 ua[3].t7 muxtest_0.x2.x2.GN1 ua[2].t12 VSS.t965 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X966 ringtest_0.drv_out.t18 ringtest_0.x3.x2.GN2 ua[1].t9 VSS.t815 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X967 VSS.t980 ringtest_0.x4._01_ a_22399_8976# VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X968 a_25336_4902# a_25168_5156# VDPWR.t349 VDPWR.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X969 VSS.t630 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t18 VSS.t629 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X970 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VSS.t842 VSS.t841 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X971 VSS.t889 VDPWR.t1267 VSS.t888 VSS.t887 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X972 VDPWR.t192 a_26808_5308# a_26735_5334# VDPWR.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X973 ringtest_0.x4.clknet_0_clk.t4 a_23879_6940# VDPWR.t796 VDPWR.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X974 VDPWR.t553 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR.t552 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X975 VDPWR.t908 VSS.t1218 VDPWR.t907 VDPWR.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X976 muxtest_0.x2.x2.GP1.t2 muxtest_0.x2.x2.GN1 VSS.t964 VSS.t963 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X977 a_21465_9294# a_21561_9116# VDPWR.t608 VDPWR.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X978 VDPWR.t905 VSS.t1219 VDPWR.t904 VDPWR.t903 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X979 ringtest_0.x4._21_ a_23809_4790# VSS.t356 VSS.t355 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X980 VSS.t374 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VSS.t371 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X981 VSS.t892 VDPWR.t1268 VSS.t891 VSS.t890 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X982 VSS.t1079 a_23879_6940# ringtest_0.x4.clknet_0_clk.t18 VSS.t1078 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X983 muxtest_0.R3R4.t3 muxtest_0.R2R3.t3 VSS.t419 sky130_fd_pr__res_high_po_1p41 l=1.75
X984 VDPWR.t294 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t3 VDPWR.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X985 a_23891_4790# ringtest_0.x4._11_.t18 a_23809_4790# VSS.t957 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X986 VDPWR.t902 VSS.t1220 VDPWR.t901 VDPWR.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X987 VDPWR.t278 a_22097_5334# a_22265_5308# VDPWR.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X988 a_22097_5334# a_21399_5340# a_21840_5308# VSS.t312 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X989 ua[3].t1 ui_in[2].t7 muxtest_0.x1.x4.A VSS.t604 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X990 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR.t518 VDPWR.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X991 VSS.t413 a_25055_3867# ringtest_0.x4.counter[5] VSS.t412 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X992 VSS.t895 VDPWR.t1269 VSS.t894 VSS.t893 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X993 VDPWR.t335 a_25761_5058# a_25677_5156# VDPWR.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X994 a_26735_5334# a_26201_5340# a_26640_5334# VDPWR.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X995 ua[1].t3 ringtest_0.x3.x2.GP1.t5 ringtest_0.ring_out.t4 VDPWR.t176 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X996 VSS.t1077 a_23879_6940# ringtest_0.x4.clknet_0_clk.t17 VSS.t1076 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X997 ringtest_0.x4._25_ a_26749_6422# VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X998 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk.t41 VSS.t128 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X999 VSS.t720 a_19289_13081.t16 ringtest_0.drv_out.t9 VSS.t719 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1000 VDPWR.t899 VSS.t1221 VDPWR.t898 VDPWR.t897 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1001 a_22201_8964# a_21981_8976# VSS.t962 VSS.t961 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1002 VSS.t897 VDPWR.t1270 VSS.t896 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1003 VSS.t900 VDPWR.t1271 VSS.t899 VSS.t898 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1004 VSS.t903 VDPWR.t1272 VSS.t902 VSS.t901 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1005 a_24135_3867# ringtest_0.x4.net6.t12 VSS.t804 VSS.t803 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1006 a_26808_4902# a_26640_5156# VSS.t510 VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1007 a_22499_4790# a_21509_4790# a_22373_5156# VSS.t744 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1008 a_12849_23648# a_13025_23980# a_12977_24040# VSS.t418 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1009 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VSS.t600 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1010 VDPWR.t326 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1011 a_22765_4478# ringtest_0.x4._11_.t19 VDPWR.t646 VDPWR.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1012 VDPWR.t896 VSS.t1222 VDPWR.t895 VDPWR.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1013 a_19842_32287# ui_in[0].t7 VDPWR.t628 VDPWR.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X1014 a_11845_23906# muxtest_0.x2.x1.nSEL0 a_12019_24012# VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1015 VDPWR.t893 VSS.t1223 VDPWR.t892 VDPWR.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1016 VDPWR.t890 VSS.t1224 VDPWR.t889 VDPWR.t888 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1017 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR.t136 VDPWR.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1018 VDPWR.t887 VSS.t1225 VDPWR.t886 VDPWR.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1019 VDPWR.t644 ringtest_0.x4.clknet_1_1__leaf_clk.t41 a_24729_4790# VDPWR.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1020 a_26367_5340# a_26201_5340# VSS.t571 VSS.t570 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1021 VDPWR.t884 VSS.t1226 VDPWR.t883 VDPWR.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1022 a_24715_5334# ringtest_0.x4._06_ VDPWR.t581 VDPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1023 muxtest_0.R4R5.t4 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A VSS.t1054 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X1024 a_23619_6788# a_23349_6422# a_23529_6422# VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1025 VSS.t628 a_25364_5878# ringtest_0.x4.clknet_1_1__leaf_clk.t17 VSS.t627 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1026 VSS.t15 ui_in[4].t16 muxtest_0.x2.x1.nSEL1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1027 a_21049_8598# ringtest_0.x4.net2.t10 VDPWR.t437 VDPWR.t436 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X1028 VSS.t915 VDPWR.t1273 VSS.t914 VSS.t913 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1029 VSS.t1122 a_21375_3867# ringtest_0.x4.counter[1] VSS.t1121 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1030 VSS.t918 VDPWR.t1274 VSS.t917 VSS.t916 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1031 VSS.t575 a_27065_5334# a_27233_5308# VSS.t574 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1032 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR.t213 VDPWR.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1033 VSS.t1020 ringtest_0.x4._21_ a_24070_5852# VSS.t1019 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1034 a_24527_5340# a_24361_5340# VDPWR.t414 VDPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1035 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP1.t7 muxtest_0.R3R4.t8 VDPWR.t662 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1036 VDPWR.t738 a_12297_23648# muxtest_0.x2.x2.GN2 VDPWR.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1037 a_27149_5334# a_26367_5340# a_27065_5334# VDPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1038 VDPWR.t673 a_25149_4220# ringtest_0.x4._22_ VDPWR.t672 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X1039 a_21767_5334# a_21233_5340# a_21672_5334# VDPWR.t1162 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1040 VSS.t524 a_21845_8816# a_21852_8720# VSS.t523 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1041 VSS.t921 VDPWR.t1275 VSS.t920 VSS.t919 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1042 ringtest_0.x4.clknet_0_clk.t3 a_23879_6940# VDPWR.t794 VDPWR.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1043 a_25364_5878# ringtest_0.x4.clknet_0_clk.t44 VSS.t733 VSS.t732 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1044 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VSS.t373 VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1045 VDPWR.t577 ringtest_0.x4.net6.t13 a_25149_4220# VDPWR.t576 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1046 VDPWR.t782 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1047 VSS.t924 VDPWR.t1276 VSS.t923 VSS.t922 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1048 VSS.t305 a_22541_5058# a_22499_4790# VSS.t304 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1049 VDPWR.t881 VSS.t1227 VDPWR.t880 VDPWR.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1050 VSS.t611 ringtest_0.drv_out.t25 a_23879_6940# VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1051 a_22486_4246# ringtest_0.x4._14_ a_22021_4220# VDPWR.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1052 VSS.t1000 a_23770_5308# ringtest_0.x4._18_ VSS.t999 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1053 VDPWR.t127 ringtest_0.x4.net10 a_25977_4220# VDPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1054 a_12297_23648# a_12473_23980# a_12425_24040# VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1055 VSS.t372 ringtest_0.ring_out.t14 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VSS.t371 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1056 ua[1].t4 ringtest_0.x3.x2.GP4.t5 ringtest_0.counter7.t4 VDPWR.t463 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1057 VDPWR.t612 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1.t1 VDPWR.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1058 ringtest_0.x4.clknet_1_0__leaf_clk.t2 a_21395_6940# VDPWR.t292 VDPWR.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1059 a_24536_6699# a_24336_6544# a_24685_6788# VSS.t833 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1060 VDPWR.t878 VSS.t1228 VDPWR.t877 VDPWR.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1061 VSS.t926 VDPWR.t1277 VSS.t925 VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1062 a_12425_24040# ui_in[3].t17 VSS.t99 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X1063 VDPWR.t599 a_27169_6641# ringtest_0.x4._08_ VDPWR.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1064 VDPWR.t624 a_20318_32213# muxtest_0.x1.x3.GN4 VDPWR.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1065 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR.t355 VDPWR.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1066 VDPWR.t792 a_23879_6940# ringtest_0.x4.clknet_0_clk.t2 VDPWR.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1067 a_24536_6699# a_24329_6640# a_24712_6422# VDPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X1068 VSS.t597 a_27815_3867# ringtest_0.x4.counter[8] VSS.t596 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1069 muxtest_0.R1R2.t4 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A VSS.t1035 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X1070 ua[1].t6 ringtest_0.x3.x2.GP2.t5 ringtest_0.drv_out.t17 VDPWR.t470 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1071 a_25421_6641# ringtest_0.x4._19_ VDPWR.t202 VDPWR.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1072 VDPWR.t875 VSS.t1229 VDPWR.t874 VDPWR.t873 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1073 a_23879_6940# ringtest_0.drv_out.t26 VSS.t613 VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1074 a_21399_5340# a_21233_5340# VSS.t1124 VSS.t1123 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1075 VSS.t1069 a_24536_6699# a_24465_6800# VSS.t1068 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1076 a_24883_6800# a_24329_6640# a_24536_6699# VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1077 muxtest_0.x2.x2.GP3 muxtest_0.x2.x2.GN3 VDPWR.t430 VDPWR.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1078 a_21395_6940# ringtest_0.x4.clknet_0_clk.t45 VDPWR.t492 VDPWR.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1079 a_26201_6788# ringtest_0.x4._11_.t20 a_26095_6788# VSS.t958 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1080 VSS.t788 a_22649_6244# a_22817_6146# VSS.t787 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1081 VSS.t928 VDPWR.t1278 VSS.t927 VSS.t916 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1082 ringtest_0.x4._07_ a_24699_6200# VSS.t829 VSS.t828 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.098625 ps=0.98 w=0.65 l=0.15
X1083 VDPWR.t524 a_21845_9116# a_21852_9416# VDPWR.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1084 a_24712_6422# a_24465_6800# VDPWR.t447 VDPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1085 VDPWR.t51 ui_in[3].t18 muxtest_0.x2.x1.nSEL0 VDPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1086 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VSS.t561 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1087 VSS.t1012 ringtest_0.x4._16_.t9 a_22765_5308# VSS.t1011 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1088 VSS.t517 a_22097_5334# a_22265_5308# VSS.t516 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1089 muxtest_0.x1.x4.A muxtest_0.x1.x3.GP3 muxtest_0.R1R2.t2 VDPWR.t711 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1090 a_16579_11759# ui_in[4].t17 VDPWR.t20 VDPWR.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X1091 VDPWR.t872 VSS.t1230 VDPWR.t871 VDPWR.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1092 VSS.t827 a_27169_6641# ringtest_0.x4._08_ VSS.t826 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1093 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR.t549 VDPWR.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1094 muxtest_0.R2R3.t1 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A VSS.t323 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X1095 a_25421_6641# ringtest_0.x4._19_ VSS.t394 VSS.t393 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1096 VDPWR.t204 a_22111_10993# ringtest_0.x4.net1 VDPWR.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1097 ringtest_0.drv_out.t1 a_19289_13081.t17 VDPWR.t469 VDPWR.t468 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X1098 ringtest_0.x3.x2.GP4.t2 ringtest_0.x3.x2.GN4 VSS.t342 VSS.t341 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1099 a_21561_8830# a_21852_8720# a_21803_8598# VDPWR.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1100 VDPWR.t869 VSS.t1231 VDPWR.t868 VDPWR.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1101 a_23993_5654# ringtest_0.x4._11_.t21 a_23899_5654# VSS.t657 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1102 VDPWR.t866 VSS.t1232 VDPWR.t865 VDPWR.t864 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1103 VSS.t296 ui_in[1].t9 a_19290_32287# VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1104 a_17377_14114# ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VSS.t495 VSS.t494 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1105 VSS.t17 ui_in[4].t18 ringtest_0.x3.x1.nSEL1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1106 a_24883_6800# a_24336_6544# a_24536_6699# VDPWR.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X1107 VDPWR.t630 ui_in[0].t8 muxtest_0.x1.x1.nSEL0 VDPWR.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1108 a_18662_32213# muxtest_0.x1.x1.nSEL1 VDPWR.t347 VDPWR.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1109 VDPWR.t863 VSS.t1233 VDPWR.t862 VDPWR.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1110 VDPWR.t860 VSS.t1234 VDPWR.t859 VDPWR.t858 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1111 VDPWR.t566 a_22649_6244# a_22817_6146# VDPWR.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1112 VDPWR.t857 VSS.t1235 VDPWR.t856 VDPWR.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1113 VSS.t1116 a_27233_5058# a_27191_4790# VSS.t1115 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1114 VDPWR.t724 a_12849_23648# muxtest_0.x2.x2.GN3 VDPWR.t723 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1115 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.ring_out.t15 VSS.t133 VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1116 ringtest_0.x4.clknet_1_1__leaf_clk.t16 a_25364_5878# VSS.t626 VSS.t625 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1117 a_24699_6200# a_24763_6143# a_24545_5878# VSS.t605 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1118 muxtest_0.x2.x2.GP2.t0 muxtest_0.x2.x2.GN2 VDPWR.t532 VDPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1119 ringtest_0.x3.x2.GP1.t0 ringtest_0.x3.x2.GN1 VDPWR.t610 VDPWR.t609 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1120 ringtest_0.x4.clknet_1_1__leaf_clk.t0 a_25364_5878# VDPWR.t379 VDPWR.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1121 VDPWR.t274 muxtest_0.x2.x1.nSEL0 a_11845_23906# VDPWR.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1122 a_21951_5878# a_21785_5878# VSS.t784 VSS.t783 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1123 VSS.t559 a_22373_5156# a_22541_5058# VSS.t558 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1124 VDPWR.t854 VSS.t1236 VDPWR.t853 VDPWR.t852 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1125 a_25975_3867# ringtest_0.x4.net8 VSS.t119 VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1126 a_21981_9142# a_21852_9416# a_21561_9116# VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1127 VSS.t931 VDPWR.t1279 VSS.t930 VSS.t929 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1128 VDPWR.t790 a_23879_6940# ringtest_0.x4.clknet_0_clk.t1 VDPWR.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1129 VSS.t934 VDPWR.t1280 VSS.t933 VSS.t932 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1130 a_21981_8976# a_21852_8720# a_21561_8830# VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1131 VDPWR.t851 VSS.t1237 VDPWR.t850 VDPWR.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1132 a_22319_6244# a_21785_5878# a_22224_6244# VDPWR.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1133 VDPWR.t343 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1.t0 VDPWR.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1134 VSS.t937 VDPWR.t1281 VSS.t936 VSS.t935 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1135 VDPWR.t686 a_19290_32287# a_19114_31955# VDPWR.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1136 VSS.t940 VDPWR.t1282 VSS.t939 VSS.t938 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1137 VDPWR.t848 VSS.t1238 VDPWR.t847 VDPWR.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1138 VSS.t943 VDPWR.t1283 VSS.t942 VSS.t941 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1139 a_21951_5878# a_21785_5878# VDPWR.t562 VDPWR.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1140 ringtest_0.x4._06_ a_24004_6128# VDPWR.t411 VDPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.18575 ps=1.415 w=1 l=0.15
X1141 VDPWR.t233 a_24968_5308# a_24895_5334# VDPWR.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1142 a_24465_6800# a_24336_6544# a_24045_6654# VSS.t832 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1143 VDPWR.t845 VSS.t1239 VDPWR.t844 VDPWR.t843 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1144 a_22390_4566# a_22164_4362# a_22021_4220# VSS.t518 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1145 VDPWR.t494 ringtest_0.x4.clknet_0_clk.t46 a_21395_6940# VDPWR.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1146 VDPWR.t694 ringtest_0.x4._18_ a_23529_6422# VDPWR.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1147 VDPWR.t773 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP4.t0 VDPWR.t772 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1148 a_12977_24040# ui_in[4].t19 VSS.t773 VSS.t772 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X1149 VDPWR.t842 VSS.t1240 VDPWR.t841 VDPWR.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1150 ringtest_0.x4._10_ a_21785_8054# VSS.t117 VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1151 VSS.t1075 a_23879_6940# ringtest_0.x4.clknet_0_clk.t16 VSS.t1074 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1152 a_23963_4790# ringtest_0.x4._15_ a_23891_4790# VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1153 VDPWR.t290 a_21395_6940# ringtest_0.x4.clknet_1_0__leaf_clk.t1 VDPWR.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1154 VSS.t946 VDPWR.t1284 VSS.t945 VSS.t944 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1155 a_24895_5334# a_24361_5340# a_24800_5334# VDPWR.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1156 a_23770_5308# ringtest_0.x4.net7 a_23899_5334# VDPWR.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1157 a_22399_9142# a_21845_9116# a_22052_9116# VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1158 a_21867_8054# ringtest_0.x4.net2.t11 a_21785_8054# VSS.t694 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1159 VDPWR.t839 VSS.t1241 VDPWR.t838 VDPWR.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1160 ringtest_0.x4._04_ a_22765_5308# VSS.t979 VSS.t978 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1161 VSS.t948 VDPWR.t1285 VSS.t947 VSS.t188 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1162 ringtest_0.x4.clknet_0_clk.t0 a_23879_6940# VDPWR.t788 VDPWR.t787 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1163 a_25364_5878# ringtest_0.x4.clknet_0_clk.t47 VSS.t731 VSS.t730 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1164 a_22399_8976# a_21845_8816# a_22052_8875# VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1165 a_20492_32319# ui_in[0].t9 VSS.t852 VSS.t851 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1166 ringtest_0.x3.x2.GP3 ringtest_0.x3.x2.GN3 VDPWR.t777 VDPWR.t776 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1167 VDPWR.t320 a_22373_5156# a_22541_5058# VDPWR.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1168 VDPWR.t836 VSS.t1242 VDPWR.t835 VDPWR.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1169 a_22052_8875# a_21845_8816# a_22228_8598# VDPWR.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X1170 a_22228_8598# a_21981_8976# VDPWR.t654 VDPWR.t653 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1171 ringtest_0.x4._01_ ringtest_0.x4._12_ VSS.t1044 VSS.t1043 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1172 VSS.t615 ringtest_0.drv_out.t27 a_23879_6940# VSS.t614 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1173 ringtest_0.x4._16_.t0 a_23381_4818# VDPWR.t256 VDPWR.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1174 a_23151_5334# ringtest_0.x4.net6.t14 VDPWR.t449 VDPWR.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1175 VDPWR.t701 VDPWR.t699 muxtest_0.x2.nselect2 VDPWR.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1176 VSS.t753 a_11845_23906# muxtest_0.x2.x2.GN1 VSS.t752 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1177 a_22295_3867# ringtest_0.x4.net4 VSS.t906 VSS.t905 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1178 VDPWR.t833 VSS.t1243 VDPWR.t832 VDPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1179 a_13025_23980# ui_in[3].t19 VDPWR.t53 VDPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X1180 VSS.t493 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B a_17377_14114# VSS.t492 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1181 VSS.t951 VDPWR.t1286 VSS.t950 VSS.t949 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1182 VDPWR.t221 a_25055_3867# ringtest_0.x4.counter[5] VDPWR.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1183 VSS.t705 ringtest_0.x4.net6.t15 a_22983_5654# VSS.t704 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1184 VDPWR.t428 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 VDPWR.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1185 ringtest_0.x4.clknet_1_0__leaf_clk.t0 a_21395_6940# VDPWR.t288 VDPWR.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 ringtest_0.x4.net2.n14 ringtest_0.x4.net2.t1 315.034
R1 ringtest_0.x4.net2.t0 ringtest_0.x4.net2.n14 265.769
R2 ringtest_0.x4.net2 ringtest_0.x4.net2.t0 262.318
R3 ringtest_0.x4.net2.n4 ringtest_0.x4.net2.t5 260.322
R4 ringtest_0.x4.net2.n9 ringtest_0.x4.net2.t10 241.536
R5 ringtest_0.x4.net2.n0 ringtest_0.x4.net2.t8 212.081
R6 ringtest_0.x4.net2.n1 ringtest_0.x4.net2.t3 212.081
R7 ringtest_0.x4.net2.n6 ringtest_0.x4.net2.t9 183.505
R8 ringtest_0.x4.net2.n4 ringtest_0.x4.net2.t2 175.169
R9 ringtest_0.x4.net2.n9 ringtest_0.x4.net2.t6 169.237
R10 ringtest_0.x4.net2.n10 ringtest_0.x4.net2.n9 159.952
R11 ringtest_0.x4.net2.n7 ringtest_0.x4.net2.n6 153.863
R12 ringtest_0.x4.net2.n3 ringtest_0.x4.net2.n2 152.698
R13 ringtest_0.x4.net2.n5 ringtest_0.x4.net2.n4 152
R14 ringtest_0.x4.net2.n0 ringtest_0.x4.net2.t7 139.78
R15 ringtest_0.x4.net2.n1 ringtest_0.x4.net2.t4 139.78
R16 ringtest_0.x4.net2.n6 ringtest_0.x4.net2.t11 114.532
R17 ringtest_0.x4.net2.n2 ringtest_0.x4.net2.n0 37.246
R18 ringtest_0.x4.net2.n8 ringtest_0.x4.net2.n5 34.4715
R19 ringtest_0.x4.net2.n2 ringtest_0.x4.net2.n1 24.1005
R20 ringtest_0.x4.net2.n12 ringtest_0.x4.net2.n3 18.9449
R21 ringtest_0.x4.net2.n13 ringtest_0.x4.net2.n12 14.916
R22 ringtest_0.x4.net2.n11 ringtest_0.x4.net2.n10 13.8005
R23 ringtest_0.x4.net2 ringtest_0.x4.net2.n7 10.8927
R24 ringtest_0.x4.net2.n14 ringtest_0.x4.net2.n13 8.72777
R25 ringtest_0.x4.net2.n8 ringtest_0.x4.net2 6.07742
R26 ringtest_0.x4.net2.n10 ringtest_0.x4.net2 3.33963
R27 ringtest_0.x4.net2.n10 ringtest_0.x4.net2 3.29747
R28 ringtest_0.x4.net2 ringtest_0.x4.net2.n13 3.29747
R29 ringtest_0.x4.net2.n11 ringtest_0.x4.net2.n8 3.19006
R30 ringtest_0.x4.net2.n3 ringtest_0.x4.net2 1.97868
R31 ringtest_0.x4.net2.n7 ringtest_0.x4.net2 1.97868
R32 ringtest_0.x4.net2.n5 ringtest_0.x4.net2 1.55726
R33 ringtest_0.x4.net2.n12 ringtest_0.x4.net2.n11 1.38649
R34 VSS.n3345 VSS.n64 4.7454e+06
R35 VSS.n318 VSS.n65 4.7454e+06
R36 VSS.n3345 VSS.n65 3.52e+06
R37 VSS.n360 VSS.n64 3.52e+06
R38 VSS.n3151 VSS.n173 3.3176e+06
R39 VSS.n3220 VSS.n3219 3.3176e+06
R40 VSS.n378 VSS.n376 2.347e+06
R41 VSS.n376 VSS.n64 2.3386e+06
R42 VSS.n3130 VSS.n173 2.3386e+06
R43 VSS.n3220 VSS.n3189 2.3386e+06
R44 VSS.n321 VSS.n66 2.15447e+06
R45 VSS.n3189 VSS.n3188 2.1446e+06
R46 VSS.n3131 VSS.n3130 2.1446e+06
R47 VSS.n3222 VSS.n3173 1.86572e+06
R48 VSS.n303 VSS.n65 1.2338e+06
R49 VSS.n334 VSS.n65 1.18072e+06
R50 VSS.n310 VSS.n309 1.1798e+06
R51 VSS.n3223 VSS.n3171 1.1798e+06
R52 VSS.n3168 VSS.n176 1.1798e+06
R53 VSS.n311 VSS.n310 1.17976e+06
R54 VSS.n3223 VSS.n3172 1.17976e+06
R55 VSS.n3168 VSS.n3167 1.17976e+06
R56 VSS.n376 VSS.t588 1.17724e+06
R57 VSS.n3189 VSS.t341 1.17707e+06
R58 VSS.n3130 VSS.t420 1.17707e+06
R59 VSS.n3344 VSS.t959 1.0027e+06
R60 VSS.n3016 VSS.n224 573621
R61 VSS.n323 VSS.n318 396385
R62 VSS.n362 VSS.n360 396385
R63 VSS.n3153 VSS.n3151 396385
R64 VSS.n3219 VSS.n3218 396385
R65 VSS.n318 VSS.n317 391216
R66 VSS.n360 VSS.n359 391216
R67 VSS.n3219 VSS.n3190 391216
R68 VSS.n3151 VSS.n3150 391216
R69 VSS.n3222 VSS.n3221 293853
R70 VSS.n3344 VSS.n66 291597
R71 VSS.n3229 VSS.n3228 86912.4
R72 VSS.n3229 VSS.n66 81673.6
R73 VSS.n3174 VSS.n67 72143.6
R74 VSS.n310 VSS.n172 66245.4
R75 VSS.n3000 VSS.n224 61252.6
R76 VSS.n3020 VSS.n172 52488.3
R77 VSS.n3228 VSS.n3227 52128.6
R78 VSS.n3333 VSS.n3332 38301.6
R79 VSS VSS.n175 35992.3
R80 VSS.n3346 VSS.n63 35421.6
R81 VSS.n3334 VSS.n3333 29605.7
R82 VSS.n3227 VSS.n173 29419.1
R83 VSS.n3227 VSS.n172 29145.5
R84 VSS.n399 VSS 25742.3
R85 VSS.n1894 VSS 23608
R86 VSS.n3343 VSS.n67 18854
R87 VSS.n3227 VSS.n3226 17410.5
R88 VSS.n341 VSS.n222 16580.9
R89 VSS.n1894 VSS.t725 13977.5
R90 VSS VSS.n173 13964.9
R91 VSS.n3170 VSS.n174 13854.2
R92 VSS.n369 VSS.n341 13333.2
R93 VSS.n3228 VSS.n74 13232.9
R94 VSS.n379 VSS.n371 11744.7
R95 VSS.n383 VSS.n371 11744.7
R96 VSS.n379 VSS.n372 11744.7
R97 VSS.n383 VSS.n372 11744.7
R98 VSS.n358 VSS.n346 11744.7
R99 VSS.n354 VSS.n346 11744.7
R100 VSS.n358 VSS.n348 11744.7
R101 VSS.n354 VSS.n348 11744.7
R102 VSS.n396 VSS.n282 11744.7
R103 VSS.n396 VSS.n388 11744.7
R104 VSS.n388 VSS.n280 11744.7
R105 VSS.n282 VSS.n280 11744.7
R106 VSS.n335 VSS.n284 11744.7
R107 VSS.n339 VSS.n284 11744.7
R108 VSS.n335 VSS.n285 11744.7
R109 VSS.n339 VSS.n285 11744.7
R110 VSS.n316 VSS.n293 11744.7
R111 VSS.n312 VSS.n293 11744.7
R112 VSS.n316 VSS.n294 11744.7
R113 VSS.n312 VSS.n294 11744.7
R114 VSS.n304 VSS.n298 11744.7
R115 VSS.n308 VSS.n298 11744.7
R116 VSS.n304 VSS.n299 11744.7
R117 VSS.n308 VSS.n299 11744.7
R118 VSS.n320 VSS.n291 11744.7
R119 VSS.n320 VSS.n292 11744.7
R120 VSS.n324 VSS.n292 11744.7
R121 VSS.n324 VSS.n291 11744.7
R122 VSS.n363 VSS.n342 11744.7
R123 VSS.n367 VSS.n342 11744.7
R124 VSS.n363 VSS.n343 11744.7
R125 VSS.n367 VSS.n343 11744.7
R126 VSS.n3187 VSS.n3175 11744.7
R127 VSS.n3182 VSS.n3175 11744.7
R128 VSS.n3187 VSS.n3177 11744.7
R129 VSS.n3182 VSS.n3177 11744.7
R130 VSS.n3205 VSS.n3202 11744.7
R131 VSS.n3205 VSS.n3203 11744.7
R132 VSS.n3207 VSS.n3202 11744.7
R133 VSS.n3207 VSS.n3203 11744.7
R134 VSS.n206 VSS.n197 11744.7
R135 VSS.n206 VSS.n199 11744.7
R136 VSS.n199 VSS.n196 11744.7
R137 VSS.n197 VSS.n196 11744.7
R138 VSS.n3149 VSS.n177 11744.7
R139 VSS.n3166 VSS.n177 11744.7
R140 VSS.n3149 VSS.n178 11744.7
R141 VSS.n3166 VSS.n178 11744.7
R142 VSS.n3133 VSS.n185 11744.7
R143 VSS.n3133 VSS.n186 11744.7
R144 VSS.n3135 VSS.n185 11744.7
R145 VSS.n3135 VSS.n186 11744.7
R146 VSS.n3154 VSS.n3143 11744.7
R147 VSS.n3154 VSS.n3147 11744.7
R148 VSS.n3144 VSS.n3143 11744.7
R149 VSS.n3147 VSS.n3144 11744.7
R150 VSS.n3330 VSS.n75 11744.7
R151 VSS.n3330 VSS.n76 11744.7
R152 VSS.n75 VSS.n73 11744.7
R153 VSS.n76 VSS.n73 11744.7
R154 VSS.n3217 VSS.n3191 11744.7
R155 VSS.n3217 VSS.n3193 11744.7
R156 VSS.n3196 VSS.n3191 11744.7
R157 VSS.n3196 VSS.n3193 11744.7
R158 VSS.n3015 VSS.n225 11744.7
R159 VSS.n3011 VSS.n226 11744.7
R160 VSS.n3015 VSS.n226 11744.7
R161 VSS.n2998 VSS.n2996 11744.7
R162 VSS.n3002 VSS.n2996 11744.7
R163 VSS.n2999 VSS.n2998 11744.7
R164 VSS.n3002 VSS.n2999 11744.7
R165 VSS.n370 VSS.n369 9554.71
R166 VSS.n3335 VSS.n3334 9243.96
R167 VSS.n3021 VSS.n3020 8452.32
R168 VSS.n3017 VSS.n222 7337.33
R169 VSS.n323 VSS.t1059 7088.89
R170 VSS.t1055 VSS.n321 7088.89
R171 VSS.n362 VSS.t1054 7088.89
R172 VSS.n368 VSS.t1056 7088.89
R173 VSS.n3153 VSS.t422 7088.89
R174 VSS.t425 VSS.n174 7088.89
R175 VSS.n3218 VSS.t345 7088.89
R176 VSS.t346 VSS.n3173 7088.89
R177 VSS.n303 VSS.t323 6925.66
R178 VSS.n309 VSS.t327 6925.66
R179 VSS.n317 VSS.t1035 6925.66
R180 VSS.n311 VSS.t1036 6925.66
R181 VSS.n3188 VSS.t816 6925.66
R182 VSS.t815 VSS.n3171 6925.66
R183 VSS.t1062 VSS.n3190 6925.66
R184 VSS.t1065 VSS.n3172 6925.66
R185 VSS.t767 VSS.n3131 6925.66
R186 VSS.t764 VSS.n176 6925.66
R187 VSS.n3150 VSS.t679 6925.66
R188 VSS.n3167 VSS.t684 6925.66
R189 VSS.n359 VSS.t1042 6925.66
R190 VSS.t1039 VSS.n283 6925.66
R191 VSS.n378 VSS.t324 6925.66
R192 VSS.n384 VSS.t330 6925.66
R193 VSS.n3020 VSS.t423 6843.4
R194 VSS.t1059 VSS.n322 6733.33
R195 VSS.n322 VSS.t1055 6733.33
R196 VSS.t1054 VSS.n361 6733.33
R197 VSS.n361 VSS.t1056 6733.33
R198 VSS.t422 VSS.n3152 6733.33
R199 VSS.n3152 VSS.t425 6733.33
R200 VSS.n3192 VSS.t345 6733.33
R201 VSS.n3192 VSS.t346 6733.33
R202 VSS.t323 VSS.n302 6578.29
R203 VSS.n302 VSS.t327 6578.29
R204 VSS.n297 VSS.t1035 6578.29
R205 VSS.t1036 VSS.n297 6578.29
R206 VSS.n3176 VSS.t816 6578.29
R207 VSS.n3176 VSS.t815 6578.29
R208 VSS.n3206 VSS.t1062 6578.29
R209 VSS.n3206 VSS.t1065 6578.29
R210 VSS.n3134 VSS.t767 6578.29
R211 VSS.n3134 VSS.t764 6578.29
R212 VSS.t679 VSS.n3148 6578.29
R213 VSS.n3148 VSS.t684 6578.29
R214 VSS.n347 VSS.t1042 6578.29
R215 VSS.n347 VSS.t1039 6578.29
R216 VSS.t324 VSS.n377 6578.29
R217 VSS.n377 VSS.t330 6578.29
R218 VSS.n334 VSS.t591 6418.9
R219 VSS.n340 VSS.t584 6418.9
R220 VSS.t591 VSS.n333 6096.95
R221 VSS.n333 VSS.t584 6096.95
R222 VSS.n386 VSS.n385 5782.24
R223 VSS.n385 VSS.n370 5742.37
R224 VSS.n479 VSS.n423 5452.27
R225 VSS.n479 VSS.n470 5452.27
R226 VSS.n423 VSS.n421 5452.27
R227 VSS.n470 VSS.n421 5452.27
R228 VSS.n467 VSS.n428 5452.27
R229 VSS.n459 VSS.n428 5452.27
R230 VSS.n467 VSS.n429 5452.27
R231 VSS.n459 VSS.n429 5452.27
R232 VSS.n489 VSS.n402 5452.27
R233 VSS.n419 VSS.n402 5452.27
R234 VSS.n489 VSS.n403 5452.27
R235 VSS.n419 VSS.n403 5452.27
R236 VSS.n434 VSS.n425 5452.27
R237 VSS.n461 VSS.n434 5452.27
R238 VSS.n437 VSS.n425 5452.27
R239 VSS.n461 VSS.n437 5452.27
R240 VSS.n413 VSS.n400 5452.27
R241 VSS.n416 VSS.n413 5452.27
R242 VSS.n414 VSS.n400 5452.27
R243 VSS.n416 VSS.n414 5452.27
R244 VSS.n439 VSS.n427 5452.27
R245 VSS.n458 VSS.n439 5452.27
R246 VSS.n440 VSS.n427 5452.27
R247 VSS.n458 VSS.n440 5452.27
R248 VSS.n481 VSS.n410 5452.27
R249 VSS.n411 VSS.n410 5452.27
R250 VSS.n481 VSS.n480 5452.27
R251 VSS.n480 VSS.n411 5452.27
R252 VSS.n451 VSS.n449 5452.27
R253 VSS.n453 VSS.n449 5452.27
R254 VSS.n452 VSS.n451 5452.27
R255 VSS.n453 VSS.n452 5452.27
R256 VSS.n1892 VSS.n1531 5434.88
R257 VSS.n1892 VSS.n1533 5434.88
R258 VSS.n1533 VSS.n1530 5434.88
R259 VSS.n1531 VSS.n1530 5434.88
R260 VSS.n3169 VSS.n3168 5417.76
R261 VSS.n3021 VSS.n3019 5047.41
R262 VSS.t194 VSS 4888.89
R263 VSS.n3019 VSS.n3018 4736.53
R264 VSS VSS.t194 4408.43
R265 VSS.n385 VSS.n384 4081.58
R266 VSS.n370 VSS.n283 4038.16
R267 VSS.t459 VSS.t468 3877.39
R268 VSS.t465 VSS.t205 3877.39
R269 VSS.n310 VSS.n222 3666.67
R270 VSS.n1540 VSS.n1537 3464.88
R271 VSS.n1543 VSS.n1537 3464.88
R272 VSS.n1540 VSS.n1538 3464.88
R273 VSS.n1543 VSS.n1538 3464.88
R274 VSS.n3169 VSS.n175 3363.82
R275 VSS VSS.t66 3346.36
R276 VSS VSS.t185 3346.36
R277 VSS VSS.t448 3346.36
R278 VSS VSS.t152 3346.36
R279 VSS VSS.t158 3346.36
R280 VSS.t898 VSS 3346.36
R281 VSS.t23 VSS 3346.36
R282 VSS.n3001 VSS.n3000 3340.87
R283 VSS.n3017 VSS.n3016 3323.88
R284 VSS.n198 VSS.n175 3119.26
R285 VSS.t959 VSS.n3343 3111.89
R286 VSS.t949 VSS.t274 3101.92
R287 VSS.t260 VSS.t867 3101.92
R288 VSS.t263 VSS.t208 3101.92
R289 VSS.n386 VSS.n224 2996.82
R290 VSS.n1359 VSS 2973.14
R291 VSS.n3223 VSS.n3222 2937.79
R292 VSS.n172 VSS.n66 2904
R293 VSS.n369 VSS.n368 2881.39
R294 VSS.t236 VSS 2857.47
R295 VSS.t474 VSS 2857.47
R296 VSS VSS.t176 2857.47
R297 VSS VSS.t941 2857.47
R298 VSS VSS.t462 2857.47
R299 VSS VSS.t58 2857.47
R300 VSS.n3224 VSS.n3223 2647.82
R301 VSS.n341 VSS.n340 2595.64
R302 VSS.n399 VSS.n398 2555.51
R303 VSS.n1209 VSS 2552.48
R304 VSS.t944 VSS.t530 2495.02
R305 VSS VSS.n572 2469.73
R306 VSS.t480 VSS 2452.87
R307 VSS.t916 VSS 2452.87
R308 VSS.t200 VSS.t215 2326.44
R309 VSS.t182 VSS.t29 2326.44
R310 VSS.t191 VSS.t35 2326.44
R311 VSS VSS.t226 2081.99
R312 VSS VSS.t179 2081.99
R313 VSS.n3018 VSS.n223 2065.3
R314 VSS.n198 VSS.t965 2053.05
R315 VSS.n3224 VSS.n3170 2012.27
R316 VSS.n207 VSS.t965 1950.07
R317 VSS.t486 VSS.n929 1938.7
R318 VSS.t968 VSS.n207 1926.65
R319 VSS.n1210 VSS.n1209 1896.67
R320 VSS.n1211 VSS.n1210 1896.67
R321 VSS.n1361 VSS.n1211 1896.67
R322 VSS.n1361 VSS.n1360 1896.67
R323 VSS.n1360 VSS.n1359 1896.67
R324 VSS.t226 VSS 1812.26
R325 VSS VSS.t949 1795.4
R326 VSS VSS.t260 1795.4
R327 VSS VSS.t263 1795.4
R328 VSS.t164 VSS 1795.4
R329 VSS.n3345 VSS.n3344 1791.03
R330 VSS.t443 VSS 1786.97
R331 VSS.t223 VSS 1786.97
R332 VSS VSS.t239 1786.97
R333 VSS VSS.t20 1702.68
R334 VSS VSS.n1528 1677.39
R335 VSS.t375 VSS.t0 1593.1
R336 VSS.t574 VSS.t314 1593.1
R337 VSS.t304 VSS.t558 1593.1
R338 VSS.t520 VSS.t523 1584.67
R339 VSS.t4 VSS.t826 1584.67
R340 VSS.t879 VSS.t355 1567.82
R341 VSS.t66 VSS.t901 1550.96
R342 VSS.t185 VSS.t236 1550.96
R343 VSS.t448 VSS.t474 1550.96
R344 VSS.t401 VSS.t8 1550.96
R345 VSS.t152 VSS.t167 1550.96
R346 VSS.t158 VSS.t266 1550.96
R347 VSS.t941 VSS.t898 1550.96
R348 VSS.t462 VSS.t23 1550.96
R349 VSS.t58 VSS.t223 1550.96
R350 VSS.n3023 VSS.t83 1550.96
R351 VSS.n3022 VSS.n3019 1530.43
R352 VSS VSS.t858 1502.01
R353 VSS.n491 VSS.n399 1445.53
R354 VSS.t606 VSS.t685 1416.09
R355 VSS.t197 VSS 1407.66
R356 VSS.t233 VSS 1407.66
R357 VSS.t41 VSS 1407.66
R358 VSS.t188 VSS 1407.66
R359 VSS VSS.t496 1407.66
R360 VSS.t173 VSS 1407.66
R361 VSS.t155 VSS 1399.23
R362 VSS.t79 VSS.t1048 1399.23
R363 VSS VSS.t2 1390.8
R364 VSS.t901 VSS 1306.51
R365 VSS.t274 VSS 1306.51
R366 VSS.t38 VSS 1306.51
R367 VSS VSS.t443 1306.51
R368 VSS.t167 VSS 1306.51
R369 VSS.t867 VSS 1306.51
R370 VSS VSS.t486 1306.51
R371 VSS VSS.t140 1306.51
R372 VSS.t266 VSS 1306.51
R373 VSS.t208 VSS 1306.51
R374 VSS VSS.t149 1306.51
R375 VSS VSS.t919 1306.51
R376 VSS VSS.t944 1306.51
R377 VSS.t471 VSS 1306.51
R378 VSS.t239 VSS 1306.51
R379 VSS.n1657 VSS.n1632 1294.86
R380 VSS.t298 VSS 1289.66
R381 VSS VSS.t104 1289.66
R382 VSS.t677 VSS 1289.66
R383 VSS.t768 VSS 1272.8
R384 VSS.n3402 VSS.t849 1229.99
R385 VSS.n3360 VSS.n3347 1198.25
R386 VSS.n3401 VSS.n3400 1198.25
R387 VSS.n3307 VSS.n86 1198.25
R388 VSS.n113 VSS.n112 1198.25
R389 VSS.n71 VSS.n68 1198.25
R390 VSS.n3342 VSS.n3341 1198.25
R391 VSS.n1529 VSS.n682 1198.25
R392 VSS.n2235 VSS.n2234 1198.25
R393 VSS.n1358 VSS.n1357 1198.25
R394 VSS.n2001 VSS.n1895 1198.25
R395 VSS.n2925 VSS.n2924 1198.25
R396 VSS.n2927 VSS.n2926 1198.25
R397 VSS.n929 VSS.n541 1196.22
R398 VSS.n2754 VSS.n572 1196.22
R399 VSS.n3403 VSS.n3402 1194.5
R400 VSS.n3129 VSS.n3128 1194.5
R401 VSS.n3033 VSS.n219 1194.5
R402 VSS.n3024 VSS.n3023 1194.5
R403 VSS.n3255 VSS.n72 1194.5
R404 VSS.n2875 VSS.n517 1194.5
R405 VSS.n1208 VSS.n1207 1194.5
R406 VSS.n2643 VSS.n640 1194.5
R407 VSS.n1065 VSS.n1064 1194.5
R408 VSS.n1528 VSS.n1527 1194.5
R409 VSS.n2442 VSS.n777 1194.5
R410 VSS.n2369 VSS.n811 1194.5
R411 VSS.n2237 VSS.n2236 1194.5
R412 VSS.t1019 VSS.t971 1188.51
R413 VSS.n3385 VSS.n38 1171.32
R414 VSS.n3114 VSS.n208 1171.32
R415 VSS.n95 VSS.n94 1171.32
R416 VSS.n2236 VSS.t337 1146.36
R417 VSS.t8 VSS 1137.93
R418 VSS.n3332 VSS.n3331 1105.32
R419 VSS VSS.t316 1104.21
R420 VSS.t1123 VSS 1078.93
R421 VSS.t121 VSS.t108 1078.93
R422 VSS.t355 VSS.t347 1078.93
R423 VSS.t734 VSS 1070.5
R424 VSS.t116 VSS 1036.78
R425 VSS.t1048 VSS 1036.78
R426 VSS.n491 VSS.n490 1032.02
R427 VSS.t176 VSS 1019.92
R428 VSS.t468 VSS 1019.92
R429 VSS.t205 VSS 1019.92
R430 VSS.t919 VSS 1019.92
R431 VSS.t608 VSS.t961 1003.07
R432 VSS.t1112 VSS 1003.07
R433 VSS.t293 VSS.t291 1003.07
R434 VSS.n1109 VSS.n1108 999.607
R435 VSS.n2709 VSS.n2708 999.607
R436 VSS.n2681 VSS.n2680 999.607
R437 VSS.t391 VSS.t1080 960.92
R438 VSS.t134 VSS.t131 952.49
R439 VSS.t522 VSS.t520 944.062
R440 VSS.t433 VSS.t498 944.062
R441 VSS.t985 VSS.t745 944.062
R442 VSS.n1208 VSS 927.203
R443 VSS VSS.n640 927.203
R444 VSS.n3402 VSS 918.774
R445 VSS VSS.t310 918.774
R446 VSS VSS.n70 918.774
R447 VSS.t215 VSS 918.774
R448 VSS VSS.n517 918.774
R449 VSS VSS.t197 918.774
R450 VSS.t29 VSS 918.774
R451 VSS VSS.t155 918.774
R452 VSS.t35 VSS 918.774
R453 VSS VSS.n1065 918.774
R454 VSS VSS.t233 918.774
R455 VSS VSS.t41 918.774
R456 VSS VSS.t188 918.774
R457 VSS VSS.t882 918.774
R458 VSS VSS.t173 918.774
R459 VSS VSS.n72 918.774
R460 VSS.t706 VSS 918.774
R461 VSS.n3023 VSS 918.774
R462 VSS.t752 VSS 918.774
R463 VSS.t496 VSS.t77 910.346
R464 VSS.t83 VSS.t673 910.346
R465 VSS VSS.n1529 901.917
R466 VSS.n2235 VSS 901.917
R467 VSS.t525 VSS.t616 893.487
R468 VSS.t751 VSS.t785 893.487
R469 VSS.n2570 VSS.n2569 870.4
R470 VSS.n1209 VSS 851.341
R471 VSS.n1210 VSS 851.341
R472 VSS.t616 VSS.t608 851.341
R473 VSS.n1211 VSS 851.341
R474 VSS VSS.n1361 851.341
R475 VSS.n1360 VSS 851.341
R476 VSS.t514 VSS.t312 851.341
R477 VSS.n1359 VSS 851.341
R478 VSS.t908 VSS 851.341
R479 VSS VSS.n3021 851.341
R480 VSS.t1021 VSS.t662 842.913
R481 VSS.n3019 VSS.n222 839.237
R482 VSS.t617 VSS.t522 834.484
R483 VSS.t961 VSS.t617 834.484
R484 VSS.t1120 VSS.t660 834.484
R485 VSS.t75 VSS.t999 834.484
R486 VSS.t750 VSS.t114 834.484
R487 VSS.t1125 VSS.t313 834.484
R488 VSS.t335 VSS.t782 834.484
R489 VSS.t791 VSS.t687 826.054
R490 VSS.t582 VSS.t302 826.054
R491 VSS.t981 VSS.t4 826.054
R492 VSS.t913 VSS.t139 826.054
R493 VSS.t291 VSS.t518 826.054
R494 VSS.t664 VSS.t1001 826.054
R495 VSS.t717 VSS.t389 826.054
R496 VSS.t772 VSS.t1013 826.054
R497 VSS.t98 VSS.t1023 826.054
R498 VSS.t958 VSS.t79 809.196
R499 VSS.t976 VSS.t768 809.196
R500 VSS.n314 VSS.n313 807.013
R501 VSS.n307 VSS.n306 807.013
R502 VSS.n319 VSS.n290 807.013
R503 VSS.n338 VSS.n337 807.013
R504 VSS.n382 VSS.n381 807.013
R505 VSS.n356 VSS.n355 807.013
R506 VSS.n366 VSS.n365 807.013
R507 VSS.n204 VSS.n203 807.013
R508 VSS.t277 VSS 805.538
R509 VSS.t0 VSS.t525 800.766
R510 VSS.t989 VSS.t12 800.766
R511 VSS.t314 VSS.t573 800.766
R512 VSS.t1115 VSS.t434 800.766
R513 VSS.t690 VSS.t295 792.337
R514 VSS.t10 VSS.t283 792.337
R515 VSS.t973 VSS.t929 792.337
R516 VSS.t671 VSS.t16 792.337
R517 VSS.t668 VSS.t14 792.337
R518 VSS.n315 VSS.n314 785.722
R519 VSS.n306 VSS.n305 785.722
R520 VSS.n325 VSS.n290 785.722
R521 VSS.n337 VSS.n336 785.722
R522 VSS.n381 VSS.n380 785.722
R523 VSS.n357 VSS.n356 785.722
R524 VSS.n365 VSS.n364 785.722
R525 VSS.n203 VSS.n202 785.722
R526 VSS.t749 VSS.t993 783.909
R527 VSS.t179 VSS.t164 775.48
R528 VSS.n3013 VSS.n3012 767.294
R529 VSS.n2997 VSS.n2995 767.294
R530 VSS.n313 VSS.n296 763.106
R531 VSS.n307 VSS.n300 763.106
R532 VSS.n319 VSS.n289 763.106
R533 VSS.n338 VSS.n286 763.106
R534 VSS.n382 VSS.n373 763.106
R535 VSS.n355 VSS.n353 763.106
R536 VSS.n366 VSS.n344 763.106
R537 VSS.n205 VSS.n204 763.106
R538 VSS.n3012 VSS.n3009 763.106
R539 VSS.n2997 VSS.n2994 763.106
R540 VSS.n394 VSS.n393 763.09
R541 VSS.n3184 VSS.n3183 763.09
R542 VSS.n3208 VSS.n3201 763.09
R543 VSS.n3165 VSS.n3164 763.09
R544 VSS.n3146 VSS.n3145 763.09
R545 VSS.n3136 VSS.n184 763.09
R546 VSS.n3328 VSS.n3327 763.09
R547 VSS.n3198 VSS.n3197 763.09
R548 VSS.t1106 VSS.t913 758.621
R549 VSS.t748 VSS.t1009 758.621
R550 VSS.t399 VSS.t697 750.192
R551 VSS.n296 VSS.n295 748.977
R552 VSS.n301 VSS.n300 748.977
R553 VSS.n332 VSS.n286 748.977
R554 VSS.n345 VSS.n344 748.977
R555 VSS.n326 VSS.n289 748.977
R556 VSS.n375 VSS.n373 748.977
R557 VSS.n353 VSS.n352 748.977
R558 VSS.n205 VSS.n201 748.977
R559 VSS.t826 VSS.t6 741.763
R560 VSS.t1016 VSS.t973 741.763
R561 VSS.t357 VSS.t631 741.763
R562 VSS.t322 VSS.t956 741.763
R563 VSS.n393 VSS.n392 732.236
R564 VSS.n3185 VSS.n3184 732.236
R565 VSS.n3209 VSS.n3208 732.236
R566 VSS.n3164 VSS.n3163 732.236
R567 VSS.n3146 VSS.n3141 732.236
R568 VSS.n3137 VSS.n3136 732.236
R569 VSS.n3327 VSS.n3326 732.236
R570 VSS.n3215 VSS.n3198 732.236
R571 VSS.t697 VSS.t710 724.904
R572 VSS.t721 VSS.t610 724.904
R573 VSS.t1082 VSS.t1104 724.904
R574 VSS.t1088 VSS.t1084 724.904
R575 VSS.t1102 VSS.t1100 724.904
R576 VSS.t1098 VSS.t1102 724.904
R577 VSS.t740 VSS.t1025 724.904
R578 VSS.t738 VSS.t740 724.904
R579 VSS.t742 VSS.t738 724.904
R580 VSS.t542 VSS.t742 724.904
R581 VSS.t548 VSS.t542 724.904
R582 VSS.t556 VSS.t552 724.904
R583 VSS.t546 VSS.t556 724.904
R584 VSS.t550 VSS.t546 724.904
R585 VSS.t554 VSS.t550 724.904
R586 VSS.t544 VSS.t554 724.904
R587 VSS.t534 VSS.t528 724.904
R588 VSS.t538 VSS.t534 724.904
R589 VSS.t540 VSS.t538 724.904
R590 VSS.t532 VSS.t540 724.904
R591 VSS.t536 VSS.t532 724.904
R592 VSS.t526 VSS.t536 724.904
R593 VSS.t635 VSS.t639 724.904
R594 VSS.t629 VSS.t633 724.904
R595 VSS.t647 VSS.t645 724.904
R596 VSS.t736 VSS.t732 724.904
R597 VSS.t732 VSS.t789 724.904
R598 VSS.t821 VSS.t578 724.904
R599 VSS.t614 VSS.t507 716.476
R600 VSS.t887 VSS.t655 716.476
R601 VSS.t971 VSS.t793 716.476
R602 VSS.t802 VSS.t1108 716.476
R603 VSS.n3331 VSS.n74 709.47
R604 VSS.t602 VSS.t1032 708.047
R605 VSS.t692 VSS.t690 708.047
R606 VSS.t18 VSS.t300 708.047
R607 VSS.t592 VSS.t85 708.047
R608 VSS.n3334 VSS.n70 708.047
R609 VSS.t132 VSS.t371 708.047
R610 VSS.t809 VSS.t811 708.047
R611 VSS.t333 VSS.t331 708.047
R612 VSS.t560 VSS.t562 708.047
R613 VSS.t566 VSS.t564 708.047
R614 VSS.t756 VSS.t754 708.047
R615 VSS.t410 VSS.t408 708.047
R616 VSS.t406 VSS.t404 708.047
R617 VSS.t841 VSS.t843 708.047
R618 VSS.n3230 VSS.n3229 708.047
R619 VSS.t695 VSS.t401 708.047
R620 VSS.t698 VSS.t695 708.047
R621 VSS.t402 VSS.t698 708.047
R622 VSS.t523 VSS.t127 708.047
R623 VSS.t2 VSS.t375 708.047
R624 VSS.t1043 VSS.t734 708.047
R625 VSS.t12 VSS.t10 708.047
R626 VSS.t361 VSS.t1021 708.047
R627 VSS.t1017 VSS.t1011 708.047
R628 VSS.t805 VSS.t1126 708.047
R629 VSS.t353 VSS.t909 708.047
R630 VSS.t440 VSS.t1123 708.047
R631 VSS.t911 VSS.t995 708.047
R632 VSS.t619 VSS.t621 708.047
R633 VSS.t435 VSS.t954 708.047
R634 VSS.t779 VSS.t794 708.047
R635 VSS.t77 VSS.t908 708.047
R636 VSS.t125 VSS.t746 708.047
R637 VSS.n3333 VSS.n72 708.047
R638 VSS.t255 VSS.t272 708.047
R639 VSS.t16 VSS.t666 708.047
R640 VSS.t102 VSS.t96 708.047
R641 VSS.t987 VSS.t90 708.047
R642 VSS.t50 VSS.t245 708.047
R643 VSS.t14 VSS.t504 708.047
R644 VSS.t715 VSS.t100 708.047
R645 VSS.t513 VSS.t308 708.047
R646 VSS.t702 VSS.t1094 699.617
R647 VSS.t1080 VSS.t414 691.188
R648 VSS.t316 VSS.t249 691.188
R649 VSS.t379 VSS.t730 691.188
R650 VSS VSS.t983 682.76
R651 VSS.n208 VSS.t257 681.482
R652 VSS.n94 VSS.t286 681.482
R653 VSS.t1076 VSS.t830 674.331
R654 VSS VSS.t647 674.331
R655 VSS.t605 VSS.t807 674.331
R656 VSS.t578 VSS.t847 674.331
R657 VSS.t758 VSS.t981 657.471
R658 VSS.t139 VSS.t997 657.471
R659 VSS.t387 VSS.t751 657.471
R660 VSS.t437 VSS.t824 657.471
R661 VSS.t483 VSS 649.043
R662 VSS.t704 VSS.t136 640.614
R663 VSS.t131 VSS.t787 640.614
R664 VSS.n3230 VSS 632.184
R665 VSS VSS.t200 632.184
R666 VSS VSS.n1208 632.184
R667 VSS VSS.n517 632.184
R668 VSS VSS.t182 632.184
R669 VSS VSS.n572 632.184
R670 VSS.n929 VSS 632.184
R671 VSS VSS.t191 632.184
R672 VSS VSS.n640 632.184
R673 VSS.n1065 VSS 632.184
R674 VSS.t20 VSS 632.184
R675 VSS.n1528 VSS 632.184
R676 VSS.t416 VSS.t1074 632.184
R677 VSS.n1529 VSS 632.184
R678 VSS VSS.t480 632.184
R679 VSS.t651 VSS.t381 632.184
R680 VSS VSS.n777 632.184
R681 VSS VSS.t916 632.184
R682 VSS VSS.n2235 632.184
R683 VSS.t349 VSS.t629 623.755
R684 VSS.t713 VSS.t625 615.327
R685 VSS.n811 VSS.t651 615.327
R686 VSS.t653 VSS.t1072 615.327
R687 VSS.t657 VSS.t123 615.327
R688 VSS.t712 VSS.t397 606.898
R689 VSS.t694 VSS.t712 606.898
R690 VSS.t530 VSS.t32 606.898
R691 VSS.t643 VSS.t572 606.898
R692 VSS.t442 VSS.t970 606.898
R693 VSS.t970 VSS.t121 606.898
R694 VSS.t347 VSS.t74 606.898
R695 VSS.t74 VSS.t957 606.898
R696 VSS.t306 VSS.t351 606.898
R697 VSS.t218 VSS.n38 606.351
R698 VSS.n70 VSS.n69 599.125
R699 VSS.n3231 VSS.n3230 599.125
R700 VSS.t1104 VSS.t430 598.467
R701 VSS.t978 VSS.t134 598.467
R702 VSS.t509 VSS.t82 598.467
R703 VSS.t594 VSS.t120 598.467
R704 VSS.t744 VSS.t1029 598.467
R705 VSS.t833 VSS.t1090 590.038
R706 VSS VSS.t758 581.61
R707 VSS.t1078 VSS.t796 581.61
R708 VSS VSS.t911 581.61
R709 VSS.t1117 VSS.t1114 573.181
R710 VSS.n3000 VSS.n175 570.136
R711 VSS VSS.t602 564.751
R712 VSS VSS.t18 564.751
R713 VSS.t85 VSS 564.751
R714 VSS.n398 VSS 564.751
R715 VSS VSS.t132 564.751
R716 VSS VSS.t809 564.751
R717 VSS VSS.t333 564.751
R718 VSS VSS.t560 564.751
R719 VSS VSS.t566 564.751
R720 VSS VSS.t756 564.751
R721 VSS VSS.t410 564.751
R722 VSS VSS.t406 564.751
R723 VSS VSS.t841 564.751
R724 VSS.n1894 VSS 564.751
R725 VSS.n1894 VSS 564.751
R726 VSS.t397 VSS 564.751
R727 VSS.n1894 VSS 564.751
R728 VSS.n1894 VSS 564.751
R729 VSS.t786 VSS.t385 564.751
R730 VSS.n1894 VSS 564.751
R731 VSS.t907 VSS 564.751
R732 VSS.n1894 VSS 564.751
R733 VSS.t272 VSS 564.751
R734 VSS.t96 VSS 564.751
R735 VSS VSS.t987 564.751
R736 VSS.n3332 VSS 564.751
R737 VSS.t670 VSS 564.751
R738 VSS.t245 VSS 564.751
R739 VSS.t100 VSS 564.751
R740 VSS VSS.t513 564.751
R741 VSS.t851 VSS.t849 563.702
R742 VSS VSS.t989 556.322
R743 VSS.t429 VSS.t1096 556.322
R744 VSS.t336 VSS.t969 556.322
R745 VSS VSS.t694 547.894
R746 VSS VSS.t1112 547.894
R747 VSS VSS.t1016 547.894
R748 VSS VSS.t1106 547.894
R749 VSS.t800 VSS.t129 547.894
R750 VSS.t999 VSS 547.894
R751 VSS.t783 VSS.t514 547.894
R752 VSS.t957 VSS 547.894
R753 VSS VSS.t1043 539.465
R754 VSS VSS.t170 539.465
R755 VSS VSS.t453 531.034
R756 VSS VSS.t459 531.034
R757 VSS VSS.t465 531.034
R758 VSS.t922 VSS 531.034
R759 VSS.t55 VSS.t395 526.468
R760 VSS.t876 VSS.t592 522.606
R761 VSS VSS.t391 522.606
R762 VSS VSS.t649 522.606
R763 VSS.t90 VSS.t280 522.606
R764 VSS.n3022 VSS.t670 522.606
R765 VSS.t308 VSS.t252 522.606
R766 VSS VSS.t116 514.177
R767 VSS.t516 VSS.t112 514.177
R768 VSS.t498 VSS 514.177
R769 VSS.t823 VSS.t1120 505.748
R770 VSS VSS.t813 505.748
R771 VSS.t552 VSS.t477 497.318
R772 VSS.t627 VSS.t358 497.318
R773 VSS.t351 VSS 497.318
R774 VSS.t114 VSS.t516 488.889
R775 VSS VSS.t988 480.461
R776 VSS.t428 VSS.t1086 480.461
R777 VSS.t570 VSS.t637 480.461
R778 VSS.t662 VSS 480.461
R779 VSS.t576 VSS 480.461
R780 VSS.t89 VSS 480.461
R781 VSS.t297 VSS 480.461
R782 VSS VSS.t47 473.495
R783 VSS VSS.t935 473.495
R784 VSS VSS.t44 473.495
R785 VSS.n1895 VSS.t63 465.17
R786 VSS VSS.t614 463.603
R787 VSS.t1086 VSS.t1052 463.603
R788 VSS.t1092 VSS.t1068 463.603
R789 VSS.t257 VSS 459.26
R790 VSS.t286 VSS 459.26
R791 VSS.t129 VSS.t426 455.173
R792 VSS.t770 VSS.t783 455.173
R793 VSS.t434 VSS 455.173
R794 VSS.t318 VSS.t433 455.173
R795 VSS.t573 VSS 446.743
R796 VSS VSS.t357 446.743
R797 VSS VSS.t1119 446.743
R798 VSS.t1110 VSS 446.743
R799 VSS.n2236 VSS.t576 446.743
R800 VSS.t781 VSS 446.743
R801 VSS.t689 VSS.t851 438.435
R802 VSS VSS.t1019 438.315
R803 VSS.t528 VSS 429.885
R804 VSS.t729 VSS.t438 429.885
R805 VSS.t359 VSS.t335 429.885
R806 VSS.t47 VSS 426.228
R807 VSS.t935 VSS 426.228
R808 VSS.t44 VSS 426.228
R809 VSS VSS.t55 426.228
R810 VSS.n3170 VSS.n3169 406.803
R811 VSS.t952 VSS 404.599
R812 VSS VSS.t106 404.599
R813 VSS VSS.t440 404.599
R814 VSS.t82 VSS.t511 404.599
R815 VSS.t511 VSS.t729 404.599
R816 VSS.t120 VSS.t580 404.599
R817 VSS.t580 VSS.t359 404.599
R818 VSS.t794 VSS 404.599
R819 VSS.t558 VSS.t991 404.599
R820 VSS VSS.t125 404.599
R821 VSS.t838 VSS.n74 403.983
R822 VSS.t310 VSS.t876 387.74
R823 VSS.t832 VSS.t1092 387.74
R824 VSS.t625 VSS.t383 387.74
R825 VSS.t280 VSS.t706 387.74
R826 VSS.t252 VSS.t752 387.74
R827 VSS.n281 VSS 384.901
R828 VSS.t63 VSS 380.899
R829 VSS.t438 VSS.t318 379.31
R830 VSS VSS.t821 379.31
R831 VSS.t882 VSS.t985 370.882
R832 VSS VSS.t680 370.37
R833 VSS.t966 VSS 370.37
R834 VSS VSS.t1063 370.37
R835 VSS.t839 VSS 370.37
R836 VSS.n1358 VSS.t853 361.798
R837 VSS.n415 VSS.n407 354.26
R838 VSS.n415 VSS.n406 354.26
R839 VSS.n418 VSS.n405 354.26
R840 VSS.n418 VSS.n417 354.26
R841 VSS.n478 VSS.n477 354.26
R842 VSS.n477 VSS.n476 354.26
R843 VSS.n445 VSS.n408 354.26
R844 VSS.n466 VSS.n430 354.26
R845 VSS.n466 VSS.n465 354.26
R846 VSS.n435 VSS.n432 354.26
R847 VSS.n436 VSS.n435 354.26
R848 VSS.n443 VSS.n442 354.26
R849 VSS.n444 VSS.n443 354.26
R850 VSS.n1891 VSS.n1534 353.13
R851 VSS.n1891 VSS.n1890 353.13
R852 VSS.n2160 VSS.n2151 352
R853 VSS VSS.t689 349.704
R854 VSS VSS.t52 341.574
R855 VSS VSS.t489 341.574
R856 VSS VSS.t864 341.574
R857 VSS.t432 VSS.n3401 337.166
R858 VSS.t1096 VSS.t832 337.166
R859 VSS.t383 VSS.t627 337.166
R860 VSS.t1119 VSS 337.166
R861 VSS.n112 VSS.t904 337.166
R862 VSS.t418 VSS.n219 337.166
R863 VSS.n3129 VSS.n187 334.815
R864 VSS.n93 VSS.n86 334.815
R865 VSS.n1890 VSS.n1889 330.486
R866 VSS.t426 VSS.t823 328.736
R867 VSS.t1011 VSS 328.736
R868 VSS VSS.t1110 328.736
R869 VSS.n3014 VSS.n3013 325.502
R870 VSS.n3003 VSS.n2995 325.502
R871 VSS.t456 VSS 325.171
R872 VSS.n1888 VSS.n1534 324.425
R873 VSS VSS.t146 323.541
R874 VSS.n3401 VSS.t687 320.307
R875 VSS VSS.t781 320.307
R876 VSS.n112 VSS.t664 320.307
R877 VSS.n219 VSS.t772 320.307
R878 VSS VSS.t779 311.877
R879 VSS.n3014 VSS.n3008 308.137
R880 VSS.n3004 VSS.n3003 308.137
R881 VSS.n3145 VSS.n3142 304.553
R882 VSS.n3197 VSS.n3195 304.553
R883 VSS.n395 VSS.n394 304.553
R884 VSS.n3183 VSS.n3181 304.553
R885 VSS.n3204 VSS.n3201 304.553
R886 VSS.n3132 VSS.n184 304.553
R887 VSS.n3165 VSS.n179 304.553
R888 VSS.n3329 VSS.n3328 304.553
R889 VSS.t997 VSS 303.449
R890 VSS.t661 VSS 303.449
R891 VSS.t991 VSS.t306 303.449
R892 VSS.n3226 VSS.n3225 299.892
R893 VSS VSS.t432 295.019
R894 VSS.t969 VSS.t594 295.019
R895 VSS.t746 VSS 295.019
R896 VSS.t904 VSS 295.019
R897 VSS VSS.t418 295.019
R898 VSS.n1538 VSS.n1535 292.5
R899 VSS.t369 VSS.n1538 292.5
R900 VSS.n1537 VSS.n1536 292.5
R901 VSS.t369 VSS.n1537 292.5
R902 VSS.t710 VSS 286.591
R903 VSS VSS.t544 286.591
R904 VSS.t81 VSS 286.591
R905 VSS.n1590 VSS.t711 281.25
R906 VSS.t371 VSS 278.161
R907 VSS.t811 VSS 278.161
R908 VSS.t331 VSS 278.161
R909 VSS.t562 VSS 278.161
R910 VSS.t564 VSS 278.161
R911 VSS.t754 VSS 278.161
R912 VSS.t408 VSS 278.161
R913 VSS.t404 VSS 278.161
R914 VSS.t843 VSS 278.161
R915 VSS.n387 VSS.t590 277.575
R916 VSS.t52 VSS 277.529
R917 VSS.t853 VSS 277.529
R918 VSS.t489 VSS 277.529
R919 VSS.t864 VSS 277.529
R920 VSS.n1118 VSS.t1211 276.531
R921 VSS.n587 VSS.t1191 276.531
R922 VSS.n623 VSS.t1192 276.531
R923 VSS.t146 VSS 276.274
R924 VSS VSS.t456 276.274
R925 VSS.n1695 VSS.t403 275.293
R926 VSS.n2443 VSS.t1012 275.293
R927 VSS.n876 VSS.t1111 275.293
R928 VSS.t1025 VSS 269.733
R929 VSS.t660 VSS.t605 269.733
R930 VSS.t385 VSS.t750 269.733
R931 VSS.n571 VSS.t1201 269.488
R932 VSS.n2836 VSS.t1162 269.445
R933 VSS.n395 VSS.n389 266.349
R934 VSS.n3181 VSS.n3178 266.349
R935 VSS.n3204 VSS.n3199 266.349
R936 VSS.n3132 VSS.n182 266.349
R937 VSS.n3161 VSS.n179 266.349
R938 VSS.n3156 VSS.n3142 266.349
R939 VSS.n3329 VSS.n77 266.349
R940 VSS.n3195 VSS.n3194 266.349
R941 VSS.n1671 VSS.t1232 265.317
R942 VSS.n744 VSS.t1152 265.317
R943 VSS.n1066 VSS.t1157 265.298
R944 VSS.n2644 VSS.t1203 265.298
R945 VSS.t585 VSS.n397 263.652
R946 VSS.n397 VSS.t590 263.652
R947 VSS.n1083 VSS.t1167 262.784
R948 VSS.n1084 VSS.t1151 262.784
R949 VSS.n1086 VSS.t1172 262.784
R950 VSS.n1107 VSS.t1212 262.784
R951 VSS.n1674 VSS.t1166 262.784
R952 VSS.n1675 VSS.t1131 262.784
R953 VSS.n591 VSS.t1206 262.784
R954 VSS.n592 VSS.t1238 262.784
R955 VSS.n594 VSS.t1146 262.784
R956 VSS.n2707 VSS.t1178 262.784
R957 VSS.n1595 VSS.t1183 262.784
R958 VSS.n1597 VSS.t1214 262.784
R959 VSS.n1006 VSS.t1187 262.784
R960 VSS.n1008 VSS.t1190 262.784
R961 VSS.n604 VSS.t1207 262.784
R962 VSS.n606 VSS.t1210 262.784
R963 VSS.n607 VSS.t1149 262.784
R964 VSS.n616 VSS.t1155 262.784
R965 VSS.n1388 VSS.t1171 262.784
R966 VSS.n1389 VSS.t1175 262.784
R967 VSS.n731 VSS.t1150 262.784
R968 VSS.n732 VSS.t1156 262.784
R969 VSS.n842 VSS.t1138 262.784
R970 VSS.n2300 VSS.t1144 262.784
R971 VSS.n2494 VSS.t1237 262.784
R972 VSS.n2495 VSS.t1243 262.784
R973 VSS.n865 VSS.t1222 262.784
R974 VSS.n867 VSS.t1227 262.784
R975 VSS.n2174 VSS.t1202 262.784
R976 VSS.n2175 VSS.t1208 262.784
R977 VSS.n1143 VSS.t1229 262.719
R978 VSS.n1183 VSS.t1196 262.719
R979 VSS.n1172 VSS.t1180 262.719
R980 VSS.n514 VSS.t1230 262.719
R981 VSS.n2880 VSS.t1193 262.719
R982 VSS.n1635 VSS.t1234 262.719
R983 VSS.n1635 VSS.t1164 262.719
R984 VSS.n2743 VSS.t1198 262.719
R985 VSS.n555 VSS.t1127 262.719
R986 VSS.n552 VSS.t1160 262.719
R987 VSS.n544 VSS.t1165 262.719
R988 VSS.n1017 VSS.t1188 262.719
R989 VSS.n1040 VSS.t1173 262.719
R990 VSS.n638 VSS.t1169 262.719
R991 VSS.n2619 VSS.t1128 262.719
R992 VSS.n661 VSS.t1241 262.719
R993 VSS.n933 VSS.t1168 262.719
R994 VSS.n960 VSS.t1133 262.719
R995 VSS.n2543 VSS.t1141 262.719
R996 VSS.n1424 VSS.t1221 262.719
R997 VSS.n1457 VSS.t1145 262.719
R998 VSS.n2098 VSS.t1215 262.719
R999 VSS.n1849 VSS.t1181 262.719
R1000 VSS.n497 VSS.t1176 262.719
R1001 VSS.n1784 VSS.t1143 262.719
R1002 VSS.n275 VSS.t1177 262.719
R1003 VSS.t295 VSS 261.303
R1004 VSS.t127 VSS 261.303
R1005 VSS.t393 VSS 261.303
R1006 VSS.t1052 VSS.t1082 261.303
R1007 VSS VSS.t471 261.303
R1008 VSS.t828 VSS.t800 261.303
R1009 VSS VSS.t922 261.303
R1010 VSS VSS.t619 261.303
R1011 VSS VSS.t708 261.303
R1012 VSS VSS.t322 261.303
R1013 VSS VSS.t1015 261.303
R1014 VSS VSS.t442 261.303
R1015 VSS VSS.t671 261.303
R1016 VSS VSS.t668 261.303
R1017 VSS.t502 VSS.t26 260.675
R1018 VSS.n2361 VSS.t1220 259.082
R1019 VSS.n2229 VSS.t1135 259.082
R1020 VSS.n2198 VSS.t1216 259.082
R1021 VSS.n1237 VSS.t1186 259.082
R1022 VSS.n1933 VSS.t1163 259.082
R1023 VSS.n1854 VSS.t1235 259.082
R1024 VSS.n1741 VSS.t1223 259.082
R1025 VSS.n2976 VSS.t1242 259.082
R1026 VSS.n245 VSS.t1233 259.082
R1027 VSS.n447 VSS.n446 255.839
R1028 VSS.n446 VSS.n445 253.365
R1029 VSS.t283 VSS 252.875
R1030 VSS.t1068 VSS.t1088 252.875
R1031 VSS VSS.t828 252.875
R1032 VSS.t106 VSS.t770 252.875
R1033 VSS.t995 VSS 252.875
R1034 VSS.n1587 VSS.t1 251
R1035 VSS.n1587 VSS.t378 251
R1036 VSS.n2449 VSS.t135 251
R1037 VSS.n2470 VSS.t386 251
R1038 VSS.n2274 VSS.t1116 251
R1039 VSS.n2216 VSS.t305 251
R1040 VSS.t680 VSS.t682 248.889
R1041 VSS.t765 VSS.t762 248.889
R1042 VSS.t963 VSS.t966 248.889
R1043 VSS.t1063 VSS.t1066 248.889
R1044 VSS.t817 VSS.t819 248.889
R1045 VSS.t836 VSS.t839 248.889
R1046 VSS.n673 VSS.t417 245.82
R1047 VSS.n2317 VSS.t315 245.82
R1048 VSS.n797 VSS.t380 245.82
R1049 VSS.n902 VSS.t577 245.82
R1050 VSS VSS.t242 244.445
R1051 VSS VSS.t38 244.445
R1052 VSS.t149 VSS 244.445
R1053 VSS.t143 VSS 244.445
R1054 VSS.t1090 VSS.t428 244.445
R1055 VSS.t170 VSS 244.445
R1056 VSS.t938 VSS 244.445
R1057 VSS VSS.t870 244.445
R1058 VSS.n1574 VSS.t521 243.028
R1059 VSS.n1574 VSS.t980 243.028
R1060 VSS.n2406 VSS.t808 243.028
R1061 VSS.n2475 VSS.t806 243.028
R1062 VSS.n2043 VSS.t769 243.028
R1063 VSS.n2249 VSS.t499 243.028
R1064 VSS.n2585 VSS.t1081 242.067
R1065 VSS.n832 VSS.t632 242.067
R1066 VSS VSS.t893 241.573
R1067 VSS.n1522 VSS.t611 240.948
R1068 VSS.n2392 VSS.t731 240.948
R1069 VSS.n16 VSS.t296 240.575
R1070 VSS.n110 VSS.t672 240.575
R1071 VSS.n1482 VSS.t1053 238.675
R1072 VSS.n2349 VSS.t350 238.675
R1073 VSS.n2512 VSS.t814 238.675
R1074 VSS.n2199 VSS.t986 238.675
R1075 VSS.n728 VSS.t531 238.44
R1076 VSS VSS.t932 238.202
R1077 VSS.n7 VSS.t299 237.327
R1078 VSS.n3037 VSS.t669 237.327
R1079 VSS.n3027 VSS.t678 237.327
R1080 VSS.n3259 VSS.t105 237.327
R1081 VSS.n2576 VSS.t1107 237.327
R1082 VSS.n1367 VSS.t1113 237.327
R1083 VSS.t633 VSS.t570 236.016
R1084 VSS.t658 VSS 236.016
R1085 VSS.t1126 VSS.t786 236.016
R1086 VSS.n979 VSS.t11 235.607
R1087 VSS.n2083 VSS.n2082 234.667
R1088 VSS.n783 VSS.t972 230.977
R1089 VSS.n890 VSS.t319 230.977
R1090 VSS.n1603 VSS.t400 229.833
R1091 VSS.n2412 VSS.n788 228.294
R1092 VSS.n2207 VSS.n2148 228.294
R1093 VSS.t269 VSS 228.09
R1094 VSS.t477 VSS.t548 227.587
R1095 VSS.t358 VSS.t643 227.587
R1096 VSS.t637 VSS.t952 227.587
R1097 VSS VSS.t798 227.587
R1098 VSS.n2766 VSS.t469 227.256
R1099 VSS.n2569 VSS.t1026 226.708
R1100 VSS.n3083 VSS.t278 225.427
R1101 VSS.n3108 VSS.t258 225.427
R1102 VSS.n3028 VSS.t871 225.427
R1103 VSS.n3047 VSS.t253 225.427
R1104 VSS.n1544 VSS.n1536 225.13
R1105 VSS.n1539 VSS.n1536 225.13
R1106 VSS.t861 VSS.t873 224.931
R1107 VSS.n2304 VSS.t1139 224.196
R1108 VSS.n1155 VSS.t1137 224.102
R1109 VSS.n644 VSS.t1197 224.102
R1110 VSS.n931 VSS.t464 223.282
R1111 VSS.n676 VSS.n675 222.691
R1112 VSS VSS.n3129 222.222
R1113 VSS.n208 VSS 222.222
R1114 VSS VSS.n86 222.222
R1115 VSS.n94 VSS 222.222
R1116 VSS.n965 VSS.t1132 221.972
R1117 VSS.n776 VSS.n774 221.804
R1118 VSS.t588 VSS.t586 221.451
R1119 VSS.n778 VSS.t1218 220.952
R1120 VSS.n779 VSS.t1224 220.952
R1121 VSS.n1060 VSS.t920 219.972
R1122 VSS.n1589 VSS.n1563 218.506
R1123 VSS.n1589 VSS.n1564 218.506
R1124 VSS.n2312 VSS.n838 218.506
R1125 VSS.n2374 VSS.n809 218.506
R1126 VSS.n763 VSS.n762 218.506
R1127 VSS.n882 VSS.n881 218.506
R1128 VSS.n2239 VSS.n900 218.506
R1129 VSS.n2142 VSS.n2132 218.506
R1130 VSS.n57 VSS.t1184 218.308
R1131 VSS.n3375 VSS.t1205 218.308
R1132 VSS.n25 VSS.t1240 218.308
R1133 VSS.n9 VSS.t1185 218.308
R1134 VSS.n212 VSS.t1159 218.308
R1135 VSS.n3106 VSS.t1154 218.308
R1136 VSS.n221 VSS.t1147 218.308
R1137 VSS.n3046 VSS.t1213 218.308
R1138 VSS.n3241 VSS.t1209 218.308
R1139 VSS.n98 VSS.t1161 218.308
R1140 VSS.n3261 VSS.t1142 218.308
R1141 VSS.n3285 VSS.t1195 218.308
R1142 VSS.n1672 VSS.t1129 218.308
R1143 VSS.n1593 VSS.t1179 218.308
R1144 VSS.n2843 VSS.t1130 218.308
R1145 VSS.n738 VSS.t1148 218.308
R1146 VSS.n2578 VSS.t1136 218.308
R1147 VSS.n877 VSS.t1219 218.308
R1148 VSS.n1268 VSS.t1239 218.308
R1149 VSS.n925 VSS.t1134 218.308
R1150 VSS.n2397 VSS.n794 218.13
R1151 VSS.n511 VSS.t449 217.977
R1152 VSS.n1167 VSS.t186 217.977
R1153 VSS.n662 VSS.t24 217.977
R1154 VSS.n656 VSS.t899 217.977
R1155 VSS.n1154 VSS.t276 217.953
R1156 VSS.n643 VSS.t210 217.953
R1157 VSS.n1175 VSS.t238 217.892
R1158 VSS.n2611 VSS.t943 217.892
R1159 VSS.n212 VSS.t279 217.78
R1160 VSS.n3106 VSS.t259 217.78
R1161 VSS.n221 VSS.t872 217.78
R1162 VSS.n3046 VSS.t254 217.78
R1163 VSS.n1409 VSS.t227 216.933
R1164 VSS.n1156 VSS.t39 216.589
R1165 VSS.n645 VSS.t150 216.589
R1166 VSS.n966 VSS.t284 216.579
R1167 VSS.n839 VSS.t250 215.992
R1168 VSS.n1155 VSS.t40 214.487
R1169 VSS.n644 VSS.t151 214.487
R1170 VSS.n8 VSS.t244 214.456
R1171 VSS.n3 VSS.t243 214.456
R1172 VSS.n58 VSS.t71 214.456
R1173 VSS.n42 VSS.t70 214.456
R1174 VSS.n3376 VSS.t220 214.456
R1175 VSS.n40 VSS.t219 214.456
R1176 VSS.n26 VSS.t878 214.456
R1177 VSS.n32 VSS.t877 214.456
R1178 VSS.n81 VSS.t892 214.456
R1179 VSS.n3244 VSS.t891 214.456
R1180 VSS.n99 VSS.t288 214.456
R1181 VSS.n97 VSS.t287 214.456
R1182 VSS.n3284 VSS.t282 214.456
R1183 VSS.n3280 VSS.t281 214.456
R1184 VSS.n3262 VSS.t940 214.456
R1185 VSS.n115 VSS.t939 214.456
R1186 VSS.n1673 VSS.t455 214.456
R1187 VSS.n1673 VSS.t445 214.456
R1188 VSS.n1683 VSS.t444 214.456
R1189 VSS.n1660 VSS.t454 214.456
R1190 VSS.n1633 VSS.t204 214.456
R1191 VSS.n519 VSS.t203 214.456
R1192 VSS.n1633 VSS.t196 214.456
R1193 VSS.n519 VSS.t195 214.456
R1194 VSS.n518 VSS.t476 214.456
R1195 VSS.n516 VSS.t450 214.456
R1196 VSS.n2899 VSS.t475 214.456
R1197 VSS.n1177 VSS.t187 214.456
R1198 VSS.n1191 VSS.t237 214.456
R1199 VSS.n1071 VSS.t275 214.456
R1200 VSS.n1150 VSS.t951 214.456
R1201 VSS.n1072 VSS.t903 214.456
R1202 VSS.n1078 VSS.t950 214.456
R1203 VSS.n1079 VSS.t68 214.456
R1204 VSS.n1082 VSS.t902 214.456
R1205 VSS.n1082 VSS.t67 214.456
R1206 VSS.n1083 VSS.t212 214.456
R1207 VSS.n1083 VSS.t211 214.456
R1208 VSS.n1084 VSS.t202 214.456
R1209 VSS.n1084 VSS.t201 214.456
R1210 VSS.n1086 VSS.t232 214.456
R1211 VSS.n1086 VSS.t231 214.456
R1212 VSS.n1107 VSS.t217 214.456
R1213 VSS.n1107 VSS.t216 214.456
R1214 VSS.n1674 VSS.t214 214.456
R1215 VSS.n1674 VSS.t213 214.456
R1216 VSS.n1675 VSS.t199 214.456
R1217 VSS.n1675 VSS.t198 214.456
R1218 VSS.n542 VSS.t207 214.456
R1219 VSS.n2823 VSS.t466 214.456
R1220 VSS.n2799 VSS.t206 214.456
R1221 VSS.n2810 VSS.t461 214.456
R1222 VSS.n553 VSS.t470 214.456
R1223 VSS.n2788 VSS.t460 214.456
R1224 VSS.n560 VSS.t178 214.456
R1225 VSS.n2760 VSS.t869 214.456
R1226 VSS.n570 VSS.t177 214.456
R1227 VSS.n576 VSS.t868 214.456
R1228 VSS.n2750 VSS.t262 214.456
R1229 VSS.n577 VSS.t169 214.456
R1230 VSS.n2721 VSS.t261 214.456
R1231 VSS.n2714 VSS.t154 214.456
R1232 VSS.n590 VSS.t168 214.456
R1233 VSS.n590 VSS.t153 214.456
R1234 VSS.n591 VSS.t886 214.456
R1235 VSS.n591 VSS.t885 214.456
R1236 VSS.n592 VSS.t184 214.456
R1237 VSS.n592 VSS.t183 214.456
R1238 VSS.n594 VSS.t62 214.456
R1239 VSS.n594 VSS.t61 214.456
R1240 VSS.n2707 VSS.t31 214.456
R1241 VSS.n2707 VSS.t30 214.456
R1242 VSS.n2844 VSS.t488 214.456
R1243 VSS.n2837 VSS.t487 214.456
R1244 VSS.n2844 VSS.t467 214.456
R1245 VSS.n1594 VSS.t142 214.456
R1246 VSS.n1605 VSS.t141 214.456
R1247 VSS.n1595 VSS.t157 214.456
R1248 VSS.n1595 VSS.t156 214.456
R1249 VSS.n1597 VSS.t230 214.456
R1250 VSS.n1597 VSS.t229 214.456
R1251 VSS.n961 VSS.t25 214.456
R1252 VSS.n941 VSS.t463 214.456
R1253 VSS.n965 VSS.t921 214.456
R1254 VSS.n985 VSS.t285 214.456
R1255 VSS.n986 VSS.t224 214.456
R1256 VSS.n1011 VSS.t60 214.456
R1257 VSS.n996 VSS.t59 214.456
R1258 VSS.n1011 VSS.t225 214.456
R1259 VSS.n1006 VSS.t248 214.456
R1260 VSS.n1006 VSS.t247 214.456
R1261 VSS.n1008 VSS.t235 214.456
R1262 VSS.n1008 VSS.t234 214.456
R1263 VSS.n2613 VSS.t900 214.456
R1264 VSS.n2627 VSS.t942 214.456
R1265 VSS.n2656 VSS.t209 214.456
R1266 VSS.n639 VSS.t265 214.456
R1267 VSS.n634 VSS.t268 214.456
R1268 VSS.n2670 VSS.t264 214.456
R1269 VSS.n619 VSS.t160 214.456
R1270 VSS.n617 VSS.t267 214.456
R1271 VSS.n617 VSS.t159 214.456
R1272 VSS.n604 VSS.t222 214.456
R1273 VSS.n604 VSS.t221 214.456
R1274 VSS.n606 VSS.t193 214.456
R1275 VSS.n606 VSS.t192 214.456
R1276 VSS.n607 VSS.t452 214.456
R1277 VSS.n607 VSS.t451 214.456
R1278 VSS.n616 VSS.t37 214.456
R1279 VSS.n616 VSS.t36 214.456
R1280 VSS.n1388 VSS.t22 214.456
R1281 VSS.n1388 VSS.t21 214.456
R1282 VSS.n1389 VSS.t290 214.456
R1283 VSS.n1389 VSS.t289 214.456
R1284 VSS.n2577 VSS.t915 214.456
R1285 VSS.n681 VSS.t914 214.456
R1286 VSS.n2536 VSS.t479 214.456
R1287 VSS.n2567 VSS.t478 214.456
R1288 VSS.n705 VSS.t33 214.456
R1289 VSS.n737 VSS.t946 214.456
R1290 VSS.n729 VSS.t945 214.456
R1291 VSS.n737 VSS.t34 214.456
R1292 VSS.n731 VSS.t447 214.456
R1293 VSS.n731 VSS.t446 214.456
R1294 VSS.n732 VSS.t43 214.456
R1295 VSS.n732 VSS.t42 214.456
R1296 VSS.n1461 VSS.t931 214.456
R1297 VSS.n1435 VSS.t930 214.456
R1298 VSS.n1434 VSS.t145 214.456
R1299 VSS.n1381 VSS.t144 214.456
R1300 VSS.n1379 VSS.t228 214.456
R1301 VSS.n2490 VSS.t172 214.456
R1302 VSS.n2486 VSS.t171 214.456
R1303 VSS.n812 VSS.t889 214.456
R1304 VSS.n2359 VSS.t888 214.456
R1305 VSS.n2321 VSS.t251 214.456
R1306 VSS.n2304 VSS.t473 214.456
R1307 VSS.n2303 VSS.t472 214.456
R1308 VSS.n842 VSS.t926 214.456
R1309 VSS.n842 VSS.t925 214.456
R1310 VSS.n2300 VSS.t482 214.456
R1311 VSS.n2300 VSS.t481 214.456
R1312 VSS.n778 VSS.t241 214.456
R1313 VSS.n778 VSS.t240 214.456
R1314 VSS.n779 VSS.t897 214.456
R1315 VSS.n779 VSS.t896 214.456
R1316 VSS.n2494 VSS.t190 214.456
R1317 VSS.n2494 VSS.t189 214.456
R1318 VSS.n2495 VSS.t948 214.456
R1319 VSS.n2495 VSS.t947 214.456
R1320 VSS.n2179 VSS.t181 214.456
R1321 VSS.n2171 VSS.t180 214.456
R1322 VSS.n2179 VSS.t166 214.456
R1323 VSS.n2163 VSS.t165 214.456
R1324 VSS.n2197 VSS.t884 214.456
R1325 VSS.n2201 VSS.t883 214.456
R1326 VSS.n2228 VSS.t485 214.456
R1327 VSS.n2124 VSS.t484 214.456
R1328 VSS.n2112 VSS.t881 214.456
R1329 VSS.n2085 VSS.t880 214.456
R1330 VSS.n878 VSS.t924 214.456
R1331 VSS.n868 VSS.t923 214.456
R1332 VSS.n865 VSS.t928 214.456
R1333 VSS.n865 VSS.t927 214.456
R1334 VSS.n867 VSS.t918 214.456
R1335 VSS.n867 VSS.t917 214.456
R1336 VSS.n2174 VSS.t857 214.456
R1337 VSS.n2174 VSS.t856 214.456
R1338 VSS.n2175 VSS.t175 214.456
R1339 VSS.n2175 VSS.t174 214.456
R1340 VSS.n1932 VSS.t28 214.456
R1341 VSS.n1930 VSS.t27 214.456
R1342 VSS.n1917 VSS.t866 214.456
R1343 VSS.n1916 VSS.t865 214.456
R1344 VSS.n1977 VSS.t65 214.456
R1345 VSS.n1897 VSS.t64 214.456
R1346 VSS.n926 VSS.t934 214.456
R1347 VSS.n2012 VSS.t933 214.456
R1348 VSS.n1324 VSS.t491 214.456
R1349 VSS.n1323 VSS.t490 214.456
R1350 VSS.n1308 VSS.t855 214.456
R1351 VSS.n1306 VSS.t854 214.456
R1352 VSS.n1294 VSS.t54 214.456
R1353 VSS.n1292 VSS.t53 214.456
R1354 VSS.n1269 VSS.t895 214.456
R1355 VSS.n1224 VSS.t894 214.456
R1356 VSS.n1230 VSS.t271 214.456
R1357 VSS.n1236 VSS.t270 214.456
R1358 VSS.n240 VSS.t863 214.456
R1359 VSS.n246 VSS.t862 214.456
R1360 VSS.n2975 VSS.t875 214.456
R1361 VSS.n2978 VSS.t874 214.456
R1362 VSS.n258 VSS.t147 214.456
R1363 VSS.n2960 VSS.t148 214.456
R1364 VSS.n277 VSS.t49 214.456
R1365 VSS.n271 VSS.t48 214.456
R1366 VSS.n1740 VSS.t163 214.456
R1367 VSS.n1739 VSS.t162 214.456
R1368 VSS.n1778 VSS.t937 214.456
R1369 VSS.n1755 VSS.t936 214.456
R1370 VSS.n495 VSS.t46 214.456
R1371 VSS.n1760 VSS.t45 214.456
R1372 VSS.n1719 VSS.t457 214.456
R1373 VSS.n1712 VSS.t458 214.456
R1374 VSS.n1850 VSS.t57 214.456
R1375 VSS.n1838 VSS.t56 214.456
R1376 VSS.n1853 VSS.t860 214.456
R1377 VSS.n1851 VSS.t859 214.456
R1378 VSS.n1539 VSS.n1535 214.409
R1379 VSS.n1545 VSS.n1544 213.911
R1380 VSS.n3340 VSS.n3339 212.78
R1381 VSS.n2406 VSS.n2405 212.317
R1382 VSS.t596 VSS.t367 211.237
R1383 VSS VSS.t907 210.728
R1384 VSS.n3226 VSS.t838 209.996
R1385 VSS.n2431 VSS.n2430 207.965
R1386 VSS.n2214 VSS.n2144 207.965
R1387 VSS.n1464 VSS.n1463 206.909
R1388 VSS.n3225 VSS.n3224 206.876
R1389 VSS.n2357 VSS.n2356 205.971
R1390 VSS.n1493 VSS.n1485 205.899
R1391 VSS.n1496 VSS.n1495 205.899
R1392 VSS.n1487 VSS.n1486 205.481
R1393 VSS.n2344 VSS.n822 205.481
R1394 VSS.n2534 VSS.n2533 205.385
R1395 VSS.n676 VSS.n674 204.692
R1396 VSS.n1503 VSS.n1502 204.692
R1397 VSS.n48 VSS.n44 204.457
R1398 VSS.n3249 VSS.n3248 204.457
R1399 VSS.n2118 VSS.n905 204.457
R1400 VSS.n2118 VSS.n906 204.457
R1401 VSS.n2134 VSS.n2133 204.457
R1402 VSS.n984 VSS.n983 204.201
R1403 VSS.n2037 VSS.n2036 204.201
R1404 VSS.n2097 VSS.n2096 204.201
R1405 VSS.n685 VSS.n684 202.724
R1406 VSS.n2555 VSS.n695 202.724
R1407 VSS.n1511 VSS.n1476 202.724
R1408 VSS.n2375 VSS.n808 202.724
R1409 VSS.n2378 VSS.n2377 202.724
R1410 VSS.t655 VSS 202.299
R1411 VSS.t785 VSS.t978 202.299
R1412 VSS.t909 VSS.t1125 202.299
R1413 VSS.t1029 VSS.t304 202.299
R1414 VSS.n704 VSS.n703 201.458
R1415 VSS.n2351 VSS.n817 201.458
R1416 VSS.n2598 VSS.n672 201.129
R1417 VSS.n2526 VSS.n708 201.129
R1418 VSS.n2528 VSS.n707 201.129
R1419 VSS.n819 VSS.n818 201.129
R1420 VSS.n2782 VSS.n2781 200.692
R1421 VSS.n2320 VSS.n2319 200.692
R1422 VSS.n1982 VSS.n1981 200.692
R1423 VSS.n2962 VSS.n2961 200.692
R1424 VSS.n1827 VSS.n1826 200.692
R1425 VSS.n2437 VSS.n2436 200.516
R1426 VSS.n886 VSS.n885 200.516
R1427 VSS.n718 VSS.n717 200.508
R1428 VSS.n699 VSS.n698 200.508
R1429 VSS.n2542 VSS.n700 200.508
R1430 VSS.n1481 VSS.n1480 200.508
R1431 VSS.n2329 VSS.n2328 200.508
R1432 VSS.n2362 VSS.n2360 200.508
R1433 VSS.n2368 VSS.n2367 200.508
R1434 VSS.n3399 VSS.n15 200.231
R1435 VSS.n3391 VSS.n21 200.231
R1436 VSS.n3268 VSS.n3267 200.231
R1437 VSS.n108 VSS.n107 200.231
R1438 VSS.n2584 VSS.n679 200.231
R1439 VSS.n776 VSS.n775 200.127
R1440 VSS.n2279 VSS.n880 200.127
R1441 VSS.n30 VSS.n24 200.105
R1442 VSS.n3048 VSS.n3045 200.105
R1443 VSS.n3077 VSS.n214 200.105
R1444 VSS.n3287 VSS.n3282 200.105
R1445 VSS.n2847 VSS.n538 199.739
R1446 VSS.n2847 VSS.n539 199.739
R1447 VSS.n1521 VSS.n1465 199.739
R1448 VSS.n790 VSS.n789 199.739
R1449 VSS.n896 VSS.n895 199.739
R1450 VSS.n1228 VSS.n1227 199.739
R1451 VSS.n1226 VSS.n1225 199.739
R1452 VSS.n1274 VSS.n1222 199.739
R1453 VSS.n1302 VSS.n1301 199.739
R1454 VSS.n1320 VSS.n1319 199.739
R1455 VSS.n2022 VSS.n919 199.739
R1456 VSS.n928 VSS.n927 199.739
R1457 VSS.n1913 VSS.n1912 199.739
R1458 VSS.n1921 VSS.n1920 199.739
R1459 VSS.n1939 VSS.n1929 199.739
R1460 VSS.n1711 VSS.n1710 199.739
R1461 VSS.n1039 VSS.n981 199.662
R1462 VSS.n1580 VSS.n1568 199.53
R1463 VSS.n1580 VSS.n1570 199.53
R1464 VSS.n1497 VSS.n1494 199.53
R1465 VSS.n2399 VSS.n2398 199.53
R1466 VSS.n2469 VSS.n764 199.53
R1467 VSS.n2047 VSS.n2046 199.53
R1468 VSS.n2267 VSS.n888 199.53
R1469 VSS.n2208 VSS.n2147 199.53
R1470 VSS.t420 VSS 198.519
R1471 VSS.t682 VSS 198.519
R1472 VSS VSS.t765 198.519
R1473 VSS VSS.t963 198.519
R1474 VSS.t341 VSS 198.519
R1475 VSS.t1066 VSS 198.519
R1476 VSS VSS.t817 198.519
R1477 VSS VSS.t836 198.519
R1478 VSS VSS.n38 197.724
R1479 VSS.n3040 VSS.n3039 197.476
R1480 VSS.n3034 VSS.n218 197.476
R1481 VSS.n1375 VSS.n1374 197.476
R1482 VSS.n1667 VSS.n1629 196.831
R1483 VSS.n2327 VSS.n831 196.589
R1484 VSS.n2477 VSS.n759 196.589
R1485 VSS.n1378 VSS.n1377 196.442
R1486 VSS.n1510 VSS.n1477 196.442
R1487 VSS.n815 VSS.n814 196.442
R1488 VSS.n2479 VSS.n2478 196.442
R1489 VSS.n2501 VSS.n2489 196.442
R1490 VSS.n308 VSS.n307 195
R1491 VSS.n309 VSS.n308 195
R1492 VSS.n305 VSS.n304 195
R1493 VSS.n304 VSS.n303 195
R1494 VSS.n313 VSS.n312 195
R1495 VSS.n312 VSS.n311 195
R1496 VSS.n316 VSS.n315 195
R1497 VSS.n317 VSS.n316 195
R1498 VSS.n320 VSS.n319 195
R1499 VSS.n321 VSS.n320 195
R1500 VSS.n325 VSS.n324 195
R1501 VSS.n324 VSS.n323 195
R1502 VSS.n367 VSS.n366 195
R1503 VSS.n368 VSS.n367 195
R1504 VSS.n364 VSS.n363 195
R1505 VSS.n363 VSS.n362 195
R1506 VSS.n339 VSS.n338 195
R1507 VSS.n340 VSS.n339 195
R1508 VSS.n336 VSS.n335 195
R1509 VSS.n335 VSS.n334 195
R1510 VSS.n391 VSS.n282 195
R1511 VSS.n282 VSS.n281 195
R1512 VSS.n3183 VSS.n3182 195
R1513 VSS.n3182 VSS.n3171 195
R1514 VSS.n3187 VSS.n3186 195
R1515 VSS.n3188 VSS.n3187 195
R1516 VSS.n3203 VSS.n3201 195
R1517 VSS.n3203 VSS.n3172 195
R1518 VSS.n3202 VSS.n3200 195
R1519 VSS.n3202 VSS.n3190 195
R1520 VSS.n3145 VSS.n3144 195
R1521 VSS.n3144 VSS.n174 195
R1522 VSS.n3155 VSS.n3154 195
R1523 VSS.n3154 VSS.n3153 195
R1524 VSS.n186 VSS.n184 195
R1525 VSS.n186 VSS.n176 195
R1526 VSS.n185 VSS.n183 195
R1527 VSS.n3131 VSS.n185 195
R1528 VSS.n3166 VSS.n3165 195
R1529 VSS.n3167 VSS.n3166 195
R1530 VSS.n3149 VSS.n180 195
R1531 VSS.n3150 VSS.n3149 195
R1532 VSS.n3328 VSS.n76 195
R1533 VSS.n3225 VSS.n76 195
R1534 VSS.n202 VSS.n197 195
R1535 VSS.n197 VSS.n187 195
R1536 VSS.n204 VSS.n199 195
R1537 VSS.n199 VSS.n198 195
R1538 VSS.n3197 VSS.n3196 195
R1539 VSS.n3196 VSS.n3173 195
R1540 VSS.n3217 VSS.n3216 195
R1541 VSS.n3218 VSS.n3217 195
R1542 VSS.n3325 VSS.n75 195
R1543 VSS.n93 VSS.n75 195
R1544 VSS.n355 VSS.n354 195
R1545 VSS.n354 VSS.n283 195
R1546 VSS.n358 VSS.n357 195
R1547 VSS.n359 VSS.n358 195
R1548 VSS.n383 VSS.n382 195
R1549 VSS.n384 VSS.n383 195
R1550 VSS.n380 VSS.n379 195
R1551 VSS.n379 VSS.n378 195
R1552 VSS.n394 VSS.n388 195
R1553 VSS.n388 VSS.n387 195
R1554 VSS.n3013 VSS.n226 195
R1555 VSS.n226 VSS.t774 195
R1556 VSS.n3009 VSS.n225 195
R1557 VSS.n2999 VSS.n2995 195
R1558 VSS.t604 VSS.n2999 195
R1559 VSS.n2996 VSS.n2994 195
R1560 VSS.t604 VSS.n2996 195
R1561 VSS.n398 VSS.t585 194.406
R1562 VSS.t112 VSS.t387 193.87
R1563 VSS.t824 VSS.t509 193.87
R1564 VSS.n2780 VSS.n2779 190.399
R1565 VSS.n836 VSS.n835 190.399
R1566 VSS.n1980 VSS.n1979 190.399
R1567 VSS.n263 VSS.n261 190.399
R1568 VSS.n1825 VSS.n1824 190.399
R1569 VSS.n2083 VSS.n2042 189.268
R1570 VSS.n2160 VSS.n2159 189.201
R1571 VSS.n3010 VSS.n225 188.968
R1572 VSS.t312 VSS.t805 185.441
R1573 VSS.t1015 VSS.t336 185.441
R1574 VSS.t673 VSS.n3022 185.441
R1575 VSS.n438 VSS.t69 179.556
R1576 VSS.t365 VSS 177.529
R1577 VSS.t412 VSS 177.529
R1578 VSS.t500 VSS 177.529
R1579 VSS.t568 VSS 177.529
R1580 VSS.t1121 VSS 177.529
R1581 VSS.t302 VSS 177.012
R1582 VSS.t123 VSS.t75 177.012
R1583 VSS.t685 VSS.t1115 177.012
R1584 VSS.t708 VSS.t437 177.012
R1585 VSS VSS.t717 177.012
R1586 VSS VSS.t98 177.012
R1587 VSS.t586 VSS 176.633
R1588 VSS.n398 VSS 176.633
R1589 VSS.n3011 VSS.n3010 174.41
R1590 VSS.t893 VSS 174.157
R1591 VSS.t932 VSS 174.157
R1592 VSS.t1074 VSS.t429 168.583
R1593 VSS.t798 VSS.t658 168.583
R1594 VSS.n387 VSS.n386 163.297
R1595 VSS.n3368 VSS.t1061 162.471
R1596 VSS.n3363 VSS.t1038 162.471
R1597 VSS.n3359 VSS.t326 162.471
R1598 VSS.n3354 VSS.t589 162.471
R1599 VSS.n3394 VSS.t691 162.471
R1600 VSS.n3315 VSS.t344 162.471
R1601 VSS.n3310 VSS.t1064 162.471
R1602 VSS.n3306 VSS.t820 162.471
R1603 VSS.n3301 VSS.t840 162.471
R1604 VSS.n3273 VSS.t17 162.471
R1605 VSS.n2925 VSS 162.179
R1606 VSS.n127 VSS.t374 162.022
R1607 VSS.n132 VSS.t812 162.022
R1608 VSS.n137 VSS.t332 162.022
R1609 VSS.n142 VSS.t601 162.022
R1610 VSS.n147 VSS.t598 162.022
R1611 VSS.n152 VSS.t755 162.022
R1612 VSS.n157 VSS.t409 162.022
R1613 VSS.n162 VSS.t405 162.022
R1614 VSS.n167 VSS.t846 162.022
R1615 VSS.n131 VSS.t133 162.022
R1616 VSS.n136 VSS.t1070 162.022
R1617 VSS.n141 VSS.t1051 162.022
R1618 VSS.n146 VSS.t561 162.022
R1619 VSS.n151 VSS.t567 162.022
R1620 VSS.n156 VSS.t761 162.022
R1621 VSS.n161 VSS.t776 162.022
R1622 VSS.n166 VSS.t778 162.022
R1623 VSS.n171 VSS.t842 162.022
R1624 VSS.n3399 VSS.t1033 160.046
R1625 VSS.n3391 VSS.t301 160.046
R1626 VSS.n3268 VSS.t256 160.046
R1627 VSS.n108 VSS.t103 160.046
R1628 VSS.n127 VSS.t372 160.017
R1629 VSS.n132 VSS.t1071 160.017
R1630 VSS.n137 VSS.t1050 160.017
R1631 VSS.n142 VSS.t563 160.017
R1632 VSS.n147 VSS.t565 160.017
R1633 VSS.n152 VSS.t760 160.017
R1634 VSS.n157 VSS.t775 160.017
R1635 VSS.n162 VSS.t777 160.017
R1636 VSS.n167 VSS.t844 160.017
R1637 VSS.n60 VSS.t1058 160.017
R1638 VSS.n3361 VSS.t1041 160.017
R1639 VSS.n3350 VSS.t329 160.017
R1640 VSS.n39 VSS.t587 160.017
R1641 VSS.n3392 VSS.t693 160.017
R1642 VSS.n22 VSS.t19 160.017
R1643 VSS.n83 VSS.t342 160.017
R1644 VSS.n3308 VSS.t1067 160.017
R1645 VSS.n89 VSS.t818 160.017
R1646 VSS.n3299 VSS.t837 160.017
R1647 VSS.n3275 VSS.t667 160.017
R1648 VSS.n3292 VSS.t97 160.017
R1649 VSS.n131 VSS.t373 160.017
R1650 VSS.n136 VSS.t810 160.017
R1651 VSS.n141 VSS.t334 160.017
R1652 VSS.n146 VSS.t600 160.017
R1653 VSS.n151 VSS.t599 160.017
R1654 VSS.n156 VSS.t757 160.017
R1655 VSS.n161 VSS.t411 160.017
R1656 VSS.n166 VSS.t407 160.017
R1657 VSS.n171 VSS.t845 160.017
R1658 VSS.n16 VSS.t603 158.534
R1659 VSS.n110 VSS.t273 158.534
R1660 VSS.t1045 VSS.n1358 157.304
R1661 VSS.n1895 VSS.t72 157.304
R1662 VSS.n3085 VSS.t424 157.291
R1663 VSS.n3087 VSS.t681 157.291
R1664 VSS.n191 VSS.t763 157.291
R1665 VSS.n192 VSS.t967 157.291
R1666 VSS.n3036 VSS.t51 157.291
R1667 VSS.n3063 VSS.t15 157.291
R1668 VSS.n3056 VSS.t716 157.291
R1669 VSS.n3095 VSS.t421 155.286
R1670 VSS.n3089 VSS.t683 155.286
R1671 VSS.n3123 VSS.t766 155.286
R1672 VSS.n3117 VSS.t964 155.286
R1673 VSS.n3068 VSS.t246 155.286
R1674 VSS.n3061 VSS.t505 155.286
R1675 VSS.n3054 VSS.t101 155.286
R1676 VSS.n2484 VSS.t910 154.131
R1677 VSS.n1045 VSS.t1044 152.381
R1678 VSS.n2513 VSS.t354 152.381
R1679 VSS.n2493 VSS.t996 152.381
R1680 VSS.n2781 VSS.n559 152
R1681 VSS.n2319 VSS.n2318 152
R1682 VSS.n1981 VSS.n1911 152
R1683 VSS.n1826 VSS.n1714 152
R1684 VSS.n2963 VSS.n2962 152
R1685 VSS.n977 VSS.t735 150.101
R1686 VSS.n2493 VSS.t912 150.101
R1687 VSS.n2926 VSS.t161 149.954
R1688 VSS VSS.n3342 144.951
R1689 VSS.n2464 VSS.t979 144.886
R1690 VSS.n2273 VSS.t686 144.886
R1691 VSS.t796 VSS.t612 143.296
R1692 VSS VSS.n777 143.296
R1693 VSS VSS.t483 143.296
R1694 VSS.n474 VSS.n473 139.727
R1695 VSS.t604 VSS.n223 137.912
R1696 VSS.n3001 VSS.t604 137.912
R1697 VSS.t960 VSS 135.415
R1698 VSS.t1094 VSS.t833 134.867
R1699 VSS.t621 VSS.t1117 134.867
R1700 VSS.t1114 VSS.t606 134.867
R1701 VSS.t782 VSS.t976 134.867
R1702 VSS.n71 VSS.t339 133.507
R1703 VSS.t430 VSS.t1078 126.438
R1704 VSS.n1632 VSS.t9 124.688
R1705 VSS.n431 VSS.n430 123.882
R1706 VSS.t26 VSS 122.472
R1707 VSS.n2490 VSS.t1231 121.927
R1708 VSS.n1917 VSS.t1228 121.927
R1709 VSS.n1324 VSS.t1158 121.927
R1710 VSS.n1308 VSS.t1225 121.927
R1711 VSS.n1294 VSS.t1170 121.927
R1712 VSS VSS.t968 121.481
R1713 VSS VSS.t835 121.481
R1714 VSS.n3018 VSS.n3017 120.984
R1715 VSS.n3016 VSS.n3015 118.285
R1716 VSS.t612 VSS 118.008
R1717 VSS.t32 VSS.t526 118.008
R1718 VSS.t572 VSS.t635 118.008
R1719 VSS.t954 VSS.t81 118.008
R1720 VSS.n452 VSS.n448 117.001
R1721 VSS.n452 VSS.t519 117.001
R1722 VSS.n449 VSS.n447 117.001
R1723 VSS.n449 VSS.t519 117.001
R1724 VSS.n480 VSS.n412 117.001
R1725 VSS.n480 VSS.t88 117.001
R1726 VSS.n410 VSS.n408 117.001
R1727 VSS.t88 VSS.n410 117.001
R1728 VSS.n444 VSS.n440 117.001
R1729 VSS.n440 VSS.t419 117.001
R1730 VSS.n442 VSS.n439 117.001
R1731 VSS.t419 VSS.n439 117.001
R1732 VSS.n414 VSS.n407 117.001
R1733 VSS.n414 VSS.t138 117.001
R1734 VSS.n413 VSS.n406 117.001
R1735 VSS.n413 VSS.t138 117.001
R1736 VSS.n437 VSS.n436 117.001
R1737 VSS.t419 VSS.n437 117.001
R1738 VSS.n434 VSS.n432 117.001
R1739 VSS.t419 VSS.n434 117.001
R1740 VSS.n405 VSS.n403 117.001
R1741 VSS.t138 VSS.n403 117.001
R1742 VSS.n417 VSS.n402 117.001
R1743 VSS.t138 VSS.n402 117.001
R1744 VSS.n465 VSS.n429 117.001
R1745 VSS.t419 VSS.n429 117.001
R1746 VSS.n430 VSS.n428 117.001
R1747 VSS.t419 VSS.n428 117.001
R1748 VSS.n476 VSS.n421 117.001
R1749 VSS.t86 VSS.n421 117.001
R1750 VSS.n479 VSS.n478 117.001
R1751 VSS.t86 VSS.n479 117.001
R1752 VSS.n2180 VSS.t1200 116.734
R1753 VSS.n1415 VSS.t1189 116.734
R1754 VSS.n2076 VSS.n2045 114.377
R1755 VSS.n1450 VSS.n1449 110.349
R1756 VSS.n898 VSS.n897 110.349
R1757 VSS.t631 VSS.t713 109.579
R1758 VSS.t649 VSS.n811 109.579
R1759 VSS.t1072 VSS.t736 109.579
R1760 VSS.t730 VSS.t661 109.579
R1761 VSS.t993 VSS.t744 109.579
R1762 VSS.n1449 VSS.t80 108.505
R1763 VSS.n2045 VSS.t360 108.505
R1764 VSS.n897 VSS.t822 108.505
R1765 VSS VSS.t343 106.942
R1766 VSS.t494 VSS.t506 102.992
R1767 VSS.t492 VSS.t675 102.992
R1768 VSS.n1079 VSS.t1140 102.353
R1769 VSS.n2714 VSS.t1226 102.353
R1770 VSS.n619 VSS.t1199 102.353
R1771 VSS.n983 VSS.t398 101.43
R1772 VSS.n2036 VSS.t122 101.43
R1773 VSS.n2096 VSS.t348 101.43
R1774 VSS.t929 VSS.t958 101.15
R1775 VSS.t639 VSS.t349 101.15
R1776 VSS.n1004 VSS.t1182 99.7825
R1777 VSS.n2172 VSS.t1204 99.7825
R1778 VSS.t320 VSS.t596 98.8769
R1779 VSS.t367 VSS.t623 98.8769
R1780 VSS.t363 VSS.t365 98.8769
R1781 VSS.t118 VSS.t1045 98.8769
R1782 VSS.t974 VSS.t412 98.8769
R1783 VSS.t803 VSS.t500 98.8769
R1784 VSS.t1027 VSS.t72 98.8769
R1785 VSS.t905 VSS.t568 98.8769
R1786 VSS.t723 VSS.t1121 98.8769
R1787 VSS.t700 VSS.t502 98.8769
R1788 VSS.t1100 VSS.t416 92.7208
R1789 VSS VSS.t641 92.7208
R1790 VSS.t381 VSS.t653 92.7208
R1791 VSS.t793 VSS.t802 92.7208
R1792 VSS.t1108 VSS.t657 92.7208
R1793 VSS.t745 VSS 92.7208
R1794 VSS.n476 VSS.n475 89.224
R1795 VSS.n465 VSS.n464 89.224
R1796 VSS.n463 VSS.n432 89.224
R1797 VSS.n436 VSS.n433 89.224
R1798 VSS.n442 VSS.n441 89.224
R1799 VSS.n456 VSS.n444 89.224
R1800 VSS.t873 VSS 88.8318
R1801 VSS.t161 VSS 88.8318
R1802 VSS.n455 VSS.n447 88.4711
R1803 VSS.t762 VSS.n187 85.9264
R1804 VSS.t819 VSS.n93 85.9264
R1805 VSS.n483 VSS.n408 84.7064
R1806 VSS.t988 VSS.t692 84.2917
R1807 VSS.t453 VSS.t402 84.2917
R1808 VSS.t666 VSS.t89 84.2917
R1809 VSS.t504 VSS.t297 84.2917
R1810 VSS VSS.t269 84.2702
R1811 VSS.n3221 VSS 83.8426
R1812 VSS.n484 VSS.n407 80.1887
R1813 VSS.n486 VSS.n406 80.1887
R1814 VSS.n487 VSS.n405 80.1887
R1815 VSS.n417 VSS.n404 80.1887
R1816 VSS.n1894 VSS 76.6073
R1817 VSS.t1009 VSS.t293 75.8626
R1818 VSS VSS.n1894 75.2814
R1819 VSS.n1568 VSS.t618 74.8666
R1820 VSS.n1570 VSS.t609 74.8666
R1821 VSS.n1494 VSS.t1069 74.8666
R1822 VSS.n831 VSS.t714 74.8666
R1823 VSS.n2398 VSS.t801 74.8666
R1824 VSS.n764 VSS.t113 74.8666
R1825 VSS.n759 VSS.t515 74.8666
R1826 VSS.n2046 VSS.t595 74.8666
R1827 VSS.n888 VSS.t510 74.8666
R1828 VSS.n2147 VSS.t292 74.8666
R1829 VSS.n24 VSS.t593 72.8576
R1830 VSS.n44 VSS.t852 72.8576
R1831 VSS.n3045 VSS.t309 72.8576
R1832 VSS.n214 VSS.t674 72.8576
R1833 VSS.n3248 VSS.t676 72.8576
R1834 VSS.n3282 VSS.t91 72.8576
R1835 VSS.n905 VSS.t78 72.8576
R1836 VSS.n906 VSS.t1031 72.8576
R1837 VSS.n2133 VSS.t352 72.8576
R1838 VSS.t419 VSS.n426 72.7469
R1839 VSS.n460 VSS.t519 72.7469
R1840 VSS.t395 VSS.t110 71.7175
R1841 VSS.t623 VSS 70.787
R1842 VSS.t423 VSS.t277 67.6928
R1843 VSS.t136 VSS.t1017 67.4335
R1844 VSS.t787 VSS.t704 67.4335
R1845 VSS.t956 VSS.t435 67.4335
R1846 VSS.n422 VSS.t138 66.396
R1847 VSS.t86 VSS.n420 66.396
R1848 VSS.n482 VSS.n409 64.8307
R1849 VSS.n3016 VSS.t774 61.6916
R1850 VSS VSS.t861 61.1229
R1851 VSS VSS.n2925 61.1229
R1852 VSS.n1532 VSS.n63 59.6152
R1853 VSS.n1541 VSS.n63 59.6152
R1854 VSS.t983 VSS.t748 59.0043
R1855 VSS.n451 VSS.n450 58.7133
R1856 VSS.n15 VSS.t688 58.5719
R1857 VSS.n21 VSS.t303 58.5719
R1858 VSS.n3039 VSS.t99 58.5719
R1859 VSS.n218 VSS.t773 58.5719
R1860 VSS.n3267 VSS.t665 58.5719
R1861 VSS.n107 VSS.t718 58.5719
R1862 VSS.n679 VSS.t998 58.5719
R1863 VSS.n1374 VSS.t982 58.5719
R1864 VSS.n3343 VSS.t960 57.2177
R1865 VSS.t506 VSS.t492 57.2177
R1866 VSS.n3333 VSS.n71 57.2177
R1867 VSS VSS.n492 56.2331
R1868 VSS.n391 VSS.n389 54.2123
R1869 VSS.n3186 VSS.n3178 54.2123
R1870 VSS.n3200 VSS.n3199 54.2123
R1871 VSS.n3161 VSS.n180 54.2123
R1872 VSS.n3156 VSS.n3155 54.2123
R1873 VSS.n183 VSS.n182 54.2123
R1874 VSS.n3325 VSS.n77 54.2123
R1875 VSS.n3216 VSS.n3194 54.2123
R1876 VSS.n1534 VSS.n1531 53.1823
R1877 VSS.n1531 VSS.t725 53.1823
R1878 VSS.n1890 VSS.n1533 53.1823
R1879 VSS.n1533 VSS.n1532 53.1823
R1880 VSS.n1544 VSS.n1543 53.1823
R1881 VSS.n1543 VSS.n1542 53.1823
R1882 VSS.n1540 VSS.n1539 53.1823
R1883 VSS.n1541 VSS.n1540 53.1823
R1884 VSS.n981 VSS.t13 52.8576
R1885 VSS.n454 VSS.n448 51.7522
R1886 VSS.t1032 VSS.t791 50.5752
R1887 VSS.t300 VSS.t582 50.5752
R1888 VSS.t830 VSS.t1098 50.5752
R1889 VSS.t641 VSS 50.5752
R1890 VSS.t1001 VSS.t255 50.5752
R1891 VSS.t389 VSS.t102 50.5752
R1892 VSS.t1013 VSS.t50 50.5752
R1893 VSS.t1023 VSS.t715 50.5752
R1894 VSS.n1532 VSS.t92 50.3004
R1895 VSS.t369 VSS.n1541 49.0584
R1896 VSS.n1542 VSS.t369 49.0584
R1897 VSS.n1889 VSS.n1530 48.7505
R1898 VSS.n1893 VSS.n1530 48.7505
R1899 VSS.n1892 VSS.n1891 48.7505
R1900 VSS.n1893 VSS.n1892 48.7505
R1901 VSS.n794 VSS.t130 48.5719
R1902 VSS.t343 VSS.n3220 47.9103
R1903 VSS.n788 VSS.t1020 47.1434
R1904 VSS.n2148 VSS.t1010 47.1434
R1905 VSS.t69 VSS 44.7453
R1906 VSS.n50 VSS 43.9579
R1907 VSS.n3079 VSS 43.9579
R1908 VSS.n3247 VSS 43.9579
R1909 VSS.n475 VSS.n474 42.1089
R1910 VSS.n488 VSS.n404 42.1089
R1911 VSS.n488 VSS.n487 42.1089
R1912 VSS.n486 VSS.n485 42.1089
R1913 VSS.n485 VSS.n484 42.1089
R1914 VSS.n483 VSS.n482 42.1089
R1915 VSS.n3342 VSS.t339 41.9598
R1916 VSS.n1568 VSS.t1034 40.0005
R1917 VSS.n1570 VSS.t962 40.0005
R1918 VSS.n981 VSS.t990 40.0005
R1919 VSS.n672 VSS.t1101 40.0005
R1920 VSS.n672 VSS.t1103 40.0005
R1921 VSS.n708 VSS.t541 40.0005
R1922 VSS.n708 VSS.t533 40.0005
R1923 VSS.n707 VSS.t535 40.0005
R1924 VSS.n707 VSS.t539 40.0005
R1925 VSS.n717 VSS.t537 40.0005
R1926 VSS.n717 VSS.t527 40.0005
R1927 VSS.n684 VSS.t741 40.0005
R1928 VSS.n684 VSS.t739 40.0005
R1929 VSS.n695 VSS.t743 40.0005
R1930 VSS.n695 VSS.t543 40.0005
R1931 VSS.n698 VSS.t549 40.0005
R1932 VSS.n698 VSS.t553 40.0005
R1933 VSS.n700 VSS.t557 40.0005
R1934 VSS.n700 VSS.t547 40.0005
R1935 VSS.n703 VSS.t551 40.0005
R1936 VSS.n703 VSS.t555 40.0005
R1937 VSS.n2533 VSS.t545 40.0005
R1938 VSS.n1485 VSS.t1089 40.0005
R1939 VSS.n1486 VSS.t1097 40.0005
R1940 VSS.n1486 VSS.t1075 40.0005
R1941 VSS.n674 VSS.t1099 40.0005
R1942 VSS.n674 VSS.t1077 40.0005
R1943 VSS.n1494 VSS.t703 40.0005
R1944 VSS.n1495 VSS.t1095 40.0005
R1945 VSS.n1495 VSS.t1085 40.0005
R1946 VSS.n1502 VSS.t1087 40.0005
R1947 VSS.n1502 VSS.t1091 40.0005
R1948 VSS.n1480 VSS.t1105 40.0005
R1949 VSS.n1480 VSS.t1083 40.0005
R1950 VSS.n1476 VSS.t613 40.0005
R1951 VSS.n1476 VSS.t1079 40.0005
R1952 VSS.n1463 VSS.t722 40.0005
R1953 VSS.n1463 VSS.t615 40.0005
R1954 VSS.n2328 VSS.t626 40.0005
R1955 VSS.n2328 VSS.t628 40.0005
R1956 VSS.n831 VSS.t384 40.0005
R1957 VSS.n822 VSS.t644 40.0005
R1958 VSS.n822 VSS.t636 40.0005
R1959 VSS.n818 VSS.t640 40.0005
R1960 VSS.n818 VSS.t630 40.0005
R1961 VSS.n817 VSS.t638 40.0005
R1962 VSS.n2356 VSS.t642 40.0005
R1963 VSS.n2356 VSS.t648 40.0005
R1964 VSS.n2360 VSS.t646 40.0005
R1965 VSS.n2360 VSS.t656 40.0005
R1966 VSS.n2367 VSS.t650 40.0005
R1967 VSS.n2367 VSS.t652 40.0005
R1968 VSS.n808 VSS.t654 40.0005
R1969 VSS.n808 VSS.t737 40.0005
R1970 VSS.n2377 VSS.t733 40.0005
R1971 VSS.n2377 VSS.t790 40.0005
R1972 VSS.n2398 VSS.t427 40.0005
R1973 VSS.n764 VSS.t115 40.0005
R1974 VSS.n759 VSS.t771 40.0005
R1975 VSS.n2046 VSS.t581 40.0005
R1976 VSS.n888 VSS.t512 40.0005
R1977 VSS.n2147 VSS.t294 40.0005
R1978 VSS.n484 VSS.n483 39.4771
R1979 VSS.n1449 VSS.t1049 38.7697
R1980 VSS.n2436 VSS.t1000 38.7697
R1981 VSS.n2045 VSS.t977 38.7697
R1982 VSS.n885 VSS.t709 38.7697
R1983 VSS.n897 VSS.t848 38.7697
R1984 VSS.n538 VSS.t128 38.5719
R1985 VSS.n538 VSS.t759 38.5719
R1986 VSS.n539 VSS.t439 38.5719
R1987 VSS.n539 VSS.t524 38.5719
R1988 VSS.n2533 VSS.t529 38.5719
R1989 VSS.n1485 VSS.t1093 38.5719
R1990 VSS.n1477 VSS.t797 38.5719
R1991 VSS.n1477 VSS.t431 38.5719
R1992 VSS.n817 VSS.t634 38.5719
R1993 VSS.n814 VSS.t571 38.5719
R1994 VSS.n814 VSS.t953 38.5719
R1995 VSS.n2405 VSS.t362 38.5719
R1996 VSS.n2405 VSS.t1022 38.5719
R1997 VSS.n789 VSS.t663 38.5719
R1998 VSS.n789 VSS.t799 38.5719
R1999 VSS.n2478 VSS.t784 38.5719
R2000 VSS.n2478 VSS.t107 38.5719
R2001 VSS.n2489 VSS.t1124 38.5719
R2002 VSS.n2489 VSS.t441 38.5719
R2003 VSS.n2042 VSS.t780 38.5719
R2004 VSS.n2042 VSS.t795 38.5719
R2005 VSS.n895 VSS.t436 38.5719
R2006 VSS.n895 VSS.t955 38.5719
R2007 VSS.n2159 VSS.t747 38.5719
R2008 VSS.n2159 VSS.t126 38.5719
R2009 VSS.n3346 VSS.t325 38.3944
R2010 VSS VSS.t1060 36.085
R2011 VSS VSS.t1037 36.085
R2012 VSS.n788 VSS.t659 35.4291
R2013 VSS.n2148 VSS.t984 35.4291
R2014 VSS.n487 VSS.n486 35.2902
R2015 VSS.n464 VSS.n431 34.659
R2016 VSS.n463 VSS.n462 34.659
R2017 VSS.n462 VSS.n433 34.659
R2018 VSS.n457 VSS.n441 34.659
R2019 VSS.n457 VSS.n456 34.659
R2020 VSS.n455 VSS.n454 34.659
R2021 VSS.n1505 VSS.n1504 34.6358
R2022 VSS.n50 VSS.n49 34.6358
R2023 VSS.n47 VSS.n2 34.6358
R2024 VSS.n3100 VSS.n3084 34.6358
R2025 VSS.n3100 VSS.n3099 34.6358
R2026 VSS.n3094 VSS.n3093 34.6358
R2027 VSS.n3128 VSS.n188 34.6358
R2028 VSS.n3128 VSS.n189 34.6358
R2029 VSS.n3122 VSS.n3121 34.6358
R2030 VSS.n3116 VSS.n3115 34.6358
R2031 VSS.n3115 VSS.n195 34.6358
R2032 VSS.n3109 VSS.n195 34.6358
R2033 VSS.n3079 VSS.n3078 34.6358
R2034 VSS.n3076 VSS.n215 34.6358
R2035 VSS.n3024 VSS.n215 34.6358
R2036 VSS.n3026 VSS.n3024 34.6358
R2037 VSS.n3029 VSS.n220 34.6358
R2038 VSS.n3033 VSS.n220 34.6358
R2039 VSS.n3053 VSS.n3042 34.6358
R2040 VSS.n3049 VSS.n3042 34.6358
R2041 VSS.n3250 VSS.n3247 34.6358
R2042 VSS.n3254 VSS.n3238 34.6358
R2043 VSS.n1617 VSS.n1616 34.6358
R2044 VSS.n1582 VSS.n1581 34.6358
R2045 VSS.n1582 VSS.n1566 34.6358
R2046 VSS.n1586 VSS.n1566 34.6358
R2047 VSS.n1575 VSS.n1571 34.6358
R2048 VSS.n1579 VSS.n1571 34.6358
R2049 VSS.n2598 VSS.n2597 34.6358
R2050 VSS.n1501 VSS.n1483 34.6358
R2051 VSS.n1509 VSS.n1478 34.6358
R2052 VSS.n2373 VSS.n810 34.6358
R2053 VSS.n2379 VSS.n2376 34.6358
R2054 VSS.n2396 VSS.n795 34.6358
R2055 VSS.n2400 VSS.n792 34.6358
R2056 VSS.n2404 VSS.n792 34.6358
R2057 VSS.n2432 VSS.n2429 34.6358
R2058 VSS.n2466 VSS.n2465 34.6358
R2059 VSS.n2471 VSS.n760 34.6358
R2060 VSS.n2514 VSS.n2485 34.6358
R2061 VSS.n2120 VSS.n2119 34.6358
R2062 VSS.n2120 VSS.n903 34.6358
R2063 VSS.n2117 VSS.n907 34.6358
R2064 VSS.n2054 VSS.n2053 34.6358
R2065 VSS.n2063 VSS.n2053 34.6358
R2066 VSS.n2064 VSS.n2063 34.6358
R2067 VSS.n2244 VSS.n2243 34.6358
R2068 VSS.n2238 VSS.n2237 34.6358
R2069 VSS.n2213 VSS.n2145 34.6358
R2070 VSS.n2209 VSS.n2145 34.6358
R2071 VSS.n2206 VSS.n2149 34.6358
R2072 VSS.n1258 VSS.n1257 34.6358
R2073 VSS.n1275 VSS.n1215 34.6358
R2074 VSS.n1335 VSS.n1334 34.6358
R2075 VSS.n2021 VSS.n920 34.6358
R2076 VSS.n1971 VSS.n1970 34.6358
R2077 VSS.n1944 VSS.n1943 34.6358
R2078 VSS.n1943 VSS.n1927 34.6358
R2079 VSS.n1722 VSS.n493 34.6358
R2080 VSS.n2780 VSS.t1236 34.2973
R2081 VSS.n835 VSS.t1194 34.2973
R2082 VSS.n1980 VSS.t1174 34.2973
R2083 VSS.n263 VSS.t1217 34.2973
R2084 VSS.n1825 VSS.t1153 34.2973
R2085 VSS.n3096 VSS.n3095 33.8829
R2086 VSS.n3090 VSS.n3089 33.8829
R2087 VSS.n3124 VSS.n3123 33.8829
R2088 VSS.n3118 VSS.n3117 33.8829
R2089 VSS.n3069 VSS.n3068 33.8829
R2090 VSS.n3062 VSS.n3061 33.8829
R2091 VSS.n3055 VSS.n3054 33.8829
R2092 VSS.n2355 VSS.n815 33.8829
R2093 VSS.n2479 VSS.n757 33.8829
R2094 VSS.t414 VSS.t1076 33.717
R2095 VSS.t789 VSS.t379 33.717
R2096 VSS.t807 VSS.t361 33.717
R2097 VSS.t313 VSS 33.717
R2098 VSS.t813 VSS.t353 33.717
R2099 VSS.t847 VSS.t337 33.717
R2100 VSS.n1377 VSS.t7 33.462
R2101 VSS.n1377 VSS.t827 33.462
R2102 VSS.n1465 VSS.t394 33.462
R2103 VSS.n1465 VSS.t508 33.462
R2104 VSS.n1227 VSS.t321 33.462
R2105 VSS.n1227 VSS.t597 33.462
R2106 VSS.n1225 VSS.t368 33.462
R2107 VSS.n1225 VSS.t624 33.462
R2108 VSS.n1222 VSS.t364 33.462
R2109 VSS.n1222 VSS.t366 33.462
R2110 VSS.n1301 VSS.t119 33.462
R2111 VSS.n1301 VSS.t1046 33.462
R2112 VSS.n1319 VSS.t975 33.462
R2113 VSS.n1319 VSS.t413 33.462
R2114 VSS.n919 VSS.t804 33.462
R2115 VSS.n919 VSS.t501 33.462
R2116 VSS.n927 VSS.t1028 33.462
R2117 VSS.n927 VSS.t73 33.462
R2118 VSS.n1912 VSS.t906 33.462
R2119 VSS.n1912 VSS.t569 33.462
R2120 VSS.n1920 VSS.t724 33.462
R2121 VSS.n1920 VSS.t1122 33.462
R2122 VSS.n1929 VSS.t701 33.462
R2123 VSS.n1929 VSS.t503 33.462
R2124 VSS.n1710 VSS.t111 33.462
R2125 VSS.n1710 VSS.t396 33.462
R2126 VSS.n3096 VSS.n3085 33.1299
R2127 VSS.n3090 VSS.n3087 33.1299
R2128 VSS.n3124 VSS.n191 33.1299
R2129 VSS.n3118 VSS.n192 33.1299
R2130 VSS.n3034 VSS.n3033 33.1299
R2131 VSS.n3069 VSS.n3036 33.1299
R2132 VSS.n3063 VSS.n3062 33.1299
R2133 VSS.n3060 VSS.n3040 33.1299
R2134 VSS.n3056 VSS.n3055 33.1299
R2135 VSS.n492 VSS.n491 32.9096
R2136 VSS.n1883 VSS.t93 32.8043
R2137 VSS.n1548 VSS.t726 32.8043
R2138 VSS VSS.t320 32.5848
R2139 VSS VSS.t363 32.5848
R2140 VSS VSS.t118 32.5848
R2141 VSS VSS.t974 32.5848
R2142 VSS VSS.t803 32.5848
R2143 VSS VSS.t1027 32.5848
R2144 VSS VSS.t905 32.5848
R2145 VSS VSS.t723 32.5848
R2146 VSS VSS.t700 32.5848
R2147 VSS.n794 VSS.t829 32.5719
R2148 VSS.n454 VSS.n453 32.5005
R2149 VSS.n453 VSS.n438 32.5005
R2150 VSS.n451 VSS.n426 32.5005
R2151 VSS.n445 VSS.n411 32.5005
R2152 VSS.n424 VSS.n411 32.5005
R2153 VSS.n482 VSS.n481 32.5005
R2154 VSS.n481 VSS.n401 32.5005
R2155 VSS.n458 VSS.n457 32.5005
R2156 VSS.n460 VSS.n458 32.5005
R2157 VSS.n443 VSS.n427 32.5005
R2158 VSS.n468 VSS.n427 32.5005
R2159 VSS.n416 VSS.n415 32.5005
R2160 VSS.n420 VSS.n416 32.5005
R2161 VSS.n485 VSS.n400 32.5005
R2162 VSS.n490 VSS.n400 32.5005
R2163 VSS.n462 VSS.n461 32.5005
R2164 VSS.n461 VSS.n460 32.5005
R2165 VSS.n435 VSS.n425 32.5005
R2166 VSS.n468 VSS.n425 32.5005
R2167 VSS.n419 VSS.n418 32.5005
R2168 VSS.n420 VSS.n419 32.5005
R2169 VSS.n489 VSS.n488 32.5005
R2170 VSS.n490 VSS.n489 32.5005
R2171 VSS.n459 VSS.n431 32.5005
R2172 VSS.n460 VSS.n459 32.5005
R2173 VSS.n467 VSS.n466 32.5005
R2174 VSS.n468 VSS.n467 32.5005
R2175 VSS.n477 VSS.n470 32.5005
R2176 VSS.n470 VSS.n469 32.5005
R2177 VSS.n474 VSS.n423 32.5005
R2178 VSS.n423 VSS.n422 32.5005
R2179 VSS.n441 VSS.n433 32.4928
R2180 VSS.n3064 VSS.n3037 32.377
R2181 VSS.n1589 VSS.n1588 32.377
R2182 VSS.n2275 VSS.n882 32.377
R2183 VSS.n2239 VSS.n2238 32.377
R2184 VSS.n2143 VSS.n2142 32.377
R2185 VSS.n2350 VSS.n2349 32.377
R2186 VSS.n2243 VSS.n898 31.624
R2187 VSS.n1588 VSS.n1587 31.2476
R2188 VSS.n2449 VSS.n2448 31.2476
R2189 VSS.n2275 VSS.n2274 31.2476
R2190 VSS.n2216 VSS.n2143 31.2476
R2191 VSS.n456 VSS.n455 30.9174
R2192 VSS.n478 VSS.n473 30.8711
R2193 VSS.n392 VSS.n391 30.8711
R2194 VSS.n3186 VSS.n3185 30.8711
R2195 VSS.n3209 VSS.n3200 30.8711
R2196 VSS.n3163 VSS.n180 30.8711
R2197 VSS.n3155 VSS.n3141 30.8711
R2198 VSS.n3137 VSS.n183 30.8711
R2199 VSS.n3326 VSS.n3325 30.8711
R2200 VSS.n3216 VSS.n3215 30.8711
R2201 VSS.n1580 VSS.n1579 30.8711
R2202 VSS.n2400 VSS.n2399 30.8711
R2203 VSS.n2075 VSS.n2047 30.8711
R2204 VSS.n2267 VSS.n2266 30.8711
R2205 VSS.n475 VSS.n404 30.7444
R2206 VSS.n2329 VSS.n821 30.4946
R2207 VSS.n2429 VSS.n783 30.4946
R2208 VSS.n2266 VSS.n890 30.4946
R2209 VSS.n1877 VSS.t370 30.3424
R2210 VSS.n1488 VSS.n673 30.1181
R2211 VSS.n2345 VSS.n819 30.1181
R2212 VSS.n2391 VSS.n797 30.1181
R2213 VSS.n2054 VSS.n902 30.1181
R2214 VSS.n3341 VSS.n3340 29.8168
R2215 VSS.t1005 VSS.t719 29.8079
R2216 VSS.t719 VSS.t94 29.8079
R2217 VSS.t1007 VSS.t727 29.8079
R2218 VSS.t1003 VSS.t1007 29.8079
R2219 VSS.t92 VSS.t1003 29.8079
R2220 VSS.n1492 VSS.n1487 29.7417
R2221 VSS.n2444 VSS.n2443 29.3652
R2222 VSS.n2586 VSS.n676 28.9887
R2223 VSS.n464 VSS.n463 28.259
R2224 VSS.n1512 VSS.n1511 27.8593
R2225 VSS.n2376 VSS.n2375 27.8593
R2226 VSS.n1575 VSS.n1574 27.4829
R2227 VSS.n2406 VSS.n2404 27.4829
R2228 VSS.n2438 VSS.n2437 27.4829
R2229 VSS.n2470 VSS.n2469 27.4829
R2230 VSS.n2475 VSS.n760 27.4829
R2231 VSS.n2077 VSS.n2076 27.4829
R2232 VSS.n2077 VSS.n2043 27.4829
R2233 VSS.n2272 VSS.n886 27.4829
R2234 VSS.n2250 VSS.n2249 27.4829
R2235 VSS.n1512 VSS.n1464 27.1064
R2236 VSS.n3385 VSS.n3384 26.9246
R2237 VSS.n3298 VSS.n95 26.9246
R2238 VSS.n2413 VSS.n2412 26.7299
R2239 VSS.n1837 VSS.n1836 26.6009
R2240 VSS.n2113 VSS.n907 26.314
R2241 VSS.n1883 VSS.n1882 26.1653
R2242 VSS.n1885 VSS.n1884 26.1653
R2243 VSS.n1548 VSS.n1547 26.1653
R2244 VSS.n469 VSS.n468 25.9813
R2245 VSS.n983 VSS.t117 25.9346
R2246 VSS.n2036 VSS.t109 25.9346
R2247 VSS.n2096 VSS.t356 25.9346
R2248 VSS.n3174 VSS.t890 25.8199
R2249 VSS.n2369 VSS.n2366 25.7355
R2250 VSS.n2227 VSS.n2125 25.7355
R2251 VSS.n2202 VSS.n2149 25.7355
R2252 VSS.n1253 VSS.n1252 25.7355
R2253 VSS.n1938 VSS.n1937 25.7355
R2254 VSS.n3403 VSS.n2 25.6926
R2255 VSS.n3255 VSS.n3254 25.6926
R2256 VSS.n1263 VSS.n1262 25.6926
R2257 VSS.n1270 VSS.n1221 25.6926
R2258 VSS.n1291 VSS.n1215 25.6926
R2259 VSS.n1334 VSS.n1321 25.6926
R2260 VSS.n2013 VSS.n920 25.6926
R2261 VSS.n2007 VSS.n2006 25.6926
R2262 VSS.n1970 VSS.n1914 25.6926
R2263 VSS.n1723 VSS.n1722 25.6926
R2264 VSS.n1616 VSS.n1590 25.6005
R2265 VSS.n2351 VSS.n2350 25.6005
R2266 VSS.n15 VSS.t792 25.4291
R2267 VSS.n21 VSS.t583 25.4291
R2268 VSS.n3039 VSS.t1024 25.4291
R2269 VSS.n218 VSS.t1014 25.4291
R2270 VSS.n3267 VSS.t1002 25.4291
R2271 VSS.n107 VSS.t390 25.4291
R2272 VSS.n679 VSS.t392 25.4291
R2273 VSS.n1374 VSS.t5 25.4291
R2274 VSS.t140 VSS.t399 25.2879
R2275 VSS.t1084 VSS.t702 25.2879
R2276 VSS.t518 VSS.t749 25.2879
R2277 VSS.n3368 VSS.n3367 25.224
R2278 VSS.n3367 VSS.n60 25.224
R2279 VSS.n3363 VSS.n3362 25.224
R2280 VSS.n3362 VSS.n3361 25.224
R2281 VSS.n3359 VSS.n3358 25.224
R2282 VSS.n3358 VSS.n3350 25.224
R2283 VSS.n3354 VSS.n3353 25.224
R2284 VSS.n3353 VSS.n39 25.224
R2285 VSS.n3394 VSS.n3393 25.224
R2286 VSS.n3393 VSS.n3392 25.224
R2287 VSS.n3390 VSS.n22 25.224
R2288 VSS.n3315 VSS.n3314 25.224
R2289 VSS.n3314 VSS.n83 25.224
R2290 VSS.n3310 VSS.n3309 25.224
R2291 VSS.n3309 VSS.n3308 25.224
R2292 VSS.n3306 VSS.n3305 25.224
R2293 VSS.n3305 VSS.n89 25.224
R2294 VSS.n3301 VSS.n3300 25.224
R2295 VSS.n3300 VSS.n3299 25.224
R2296 VSS.n3274 VSS.n3273 25.224
R2297 VSS.n3275 VSS.n3274 25.224
R2298 VSS.n3292 VSS.n3279 25.224
R2299 VSS.n127 VSS.n125 25.224
R2300 VSS.n131 VSS.n125 25.224
R2301 VSS.n132 VSS.n124 25.224
R2302 VSS.n136 VSS.n124 25.224
R2303 VSS.n137 VSS.n123 25.224
R2304 VSS.n141 VSS.n123 25.224
R2305 VSS.n142 VSS.n122 25.224
R2306 VSS.n146 VSS.n122 25.224
R2307 VSS.n147 VSS.n121 25.224
R2308 VSS.n151 VSS.n121 25.224
R2309 VSS.n152 VSS.n120 25.224
R2310 VSS.n156 VSS.n120 25.224
R2311 VSS.n157 VSS.n119 25.224
R2312 VSS.n161 VSS.n119 25.224
R2313 VSS.n162 VSS.n118 25.224
R2314 VSS.n166 VSS.n118 25.224
R2315 VSS.n167 VSS.n117 25.224
R2316 VSS.n171 VSS.n117 25.224
R2317 VSS.n2344 VSS.n821 25.224
R2318 VSS.n2345 VSS.n2344 25.224
R2319 VSS.n1976 VSS.n1975 24.9894
R2320 VSS.n1832 VSS.n1831 24.9894
R2321 VSS.n3083 VSS.n3082 24.9767
R2322 VSS.n3108 VSS.n3107 24.9767
R2323 VSS.n3047 VSS.n3044 24.9767
R2324 VSS.n2846 VSS.n2845 24.968
R2325 VSS.n3339 VSS.t495 24.9236
R2326 VSS.n3339 VSS.t493 24.9236
R2327 VSS.n1629 VSS.t696 24.9236
R2328 VSS.n1629 VSS.t699 24.9236
R2329 VSS.n1564 VSS.t376 24.9236
R2330 VSS.n1564 VSS.t377 24.9236
R2331 VSS.n1563 VSS.t834 24.9236
R2332 VSS.n1563 VSS.t3 24.9236
R2333 VSS.n675 VSS.t831 24.9236
R2334 VSS.n675 VSS.t415 24.9236
R2335 VSS.n838 VSS.t317 24.9236
R2336 VSS.n838 VSS.t575 24.9236
R2337 VSS.n809 VSS.t382 24.9236
R2338 VSS.n809 VSS.t1073 24.9236
R2339 VSS.n2430 VSS.t1109 24.9236
R2340 VSS.n2430 VSS.t124 24.9236
R2341 VSS.n2436 VSS.t76 24.9236
R2342 VSS.n775 VSS.t1018 24.9236
R2343 VSS.n775 VSS.t705 24.9236
R2344 VSS.n774 VSS.t137 24.9236
R2345 VSS.n774 VSS.t788 24.9236
R2346 VSS.n762 VSS.t388 24.9236
R2347 VSS.n762 VSS.t517 24.9236
R2348 VSS.n880 VSS.t620 24.9236
R2349 VSS.n880 VSS.t622 24.9236
R2350 VSS.n881 VSS.t1118 24.9236
R2351 VSS.n881 VSS.t607 24.9236
R2352 VSS.n885 VSS.t825 24.9236
R2353 VSS.n900 VSS.t579 24.9236
R2354 VSS.n900 VSS.t338 24.9236
R2355 VSS.n2132 VSS.t307 24.9236
R2356 VSS.n2132 VSS.t559 24.9236
R2357 VSS.n2144 VSS.t1030 24.9236
R2358 VSS.n2144 VSS.t994 24.9236
R2359 VSS VSS.t494 24.7946
R2360 VSS.n2327 VSS.n2326 24.4711
R2361 VSS.n2477 VSS.n2476 24.4711
R2362 VSS.n2432 VSS.n2431 24.4711
R2363 VSS.n2484 VSS.n757 24.4711
R2364 VSS.n2485 VSS.n2484 24.4711
R2365 VSS.n2214 VSS.n2213 24.4711
R2366 VSS.t1060 VSS.t1057 24.2493
R2367 VSS.t1037 VSS.t1040 24.2493
R2368 VSS.t325 VSS.t328 24.2493
R2369 VSS.n3398 VSS.n16 24.0946
R2370 VSS.n3269 VSS.n110 24.0946
R2371 VSS.n281 VSS.t218 23.7273
R2372 VSS.n2442 VSS.n780 23.7181
R2373 VSS.n1397 VSS.n1382 23.7181
R2374 VSS.n1408 VSS.n1382 23.7181
R2375 VSS.n2571 VSS.n682 23.7181
R2376 VSS.n2571 VSS.n2570 23.7181
R2377 VSS.n2392 VSS.n795 23.7181
R2378 VSS.n2438 VSS.n780 23.7181
R2379 VSS.n2464 VSS.n766 23.7181
R2380 VSS.n2465 VSS.n2464 23.7181
R2381 VSS.n2234 VSS.n903 23.7181
R2382 VSS.n2273 VSS.n2272 23.7181
R2383 VSS.n1300 VSS.n1213 23.7181
R2384 VSS.n1357 VSS.n1212 23.7181
R2385 VSS.n1340 VSS.n1339 23.7181
R2386 VSS.n1327 VSS.n918 23.7181
R2387 VSS.n2002 VSS.n2001 23.7181
R2388 VSS.n1963 VSS.n1962 23.7181
R2389 VSS.n2924 VSS.n493 23.7181
R2390 VSS.t110 VSS 23.6345
R2391 VSS.n2512 VSS.n2511 23.4338
R2392 VSS.n1481 VSS.n1478 23.3417
R2393 VSS.n2368 VSS.n810 23.3417
R2394 VSS.n450 VSS.n448 23.2076
R2395 VSS.n3115 VSS.n3114 23.1729
R2396 VSS.n2847 VSS.n537 22.9652
R2397 VSS.n1574 VSS.n537 22.9652
R2398 VSS.n2407 VSS.n2406 22.9652
R2399 VSS.n2407 VSS.n790 22.9652
R2400 VSS.n2448 VSS.n776 22.9652
R2401 VSS.n2476 VSS.n2475 22.9652
R2402 VSS.n2081 VSS.n2043 22.9652
R2403 VSS.n2082 VSS.n2081 22.9652
R2404 VSS.n2279 VSS.n2278 22.9652
R2405 VSS.n2249 VSS.n2248 22.9652
R2406 VSS.n2248 VSS.n896 22.9652
R2407 VSS.n2208 VSS.n2207 22.9652
R2408 VSS.n3221 VSS.n3174 22.9387
R2409 VSS.n3332 VSS.t835 22.8805
R2410 VSS.n2392 VSS.n2391 22.5887
R2411 VSS.n24 VSS.t311 22.3257
R2412 VSS.n44 VSS.t850 22.3257
R2413 VSS.n3045 VSS.t753 22.3257
R2414 VSS.n214 VSS.t84 22.3257
R2415 VSS.n3248 VSS.t340 22.3257
R2416 VSS.n3282 VSS.t707 22.3257
R2417 VSS.n905 VSS.t497 22.3257
R2418 VSS.n906 VSS.t1047 22.3257
R2419 VSS.n2133 VSS.t992 22.3257
R2420 VSS.n1587 VSS.n1586 22.2123
R2421 VSS.n2449 VSS.n766 22.2123
R2422 VSS.n2471 VSS.n2470 22.2123
R2423 VSS.n2216 VSS.n2215 22.2123
R2424 VSS.n1253 VSS.n1228 22.2123
R2425 VSS.n1257 VSS.n1228 22.2123
R2426 VSS.n1258 VSS.n1226 22.2123
R2427 VSS.n1262 VSS.n1226 22.2123
R2428 VSS.n1274 VSS.n1221 22.2123
R2429 VSS.n1275 VSS.n1274 22.2123
R2430 VSS.n1302 VSS.n1300 22.2123
R2431 VSS.n1302 VSS.n1212 22.2123
R2432 VSS.n1339 VSS.n1320 22.2123
R2433 VSS.n1335 VSS.n1320 22.2123
R2434 VSS.n2022 VSS.n918 22.2123
R2435 VSS.n2022 VSS.n2021 22.2123
R2436 VSS.n2006 VSS.n928 22.2123
R2437 VSS.n2002 VSS.n928 22.2123
R2438 VSS.n1975 VSS.n1913 22.2123
R2439 VSS.n1971 VSS.n1913 22.2123
R2440 VSS.n1962 VSS.n1921 22.2123
R2441 VSS.n1944 VSS.n1921 22.2123
R2442 VSS.n1939 VSS.n1927 22.2123
R2443 VSS.n1939 VSS.n1938 22.2123
R2444 VSS.n1836 VSS.n1711 22.2123
R2445 VSS.n1832 VSS.n1711 22.2123
R2446 VSS.n446 VSS.n412 21.6752
R2447 VSS.n3347 VSS 21.6512
R2448 VSS.n3399 VSS.n3398 21.4593
R2449 VSS.n3391 VSS.n3390 21.4593
R2450 VSS.n3269 VSS.n3268 21.4593
R2451 VSS.n3279 VSS.n108 21.4593
R2452 VSS.n2847 VSS.n2846 21.4593
R2453 VSS.n2411 VSS.n790 21.4593
R2454 VSS.n2444 VSS.n776 21.4593
R2455 VSS.n2076 VSS.n2075 21.4593
R2456 VSS.n2244 VSS.n896 21.4593
R2457 VSS.n2322 VSS.n832 20.8482
R2458 VSS.n1488 VSS.n1487 20.7064
R2459 VSS.n2597 VSS.n676 20.7064
R2460 VSS.n3363 VSS.n60 20.3299
R2461 VSS.n3354 VSS.n3350 20.3299
R2462 VSS.n3310 VSS.n83 20.3299
R2463 VSS.n3301 VSS.n89 20.3299
R2464 VSS.t1057 VSS 19.3418
R2465 VSS.t1040 VSS 19.3418
R2466 VSS.t328 VSS 19.3418
R2467 VSS.n3369 VSS.n3368 19.2926
R2468 VSS.n3316 VSS.n3315 19.2926
R2469 VSS.n1894 VSS.t1005 19.2511
R2470 VSS.t675 VSS 19.0729
R2471 VSS.n3077 VSS.n3076 18.824
R2472 VSS.n132 VSS.n131 18.824
R2473 VSS.n137 VSS.n136 18.824
R2474 VSS.n142 VSS.n141 18.824
R2475 VSS.n147 VSS.n146 18.824
R2476 VSS.n152 VSS.n151 18.824
R2477 VSS.n157 VSS.n156 18.824
R2478 VSS.n162 VSS.n161 18.824
R2479 VSS.n167 VSS.n166 18.824
R2480 VSS.n1035 VSS.n1034 18.2791
R2481 VSS.n1437 VSS.n1436 18.2791
R2482 VSS.n1777 VSS.n1776 18.2791
R2483 VSS.n33 VSS.n22 17.7867
R2484 VSS.n3292 VSS.n3291 17.7867
R2485 VSS.n1754 VSS.n1735 17.7007
R2486 VSS.n1859 VSS.n1858 17.4137
R2487 VSS.n3360 VSS.n3359 17.3181
R2488 VSS.n3084 VSS.n3083 17.3181
R2489 VSS.n3109 VSS.n3108 17.3181
R2490 VSS.n3029 VSS.n3028 17.3181
R2491 VSS.n3307 VSS.n3306 17.3181
R2492 VSS.n2585 VSS.n2584 17.3181
R2493 VSS.n2872 VSS.n2871 17.195
R2494 VSS.n1061 VSS.n1060 16.9936
R2495 VSS.n2959 VSS.n264 16.9545
R2496 VSS.n2437 VSS.n781 16.9417
R2497 VSS.n2268 VSS.n886 16.9417
R2498 VSS.t242 VSS.t298 16.8587
R2499 VSS.t6 VSS.t143 16.8587
R2500 VSS.t249 VSS.t574 16.8587
R2501 VSS.t108 VSS.t879 16.8587
R2502 VSS.t104 VSS.t938 16.8587
R2503 VSS.t870 VSS.t677 16.8587
R2504 VSS.n2979 VSS.n255 16.8353
R2505 VSS.n2974 VSS.n256 16.7924
R2506 VSS.n1659 VSS.n1632 16.763
R2507 VSS.n1542 VSS.n67 16.4566
R2508 VSS.n1493 VSS.n1492 16.1887
R2509 VSS.n2586 VSS.n2585 16.1887
R2510 VSS.n2326 VSS.n832 16.1887
R2511 VSS.n3361 VSS.n3360 15.8123
R2512 VSS.n3384 VSS.n39 15.8123
R2513 VSS.n3078 VSS.n3077 15.8123
R2514 VSS.n3049 VSS.n3048 15.8123
R2515 VSS.n3308 VSS.n3307 15.8123
R2516 VSS.n3299 VSS.n3298 15.8123
R2517 VSS.n127 VSS.n69 15.8123
R2518 VSS.n3231 VSS.n171 15.8123
R2519 VSS.n1523 VSS.n1522 15.3963
R2520 VSS.n2924 VSS.n2923 15.3963
R2521 VSS.n2928 VSS.n2927 15.3963
R2522 VSS.n3028 VSS.n3027 15.0593
R2523 VSS.t94 VSS.n1893 14.9042
R2524 VSS.n1893 VSS.t727 14.9042
R2525 VSS.n2234 VSS.n2233 14.8179
R2526 VSS.n2927 VSS.n278 14.8179
R2527 VSS.n3384 VSS.n3383 14.775
R2528 VSS.n3400 VSS.n4 14.775
R2529 VSS.n3298 VSS.n92 14.775
R2530 VSS.n3263 VSS.n113 14.775
R2531 VSS.n1599 VSS.n1598 14.775
R2532 VSS.n2575 VSS.n682 14.775
R2533 VSS.n2302 VSS.n2301 14.775
R2534 VSS.n2288 VSS.n2287 14.775
R2535 VSS.n1357 VSS.n1356 14.775
R2536 VSS.n2001 VSS.n2000 14.775
R2537 VSS.n1657 VSS.n1656 14.2735
R2538 VSS.n2196 VSS.n2151 14.065
R2539 VSS.n1678 VSS.n1677 14.0503
R2540 VSS.n1010 VSS.n1009 14.0503
R2541 VSS.n736 VSS.n733 14.0503
R2542 VSS.n2413 VSS.n783 13.9299
R2543 VSS.n2250 VSS.n890 13.9299
R2544 VSS.n2178 VSS.n2177 13.8859
R2545 VSS.n3394 VSS.n16 13.5534
R2546 VSS.n3273 VSS.n110 13.5534
R2547 VSS.n3335 VSS.n69 12.8005
R2548 VSS.n3335 VSS.n68 12.8005
R2549 VSS.n3341 VSS.n68 12.8005
R2550 VSS.n1108 VSS.n1085 12.8005
R2551 VSS.n2708 VSS.n593 12.8005
R2552 VSS.n2682 VSS.n2681 12.8005
R2553 VSS.n2498 VSS.n2497 12.8005
R2554 VSS.n2280 VSS.n2279 12.5161
R2555 VSS.n3009 VSS.n3008 12.424
R2556 VSS.n3004 VSS.n2994 12.424
R2557 VSS.n1061 VSS.n931 12.1384
R2558 VSS.n2357 VSS.n2355 11.9309
R2559 VSS.n3082 VSS.n3081 11.3835
R2560 VSS.n2369 VSS.n2368 11.2946
R2561 VSS.n2274 VSS.n2273 11.2946
R2562 VSS.n53 VSS.n52 11.2844
R2563 VSS.n3246 VSS.n3245 11.2844
R2564 VSS.n306 VSS.n299 11.0382
R2565 VSS.n302 VSS.n299 11.0382
R2566 VSS.n300 VSS.n298 11.0382
R2567 VSS.n302 VSS.n298 11.0382
R2568 VSS.n314 VSS.n294 11.0382
R2569 VSS.n297 VSS.n294 11.0382
R2570 VSS.n296 VSS.n293 11.0382
R2571 VSS.n297 VSS.n293 11.0382
R2572 VSS.n291 VSS.n289 11.0382
R2573 VSS.n322 VSS.n291 11.0382
R2574 VSS.n292 VSS.n290 11.0382
R2575 VSS.n322 VSS.n292 11.0382
R2576 VSS.n365 VSS.n343 11.0382
R2577 VSS.n361 VSS.n343 11.0382
R2578 VSS.n344 VSS.n342 11.0382
R2579 VSS.n361 VSS.n342 11.0382
R2580 VSS.n337 VSS.n285 11.0382
R2581 VSS.n333 VSS.n285 11.0382
R2582 VSS.n286 VSS.n284 11.0382
R2583 VSS.n333 VSS.n284 11.0382
R2584 VSS.n3184 VSS.n3177 11.0382
R2585 VSS.n3177 VSS.n3176 11.0382
R2586 VSS.n3181 VSS.n3175 11.0382
R2587 VSS.n3176 VSS.n3175 11.0382
R2588 VSS.n3208 VSS.n3207 11.0382
R2589 VSS.n3207 VSS.n3206 11.0382
R2590 VSS.n3205 VSS.n3204 11.0382
R2591 VSS.n3206 VSS.n3205 11.0382
R2592 VSS.n3147 VSS.n3146 11.0382
R2593 VSS.n3152 VSS.n3147 11.0382
R2594 VSS.n3143 VSS.n3142 11.0382
R2595 VSS.n3152 VSS.n3143 11.0382
R2596 VSS.n3136 VSS.n3135 11.0382
R2597 VSS.n3135 VSS.n3134 11.0382
R2598 VSS.n3133 VSS.n3132 11.0382
R2599 VSS.n3134 VSS.n3133 11.0382
R2600 VSS.n3164 VSS.n178 11.0382
R2601 VSS.n3148 VSS.n178 11.0382
R2602 VSS.n179 VSS.n177 11.0382
R2603 VSS.n3148 VSS.n177 11.0382
R2604 VSS.n203 VSS.n196 11.0382
R2605 VSS.n207 VSS.n196 11.0382
R2606 VSS.n206 VSS.n205 11.0382
R2607 VSS.n207 VSS.n206 11.0382
R2608 VSS.n3198 VSS.n3193 11.0382
R2609 VSS.n3193 VSS.n3192 11.0382
R2610 VSS.n3195 VSS.n3191 11.0382
R2611 VSS.n3192 VSS.n3191 11.0382
R2612 VSS.n3327 VSS.n73 11.0382
R2613 VSS.n3331 VSS.n73 11.0382
R2614 VSS.n3330 VSS.n3329 11.0382
R2615 VSS.n3331 VSS.n3330 11.0382
R2616 VSS.n356 VSS.n348 11.0382
R2617 VSS.n348 VSS.n347 11.0382
R2618 VSS.n353 VSS.n346 11.0382
R2619 VSS.n347 VSS.n346 11.0382
R2620 VSS.n381 VSS.n372 11.0382
R2621 VSS.n377 VSS.n372 11.0382
R2622 VSS.n373 VSS.n371 11.0382
R2623 VSS.n377 VSS.n371 11.0382
R2624 VSS.n393 VSS.n280 11.0382
R2625 VSS.n397 VSS.n280 11.0382
R2626 VSS.n396 VSS.n395 11.0382
R2627 VSS.n397 VSS.n396 11.0382
R2628 VSS.n3015 VSS.n3014 11.0382
R2629 VSS.n3012 VSS.n3011 11.0382
R2630 VSS.n3003 VSS.n3002 11.0382
R2631 VSS.n3002 VSS.n3001 11.0382
R2632 VSS.n2998 VSS.n2997 11.0382
R2633 VSS.n2998 VSS.n223 11.0382
R2634 VSS.n2761 VSS.n561 10.9091
R2635 VSS.n2569 VSS.n2568 10.8805
R2636 VSS.n471 VSS.t87 10.6509
R2637 VSS.n3005 VSS.n3004 10.6195
R2638 VSS.n3008 VSS.n3007 10.6189
R2639 VSS.n1409 VSS.n1408 10.5983
R2640 VSS.n1581 VSS.n1580 10.5417
R2641 VSS.n1497 VSS.n1493 10.5417
R2642 VSS.n2064 VSS.n2047 10.5417
R2643 VSS.n2268 VSS.n2267 10.5417
R2644 VSS.n2209 VSS.n2208 10.5417
R2645 VSS.n392 VSS.n390 10.4476
R2646 VSS.n3185 VSS.n3180 10.4476
R2647 VSS.n3210 VSS.n3209 10.4476
R2648 VSS.n3163 VSS.n3162 10.4476
R2649 VSS.n3157 VSS.n3141 10.4476
R2650 VSS.n3138 VSS.n3137 10.4476
R2651 VSS.n3326 VSS.n3324 10.4476
R2652 VSS.n3215 VSS.n3214 10.4476
R2653 VSS.n3392 VSS.n3391 10.1652
R2654 VSS.n3275 VSS.n108 10.1652
R2655 VSS.n1522 VSS.n1521 10.1652
R2656 VSS.n1521 VSS.n1464 10.1652
R2657 VSS.n2330 VSS.n2327 10.1652
R2658 VSS.n2431 VSS.n781 10.1652
R2659 VSS.n2480 VSS.n2477 10.1652
R2660 VSS.n2215 VSS.n2214 10.1652
R2661 VSS.n1606 VSS.n1590 9.88085
R2662 VSS.n1236 VSS.n1235 9.7205
R2663 VSS.n247 VSS.n246 9.7205
R2664 VSS.n1932 VSS.n1931 9.71789
R2665 VSS.n1853 VSS.n1852 9.71789
R2666 VSS.n53 VSS.n42 9.70901
R2667 VSS.n3377 VSS.n3376 9.70901
R2668 VSS.n27 VSS.n26 9.70901
R2669 VSS.n3245 VSS.n3244 9.70901
R2670 VSS.n100 VSS.n99 9.70901
R2671 VSS.n3284 VSS.n3283 9.70901
R2672 VSS.n48 VSS.n47 9.41227
R2673 VSS.n3249 VSS.n3238 9.41227
R2674 VSS.n2399 VSS.n2397 9.41227
R2675 VSS.n2118 VSS.n2117 9.41227
R2676 VSS.n2141 VSS.n2134 9.41227
R2677 VSS.n1090 VSS.n1085 9.3031
R2678 VSS.n2690 VSS.n593 9.3031
R2679 VSS.n2682 VSS.n601 9.3031
R2680 VSS.n1397 VSS.n1396 9.3031
R2681 VSS.n2301 VSS.n2299 9.3031
R2682 VSS.n2288 VSS.n862 9.3031
R2683 VSS.n3386 VSS.n3385 9.3005
R2684 VSS.n3379 VSS.n3378 9.3005
R2685 VSS.n3381 VSS.n3380 9.3005
R2686 VSS.n3383 VSS.n3382 9.3005
R2687 VSS.n3384 VSS.n36 9.3005
R2688 VSS.n55 VSS.n54 9.3005
R2689 VSS.n56 VSS.n41 9.3005
R2690 VSS.n3370 VSS.n3369 9.3005
R2691 VSS.n3368 VSS.n59 9.3005
R2692 VSS.n3367 VSS.n3366 9.3005
R2693 VSS.n3365 VSS.n60 9.3005
R2694 VSS.n3364 VSS.n3363 9.3005
R2695 VSS.n3362 VSS.n61 9.3005
R2696 VSS.n3361 VSS.n62 9.3005
R2697 VSS.n3360 VSS.n3348 9.3005
R2698 VSS.n3359 VSS.n3349 9.3005
R2699 VSS.n3358 VSS.n3357 9.3005
R2700 VSS.n3356 VSS.n3350 9.3005
R2701 VSS.n3355 VSS.n3354 9.3005
R2702 VSS.n3353 VSS.n3352 9.3005
R2703 VSS.n3351 VSS.n39 9.3005
R2704 VSS.n29 VSS.n28 9.3005
R2705 VSS.n31 VSS.n23 9.3005
R2706 VSS.n34 VSS.n33 9.3005
R2707 VSS.n3400 VSS.n13 9.3005
R2708 VSS.n3399 VSS.n14 9.3005
R2709 VSS.n3398 VSS.n3397 9.3005
R2710 VSS.n3396 VSS.n16 9.3005
R2711 VSS.n3395 VSS.n3394 9.3005
R2712 VSS.n3393 VSS.n18 9.3005
R2713 VSS.n3392 VSS.n19 9.3005
R2714 VSS.n3391 VSS.n20 9.3005
R2715 VSS.n3390 VSS.n3389 9.3005
R2716 VSS.n35 VSS.n22 9.3005
R2717 VSS.n51 VSS.n50 9.3005
R2718 VSS.n49 VSS.n43 9.3005
R2719 VSS.n47 VSS.n46 9.3005
R2720 VSS.n45 VSS.n2 9.3005
R2721 VSS.n3404 VSS.n3403 9.3005
R2722 VSS.n6 VSS.n5 9.3005
R2723 VSS.n11 VSS.n10 9.3005
R2724 VSS.n12 VSS.n4 9.3005
R2725 VSS.n3050 VSS.n3049 9.3005
R2726 VSS.n3051 VSS.n3042 9.3005
R2727 VSS.n3080 VSS.n3079 9.3005
R2728 VSS.n3078 VSS.n213 9.3005
R2729 VSS.n3076 VSS.n3075 9.3005
R2730 VSS.n3074 VSS.n215 9.3005
R2731 VSS.n3024 VSS.n216 9.3005
R2732 VSS.n3026 VSS.n3025 9.3005
R2733 VSS.n3030 VSS.n3029 9.3005
R2734 VSS.n3031 VSS.n220 9.3005
R2735 VSS.n3033 VSS.n3032 9.3005
R2736 VSS.n3035 VSS.n217 9.3005
R2737 VSS.n3070 VSS.n3069 9.3005
R2738 VSS.n3067 VSS.n3066 9.3005
R2739 VSS.n3065 VSS.n3064 9.3005
R2740 VSS.n3062 VSS.n3038 9.3005
R2741 VSS.n3060 VSS.n3059 9.3005
R2742 VSS.n3058 VSS.n3057 9.3005
R2743 VSS.n3055 VSS.n3041 9.3005
R2744 VSS.n3053 VSS.n3052 9.3005
R2745 VSS.n3114 VSS.n3113 9.3005
R2746 VSS.n3110 VSS.n3109 9.3005
R2747 VSS.n3111 VSS.n195 9.3005
R2748 VSS.n3115 VSS.n194 9.3005
R2749 VSS.n3084 VSS.n211 9.3005
R2750 VSS.n3101 VSS.n3100 9.3005
R2751 VSS.n3099 VSS.n3098 9.3005
R2752 VSS.n3097 VSS.n3096 9.3005
R2753 VSS.n3094 VSS.n3086 9.3005
R2754 VSS.n3093 VSS.n3092 9.3005
R2755 VSS.n3091 VSS.n3090 9.3005
R2756 VSS.n3088 VSS.n188 9.3005
R2757 VSS.n3128 VSS.n3127 9.3005
R2758 VSS.n3126 VSS.n189 9.3005
R2759 VSS.n3125 VSS.n3124 9.3005
R2760 VSS.n3122 VSS.n190 9.3005
R2761 VSS.n3121 VSS.n3120 9.3005
R2762 VSS.n3119 VSS.n3118 9.3005
R2763 VSS.n3116 VSS.n193 9.3005
R2764 VSS.n3295 VSS.n95 9.3005
R2765 VSS.n102 VSS.n101 9.3005
R2766 VSS.n104 VSS.n103 9.3005
R2767 VSS.n105 VSS.n92 9.3005
R2768 VSS.n3298 VSS.n3297 9.3005
R2769 VSS.n3243 VSS.n3240 9.3005
R2770 VSS.n3242 VSS.n80 9.3005
R2771 VSS.n3317 VSS.n3316 9.3005
R2772 VSS.n3315 VSS.n82 9.3005
R2773 VSS.n3314 VSS.n3313 9.3005
R2774 VSS.n3312 VSS.n83 9.3005
R2775 VSS.n3311 VSS.n3310 9.3005
R2776 VSS.n3309 VSS.n84 9.3005
R2777 VSS.n3308 VSS.n85 9.3005
R2778 VSS.n3307 VSS.n87 9.3005
R2779 VSS.n3306 VSS.n88 9.3005
R2780 VSS.n3305 VSS.n3304 9.3005
R2781 VSS.n3303 VSS.n89 9.3005
R2782 VSS.n3302 VSS.n3301 9.3005
R2783 VSS.n3300 VSS.n90 9.3005
R2784 VSS.n3299 VSS.n91 9.3005
R2785 VSS.n3286 VSS.n3281 9.3005
R2786 VSS.n3289 VSS.n3288 9.3005
R2787 VSS.n3291 VSS.n3290 9.3005
R2788 VSS.n3247 VSS.n3239 9.3005
R2789 VSS.n3251 VSS.n3250 9.3005
R2790 VSS.n3252 VSS.n3238 9.3005
R2791 VSS.n3254 VSS.n3253 9.3005
R2792 VSS.n3256 VSS.n3255 9.3005
R2793 VSS.n3258 VSS.n3257 9.3005
R2794 VSS.n3260 VSS.n114 9.3005
R2795 VSS.n3264 VSS.n3263 9.3005
R2796 VSS.n3265 VSS.n113 9.3005
R2797 VSS.n3268 VSS.n3266 9.3005
R2798 VSS.n3270 VSS.n3269 9.3005
R2799 VSS.n3271 VSS.n110 9.3005
R2800 VSS.n3273 VSS.n3272 9.3005
R2801 VSS.n3274 VSS.n109 9.3005
R2802 VSS.n3276 VSS.n3275 9.3005
R2803 VSS.n3277 VSS.n108 9.3005
R2804 VSS.n3279 VSS.n3278 9.3005
R2805 VSS.n3293 VSS.n3292 9.3005
R2806 VSS.n3232 VSS.n3231 9.3005
R2807 VSS.n171 VSS.n170 9.3005
R2808 VSS.n3341 VSS.n3338 9.3005
R2809 VSS.n3337 VSS.n68 9.3005
R2810 VSS.n3336 VSS.n3335 9.3005
R2811 VSS.n126 VSS.n69 9.3005
R2812 VSS.n128 VSS.n127 9.3005
R2813 VSS.n129 VSS.n125 9.3005
R2814 VSS.n131 VSS.n130 9.3005
R2815 VSS.n133 VSS.n132 9.3005
R2816 VSS.n134 VSS.n124 9.3005
R2817 VSS.n136 VSS.n135 9.3005
R2818 VSS.n138 VSS.n137 9.3005
R2819 VSS.n139 VSS.n123 9.3005
R2820 VSS.n141 VSS.n140 9.3005
R2821 VSS.n143 VSS.n142 9.3005
R2822 VSS.n144 VSS.n122 9.3005
R2823 VSS.n146 VSS.n145 9.3005
R2824 VSS.n148 VSS.n147 9.3005
R2825 VSS.n149 VSS.n121 9.3005
R2826 VSS.n151 VSS.n150 9.3005
R2827 VSS.n153 VSS.n152 9.3005
R2828 VSS.n154 VSS.n120 9.3005
R2829 VSS.n156 VSS.n155 9.3005
R2830 VSS.n158 VSS.n157 9.3005
R2831 VSS.n159 VSS.n119 9.3005
R2832 VSS.n161 VSS.n160 9.3005
R2833 VSS.n163 VSS.n162 9.3005
R2834 VSS.n164 VSS.n118 9.3005
R2835 VSS.n166 VSS.n165 9.3005
R2836 VSS.n168 VSS.n167 9.3005
R2837 VSS.n169 VSS.n117 9.3005
R2838 VSS.n1679 VSS.n1678 9.3005
R2839 VSS.n1681 VSS.n1680 9.3005
R2840 VSS.n1682 VSS.n1670 9.3005
R2841 VSS.n1685 VSS.n1684 9.3005
R2842 VSS.n1686 VSS.n1668 9.3005
R2843 VSS.n1694 VSS.n1693 9.3005
R2844 VSS.n1697 VSS.n1696 9.3005
R2845 VSS.n1666 VSS.n1627 9.3005
R2846 VSS.n1665 VSS.n1664 9.3005
R2847 VSS.n1663 VSS.n1630 9.3005
R2848 VSS.n1662 VSS.n1661 9.3005
R2849 VSS.n1658 VSS.n1631 9.3005
R2850 VSS.n1096 VSS.n1085 9.3005
R2851 VSS.n1098 VSS.n1085 9.3005
R2852 VSS.n1110 VSS.n1109 9.3005
R2853 VSS.n1112 VSS.n1111 9.3005
R2854 VSS.n1113 VSS.n1081 9.3005
R2855 VSS.n1115 VSS.n1114 9.3005
R2856 VSS.n1120 VSS.n1119 9.3005
R2857 VSS.n1126 VSS.n1125 9.3005
R2858 VSS.n1128 VSS.n1127 9.3005
R2859 VSS.n1137 VSS.n1136 9.3005
R2860 VSS.n1139 VSS.n1138 9.3005
R2861 VSS.n1141 VSS.n1140 9.3005
R2862 VSS.n1142 VSS.n1070 9.3005
R2863 VSS.n1145 VSS.n1144 9.3005
R2864 VSS.n1146 VSS.n1069 9.3005
R2865 VSS.n1148 VSS.n1147 9.3005
R2866 VSS.n1149 VSS.n1068 9.3005
R2867 VSS.n1152 VSS.n1151 9.3005
R2868 VSS.n1207 VSS.n1206 9.3005
R2869 VSS.n1205 VSS.n1067 9.3005
R2870 VSS.n1204 VSS.n1203 9.3005
R2871 VSS.n1203 VSS.n1202 9.3005
R2872 VSS.n1166 VSS.n1157 9.3005
R2873 VSS.n1166 VSS.n1165 9.3005
R2874 VSS.n1193 VSS.n1192 9.3005
R2875 VSS.n1190 VSS.n1162 9.3005
R2876 VSS.n1189 VSS.n1188 9.3005
R2877 VSS.n1187 VSS.n1168 9.3005
R2878 VSS.n1186 VSS.n1185 9.3005
R2879 VSS.n1184 VSS.n1169 9.3005
R2880 VSS.n1182 VSS.n1181 9.3005
R2881 VSS.n1180 VSS.n1170 9.3005
R2882 VSS.n1179 VSS.n1178 9.3005
R2883 VSS.n1176 VSS.n1171 9.3005
R2884 VSS.n2901 VSS.n2900 9.3005
R2885 VSS.n2898 VSS.n2897 9.3005
R2886 VSS.n2889 VSS.n512 9.3005
R2887 VSS.n2888 VSS.n2887 9.3005
R2888 VSS.n2886 VSS.n513 9.3005
R2889 VSS.n2885 VSS.n2884 9.3005
R2890 VSS.n2883 VSS.n2882 9.3005
R2891 VSS.n2881 VSS.n515 9.3005
R2892 VSS.n2879 VSS.n2878 9.3005
R2893 VSS.n2877 VSS.n2876 9.3005
R2894 VSS.n2875 VSS.n2874 9.3005
R2895 VSS.n2873 VSS.n2872 9.3005
R2896 VSS.n2871 VSS.n2870 9.3005
R2897 VSS.n2869 VSS.n2868 9.3005
R2898 VSS.n2867 VSS.n2866 9.3005
R2899 VSS.n1640 VSS.n521 9.3005
R2900 VSS.n1638 VSS.n1637 9.3005
R2901 VSS.n1646 VSS.n1645 9.3005
R2902 VSS.n1647 VSS.n1636 9.3005
R2903 VSS.n1649 VSS.n1648 9.3005
R2904 VSS.n1651 VSS.n1650 9.3005
R2905 VSS.n1652 VSS.n1634 9.3005
R2906 VSS.n1654 VSS.n1653 9.3005
R2907 VSS.n1656 VSS.n1655 9.3005
R2908 VSS.n2834 VSS.n2833 9.3005
R2909 VSS.n2831 VSS.n2830 9.3005
R2910 VSS.n2829 VSS.n543 9.3005
R2911 VSS.n2828 VSS.n2827 9.3005
R2912 VSS.n2826 VSS.n2825 9.3005
R2913 VSS.n2824 VSS.n545 9.3005
R2914 VSS.n2822 VSS.n2821 9.3005
R2915 VSS.n2832 VSS.n541 9.3005
R2916 VSS.n2839 VSS.n2838 9.3005
R2917 VSS.n2840 VSS.n540 9.3005
R2918 VSS.n2842 VSS.n2841 9.3005
R2919 VSS.n2845 VSS.n533 9.3005
R2920 VSS.n2848 VSS.n2847 9.3005
R2921 VSS.n1574 VSS.n1573 9.3005
R2922 VSS.n1608 VSS.n1590 9.3005
R2923 VSS.n1602 VSS.n1601 9.3005
R2924 VSS.n1600 VSS.n1599 9.3005
R2925 VSS.n1604 VSS.n1592 9.3005
R2926 VSS.n1607 VSS.n1606 9.3005
R2927 VSS.n1616 VSS.n1615 9.3005
R2928 VSS.n1618 VSS.n1617 9.3005
R2929 VSS.n1588 VSS.n1561 9.3005
R2930 VSS.n1587 VSS.n1565 9.3005
R2931 VSS.n1586 VSS.n1585 9.3005
R2932 VSS.n1584 VSS.n1566 9.3005
R2933 VSS.n1583 VSS.n1582 9.3005
R2934 VSS.n1581 VSS.n1567 9.3005
R2935 VSS.n1580 VSS.n1569 9.3005
R2936 VSS.n1579 VSS.n1578 9.3005
R2937 VSS.n1577 VSS.n1571 9.3005
R2938 VSS.n1576 VSS.n1575 9.3005
R2939 VSS.n1572 VSS.n537 9.3005
R2940 VSS.n2846 VSS.n534 9.3005
R2941 VSS.n2820 VSS.n546 9.3005
R2942 VSS.n2812 VSS.n2811 9.3005
R2943 VSS.n2809 VSS.n551 9.3005
R2944 VSS.n2808 VSS.n2807 9.3005
R2945 VSS.n2801 VSS.n2800 9.3005
R2946 VSS.n2697 VSS.n593 9.3005
R2947 VSS.n2693 VSS.n593 9.3005
R2948 VSS.n2710 VSS.n2709 9.3005
R2949 VSS.n2712 VSS.n2711 9.3005
R2950 VSS.n2713 VSS.n589 9.3005
R2951 VSS.n2717 VSS.n2716 9.3005
R2952 VSS.n2720 VSS.n2719 9.3005
R2953 VSS.n2722 VSS.n586 9.3005
R2954 VSS.n2724 VSS.n2723 9.3005
R2955 VSS.n2737 VSS.n2736 9.3005
R2956 VSS.n2739 VSS.n2738 9.3005
R2957 VSS.n2741 VSS.n2740 9.3005
R2958 VSS.n2742 VSS.n575 9.3005
R2959 VSS.n2745 VSS.n2744 9.3005
R2960 VSS.n2746 VSS.n574 9.3005
R2961 VSS.n2748 VSS.n2747 9.3005
R2962 VSS.n2749 VSS.n573 9.3005
R2963 VSS.n2752 VSS.n2751 9.3005
R2964 VSS.n2754 VSS.n2753 9.3005
R2965 VSS.n2757 VSS.n2756 9.3005
R2966 VSS.n2759 VSS.n2758 9.3005
R2967 VSS.n2762 VSS.n2761 9.3005
R2968 VSS.n2767 VSS.n2766 9.3005
R2969 VSS.n2777 VSS.n2776 9.3005
R2970 VSS.n2778 VSS.n558 9.3005
R2971 VSS.n2784 VSS.n2783 9.3005
R2972 VSS.n2785 VSS.n557 9.3005
R2973 VSS.n2787 VSS.n2786 9.3005
R2974 VSS.n2789 VSS.n556 9.3005
R2975 VSS.n2791 VSS.n2790 9.3005
R2976 VSS.n2793 VSS.n2792 9.3005
R2977 VSS.n2794 VSS.n554 9.3005
R2978 VSS.n2796 VSS.n2795 9.3005
R2979 VSS.n2798 VSS.n2797 9.3005
R2980 VSS.n964 VSS.n930 9.3005
R2981 VSS.n963 VSS.n962 9.3005
R2982 VSS.n959 VSS.n932 9.3005
R2983 VSS.n958 VSS.n957 9.3005
R2984 VSS.n956 VSS.n955 9.3005
R2985 VSS.n954 VSS.n934 9.3005
R2986 VSS.n953 VSS.n952 9.3005
R2987 VSS.n951 VSS.n935 9.3005
R2988 VSS.n943 VSS.n942 9.3005
R2989 VSS.n940 VSS.n939 9.3005
R2990 VSS.n1064 VSS.n1063 9.3005
R2991 VSS.n1062 VSS.n1061 9.3005
R2992 VSS.n1058 VSS.n1057 9.3005
R2993 VSS.n977 VSS.n976 9.3005
R2994 VSS.n978 VSS.n973 9.3005
R2995 VSS.n1047 VSS.n1046 9.3005
R2996 VSS.n1044 VSS.n1043 9.3005
R2997 VSS.n1042 VSS.n1041 9.3005
R2998 VSS.n1039 VSS.n980 9.3005
R2999 VSS.n1038 VSS 9.3005
R3000 VSS.n1037 VSS.n982 9.3005
R3001 VSS.n1036 VSS.n1035 9.3005
R3002 VSS.n1034 VSS.n1033 9.3005
R3003 VSS.n1032 VSS.n1031 9.3005
R3004 VSS.n1030 VSS.n987 9.3005
R3005 VSS.n1029 VSS.n1028 9.3005
R3006 VSS.n989 VSS.n988 9.3005
R3007 VSS.n1002 VSS.n1001 9.3005
R3008 VSS.n1003 VSS.n994 9.3005
R3009 VSS.n1019 VSS.n1018 9.3005
R3010 VSS.n1016 VSS.n995 9.3005
R3011 VSS.n1015 VSS.n1014 9.3005
R3012 VSS.n1013 VSS.n1012 9.3005
R3013 VSS.n1010 VSS.n1005 9.3005
R3014 VSS.n2683 VSS.n2682 9.3005
R3015 VSS.n2682 VSS.n605 9.3005
R3016 VSS.n2680 VSS.n2679 9.3005
R3017 VSS.n2678 VSS.n2677 9.3005
R3018 VSS.n2676 VSS.n618 9.3005
R3019 VSS.n2675 VSS.n2674 9.3005
R3020 VSS.n2672 VSS.n2671 9.3005
R3021 VSS.n2669 VSS.n2668 9.3005
R3022 VSS.n630 VSS.n624 9.3005
R3023 VSS.n635 VSS.n632 9.3005
R3024 VSS.n2658 VSS.n2657 9.3005
R3025 VSS.n2655 VSS.n633 9.3005
R3026 VSS.n2654 VSS.n2653 9.3005
R3027 VSS.n2652 VSS.n636 9.3005
R3028 VSS.n2651 VSS.n2650 9.3005
R3029 VSS.n2649 VSS.n637 9.3005
R3030 VSS.n2648 VSS.n2647 9.3005
R3031 VSS.n2646 VSS.n2645 9.3005
R3032 VSS.n2643 VSS.n2642 9.3005
R3033 VSS.n2641 VSS.n641 9.3005
R3034 VSS.n2640 VSS.n2639 9.3005
R3035 VSS.n2639 VSS.n2638 9.3005
R3036 VSS.n655 VSS.n646 9.3005
R3037 VSS.n655 VSS.n654 9.3005
R3038 VSS.n2629 VSS.n2628 9.3005
R3039 VSS.n2626 VSS.n651 9.3005
R3040 VSS.n2625 VSS.n2624 9.3005
R3041 VSS.n2623 VSS.n657 9.3005
R3042 VSS.n2622 VSS.n2621 9.3005
R3043 VSS.n2620 VSS.n658 9.3005
R3044 VSS.n2618 VSS.n2617 9.3005
R3045 VSS.n2616 VSS.n659 9.3005
R3046 VSS.n2615 VSS.n2614 9.3005
R3047 VSS.n2612 VSS.n660 9.3005
R3048 VSS.n1521 VSS.n1520 9.3005
R3049 VSS.n1509 VSS.n1508 9.3005
R3050 VSS.n1506 VSS.n1505 9.3005
R3051 VSS.n2584 VSS.n2583 9.3005
R3052 VSS.n2575 VSS.n2574 9.3005
R3053 VSS.n686 VSS.n683 9.3005
R3054 VSS.n2566 VSS.n2565 9.3005
R3055 VSS.n694 VSS.n687 9.3005
R3056 VSS.n2557 VSS.n2556 9.3005
R3057 VSS.n2554 VSS.n2553 9.3005
R3058 VSS.n2547 VSS.n696 9.3005
R3059 VSS.n2546 VSS.n2545 9.3005
R3060 VSS.n2544 VSS.n697 9.3005
R3061 VSS.n2541 VSS.n2540 9.3005
R3062 VSS.n2539 VSS.n701 9.3005
R3063 VSS.n2538 VSS.n2537 9.3005
R3064 VSS.n2535 VSS.n702 9.3005
R3065 VSS.n2532 VSS.n2531 9.3005
R3066 VSS.n2530 VSS.n2529 9.3005
R3067 VSS.n2527 VSS.n706 9.3005
R3068 VSS.n2526 VSS.n2525 9.3005
R3069 VSS.n710 VSS.n709 9.3005
R3070 VSS.n726 VSS.n725 9.3005
R3071 VSS.n727 VSS.n716 9.3005
R3072 VSS.n746 VSS.n745 9.3005
R3073 VSS.n743 VSS.n742 9.3005
R3074 VSS.n741 VSS.n740 9.3005
R3075 VSS.n739 VSS.n730 9.3005
R3076 VSS.n736 VSS.n735 9.3005
R3077 VSS.n2572 VSS.n2571 9.3005
R3078 VSS.n2573 VSS.n682 9.3005
R3079 VSS.n2579 VSS.n680 9.3005
R3080 VSS.n2581 VSS.n2580 9.3005
R3081 VSS.n2582 VSS.n678 9.3005
R3082 VSS.n2585 VSS.n677 9.3005
R3083 VSS.n2587 VSS.n2586 9.3005
R3084 VSS.n2588 VSS.n676 9.3005
R3085 VSS.n2597 VSS.n2596 9.3005
R3086 VSS.n2599 VSS.n2598 9.3005
R3087 VSS.n1489 VSS.n1488 9.3005
R3088 VSS.n1490 VSS.n1487 9.3005
R3089 VSS.n1492 VSS.n1491 9.3005
R3090 VSS.n1493 VSS.n1484 9.3005
R3091 VSS.n1498 VSS.n1497 9.3005
R3092 VSS.n1499 VSS.n1483 9.3005
R3093 VSS.n1501 VSS.n1500 9.3005
R3094 VSS.n1504 VSS.n1479 9.3005
R3095 VSS.n1507 VSS.n1478 9.3005
R3096 VSS.n1513 VSS.n1512 9.3005
R3097 VSS.n1475 VSS.n1464 9.3005
R3098 VSS.n1522 VSS.n1462 9.3005
R3099 VSS.n1524 VSS.n1523 9.3005
R3100 VSS.n1525 VSS.n1363 9.3005
R3101 VSS.n1527 VSS.n1526 9.3005
R3102 VSS.n1460 VSS.n1362 9.3005
R3103 VSS.n1459 VSS.n1458 9.3005
R3104 VSS.n1456 VSS.n1364 9.3005
R3105 VSS.n1455 VSS.n1454 9.3005
R3106 VSS.n1453 VSS.n1365 9.3005
R3107 VSS.n1452 VSS.n1451 9.3005
R3108 VSS.n1448 VSS.n1366 9.3005
R3109 VSS.n1447 VSS.n1446 9.3005
R3110 VSS.n1436 VSS.n1368 9.3005
R3111 VSS.n1397 VSS.n1386 9.3005
R3112 VSS.n1398 VSS.n1397 9.3005
R3113 VSS.n1406 VSS.n1382 9.3005
R3114 VSS.n1408 VSS.n1407 9.3005
R3115 VSS.n1411 VSS.n1410 9.3005
R3116 VSS.n1413 VSS.n1412 9.3005
R3117 VSS.n1414 VSS.n1380 9.3005
R3118 VSS.n1416 VSS.n1415 9.3005
R3119 VSS.n1418 VSS.n1417 9.3005
R3120 VSS.n1420 VSS.n1419 9.3005
R3121 VSS.n1421 VSS.n1378 9.3005
R3122 VSS.n1423 VSS.n1422 9.3005
R3123 VSS.n1425 VSS.n1376 9.3005
R3124 VSS.n1427 VSS.n1426 9.3005
R3125 VSS.n1433 VSS.n1432 9.3005
R3126 VSS.n1438 VSS.n1437 9.3005
R3127 VSS.n2301 VSS.n844 9.3005
R3128 VSS.n2301 VSS.n843 9.3005
R3129 VSS.n2302 VSS.n841 9.3005
R3130 VSS.n2307 VSS.n2306 9.3005
R3131 VSS.n2310 VSS.n2309 9.3005
R3132 VSS.n2311 VSS.n837 9.3005
R3133 VSS.n2314 VSS.n2313 9.3005
R3134 VSS.n2316 VSS.n2315 9.3005
R3135 VSS.n834 VSS.n833 9.3005
R3136 VSS.n2323 VSS.n2322 9.3005
R3137 VSS.n2324 VSS.n832 9.3005
R3138 VSS.n2326 VSS.n2325 9.3005
R3139 VSS.n2331 VSS.n2330 9.3005
R3140 VSS.n823 VSS.n821 9.3005
R3141 VSS.n2344 VSS.n2343 9.3005
R3142 VSS.n2346 VSS.n2345 9.3005
R3143 VSS.n2348 VSS.n2347 9.3005
R3144 VSS.n2350 VSS.n816 9.3005
R3145 VSS.n2353 VSS.n2352 9.3005
R3146 VSS.n2355 VSS.n2354 9.3005
R3147 VSS.n2358 VSS.n813 9.3005
R3148 VSS.n2364 VSS.n2363 9.3005
R3149 VSS.n2366 VSS.n2365 9.3005
R3150 VSS.n2370 VSS.n2369 9.3005
R3151 VSS.n2371 VSS.n810 9.3005
R3152 VSS.n2373 VSS.n2372 9.3005
R3153 VSS.n2376 VSS.n807 9.3005
R3154 VSS.n2380 VSS.n2379 9.3005
R3155 VSS.n2391 VSS.n2390 9.3005
R3156 VSS.n2393 VSS.n2392 9.3005
R3157 VSS.n2394 VSS.n795 9.3005
R3158 VSS.n2396 VSS.n2395 9.3005
R3159 VSS.n2399 VSS.n793 9.3005
R3160 VSS.n2401 VSS.n2400 9.3005
R3161 VSS.n2402 VSS.n792 9.3005
R3162 VSS.n2404 VSS.n2403 9.3005
R3163 VSS.n2406 VSS.n791 9.3005
R3164 VSS.n2408 VSS.n2407 9.3005
R3165 VSS.n2409 VSS.n790 9.3005
R3166 VSS.n2411 VSS.n2410 9.3005
R3167 VSS.n2414 VSS.n2413 9.3005
R3168 VSS.n2416 VSS.n783 9.3005
R3169 VSS.n2429 VSS.n2428 9.3005
R3170 VSS.n2433 VSS.n2432 9.3005
R3171 VSS.n2434 VSS.n781 9.3005
R3172 VSS.n2437 VSS.n2435 9.3005
R3173 VSS.n2439 VSS.n2438 9.3005
R3174 VSS.n2442 VSS.n2441 9.3005
R3175 VSS.n2445 VSS.n2444 9.3005
R3176 VSS.n2446 VSS.n776 9.3005
R3177 VSS.n2448 VSS.n2447 9.3005
R3178 VSS.n2450 VSS.n2449 9.3005
R3179 VSS.n2451 VSS.n766 9.3005
R3180 VSS.n2464 VSS.n2463 9.3005
R3181 VSS.n2465 VSS.n765 9.3005
R3182 VSS.n2467 VSS.n2466 9.3005
R3183 VSS.n2469 VSS.n2468 9.3005
R3184 VSS.n2470 VSS.n761 9.3005
R3185 VSS.n2472 VSS.n2471 9.3005
R3186 VSS.n2473 VSS.n760 9.3005
R3187 VSS.n2475 VSS.n2474 9.3005
R3188 VSS.n2476 VSS.n758 9.3005
R3189 VSS.n2481 VSS.n2480 9.3005
R3190 VSS.n2482 VSS.n757 9.3005
R3191 VSS.n2484 VSS.n2483 9.3005
R3192 VSS.n2485 VSS.n755 9.3005
R3193 VSS.n2515 VSS.n2514 9.3005
R3194 VSS.n2511 VSS.n2510 9.3005
R3195 VSS.n2503 VSS.n2502 9.3005
R3196 VSS.n2500 VSS.n2488 9.3005
R3197 VSS.n2498 VSS.n2492 9.3005
R3198 VSS.n2289 VSS.n2288 9.3005
R3199 VSS.n2288 VSS.n866 9.3005
R3200 VSS.n2287 VSS.n2286 9.3005
R3201 VSS.n2285 VSS.n2284 9.3005
R3202 VSS.n2283 VSS.n2282 9.3005
R3203 VSS.n2281 VSS.n2280 9.3005
R3204 VSS.n2279 VSS.n879 9.3005
R3205 VSS.n2278 VSS.n2277 9.3005
R3206 VSS.n2276 VSS.n2275 9.3005
R3207 VSS.n2274 VSS.n883 9.3005
R3208 VSS.n2273 VSS.n884 9.3005
R3209 VSS.n2272 VSS.n2271 9.3005
R3210 VSS.n2270 VSS.n886 9.3005
R3211 VSS.n2269 VSS.n2268 9.3005
R3212 VSS.n2267 VSS.n889 9.3005
R3213 VSS.n2266 VSS.n2265 9.3005
R3214 VSS.n892 VSS.n890 9.3005
R3215 VSS.n2251 VSS.n2250 9.3005
R3216 VSS.n2249 VSS.n894 9.3005
R3217 VSS.n2248 VSS.n2247 9.3005
R3218 VSS.n2246 VSS.n896 9.3005
R3219 VSS.n2245 VSS.n2244 9.3005
R3220 VSS.n2243 VSS.n2242 9.3005
R3221 VSS.n2241 VSS.n2240 9.3005
R3222 VSS.n2238 VSS.n899 9.3005
R3223 VSS.n2237 VSS.n901 9.3005
R3224 VSS.n2055 VSS.n2054 9.3005
R3225 VSS.n2056 VSS.n2053 9.3005
R3226 VSS.n2063 VSS.n2062 9.3005
R3227 VSS.n2065 VSS.n2064 9.3005
R3228 VSS.n2048 VSS.n2047 9.3005
R3229 VSS.n2075 VSS.n2074 9.3005
R3230 VSS.n2076 VSS.n2044 9.3005
R3231 VSS.n2078 VSS.n2077 9.3005
R3232 VSS.n2079 VSS.n2043 9.3005
R3233 VSS.n2081 VSS.n2080 9.3005
R3234 VSS.n2041 VSS.n2040 9.3005
R3235 VSS.n2087 VSS.n2086 9.3005
R3236 VSS.n2088 VSS.n2039 9.3005
R3237 VSS.n2090 VSS.n2089 9.3005
R3238 VSS.n2091 VSS.n2038 9.3005
R3239 VSS.n2093 VSS.n2092 9.3005
R3240 VSS.n2095 VSS.n2094 9.3005
R3241 VSS.n2100 VSS.n2099 9.3005
R3242 VSS.n2032 VSS.n909 9.3005
R3243 VSS.n2110 VSS.n2109 9.3005
R3244 VSS.n2111 VSS.n908 9.3005
R3245 VSS.n2114 VSS.n2113 9.3005
R3246 VSS.n2115 VSS.n907 9.3005
R3247 VSS.n2117 VSS.n2116 9.3005
R3248 VSS.n2119 VSS.n904 9.3005
R3249 VSS.n2121 VSS.n2120 9.3005
R3250 VSS.n2122 VSS.n903 9.3005
R3251 VSS.n2234 VSS.n2123 9.3005
R3252 VSS.n2233 VSS.n2232 9.3005
R3253 VSS.n2231 VSS.n2230 9.3005
R3254 VSS.n2227 VSS.n2226 9.3005
R3255 VSS.n2135 VSS.n2125 9.3005
R3256 VSS.n2141 VSS.n2140 9.3005
R3257 VSS.n2143 VSS.n2130 9.3005
R3258 VSS.n2217 VSS.n2216 9.3005
R3259 VSS.n2215 VSS.n2131 9.3005
R3260 VSS.n2213 VSS.n2212 9.3005
R3261 VSS.n2211 VSS.n2145 9.3005
R3262 VSS.n2210 VSS.n2209 9.3005
R3263 VSS.n2208 VSS.n2146 9.3005
R3264 VSS.n2206 VSS.n2205 9.3005
R3265 VSS.n2204 VSS.n2149 9.3005
R3266 VSS.n2203 VSS.n2202 9.3005
R3267 VSS.n2200 VSS.n2150 9.3005
R3268 VSS.n2196 VSS.n2195 9.3005
R3269 VSS.n2161 VSS.n2152 9.3005
R3270 VSS.n2169 VSS.n2168 9.3005
R3271 VSS.n2170 VSS.n2157 9.3005
R3272 VSS.n2186 VSS.n2185 9.3005
R3273 VSS.n2184 VSS.n2158 9.3005
R3274 VSS.n2183 VSS.n2182 9.3005
R3275 VSS.n2181 VSS.n2180 9.3005
R3276 VSS.n2178 VSS.n2173 9.3005
R3277 VSS.n1935 VSS.n1934 9.3005
R3278 VSS.n1937 VSS.n1936 9.3005
R3279 VSS.n1239 VSS.n1238 9.3005
R3280 VSS.n1252 VSS.n1251 9.3005
R3281 VSS.n1254 VSS.n1253 9.3005
R3282 VSS.n1255 VSS.n1228 9.3005
R3283 VSS.n1257 VSS.n1256 9.3005
R3284 VSS.n1259 VSS.n1258 9.3005
R3285 VSS.n1260 VSS.n1226 9.3005
R3286 VSS.n1262 VSS.n1261 9.3005
R3287 VSS.n1264 VSS.n1263 9.3005
R3288 VSS.n1266 VSS.n1265 9.3005
R3289 VSS.n1267 VSS.n1223 9.3005
R3290 VSS.n1271 VSS.n1270 9.3005
R3291 VSS.n1272 VSS.n1221 9.3005
R3292 VSS.n1274 VSS.n1273 9.3005
R3293 VSS.n1276 VSS.n1275 9.3005
R3294 VSS.n1278 VSS.n1215 9.3005
R3295 VSS.n1291 VSS.n1290 9.3005
R3296 VSS.n1293 VSS.n1214 9.3005
R3297 VSS.n1297 VSS.n1296 9.3005
R3298 VSS.n1300 VSS.n1299 9.3005
R3299 VSS.n1303 VSS.n1302 9.3005
R3300 VSS.n1304 VSS.n1212 9.3005
R3301 VSS.n1357 VSS.n1305 9.3005
R3302 VSS.n1356 VSS.n1355 9.3005
R3303 VSS.n1354 VSS.n1353 9.3005
R3304 VSS.n1352 VSS.n1351 9.3005
R3305 VSS.n1340 VSS.n1310 9.3005
R3306 VSS.n1340 VSS.n1318 9.3005
R3307 VSS.n1341 VSS.n1340 9.3005
R3308 VSS.n1339 VSS.n1338 9.3005
R3309 VSS.n1337 VSS.n1320 9.3005
R3310 VSS.n1336 VSS.n1335 9.3005
R3311 VSS.n1334 VSS.n1333 9.3005
R3312 VSS.n1332 VSS.n1321 9.3005
R3313 VSS.n1331 VSS.n1330 9.3005
R3314 VSS.n1329 VSS.n1322 9.3005
R3315 VSS.n1325 VSS.n918 9.3005
R3316 VSS.n2023 VSS.n2022 9.3005
R3317 VSS.n2021 VSS.n2020 9.3005
R3318 VSS.n2015 VSS.n920 9.3005
R3319 VSS.n2014 VSS.n2013 9.3005
R3320 VSS.n2011 VSS.n924 9.3005
R3321 VSS.n2010 VSS.n2009 9.3005
R3322 VSS.n2008 VSS.n2007 9.3005
R3323 VSS.n2006 VSS.n2005 9.3005
R3324 VSS.n2004 VSS.n928 9.3005
R3325 VSS.n2003 VSS.n2002 9.3005
R3326 VSS.n2001 VSS.n1896 9.3005
R3327 VSS.n2000 VSS.n1999 9.3005
R3328 VSS.n1998 VSS.n1997 9.3005
R3329 VSS.n1996 VSS.n1898 9.3005
R3330 VSS.n1995 VSS.n1994 9.3005
R3331 VSS.n1907 VSS.n1899 9.3005
R3332 VSS.n1978 VSS.n1909 9.3005
R3333 VSS.n1984 VSS.n1983 9.3005
R3334 VSS.n1976 VSS.n1910 9.3005
R3335 VSS.n1975 VSS.n1974 9.3005
R3336 VSS.n1973 VSS.n1913 9.3005
R3337 VSS.n1972 VSS.n1971 9.3005
R3338 VSS.n1970 VSS.n1969 9.3005
R3339 VSS.n1968 VSS.n1914 9.3005
R3340 VSS.n1967 VSS.n1966 9.3005
R3341 VSS.n1965 VSS.n1915 9.3005
R3342 VSS.n1963 VSS.n1918 9.3005
R3343 VSS.n1962 VSS.n1961 9.3005
R3344 VSS.n1926 VSS.n1921 9.3005
R3345 VSS.n1945 VSS.n1944 9.3005
R3346 VSS.n1943 VSS.n1942 9.3005
R3347 VSS.n1941 VSS.n1927 9.3005
R3348 VSS.n1940 VSS.n1939 9.3005
R3349 VSS.n1938 VSS.n1928 9.3005
R3350 VSS.n244 VSS.n241 9.3005
R3351 VSS.n255 VSS.n254 9.3005
R3352 VSS.n2980 VSS.n2979 9.3005
R3353 VSS.n2977 VSS.n239 9.3005
R3354 VSS.n2974 VSS.n2973 9.3005
R3355 VSS.n2972 VSS.n256 9.3005
R3356 VSS.n2971 VSS.n2970 9.3005
R3357 VSS.n2969 VSS.n257 9.3005
R3358 VSS.n2968 VSS.n2967 9.3005
R3359 VSS.n2966 VSS.n259 9.3005
R3360 VSS.n2965 VSS.n2964 9.3005
R3361 VSS.n262 VSS.n260 9.3005
R3362 VSS.n2959 VSS.n2958 9.3005
R3363 VSS.n2957 VSS.n264 9.3005
R3364 VSS.n272 VSS.n265 9.3005
R3365 VSS.n2949 VSS.n2948 9.3005
R3366 VSS.n2947 VSS.n2946 9.3005
R3367 VSS.n2940 VSS.n273 9.3005
R3368 VSS.n2939 VSS.n2938 9.3005
R3369 VSS.n2937 VSS.n274 9.3005
R3370 VSS.n2936 VSS.n2935 9.3005
R3371 VSS.n2934 VSS.n2933 9.3005
R3372 VSS.n2932 VSS.n276 9.3005
R3373 VSS.n2931 VSS.n2930 9.3005
R3374 VSS.n2929 VSS.n2928 9.3005
R3375 VSS.n2927 VSS.n279 9.3005
R3376 VSS.n1738 VSS.n278 9.3005
R3377 VSS.n1743 VSS.n1742 9.3005
R3378 VSS.n1745 VSS.n1735 9.3005
R3379 VSS.n1754 VSS.n1753 9.3005
R3380 VSS.n1756 VSS.n1733 9.3005
R3381 VSS.n1793 VSS.n1792 9.3005
R3382 VSS.n1791 VSS.n1734 9.3005
R3383 VSS.n1790 VSS.n1789 9.3005
R3384 VSS.n1788 VSS.n1757 9.3005
R3385 VSS.n1787 VSS.n1786 9.3005
R3386 VSS.n1785 VSS.n1758 9.3005
R3387 VSS.n1783 VSS.n1782 9.3005
R3388 VSS.n1781 VSS.n1759 9.3005
R3389 VSS.n1780 VSS.n1779 9.3005
R3390 VSS.n1777 VSS 9.3005
R3391 VSS.n1776 VSS.n1775 9.3005
R3392 VSS.n1774 VSS.n1773 9.3005
R3393 VSS.n1772 VSS.n1771 9.3005
R3394 VSS.n1764 VSS.n1762 9.3005
R3395 VSS.n2911 VSS.n499 9.3005
R3396 VSS.n2913 VSS.n2912 9.3005
R3397 VSS.n2914 VSS.n498 9.3005
R3398 VSS.n2916 VSS.n2915 9.3005
R3399 VSS.n2918 VSS.n2917 9.3005
R3400 VSS.n2919 VSS.n496 9.3005
R3401 VSS.n2921 VSS.n2920 9.3005
R3402 VSS.n2923 VSS.n2922 9.3005
R3403 VSS.n2924 VSS.n494 9.3005
R3404 VSS.n1720 VSS.n493 9.3005
R3405 VSS.n1722 VSS.n1721 9.3005
R3406 VSS.n1724 VSS.n1723 9.3005
R3407 VSS.n1814 VSS.n1813 9.3005
R3408 VSS.n1816 VSS.n1815 9.3005
R3409 VSS.n1716 VSS.n1715 9.3005
R3410 VSS.n1822 VSS.n1821 9.3005
R3411 VSS.n1823 VSS.n1713 9.3005
R3412 VSS.n1829 VSS.n1828 9.3005
R3413 VSS.n1831 VSS.n1830 9.3005
R3414 VSS.n1833 VSS.n1832 9.3005
R3415 VSS.n1834 VSS.n1711 9.3005
R3416 VSS.n1836 VSS.n1835 9.3005
R3417 VSS.n1837 VSS.n1709 9.3005
R3418 VSS.n1840 VSS.n1839 9.3005
R3419 VSS.n1841 VSS.n1708 9.3005
R3420 VSS.n1843 VSS.n1842 9.3005
R3421 VSS.n1844 VSS.n1705 9.3005
R3422 VSS.n1871 VSS.n1870 9.3005
R3423 VSS.n1869 VSS.n1868 9.3005
R3424 VSS.n1866 VSS.n1845 9.3005
R3425 VSS.n1865 VSS.n1864 9.3005
R3426 VSS.n1863 VSS.n1848 9.3005
R3427 VSS.n1862 VSS.n1861 9.3005
R3428 VSS.n1860 VSS.n1859 9.3005
R3429 VSS.n1858 VSS.n1857 9.3005
R3430 VSS.n1856 VSS.n1855 9.3005
R3431 VSS.n2584 VSS.n678 9.12791
R3432 VSS.n1504 VSS.n1503 9.03579
R3433 VSS.n1482 VSS.n1481 9.03579
R3434 VSS.n2352 VSS.n2351 9.03579
R3435 VSS.n2534 VSS.n2532 8.9684
R3436 VSS.n328 VSS.n327 8.44328
R3437 VSS.n350 VSS.n349 8.44328
R3438 VSS.n3159 VSS.n3158 8.44328
R3439 VSS.n3213 VSS.n3212 8.44328
R3440 VSS.t610 VSS.t393 8.42962
R3441 VSS.t507 VSS.t721 8.42962
R3442 VSS.t645 VSS.t887 8.42962
R3443 VSS VSS.n3345 8.3721
R3444 VSS.n331 VSS.n330 8.33966
R3445 VSS.n3323 VSS.n3322 8.33966
R3446 VSS.n200 VSS.n181 8.31061
R3447 VSS.n2993 VSS.n227 8.30267
R3448 VSS.n2469 VSS.n763 8.28285
R3449 VSS.n1207 VSS.n1067 8.23546
R3450 VSS.n1661 VSS.n1630 8.23546
R3451 VSS.n1665 VSS.n1630 8.23546
R3452 VSS.n1666 VSS.n1665 8.23546
R3453 VSS.n1694 VSS.n1668 8.23546
R3454 VSS.n1031 VSS.n1030 8.23546
R3455 VSS.n1030 VSS.n1029 8.23546
R3456 VSS.n978 VSS.n977 8.23546
R3457 VSS.n1046 VSS.n978 8.23546
R3458 VSS.n1039 VSS.n1038 8.23546
R3459 VSS.n1038 VSS.n982 8.23546
R3460 VSS.n2643 VSS.n641 8.23546
R3461 VSS.n2527 VSS.n2526 8.23546
R3462 VSS.n2526 VSS.n709 8.23546
R3463 VSS.n727 VSS.n726 8.23546
R3464 VSS.n2556 VSS.n694 8.23546
R3465 VSS.n2554 VSS.n696 8.23546
R3466 VSS.n2545 VSS.n2544 8.23546
R3467 VSS.n2541 VSS.n701 8.23546
R3468 VSS.n1419 VSS.n1378 8.23546
R3469 VSS.n1423 VSS.n1378 8.23546
R3470 VSS.n1426 VSS.n1425 8.23546
R3471 VSS.n1448 VSS.n1447 8.23546
R3472 VSS.n1451 VSS.n1448 8.23546
R3473 VSS.n1455 VSS.n1365 8.23546
R3474 VSS.n1456 VSS.n1455 8.23546
R3475 VSS.n1458 VSS.n1456 8.23546
R3476 VSS.n1527 VSS.n1362 8.23546
R3477 VSS.n1527 VSS.n1363 8.23546
R3478 VSS.n2086 VSS.n2039 8.23546
R3479 VSS.n2090 VSS.n2039 8.23546
R3480 VSS.n2091 VSS.n2090 8.23546
R3481 VSS.n2092 VSS.n2091 8.23546
R3482 VSS.n2099 VSS.n2095 8.23546
R3483 VSS.n2110 VSS.n909 8.23546
R3484 VSS.n2111 VSS.n2110 8.23546
R3485 VSS.n1839 VSS.n1708 8.23546
R3486 VSS.n1843 VSS.n1708 8.23546
R3487 VSS.n1844 VSS.n1843 8.23546
R3488 VSS.n1870 VSS.n1844 8.23546
R3489 VSS.n1870 VSS.n1869 8.23546
R3490 VSS.n1869 VSS.n1845 8.23546
R3491 VSS.n1864 VSS.n1863 8.23546
R3492 VSS.n1863 VSS.n1862 8.23546
R3493 VSS.n1773 VSS.n1772 8.23546
R3494 VSS.n1772 VSS.n1762 8.23546
R3495 VSS.n1762 VSS.n499 8.23546
R3496 VSS.n2913 VSS.n499 8.23546
R3497 VSS.n2914 VSS.n2913 8.23546
R3498 VSS.n2915 VSS.n2914 8.23546
R3499 VSS.n2919 VSS.n2918 8.23546
R3500 VSS.n2920 VSS.n2919 8.23546
R3501 VSS.n1792 VSS.n1756 8.23546
R3502 VSS.n1792 VSS.n1791 8.23546
R3503 VSS.n1791 VSS.n1790 8.23546
R3504 VSS.n1790 VSS.n1757 8.23546
R3505 VSS.n1786 VSS.n1757 8.23546
R3506 VSS.n1786 VSS.n1785 8.23546
R3507 VSS.n1783 VSS.n1759 8.23546
R3508 VSS.n1779 VSS.n1759 8.23546
R3509 VSS.n2948 VSS.n272 8.23546
R3510 VSS.n2948 VSS.n2947 8.23546
R3511 VSS.n2947 VSS.n273 8.23546
R3512 VSS.n2938 VSS.n273 8.23546
R3513 VSS.n2938 VSS.n2937 8.23546
R3514 VSS.n2937 VSS.n2936 8.23546
R3515 VSS.n2933 VSS.n2932 8.23546
R3516 VSS.n2932 VSS.n2931 8.23546
R3517 VSS.n1045 VSS.n1044 8.14595
R3518 VSS.n1696 VSS.n1667 8.05644
R3519 VSS.n329 VSS.n287 7.97888
R3520 VSS.n374 VSS.n228 7.97888
R3521 VSS.n3179 VSS.n78 7.97888
R3522 VSS.n3140 VSS.n3139 7.97888
R3523 VSS.n328 VSS.n288 7.97601
R3524 VSS.n351 VSS.n350 7.97601
R3525 VSS.n3212 VSS.n3211 7.97601
R3526 VSS.n3160 VSS.n3159 7.97601
R3527 VSS.n1497 VSS.n1496 7.90638
R3528 VSS.n2412 VSS.n2411 7.90638
R3529 VSS.n2207 VSS.n2206 7.90638
R3530 VSS.n1433 VSS.n1375 7.78791
R3531 VSS.n2084 VSS.n2083 7.72113
R3532 VSS.n2875 VSS.n518 7.6984
R3533 VSS.n1661 VSS.n1660 7.6984
R3534 VSS.n1031 VSS.n986 7.6984
R3535 VSS.n1041 VSS.n979 7.6984
R3536 VSS.n2529 VSS.n705 7.6984
R3537 VSS.n2567 VSS.n2566 7.6984
R3538 VSS.n2566 VSS.n685 7.6984
R3539 VSS.n2537 VSS.n2536 7.6984
R3540 VSS.n1434 VSS.n1433 7.6984
R3541 VSS.n1461 VSS.n1363 7.6984
R3542 VSS.n2086 VSS.n2085 7.6984
R3543 VSS.n2112 VSS.n2111 7.6984
R3544 VSS.n1839 VSS.n1838 7.6984
R3545 VSS.n1862 VSS.n1850 7.6984
R3546 VSS.n1773 VSS.n1760 7.6984
R3547 VSS.n2920 VSS.n495 7.6984
R3548 VSS.n1756 VSS.n1755 7.6984
R3549 VSS.n1779 VSS.n1778 7.6984
R3550 VSS.n272 VSS.n271 7.6984
R3551 VSS.n2931 VSS.n277 7.6984
R3552 VSS.n3083 VSS.n212 7.64725
R3553 VSS.n3108 VSS.n3106 7.64725
R3554 VSS.n3028 VSS.n221 7.64725
R3555 VSS.n3047 VSS.n3046 7.64725
R3556 VSS.n2162 VSS.n2160 7.6005
R3557 VSS.n1450 VSS.n1365 7.51938
R3558 VSS.n984 VSS.n982 7.34036
R3559 VSS.n2095 VSS.n2037 7.34036
R3560 VSS.n718 VSS.n709 7.25085
R3561 VSS.n1435 VSS.n1367 7.25085
R3562 VSS.n390 VSS.n227 7.16724
R3563 VSS.n3180 VSS.n3179 7.16724
R3564 VSS.n3211 VSS.n3210 7.16724
R3565 VSS.n3162 VSS.n3160 7.16724
R3566 VSS.n3158 VSS.n3157 7.16724
R3567 VSS.n3139 VSS.n3138 7.16724
R3568 VSS.n3324 VSS.n3323 7.16724
R3569 VSS.n3214 VSS.n3213 7.16724
R3570 VSS.n2528 VSS.n2527 7.16134
R3571 VSS.n3400 VSS.n3399 7.15344
R3572 VSS.n3268 VSS.n113 7.15344
R3573 VSS.n2876 VSS.n2875 7.11268
R3574 VSS.n1064 VSS.n930 7.11268
R3575 VSS.n1696 VSS.n1695 6.98232
R3576 VSS.n1029 VSS.n988 6.88949
R3577 VSS.n1419 VSS.n1418 6.88949
R3578 VSS.n2556 VSS.n2555 6.62428
R3579 VSS.n1166 VSS.n1156 6.61527
R3580 VSS.n655 VSS.n645 6.61527
R3581 VSS.n1882 VSS.t1008 6.6005
R3582 VSS.n1882 VSS.t1004 6.6005
R3583 VSS.n1884 VSS.t95 6.6005
R3584 VSS.n1884 VSS.t728 6.6005
R3585 VSS.n1547 VSS.t1006 6.6005
R3586 VSS.n1547 VSS.t720 6.6005
R3587 VSS.n1203 VSS.n1156 6.57117
R3588 VSS.n2639 VSS.n645 6.57117
R3589 VSS.n840 VSS.n839 6.57117
R3590 VSS.n2305 VSS.n840 6.57117
R3591 VSS.n728 VSS.n727 6.53477
R3592 VSS.n3388 VSS.n3387 6.50373
R3593 VSS.n3043 VSS.n209 6.50373
R3594 VSS.n3296 VSS.n3294 6.50373
R3595 VSS.n49 VSS.n48 6.4005
R3596 VSS.n3250 VSS.n3249 6.4005
R3597 VSS.n2119 VSS.n2118 6.4005
R3598 VSS.n2134 VSS.n2125 6.4005
R3599 VSS.n56 VSS.n55 6.26433
R3600 VSS.n3380 VSS.n3379 6.26433
R3601 VSS.n3243 VSS.n3242 6.26433
R3602 VSS.n103 VSS.n102 6.26433
R3603 VSS.n2580 VSS.n2579 6.26433
R3604 VSS.n2311 VSS.n2310 6.26433
R3605 VSS.n2284 VSS.n2283 6.26433
R3606 VSS.n1267 VSS.n1266 6.26433
R3607 VSS.n1296 VSS.n1293 6.26433
R3608 VSS.n1353 VSS.n1352 6.26433
R3609 VSS.n1330 VSS.n1329 6.26433
R3610 VSS.n2011 VSS.n2010 6.26433
R3611 VSS.n1997 VSS.n1996 6.26433
R3612 VSS.n1996 VSS.n1995 6.26433
R3613 VSS.n1966 VSS.n1965 6.26433
R3614 VSS.n1815 VSS.n1814 6.26433
R3615 VSS.n1815 VSS.n1715 6.26433
R3616 VSS.n2970 VSS.n2969 6.26433
R3617 VSS.n2969 VSS.n2968 6.26433
R3618 VSS.n2501 VSS.n2500 6.12816
R3619 VSS.n1604 VSS.n1603 6.06007
R3620 VSS.n315 VSS.n295 6.05269
R3621 VSS.n305 VSS.n301 6.05269
R3622 VSS.n326 VSS.n325 6.05269
R3623 VSS.n336 VSS.n332 6.05269
R3624 VSS.n380 VSS.n375 6.05269
R3625 VSS.n357 VSS.n352 6.05269
R3626 VSS.n364 VSS.n345 6.05269
R3627 VSS.n202 VSS.n201 6.05269
R3628 VSS.n1138 VSS.n1137 6.02861
R3629 VSS.n2738 VSS.n2737 6.02861
R3630 VSS.n2800 VSS.n2798 6.02861
R3631 VSS.n2822 VSS.n546 6.02861
R3632 VSS.n2657 VSS.n635 6.02861
R3633 VSS.n1503 VSS.n1501 6.02403
R3634 VSS.n1511 VSS.n1510 6.02403
R3635 VSS.n2363 VSS.n2359 5.98311
R3636 VSS.n2230 VSS.n2124 5.98311
R3637 VSS.n2201 VSS.n2200 5.98311
R3638 VSS.n1238 VSS.n1230 5.98311
R3639 VSS.n1934 VSS.n1930 5.98311
R3640 VSS.n1855 VSS.n1851 5.98311
R3641 VSS.n1742 VSS.n1739 5.98311
R3642 VSS.n2978 VSS.n2977 5.98311
R3643 VSS.n244 VSS.n240 5.98311
R3644 VSS.n55 VSS.n42 5.85582
R3645 VSS.n3380 VSS.n40 5.85582
R3646 VSS.n32 VSS.n31 5.85582
R3647 VSS.n6 VSS.n3 5.85582
R3648 VSS.n10 VSS.n7 5.85582
R3649 VSS.n3244 VSS.n3243 5.85582
R3650 VSS.n103 VSS.n97 5.85582
R3651 VSS.n3258 VSS.n115 5.85582
R3652 VSS.n3260 VSS.n3259 5.85582
R3653 VSS.n3288 VSS.n3280 5.85582
R3654 VSS.n1605 VSS.n1604 5.85582
R3655 VSS.n2580 VSS.n681 5.85582
R3656 VSS.n2306 VSS.n2303 5.85582
R3657 VSS.n2502 VSS.n2486 5.85582
R3658 VSS.n2284 VSS.n868 5.85582
R3659 VSS.n2169 VSS.n2163 5.85582
R3660 VSS.n1266 VSS.n1224 5.85582
R3661 VSS.n1293 VSS.n1292 5.85582
R3662 VSS.n1353 VSS.n1306 5.85582
R3663 VSS.n1330 VSS.n1323 5.85582
R3664 VSS.n2012 VSS.n2011 5.85582
R3665 VSS.n1997 VSS.n1897 5.85582
R3666 VSS.n1966 VSS.n1916 5.85582
R3667 VSS.n1814 VSS.n1719 5.85582
R3668 VSS.n2970 VSS.n258 5.85582
R3669 VSS.n1995 VSS.n1899 5.65809
R3670 VSS.n1822 VSS.n1715 5.65809
R3671 VSS.n2968 VSS.n259 5.65809
R3672 VSS.n1154 VSS.n1067 5.63966
R3673 VSS.n977 VSS.n966 5.63966
R3674 VSS.n1064 VSS.n931 5.63966
R3675 VSS.n643 VSS.n641 5.63966
R3676 VSS.n2835 VSS.n541 5.5878
R3677 VSS.n699 VSS.n696 5.55015
R3678 VSS.n2755 VSS.n2754 5.48621
R3679 VSS.n2787 VSS.n557 5.48128
R3680 VSS.n2170 VSS.n2169 5.37524
R3681 VSS.n2443 VSS.n2442 5.27109
R3682 VSS.n2313 VSS.n2312 5.24958
R3683 VSS.n1085 VSS.n1083 5.13108
R3684 VSS.n1085 VSS.n1084 5.13108
R3685 VSS.n1108 VSS.n1086 5.13108
R3686 VSS.n1108 VSS.n1107 5.13108
R3687 VSS.n1677 VSS.n1674 5.13108
R3688 VSS.n1677 VSS.n1675 5.13108
R3689 VSS.n593 VSS.n591 5.13108
R3690 VSS.n593 VSS.n592 5.13108
R3691 VSS.n2708 VSS.n594 5.13108
R3692 VSS.n2708 VSS.n2707 5.13108
R3693 VSS.n1598 VSS.n1595 5.13108
R3694 VSS.n1598 VSS.n1597 5.13108
R3695 VSS.n1009 VSS.n1006 5.13108
R3696 VSS.n1009 VSS.n1008 5.13108
R3697 VSS.n2682 VSS.n604 5.13108
R3698 VSS.n2682 VSS.n606 5.13108
R3699 VSS.n2681 VSS.n607 5.13108
R3700 VSS.n2681 VSS.n616 5.13108
R3701 VSS.n1397 VSS.n1388 5.13108
R3702 VSS.n1397 VSS.n1389 5.13108
R3703 VSS.n733 VSS.n731 5.13108
R3704 VSS.n733 VSS.n732 5.13108
R3705 VSS.n2301 VSS.n842 5.13108
R3706 VSS.n2301 VSS.n2300 5.13108
R3707 VSS.n2497 VSS.n2494 5.13108
R3708 VSS.n2497 VSS.n2495 5.13108
R3709 VSS.n2288 VSS.n865 5.13108
R3710 VSS.n2288 VSS.n867 5.13108
R3711 VSS.n2177 VSS.n2174 5.13108
R3712 VSS.n2177 VSS.n2175 5.13108
R3713 VSS.n2537 VSS.n704 4.92358
R3714 VSS.n2926 VSS.n492 4.89029
R3715 VSS.n2781 VSS.n2780 4.85762
R3716 VSS.n2319 VSS.n835 4.85762
R3717 VSS.n1981 VSS.n1980 4.85762
R3718 VSS.n2962 VSS.n263 4.85762
R3719 VSS.n1826 VSS.n1825 4.85762
R3720 VSS.n2230 VSS.n2229 4.8005
R3721 VSS.n1238 VSS.n1237 4.8005
R3722 VSS.n1934 VSS.n1933 4.8005
R3723 VSS.n1855 VSS.n1854 4.8005
R3724 VSS.n1742 VSS.n1741 4.8005
R3725 VSS.n2977 VSS.n2976 4.8005
R3726 VSS.n245 VSS.n244 4.8005
R3727 VSS.n3387 VSS.n36 4.788
R3728 VSS.n209 VSS.n194 4.788
R3729 VSS.n3297 VSS.n3296 4.788
R3730 VSS.n1175 VSS.n1174 4.72533
R3731 VSS.n2611 VSS.n2610 4.72533
R3732 VSS.n1127 VSS.n1126 4.67352
R3733 VSS.n1142 VSS.n1141 4.67352
R3734 VSS.n1144 VSS.n1142 4.67352
R3735 VSS.n1148 VSS.n1069 4.67352
R3736 VSS.n1149 VSS.n1148 4.67352
R3737 VSS.n1190 VSS.n1189 4.67352
R3738 VSS.n1189 VSS.n1168 4.67352
R3739 VSS.n1185 VSS.n1168 4.67352
R3740 VSS.n1185 VSS.n1184 4.67352
R3741 VSS.n1182 VSS.n1170 4.67352
R3742 VSS.n2898 VSS.n512 4.67352
R3743 VSS.n2887 VSS.n512 4.67352
R3744 VSS.n2887 VSS.n2886 4.67352
R3745 VSS.n2886 VSS.n2885 4.67352
R3746 VSS.n2882 VSS.n2881 4.67352
R3747 VSS.n2868 VSS.n2867 4.67352
R3748 VSS.n2867 VSS.n521 4.67352
R3749 VSS.n1637 VSS.n521 4.67352
R3750 VSS.n1646 VSS.n1637 4.67352
R3751 VSS.n1647 VSS.n1646 4.67352
R3752 VSS.n1648 VSS.n1647 4.67352
R3753 VSS.n1652 VSS.n1651 4.67352
R3754 VSS.n1653 VSS.n1652 4.67352
R3755 VSS.n2723 VSS.n2722 4.67352
R3756 VSS.n2742 VSS.n2741 4.67352
R3757 VSS.n2744 VSS.n2742 4.67352
R3758 VSS.n2748 VSS.n574 4.67352
R3759 VSS.n2749 VSS.n2748 4.67352
R3760 VSS.n2790 VSS.n2789 4.67352
R3761 VSS.n2794 VSS.n2793 4.67352
R3762 VSS.n2795 VSS.n2794 4.67352
R3763 VSS.n2809 VSS.n2808 4.67352
R3764 VSS.n2811 VSS.n2809 4.67352
R3765 VSS.n2825 VSS.n2824 4.67352
R3766 VSS.n2829 VSS.n2828 4.67352
R3767 VSS.n2830 VSS.n2829 4.67352
R3768 VSS.n2669 VSS.n624 4.67352
R3769 VSS.n2655 VSS.n2654 4.67352
R3770 VSS.n2654 VSS.n636 4.67352
R3771 VSS.n2650 VSS.n2649 4.67352
R3772 VSS.n2649 VSS.n2648 4.67352
R3773 VSS.n2626 VSS.n2625 4.67352
R3774 VSS.n2625 VSS.n657 4.67352
R3775 VSS.n2621 VSS.n657 4.67352
R3776 VSS.n2621 VSS.n2620 4.67352
R3777 VSS.n2618 VSS.n659 4.67352
R3778 VSS.n942 VSS.n935 4.67352
R3779 VSS.n953 VSS.n935 4.67352
R3780 VSS.n954 VSS.n953 4.67352
R3781 VSS.n955 VSS.n954 4.67352
R3782 VSS.n959 VSS.n958 4.67352
R3783 VSS.n1167 VSS.n1166 4.63943
R3784 VSS.n1174 VSS.n511 4.63943
R3785 VSS.n656 VSS.n655 4.63943
R3786 VSS.n2610 VSS.n662 4.63943
R3787 VSS.n2498 VSS.n2491 4.62124
R3788 VSS.n1963 VSS.n1919 4.62124
R3789 VSS.n1174 VSS.n1173 4.62124
R3790 VSS.n1058 VSS.n967 4.62124
R3791 VSS.n2610 VSS.n2609 4.62124
R3792 VSS.n2308 VSS.n840 4.62124
R3793 VSS.n1203 VSS.n1154 4.6085
R3794 VSS.n2639 VSS.n643 4.6085
R3795 VSS.n1176 VSS.n1175 4.60638
R3796 VSS.n2612 VSS.n2611 4.60638
R3797 VSS.n473 VSS.n472 4.5578
R3798 VSS.n1192 VSS.n1167 4.55559
R3799 VSS.n2900 VSS.n511 4.55559
R3800 VSS.n2628 VSS.n656 4.55559
R3801 VSS.n940 VSS.n662 4.55559
R3802 VSS.n2598 VSS.n673 4.51815
R3803 VSS.n1496 VSS.n1483 4.51815
R3804 VSS.n2348 VSS.n819 4.51815
R3805 VSS.n2375 VSS.n2374 4.51815
R3806 VSS.n2237 VSS.n902 4.51815
R3807 VSS.n1726 VSS.n1725 4.51401
R3808 VSS.n1820 VSS.n1819 4.51401
R3809 VSS.n247 VSS.n243 4.51401
R3810 VSS.n2982 VSS.n2981 4.51401
R3811 VSS.n1744 VSS.n1737 4.51401
R3812 VSS.n1795 VSS.n1794 4.51401
R3813 VSS.n1765 VSS.n1761 4.51401
R3814 VSS.n2910 VSS.n2909 4.51401
R3815 VSS.n1396 VSS.n1395 4.51401
R3816 VSS.n1405 VSS.n1404 4.51401
R3817 VSS.n2524 VSS.n2523 4.51401
R3818 VSS.n748 VSS.n747 4.51401
R3819 VSS.n2904 VSS.n508 4.51401
R3820 VSS.n2894 VSS.n2890 4.51401
R3821 VSS.n1158 VSS.n1153 4.51401
R3822 VSS.n1194 VSS 4.51401
R3823 VSS.n1124 VSS.n1123 4.51401
R3824 VSS.n1135 VSS.n1134 4.51401
R3825 VSS.n1093 VSS.n1090 4.51401
R3826 VSS.n1105 VSS.n1104 4.51401
R3827 VSS.n1700 VSS.n1625 4.51401
R3828 VSS.n1692 VSS.n1691 4.51401
R3829 VSS.n523 VSS.n520 4.51401
R3830 VSS.n1644 VSS.n1643 4.51401
R3831 VSS.n2730 VSS.n584 4.51401
R3832 VSS.n2735 VSS.n2734 4.51401
R3833 VSS.n2700 VSS.n2690 4.51401
R3834 VSS.n2705 VSS.n2704 4.51401
R3835 VSS.n1621 VSS.n1559 4.51401
R3836 VSS.n1614 VSS.n1613 4.51401
R3837 VSS.n2806 VSS.n2805 4.51401
R3838 VSS.n2819 VSS.n2818 4.51401
R3839 VSS.n2770 VSS.n568 4.51401
R3840 VSS.n2775 VSS.n2774 4.51401
R3841 VSS.n2857 VSS.n531 4.51401
R3842 VSS.n536 VSS.n535 4.51401
R3843 VSS.n626 VSS.n622 4.51401
R3844 VSS.n2660 VSS.n2659 4.51401
R3845 VSS.n2686 VSS.n601 4.51401
R3846 VSS.n614 VSS.n613 4.51401
R3847 VSS.n1027 VSS.n1026 4.51401
R3848 VSS.n1021 VSS.n1020 4.51401
R3849 VSS.n2608 VSS.n2607 4.51401
R3850 VSS.n950 VSS.n949 4.51401
R3851 VSS.n647 VSS.n642 4.51401
R3852 VSS.n2630 VSS 4.51401
R3853 VSS.n969 VSS.n968 4.51401
R3854 VSS.n1049 VSS.n1048 4.51401
R3855 VSS.n2457 VSS.n772 4.51401
R3856 VSS.n2462 VSS.n2461 4.51401
R3857 VSS.n2225 VSS.n2224 4.51401
R3858 VSS.n2219 VSS.n2218 4.51401
R3859 VSS.n1902 VSS.n1900 4.51401
R3860 VSS.n1986 VSS.n1985 4.51401
R3861 VSS.n2564 VSS.n2563 4.51401
R3862 VSS.n2552 VSS.n2551 4.51401
R3863 VSS.n1472 VSS.n1470 4.51401
R3864 VSS.n1514 VSS 4.51401
R3865 VSS.n1431 VSS.n1430 4.51401
R3866 VSS.n1445 VSS.n1444 4.51401
R3867 VSS.n2602 VSS.n669 4.51401
R3868 VSS.n2593 VSS.n2589 4.51401
R3869 VSS.n2103 VSS.n2030 4.51401
R3870 VSS.n2108 VSS.n2107 4.51401
R3871 VSS.n2026 VSS.n915 4.51401
R3872 VSS.n2017 VSS.n2016 4.51401
R3873 VSS.n2415 VSS.n787 4.51401
R3874 VSS.n2425 VSS.n782 4.51401
R3875 VSS.n2336 VSS.n829 4.51401
R3876 VSS.n2340 VSS.n820 4.51401
R3877 VSS.n2299 VSS.n2298 4.51401
R3878 VSS.n856 VSS.n855 4.51401
R3879 VSS.n2518 VSS.n753 4.51401
R3880 VSS.n2509 VSS.n2508 4.51401
R3881 VSS.n2383 VSS.n804 4.51401
R3882 VSS.n2387 VSS.n796 4.51401
R3883 VSS.n1311 VSS.n1307 4.51401
R3884 VSS.n1343 VSS.n1342 4.51401
R3885 VSS.n2061 VSS.n2060 4.51401
R3886 VSS.n2073 VSS.n2072 4.51401
R3887 VSS.n2292 VSS.n862 4.51401
R3888 VSS.n875 VSS.n874 4.51401
R3889 VSS.n2194 VSS.n2193 4.51401
R3890 VSS.n2188 VSS.n2187 4.51401
R3891 VSS.n2257 VSS.n887 4.51401
R3892 VSS.n2262 VSS.n2252 4.51401
R3893 VSS.n1284 VSS.n1219 4.51401
R3894 VSS.n1289 VSS.n1288 4.51401
R3895 VSS.n1235 VSS.n1234 4.51401
R3896 VSS.n1248 VSS.n1229 4.51401
R3897 VSS.n1952 VSS.n1949 4.51401
R3898 VSS.n1947 VSS.n1946 4.51401
R3899 VSS.n1874 VSS.n1704 4.51401
R3900 VSS.n1867 VSS.n1552 4.51401
R3901 VSS.n2956 VSS.n2955 4.51401
R3902 VSS.n2945 VSS.n2944 4.51401
R3903 VSS.n3387 VSS.n3386 4.50726
R3904 VSS.n3113 VSS.n209 4.50726
R3905 VSS.n3296 VSS.n3295 4.50726
R3906 VSS.n1699 VSS.n1698 4.5005
R3907 VSS.n1687 VSS.n1628 4.5005
R3908 VSS.n1690 VSS.n1669 4.5005
R3909 VSS.n1095 VSS.n1094 4.5005
R3910 VSS.n1100 VSS.n1099 4.5005
R3911 VSS.n1097 VSS.n1087 4.5005
R3912 VSS.n1121 VSS.n1077 4.5005
R3913 VSS.n1130 VSS.n1129 4.5005
R3914 VSS.n1074 VSS.n1073 4.5005
R3915 VSS.n1201 VSS.n1200 4.5005
R3916 VSS.n1163 VSS.n1159 4.5005
R3917 VSS.n1164 VSS.n1161 4.5005
R3918 VSS.n2903 VSS.n2902 4.5005
R3919 VSS.n2891 VSS.n510 4.5005
R3920 VSS.n2896 VSS.n2895 4.5005
R3921 VSS.n2865 VSS.n2864 4.5005
R3922 VSS.n524 VSS.n522 4.5005
R3923 VSS.n1642 VSS.n1641 4.5005
R3924 VSS.n563 VSS.n562 4.5005
R3925 VSS.n2803 VSS.n2802 4.5005
R3926 VSS.n2814 VSS.n2813 4.5005
R3927 VSS.n548 VSS.n547 4.5005
R3928 VSS.n1620 VSS.n1619 4.5005
R3929 VSS.n1609 VSS.n1562 4.5005
R3930 VSS.n1612 VSS.n1591 4.5005
R3931 VSS.n2699 VSS.n2698 4.5005
R3932 VSS.n2696 VSS.n2695 4.5005
R3933 VSS.n2692 VSS.n595 4.5005
R3934 VSS.n2729 VSS.n2728 4.5005
R3935 VSS.n2727 VSS.n2726 4.5005
R3936 VSS.n579 VSS.n578 4.5005
R3937 VSS.n2769 VSS.n2768 4.5005
R3938 VSS.n2765 VSS.n2764 4.5005
R3939 VSS.n2856 VSS.n2855 4.5005
R3940 VSS.n2854 VSS.n2853 4.5005
R3941 VSS.n2850 VSS.n2849 4.5005
R3942 VSS.n653 VSS.n650 4.5005
R3943 VSS.n938 VSS.n663 4.5005
R3944 VSS.n945 VSS.n944 4.5005
R3945 VSS.n948 VSS.n936 4.5005
R3946 VSS.n997 VSS.n990 4.5005
R3947 VSS.n1000 VSS.n999 4.5005
R3948 VSS.n998 VSS.n993 4.5005
R3949 VSS.n2685 VSS.n2684 4.5005
R3950 VSS.n608 VSS.n603 4.5005
R3951 VSS.n612 VSS.n611 4.5005
R3952 VSS.n2667 VSS.n2666 4.5005
R3953 VSS.n627 VSS.n625 4.5005
R3954 VSS.n631 VSS.n629 4.5005
R3955 VSS.n2637 VSS.n2636 4.5005
R3956 VSS.n652 VSS.n648 4.5005
R3957 VSS.n1056 VSS.n1055 4.5005
R3958 VSS.n974 VSS.n970 4.5005
R3959 VSS.n975 VSS.n972 4.5005
R3960 VSS.n1471 VSS.n1466 4.5005
R3961 VSS.n1519 VSS.n1518 4.5005
R3962 VSS.n1469 VSS.n1467 4.5005
R3963 VSS.n692 VSS.n688 4.5005
R3964 VSS.n2559 VSS.n2558 4.5005
R3965 VSS.n2548 VSS.n693 4.5005
R3966 VSS.n719 VSS.n711 4.5005
R3967 VSS.n724 VSS.n723 4.5005
R3968 VSS.n720 VSS.n715 4.5005
R3969 VSS.n1391 VSS.n1390 4.5005
R3970 VSS.n1400 VSS.n1399 4.5005
R3971 VSS.n1387 VSS.n1383 4.5005
R3972 VSS.n1428 VSS.n1372 4.5005
R3973 VSS.n1440 VSS.n1439 4.5005
R3974 VSS.n1373 VSS.n1369 4.5005
R3975 VSS.n2601 VSS.n2600 4.5005
R3976 VSS.n2590 VSS.n671 4.5005
R3977 VSS.n2595 VSS.n2594 4.5005
R3978 VSS.n2507 VSS.n2487 4.5005
R3979 VSS.n846 VSS.n845 4.5005
R3980 VSS.n851 VSS.n850 4.5005
R3981 VSS.n854 VSS.n853 4.5005
R3982 VSS.n2335 VSS.n2334 4.5005
R3983 VSS.n2333 VSS.n2332 4.5005
R3984 VSS.n2342 VSS.n2341 4.5005
R3985 VSS.n2418 VSS.n2417 4.5005
R3986 VSS.n2419 VSS.n784 4.5005
R3987 VSS.n2427 VSS.n2426 4.5005
R3988 VSS.n2456 VSS.n2455 4.5005
R3989 VSS.n2454 VSS.n2453 4.5005
R3990 VSS.n768 VSS.n767 4.5005
R3991 VSS.n2517 VSS.n2516 4.5005
R3992 VSS.n2504 VSS.n756 4.5005
R3993 VSS.n2382 VSS.n2381 4.5005
R3994 VSS.n805 VSS.n798 4.5005
R3995 VSS.n2389 VSS.n2388 4.5005
R3996 VSS.n2165 VSS.n2156 4.5005
R3997 VSS.n2291 VSS.n2290 4.5005
R3998 VSS.n869 VSS.n864 4.5005
R3999 VSS.n873 VSS.n872 4.5005
R4000 VSS.n2057 VSS.n2052 4.5005
R4001 VSS.n2068 VSS.n2067 4.5005
R4002 VSS.n2066 VSS.n2049 4.5005
R4003 VSS.n2102 VSS.n2101 4.5005
R4004 VSS.n2035 VSS.n2034 4.5005
R4005 VSS.n911 VSS.n910 4.5005
R4006 VSS.n2136 VSS.n2126 4.5005
R4007 VSS.n2138 VSS.n2137 4.5005
R4008 VSS.n2139 VSS.n2129 4.5005
R4009 VSS.n2164 VSS.n2153 4.5005
R4010 VSS.n2167 VSS.n2166 4.5005
R4011 VSS.n2256 VSS.n2255 4.5005
R4012 VSS.n2253 VSS.n891 4.5005
R4013 VSS.n2264 VSS.n2263 4.5005
R4014 VSS.n1241 VSS.n1240 4.5005
R4015 VSS.n1242 VSS.n1231 4.5005
R4016 VSS.n1250 VSS.n1249 4.5005
R4017 VSS.n1283 VSS.n1282 4.5005
R4018 VSS.n1281 VSS.n1280 4.5005
R4019 VSS.n1277 VSS.n1216 4.5005
R4020 VSS.n1350 VSS.n1349 4.5005
R4021 VSS.n1316 VSS.n1312 4.5005
R4022 VSS.n1317 VSS.n1315 4.5005
R4023 VSS.n2025 VSS.n2024 4.5005
R4024 VSS.n921 VSS.n917 4.5005
R4025 VSS.n2019 VSS.n2018 4.5005
R4026 VSS.n1993 VSS.n1992 4.5005
R4027 VSS.n1903 VSS.n1901 4.5005
R4028 VSS.n1908 VSS.n1906 4.5005
R4029 VSS.n1925 VSS.n1923 4.5005
R4030 VSS.n1951 VSS.n1950 4.5005
R4031 VSS.n1960 VSS.n1959 4.5005
R4032 VSS.n1847 VSS.n1846 4.5005
R4033 VSS.n249 VSS.n248 4.5005
R4034 VSS.n252 VSS.n251 4.5005
R4035 VSS.n253 VSS.n238 4.5005
R4036 VSS.n1747 VSS.n1746 4.5005
R4037 VSS.n1752 VSS.n1751 4.5005
R4038 VSS.n1736 VSS.n1732 4.5005
R4039 VSS.n1766 VSS.n1763 4.5005
R4040 VSS.n1770 VSS.n1769 4.5005
R4041 VSS.n501 VSS.n500 4.5005
R4042 VSS.n1812 VSS.n1811 4.5005
R4043 VSS.n1727 VSS.n1718 4.5005
R4044 VSS.n1818 VSS.n1817 4.5005
R4045 VSS.n1873 VSS.n1872 4.5005
R4046 VSS.n1707 VSS.n1706 4.5005
R4047 VSS.n269 VSS.n266 4.5005
R4048 VSS.n2951 VSS.n2950 4.5005
R4049 VSS.n2941 VSS.n270 4.5005
R4050 VSS.n1889 VSS.n1888 4.4805
R4051 VSS.n2199 VSS.n2198 4.38311
R4052 VSS.n1126 VSS.n1078 4.36875
R4053 VSS.n1127 VSS.n1072 4.36875
R4054 VSS.n1141 VSS.n1071 4.36875
R4055 VSS.n1150 VSS.n1149 4.36875
R4056 VSS.n1191 VSS.n1190 4.36875
R4057 VSS.n1178 VSS.n1177 4.36875
R4058 VSS.n2899 VSS.n2898 4.36875
R4059 VSS.n2879 VSS.n516 4.36875
R4060 VSS.n2868 VSS.n519 4.36875
R4061 VSS.n1653 VSS.n1633 4.36875
R4062 VSS.n2722 VSS.n2721 4.36875
R4063 VSS.n2723 VSS.n577 4.36875
R4064 VSS.n2741 VSS.n576 4.36875
R4065 VSS.n2750 VSS.n2749 4.36875
R4066 VSS.n2789 VSS.n2788 4.36875
R4067 VSS.n2795 VSS.n553 4.36875
R4068 VSS.n2811 VSS.n2810 4.36875
R4069 VSS.n2824 VSS.n2823 4.36875
R4070 VSS.n2830 VSS.n542 4.36875
R4071 VSS.n2670 VSS.n2669 4.36875
R4072 VSS.n634 VSS.n624 4.36875
R4073 VSS.n2656 VSS.n2655 4.36875
R4074 VSS.n2648 VSS.n639 4.36875
R4075 VSS.n2627 VSS.n2626 4.36875
R4076 VSS.n2614 VSS.n2613 4.36875
R4077 VSS.n942 VSS.n941 4.36875
R4078 VSS.n962 VSS.n961 4.36875
R4079 VSS.n2306 VSS.n2305 4.28986
R4080 VSS.n2310 VSS.n839 4.28986
R4081 VSS.n2500 VSS.n2499 4.28986
R4082 VSS.n1296 VSS.n1295 4.28986
R4083 VSS.n1352 VSS.n1309 4.28986
R4084 VSS.n1329 VSS.n1328 4.28986
R4085 VSS.n1965 VSS.n1964 4.28986
R4086 VSS.n2330 VSS.n2329 4.14168
R4087 VSS.n1041 VSS.n1040 4.11798
R4088 VSS.n1040 VSS.n1039 4.11798
R4089 VSS.n2544 VSS.n2543 4.11798
R4090 VSS.n1424 VSS.n1423 4.11798
R4091 VSS.n1425 VSS.n1424 4.11798
R4092 VSS.n1458 VSS.n1457 4.11798
R4093 VSS.n1457 VSS.n1362 4.11798
R4094 VSS.n2099 VSS.n2098 4.11798
R4095 VSS.n1849 VSS.n1845 4.11798
R4096 VSS.n1864 VSS.n1849 4.11798
R4097 VSS.n2915 VSS.n497 4.11798
R4098 VSS.n2918 VSS.n497 4.11798
R4099 VSS.n1785 VSS.n1784 4.11798
R4100 VSS.n1784 VSS.n1783 4.11798
R4101 VSS.n2936 VSS.n275 4.11798
R4102 VSS.n2933 VSS.n275 4.11798
R4103 VSS.n1059 VSS.n1058 4.09013
R4104 VSS.n2499 VSS.n2498 4.07323
R4105 VSS.n1295 VSS.n1213 4.07323
R4106 VSS.n1340 VSS.n1309 4.07323
R4107 VSS.n1328 VSS.n1327 4.07323
R4108 VSS.n1964 VSS.n1963 4.07323
R4109 VSS.n1671 VSS.n1668 4.03876
R4110 VSS.n745 VSS.n744 4.03876
R4111 VSS.n2992 VSS 4.02175
R4112 VSS.n230 VSS 4.02175
R4113 VSS.n3321 VSS 4.02175
R4114 VSS.n231 VSS 4.02175
R4115 VSS.n1207 VSS.n1066 3.97459
R4116 VSS.n2644 VSS.n2643 3.97459
R4117 VSS.n1113 VSS.n1112 3.96548
R4118 VSS.n1114 VSS.n1113 3.96548
R4119 VSS.n1682 VSS.n1681 3.96548
R4120 VSS.n2713 VSS.n2712 3.96548
R4121 VSS.n2716 VSS.n2713 3.96548
R4122 VSS.n2842 VSS.n540 3.96548
R4123 VSS.n1003 VSS.n1002 3.96548
R4124 VSS.n1018 VSS.n1003 3.96548
R4125 VSS.n1016 VSS.n1015 3.96548
R4126 VSS.n2677 VSS.n2676 3.96548
R4127 VSS.n2676 VSS.n2675 3.96548
R4128 VSS.n740 VSS.n739 3.96548
R4129 VSS.n1414 VSS.n1413 3.96548
R4130 VSS.n1415 VSS.n1414 3.96548
R4131 VSS.n780 VSS.n778 3.90948
R4132 VSS.n780 VSS.n779 3.90948
R4133 VSS.n390 VSS.n389 3.78485
R4134 VSS.n3180 VSS.n3178 3.78485
R4135 VSS.n3210 VSS.n3199 3.78485
R4136 VSS.n3162 VSS.n3161 3.78485
R4137 VSS.n3157 VSS.n3156 3.78485
R4138 VSS.n3138 VSS.n182 3.78485
R4139 VSS.n3324 VSS.n77 3.78485
R4140 VSS.n3214 VSS.n3194 3.78485
R4141 VSS.n2542 VSS.n2541 3.75994
R4142 VSS.n412 VSS.n409 3.75517
R4143 VSS.n1112 VSS.n1082 3.7069
R4144 VSS.n1683 VSS.n1682 3.7069
R4145 VSS.n2712 VSS.n590 3.7069
R4146 VSS.n2837 VSS.n540 3.7069
R4147 VSS.n2759 VSS.n570 3.7069
R4148 VSS.n2760 VSS.n2759 3.7069
R4149 VSS.n1002 VSS.n996 3.7069
R4150 VSS.n1012 VSS.n1011 3.7069
R4151 VSS.n2677 VSS.n617 3.7069
R4152 VSS.n740 VSS.n729 3.7069
R4153 VSS.n1413 VSS.n1381 3.7069
R4154 VSS.n1415 VSS.n1379 3.7069
R4155 VSS.n2316 VSS.n836 3.50735
R4156 VSS.n1979 VSS.n1978 3.50735
R4157 VSS.n1824 VSS.n1823 3.50735
R4158 VSS.n2964 VSS.n261 3.50735
R4159 VSS.n490 VSS.n401 3.46461
R4160 VSS.n422 VSS.n401 3.46461
R4161 VSS.t88 VSS.t138 3.46461
R4162 VSS.t88 VSS.t86 3.46461
R4163 VSS.n424 VSS.n420 3.46461
R4164 VSS.n469 VSS.n424 3.46461
R4165 VSS.n2185 VSS.n2184 3.44377
R4166 VSS.n2184 VSS.n2183 3.44377
R4167 VSS.n1953 VSS.n1952 3.43942
R4168 VSS.n749 VSS.n748 3.43925
R4169 VSS.n2523 VSS.n2522 3.43925
R4170 VSS.n2894 VSS.n505 3.43925
R4171 VSS.n2905 VSS.n2904 3.43925
R4172 VSS.n1195 VSS.n1194 3.43925
R4173 VSS.n1197 VSS.n1158 3.43925
R4174 VSS.n1134 VSS.n1133 3.43925
R4175 VSS.n1123 VSS.n1122 3.43925
R4176 VSS.n1691 VSS.n1556 3.43925
R4177 VSS.n1701 VSS.n1700 3.43925
R4178 VSS.n1643 VSS.n527 3.43925
R4179 VSS.n2861 VSS.n523 3.43925
R4180 VSS.n2734 VSS.n2733 3.43925
R4181 VSS.n2731 VSS.n2730 3.43925
R4182 VSS.n2704 VSS.n2703 3.43925
R4183 VSS.n2701 VSS.n2700 3.43925
R4184 VSS.n1613 VSS.n1557 3.43925
R4185 VSS.n1622 VSS.n1621 3.43925
R4186 VSS.n2818 VSS.n2817 3.43925
R4187 VSS.n2805 VSS.n2804 3.43925
R4188 VSS.n2774 VSS.n2773 3.43925
R4189 VSS.n2771 VSS.n2770 3.43925
R4190 VSS.n535 VSS.n528 3.43925
R4191 VSS.n2858 VSS.n2857 3.43925
R4192 VSS.n2661 VSS.n2660 3.43925
R4193 VSS.n2663 VSS.n626 3.43925
R4194 VSS.n613 VSS.n598 3.43925
R4195 VSS.n2687 VSS.n2686 3.43925
R4196 VSS.n1022 VSS.n1021 3.43925
R4197 VSS.n1026 VSS.n1025 3.43925
R4198 VSS.n949 VSS.n665 3.43925
R4199 VSS.n2607 VSS.n2606 3.43925
R4200 VSS.n2631 VSS.n2630 3.43925
R4201 VSS.n2633 VSS.n647 3.43925
R4202 VSS.n1050 VSS.n1049 3.43925
R4203 VSS.n1052 VSS.n969 3.43925
R4204 VSS.n2461 VSS.n2460 3.43925
R4205 VSS.n2458 VSS.n2457 3.43925
R4206 VSS.n2220 VSS.n2219 3.43925
R4207 VSS.n2224 VSS.n2223 3.43925
R4208 VSS.n1987 VSS.n1986 3.43925
R4209 VSS.n1989 VSS.n1902 3.43925
R4210 VSS.n1515 VSS.n1514 3.43925
R4211 VSS.n1473 VSS.n1472 3.43925
R4212 VSS.n1444 VSS.n1443 3.43925
R4213 VSS.n1430 VSS.n1429 3.43925
R4214 VSS.n2593 VSS.n666 3.43925
R4215 VSS.n2603 VSS.n2602 3.43925
R4216 VSS.n2107 VSS.n2106 3.43925
R4217 VSS.n2104 VSS.n2103 3.43925
R4218 VSS.n2017 VSS.n913 3.43925
R4219 VSS.n2027 VSS.n2026 3.43925
R4220 VSS.n2340 VSS.n2339 3.43925
R4221 VSS.n2337 VSS.n2336 3.43925
R4222 VSS.n857 VSS.n856 3.43925
R4223 VSS.n2298 VSS.n2297 3.43925
R4224 VSS.n2508 VSS.n750 3.43925
R4225 VSS.n2519 VSS.n2518 3.43925
R4226 VSS.n2387 VSS.n2386 3.43925
R4227 VSS.n2384 VSS.n2383 3.43925
R4228 VSS.n1344 VSS.n1343 3.43925
R4229 VSS.n1346 VSS.n1311 3.43925
R4230 VSS.n2189 VSS.n2188 3.43925
R4231 VSS.n2193 VSS.n2192 3.43925
R4232 VSS.n2262 VSS.n2261 3.43925
R4233 VSS.n2258 VSS.n2257 3.43925
R4234 VSS.n1288 VSS.n1287 3.43925
R4235 VSS.n1285 VSS.n1284 3.43925
R4236 VSS.n2983 VSS.n2982 3.41839
R4237 VSS.n243 VSS.n242 3.41839
R4238 VSS.n2944 VSS.n2943 3.41636
R4239 VSS.n2955 VSS.n2954 3.41636
R4240 VSS.n1796 VSS.n1795 3.41624
R4241 VSS.n1737 VSS.n1730 3.41624
R4242 VSS.n2909 VSS.n2908 3.41605
R4243 VSS.n1765 VSS.n504 3.41605
R4244 VSS.n1404 VSS.n1403 3.41514
R4245 VSS.n1104 VSS.n1103 3.41514
R4246 VSS.n874 VSS.n858 3.41514
R4247 VSS.n250 VSS.n235 3.4105
R4248 VSS.n2984 VSS.n236 3.4105
R4249 VSS.n1749 VSS.n1748 3.4105
R4250 VSS.n1750 VSS.n1731 3.4105
R4251 VSS.n1767 VSS.n1728 3.4105
R4252 VSS.n1768 VSS.n502 3.4105
R4253 VSS.n1395 VSS.n1394 3.4105
R4254 VSS.n1385 VSS.n1384 3.4105
R4255 VSS.n1402 VSS.n1401 3.4105
R4256 VSS.n721 VSS.n712 3.4105
R4257 VSS.n722 VSS.n714 3.4105
R4258 VSS.n509 VSS.n507 3.4105
R4259 VSS.n2893 VSS.n2892 3.4105
R4260 VSS.n1199 VSS.n1198 3.4105
R4261 VSS.n1196 VSS.n1160 3.4105
R4262 VSS.n1076 VSS.n1075 3.4105
R4263 VSS.n1132 VSS.n1131 3.4105
R4264 VSS.n1093 VSS.n1092 3.4105
R4265 VSS.n1089 VSS.n1088 3.4105
R4266 VSS.n1102 VSS.n1101 3.4105
R4267 VSS.n1626 VSS.n1624 3.4105
R4268 VSS.n1689 VSS.n1688 3.4105
R4269 VSS.n2863 VSS.n2862 3.4105
R4270 VSS.n1639 VSS.n525 3.4105
R4271 VSS.n585 VSS.n583 3.4105
R4272 VSS.n2725 VSS.n580 3.4105
R4273 VSS.n2691 VSS.n2689 3.4105
R4274 VSS.n2694 VSS.n596 3.4105
R4275 VSS.n1560 VSS.n1558 3.4105
R4276 VSS.n1611 VSS.n1610 3.4105
R4277 VSS.n550 VSS.n549 3.4105
R4278 VSS.n2816 VSS.n2815 3.4105
R4279 VSS.n569 VSS.n567 3.4105
R4280 VSS.n2763 VSS.n564 3.4105
R4281 VSS.n532 VSS.n530 3.4105
R4282 VSS.n2852 VSS.n2851 3.4105
R4283 VSS.n2665 VSS.n2664 3.4105
R4284 VSS.n2662 VSS.n628 3.4105
R4285 VSS.n602 VSS.n600 3.4105
R4286 VSS.n610 VSS.n609 3.4105
R4287 VSS.n1024 VSS.n991 3.4105
R4288 VSS.n1023 VSS.n992 3.4105
R4289 VSS.n937 VSS.n664 3.4105
R4290 VSS.n947 VSS.n946 3.4105
R4291 VSS.n2635 VSS.n2634 3.4105
R4292 VSS.n2632 VSS.n649 3.4105
R4293 VSS.n1054 VSS.n1053 3.4105
R4294 VSS.n1051 VSS.n971 3.4105
R4295 VSS.n773 VSS.n771 3.4105
R4296 VSS.n2452 VSS.n769 3.4105
R4297 VSS.n2222 VSS.n2127 3.4105
R4298 VSS.n2221 VSS.n2128 3.4105
R4299 VSS.n1991 VSS.n1990 3.4105
R4300 VSS.n1905 VSS.n1904 3.4105
R4301 VSS.n2550 VSS.n689 3.4105
R4302 VSS.n2562 VSS.n689 3.4105
R4303 VSS.n2551 VSS.n2550 3.4105
R4304 VSS.n2563 VSS.n2562 3.4105
R4305 VSS.n2561 VSS.n2560 3.4105
R4306 VSS.n2549 VSS.n691 3.4105
R4307 VSS.n1474 VSS.n1468 3.4105
R4308 VSS.n1517 VSS.n1516 3.4105
R4309 VSS.n1371 VSS.n1370 3.4105
R4310 VSS.n1442 VSS.n1441 3.4105
R4311 VSS.n670 VSS.n668 3.4105
R4312 VSS.n2592 VSS.n2591 3.4105
R4313 VSS.n2031 VSS.n2029 3.4105
R4314 VSS.n2033 VSS.n912 3.4105
R4315 VSS.n916 VSS.n914 3.4105
R4316 VSS.n923 VSS.n922 3.4105
R4317 VSS.n2424 VSS.n667 3.4105
R4318 VSS.n786 VSS.n667 3.4105
R4319 VSS.n2425 VSS.n2424 3.4105
R4320 VSS.n787 VSS.n786 3.4105
R4321 VSS.n2421 VSS.n2420 3.4105
R4322 VSS.n2423 VSS.n785 3.4105
R4323 VSS.n830 VSS.n828 3.4105
R4324 VSS.n825 VSS.n824 3.4105
R4325 VSS.n849 VSS.n847 3.4105
R4326 VSS.n852 VSS.n848 3.4105
R4327 VSS.n754 VSS.n752 3.4105
R4328 VSS.n2506 VSS.n2505 3.4105
R4329 VSS.n806 VSS.n803 3.4105
R4330 VSS.n800 VSS.n799 3.4105
R4331 VSS.n1348 VSS.n1347 3.4105
R4332 VSS.n1314 VSS.n1313 3.4105
R4333 VSS.n2071 VSS.n802 3.4105
R4334 VSS.n2059 VSS.n802 3.4105
R4335 VSS.n2072 VSS.n2071 3.4105
R4336 VSS.n2060 VSS.n2059 3.4105
R4337 VSS.n2058 VSS.n2051 3.4105
R4338 VSS.n2070 VSS.n2069 3.4105
R4339 VSS.n2293 VSS.n2292 3.4105
R4340 VSS.n863 VSS.n860 3.4105
R4341 VSS.n871 VSS.n870 3.4105
R4342 VSS.n2191 VSS.n2154 3.4105
R4343 VSS.n2190 VSS.n2155 3.4105
R4344 VSS.n2259 VSS.n2254 3.4105
R4345 VSS.n2260 VSS.n893 3.4105
R4346 VSS.n1220 VSS.n1218 3.4105
R4347 VSS.n1279 VSS.n1217 3.4105
R4348 VSS.n1247 VSS.n859 3.4105
R4349 VSS.n1233 VSS.n859 3.4105
R4350 VSS.n1248 VSS.n1247 3.4105
R4351 VSS.n1234 VSS.n1233 3.4105
R4352 VSS.n1244 VSS.n1243 3.4105
R4353 VSS.n1246 VSS.n1232 3.4105
R4354 VSS.n1948 VSS.n1947 3.4105
R4355 VSS.n1924 VSS.n1922 3.4105
R4356 VSS.n1958 VSS.n1957 3.4105
R4357 VSS.n1955 VSS.n1948 3.4105
R4358 VSS.n1957 VSS.n1956 3.4105
R4359 VSS.n1875 VSS.n1874 3.4105
R4360 VSS.n2953 VSS.n2952 3.4105
R4361 VSS.n2942 VSS.n268 3.4105
R4362 VSS.n1819 VSS.n1549 3.4105
R4363 VSS.n1805 VSS.n1726 3.4105
R4364 VSS.n1810 VSS.n1809 3.4105
R4365 VSS.n1808 VSS.n1717 3.4105
R4366 VSS.n1875 VSS.n1552 3.4105
R4367 VSS.n1875 VSS.n1551 3.4105
R4368 VSS.n1875 VSS.n1550 3.4105
R4369 VSS.n30 VSS.n29 3.40476
R4370 VSS.n3287 VSS.n3286 3.40476
R4371 VSS.n704 VSS.n701 3.31239
R4372 VSS.n2098 VSS.n2097 3.22288
R4373 VSS.n2185 VSS.n2171 3.21921
R4374 VSS.n2180 VSS.n2179 3.21921
R4375 VSS.n2318 VSS.n834 3.2005
R4376 VSS.n1983 VSS.n1911 3.2005
R4377 VSS.n1828 VSS.n1714 3.2005
R4378 VSS.n2963 VSS.n262 3.2005
R4379 VSS.n57 VSS.n56 3.13241
R4380 VSS.n3379 VSS.n3375 3.13241
R4381 VSS.n29 VSS.n25 3.13241
R4382 VSS.n10 VSS.n9 3.13241
R4383 VSS.n3242 VSS.n3241 3.13241
R4384 VSS.n102 VSS.n98 3.13241
R4385 VSS.n3261 VSS.n3260 3.13241
R4386 VSS.n3286 VSS.n3285 3.13241
R4387 VSS.n1602 VSS.n1593 3.13241
R4388 VSS.n2579 VSS.n2578 3.13241
R4389 VSS.n1268 VSS.n1267 3.13241
R4390 VSS.n2010 VSS.n925 3.13241
R4391 VSS.n1546 VSS.n1545 3.1005
R4392 VSS.n2766 VSS.n561 3.09945
R4393 VSS.n1151 VSS.n1066 3.05276
R4394 VSS.n2645 VSS.n2644 3.05276
R4395 VSS.n1677 VSS.n1676 3.04861
R4396 VSS.n1108 VSS.n1106 3.04861
R4397 VSS.n1598 VSS.n1596 3.04861
R4398 VSS.n2708 VSS.n2706 3.04861
R4399 VSS.n1009 VSS.n1007 3.04861
R4400 VSS.n2681 VSS.n615 3.04861
R4401 VSS.n734 VSS.n733 3.04861
R4402 VSS.n2497 VSS.n2496 3.04861
R4403 VSS.n2177 VSS.n2176 3.04861
R4404 VSS.n1298 VSS.n1213 3.04861
R4405 VSS.n1327 VSS.n1326 3.04861
R4406 VSS.n2240 VSS.n898 3.01226
R4407 VSS.n2363 VSS.n2362 2.92224
R4408 VSS.n1058 VSS.n966 2.92166
R4409 VSS.n3407 VSS.n3406 2.90519
R4410 VSS.n3010 VSS.t774 2.89674
R4411 VSS.n1114 VSS.n1080 2.88804
R4412 VSS.n2716 VSS.n2715 2.88804
R4413 VSS.n2675 VSS.n620 2.88804
R4414 VSS.n3073 VSS.n3072 2.88636
R4415 VSS.n31 VSS.n30 2.86007
R4416 VSS.n3288 VSS.n3287 2.86007
R4417 VSS.n1080 VSS.n1079 2.79323
R4418 VSS.n2715 VSS.n2714 2.79323
R4419 VSS.n620 VSS.n619 2.79323
R4420 VSS.n1684 VSS.n1671 2.77203
R4421 VSS.n744 VSS.n743 2.77203
R4422 VSS.n58 VSS.n57 2.7239
R4423 VSS.n3376 VSS.n3375 2.7239
R4424 VSS.n26 VSS.n25 2.7239
R4425 VSS.n9 VSS.n8 2.7239
R4426 VSS.n3241 VSS.n81 2.7239
R4427 VSS.n99 VSS.n98 2.7239
R4428 VSS.n3262 VSS.n3261 2.7239
R4429 VSS.n3285 VSS.n3284 2.7239
R4430 VSS.n1594 VSS.n1593 2.7239
R4431 VSS.n2578 VSS.n2577 2.7239
R4432 VSS.n878 VSS.n877 2.7239
R4433 VSS.n1269 VSS.n1268 2.7239
R4434 VSS.n926 VSS.n925 2.7239
R4435 VSS.n2545 VSS.n699 2.68581
R4436 VSS.n3406 VSS.n3405 2.63717
R4437 VSS.n3237 VSS.n3236 2.63717
R4438 VSS.n2321 VSS.n2320 2.63064
R4439 VSS.n1982 VSS.n1977 2.63064
R4440 VSS.n1827 VSS.n1712 2.63064
R4441 VSS.n2961 VSS.n2960 2.63064
R4442 VSS.n3347 VSS.n3346 2.59858
R4443 VSS VSS.n229 2.56738
R4444 VSS.n2779 VSS.n2778 2.55412
R4445 VSS.n1658 VSS.n1657 2.50679
R4446 VSS.n2570 VSS.n683 2.50679
R4447 VSS.n2082 VSS.n2041 2.50679
R4448 VSS.n1060 VSS.n1059 2.38348
R4449 VSS.n1144 VSS.n1143 2.33701
R4450 VSS.n1143 VSS.n1069 2.33701
R4451 VSS.n1184 VSS.n1183 2.33701
R4452 VSS.n1183 VSS.n1182 2.33701
R4453 VSS.n1172 VSS.n1170 2.33701
R4454 VSS.n1178 VSS.n1172 2.33701
R4455 VSS.n2885 VSS.n514 2.33701
R4456 VSS.n2882 VSS.n514 2.33701
R4457 VSS.n2881 VSS.n2880 2.33701
R4458 VSS.n2880 VSS.n2879 2.33701
R4459 VSS.n1648 VSS.n1635 2.33701
R4460 VSS.n1651 VSS.n1635 2.33701
R4461 VSS.n2744 VSS.n2743 2.33701
R4462 VSS.n2743 VSS.n574 2.33701
R4463 VSS.n2790 VSS.n555 2.33701
R4464 VSS.n2793 VSS.n555 2.33701
R4465 VSS.n2808 VSS.n552 2.33701
R4466 VSS.n2825 VSS.n544 2.33701
R4467 VSS.n2828 VSS.n544 2.33701
R4468 VSS.n638 VSS.n636 2.33701
R4469 VSS.n2650 VSS.n638 2.33701
R4470 VSS.n2620 VSS.n2619 2.33701
R4471 VSS.n2619 VSS.n2618 2.33701
R4472 VSS.n661 VSS.n659 2.33701
R4473 VSS.n2614 VSS.n661 2.33701
R4474 VSS.n955 VSS.n933 2.33701
R4475 VSS.n958 VSS.n933 2.33701
R4476 VSS.n960 VSS.n959 2.33701
R4477 VSS.n962 VSS.n960 2.33701
R4478 VSS.n2783 VSS.n559 2.33067
R4479 VSS.n295 VSS.n288 2.3255
R4480 VSS.n301 VSS.n287 2.3255
R4481 VSS.n327 VSS.n326 2.3255
R4482 VSS.n332 VSS.n331 2.3255
R4483 VSS.n375 VSS.n374 2.3255
R4484 VSS.n352 VSS.n351 2.3255
R4485 VSS.n349 VSS.n345 2.3255
R4486 VSS.n201 VSS.n200 2.3255
R4487 VSS.n3027 VSS.n3026 2.25932
R4488 VSS.n3067 VSS.n3037 2.25932
R4489 VSS.n1617 VSS.n1589 2.25932
R4490 VSS.n1505 VSS.n1482 2.25932
R4491 VSS.n2349 VSS.n2348 2.25932
R4492 VSS.n2374 VSS.n2373 2.25932
R4493 VSS.n2379 VSS.n2378 2.25932
R4494 VSS.n2378 VSS.n797 2.25932
R4495 VSS.n2466 VSS.n763 2.25932
R4496 VSS.n2278 VSS.n882 2.25932
R4497 VSS.n2240 VSS.n2239 2.25932
R4498 VSS.n2142 VSS.n2141 2.25932
R4499 VSS.n1117 VSS.n1116 2.25312
R4500 VSS.n2718 VSS.n588 2.25312
R4501 VSS.n2673 VSS.n621 2.25312
R4502 VSS.n2440 VSS.n780 2.25293
R4503 VSS.n2989 VSS.n2988 2.23999
R4504 VSS.n1118 VSS.n1117 2.2228
R4505 VSS.n588 VSS.n587 2.2228
R4506 VSS.n623 VSS.n621 2.2228
R4507 VSS.n877 VSS.n876 2.17922
R4508 VSS.n3234 VSS.n3233 2.14347
R4509 VSS.n2305 VSS.n2304 2.13383
R4510 VSS.n1156 VSS.n1155 2.11085
R4511 VSS.n645 VSS.n644 2.11085
R4512 VSS.n1015 VSS.n1004 2.06919
R4513 VSS.n3006 VSS.n3005 2.03479
R4514 VSS.n2799 VSS.n552 2.03225
R4515 VSS.n1681 VSS.n1672 1.98299
R4516 VSS.n2843 VSS.n2842 1.98299
R4517 VSS.n1018 VSS.n1017 1.98299
R4518 VSS.n1017 VSS.n1016 1.98299
R4519 VSS.n739 VSS.n738 1.98299
R4520 VSS.n2161 VSS.n2151 1.97497
R4521 VSS VSS.n3431 1.92557
R4522 VSS.n2782 VSS.n560 1.91571
R4523 VSS.n1012 VSS.n1004 1.8968
R4524 VSS.n2513 VSS.n2512 1.88285
R4525 VSS.n2362 VSS.n2361 1.87876
R4526 VSS.n2183 VSS.n2172 1.79699
R4527 VSS.n3007 VSS.n3006 1.77326
R4528 VSS.n2535 VSS.n2534 1.75824
R4529 VSS.n3374 VSS.n3373 1.753
R4530 VSS.n3372 VSS.n3371 1.753
R4531 VSS.n3105 VSS.n3104 1.753
R4532 VSS.n3103 VSS.n3102 1.753
R4533 VSS.n96 VSS.n79 1.753
R4534 VSS.n3319 VSS.n3318 1.753
R4535 VSS.n2358 VSS.n2357 1.7528
R4536 VSS.n1673 VSS.n1672 1.72441
R4537 VSS.n2844 VSS.n2843 1.72441
R4538 VSS.n738 VSS.n737 1.72441
R4539 VSS.n1954 VSS.n1953 1.72315
R4540 VSS.n1807 VSS.n526 1.70468
R4541 VSS.n1806 VSS.n526 1.70468
R4542 VSS.n2295 VSS.n858 1.70393
R4543 VSS.n2295 VSS.n2294 1.70393
R4544 VSS.n1403 VSS.n599 1.70393
R4545 VSS.n1393 VSS.n599 1.70393
R4546 VSS.n1103 VSS.n597 1.70393
R4547 VSS.n1091 VSS.n597 1.70393
R4548 VSS.n2908 VSS.n2907 1.70348
R4549 VSS.n2907 VSS.n504 1.70348
R4550 VSS.n1797 VSS.n1796 1.70338
R4551 VSS.n1797 VSS.n1730 1.70338
R4552 VSS.n2943 VSS.n267 1.70332
R4553 VSS.n2954 VSS.n267 1.70332
R4554 VSS.n2983 VSS.n237 1.70231
R4555 VSS.n242 VSS.n237 1.70231
R4556 VSS.n745 VSS.n728 1.7012
R4557 VSS.n1988 VSS.n1987 1.69188
R4558 VSS.n1989 VSS.n1988 1.69188
R4559 VSS.n2220 VSS.n770 1.69188
R4560 VSS.n2223 VSS.n770 1.69188
R4561 VSS.n2460 VSS.n2459 1.69188
R4562 VSS.n2459 VSS.n2458 1.69188
R4563 VSS.n1050 VSS.n529 1.69188
R4564 VSS.n1052 VSS.n529 1.69188
R4565 VSS.n2859 VSS.n528 1.69188
R4566 VSS.n2859 VSS.n2858 1.69188
R4567 VSS.n2860 VSS.n527 1.69188
R4568 VSS.n2861 VSS.n2860 1.69188
R4569 VSS.n690 VSS.n689 1.69188
R4570 VSS.n2028 VSS.n913 1.69188
R4571 VSS.n2028 VSS.n2027 1.69188
R4572 VSS.n2106 VSS.n2105 1.69188
R4573 VSS.n2105 VSS.n2104 1.69188
R4574 VSS.n2604 VSS.n666 1.69188
R4575 VSS.n2604 VSS.n2603 1.69188
R4576 VSS.n2605 VSS.n665 1.69188
R4577 VSS.n2606 VSS.n2605 1.69188
R4578 VSS.n2817 VSS.n506 1.69188
R4579 VSS.n2804 VSS.n506 1.69188
R4580 VSS.n2906 VSS.n505 1.69188
R4581 VSS.n2906 VSS.n2905 1.69188
R4582 VSS.n2422 VSS.n667 1.69188
R4583 VSS.n1345 VSS.n1344 1.69188
R4584 VSS.n1346 VSS.n1345 1.69188
R4585 VSS.n2386 VSS.n2385 1.69188
R4586 VSS.n2385 VSS.n2384 1.69188
R4587 VSS.n1515 VSS.n801 1.69188
R4588 VSS.n1473 VSS.n801 1.69188
R4589 VSS.n2631 VSS.n566 1.69188
R4590 VSS.n2633 VSS.n566 1.69188
R4591 VSS.n2773 VSS.n2772 1.69188
R4592 VSS.n2772 VSS.n2771 1.69188
R4593 VSS.n1195 VSS.n565 1.69188
R4594 VSS.n1197 VSS.n565 1.69188
R4595 VSS.n2050 VSS.n802 1.69188
R4596 VSS.n1287 VSS.n1286 1.69188
R4597 VSS.n1286 VSS.n1285 1.69188
R4598 VSS.n2261 VSS.n827 1.69188
R4599 VSS.n2258 VSS.n827 1.69188
R4600 VSS.n2339 VSS.n2338 1.69188
R4601 VSS.n2338 VSS.n2337 1.69188
R4602 VSS.n1443 VSS.n826 1.69188
R4603 VSS.n1429 VSS.n826 1.69188
R4604 VSS.n2661 VSS.n582 1.69188
R4605 VSS.n2663 VSS.n582 1.69188
R4606 VSS.n2733 VSS.n2732 1.69188
R4607 VSS.n2732 VSS.n2731 1.69188
R4608 VSS.n1133 VSS.n581 1.69188
R4609 VSS.n1122 VSS.n581 1.69188
R4610 VSS.n2296 VSS.n857 1.69188
R4611 VSS.n2297 VSS.n2296 1.69188
R4612 VSS.n2688 VSS.n598 1.69188
R4613 VSS.n2688 VSS.n2687 1.69188
R4614 VSS.n2703 VSS.n2702 1.69188
R4615 VSS.n2702 VSS.n2701 1.69188
R4616 VSS.n1245 VSS.n859 1.69188
R4617 VSS.n2189 VSS.n751 1.69188
R4618 VSS.n2192 VSS.n751 1.69188
R4619 VSS.n2520 VSS.n750 1.69188
R4620 VSS.n2520 VSS.n2519 1.69188
R4621 VSS.n2521 VSS.n749 1.69188
R4622 VSS.n2522 VSS.n2521 1.69188
R4623 VSS.n1022 VSS.n713 1.69188
R4624 VSS.n1025 VSS.n713 1.69188
R4625 VSS.n1623 VSS.n1557 1.69188
R4626 VSS.n1623 VSS.n1622 1.69188
R4627 VSS.n1702 VSS.n1556 1.69188
R4628 VSS.n1702 VSS.n1701 1.69188
R4629 VSS.n2180 VSS.n2172 1.64728
R4630 VSS.n2555 VSS.n2554 1.61169
R4631 VSS.n3340 VSS 1.54822
R4632 VSS.n3099 VSS.n3085 1.50638
R4633 VSS.n3093 VSS.n3087 1.50638
R4634 VSS.n191 VSS.n189 1.50638
R4635 VSS.n3121 VSS.n192 1.50638
R4636 VSS.n3035 VSS.n3034 1.50638
R4637 VSS.n3036 VSS.n3035 1.50638
R4638 VSS.n3064 VSS.n3063 1.50638
R4639 VSS.n3057 VSS.n3040 1.50638
R4640 VSS.n3057 VSS.n3056 1.50638
R4641 VSS.n3048 VSS.n3047 1.50638
R4642 VSS.n2835 VSS.n2834 1.47352
R4643 VSS.n3006 VSS.n2993 1.44312
R4644 VSS.n2751 VSS.n571 1.34658
R4645 VSS.n2991 VSS.n229 1.3415
R4646 VSS.n1059 VSS.n965 1.3283
R4647 VSS.n2990 VSS.n2989 1.31337
R4648 VSS.n1119 VSS.n1118 1.29527
R4649 VSS.n2720 VSS.n587 1.29527
R4650 VSS.n2671 VSS.n623 1.29527
R4651 VSS.n1695 VSS.n1694 1.25365
R4652 VSS.n2756 VSS.n2755 1.25033
R4653 VSS.n17 VSS.n1 1.21169
R4654 VSS.n3072 VSS.n3071 1.21169
R4655 VSS.n3235 VSS.n111 1.21169
R4656 VSS.n1410 VSS.n1409 1.20723
R4657 VSS.n2361 VSS.n812 1.18311
R4658 VSS.n2229 VSS.n2228 1.18311
R4659 VSS.n2198 VSS.n2197 1.18311
R4660 VSS.n1237 VSS.n1236 1.18311
R4661 VSS.n1933 VSS.n1932 1.18311
R4662 VSS.n1854 VSS.n1853 1.18311
R4663 VSS.n1741 VSS.n1740 1.18311
R4664 VSS.n2976 VSS.n2975 1.18311
R4665 VSS.n246 VSS.n245 1.18311
R4666 VSS.n450 VSS.n409 1.15795
R4667 VSS.n2320 VSS.n834 1.14023
R4668 VSS.n1983 VSS.n1982 1.14023
R4669 VSS.n1828 VSS.n1827 1.14023
R4670 VSS.n2961 VSS.n262 1.14023
R4671 VSS.n2397 VSS.n2396 1.12991
R4672 VSS.n2838 VSS.n2836 1.12954
R4673 VSS.n1799 VSS 1.12383
R4674 VSS.n1798 VSS 1.11689
R4675 VSS.n2989 VSS.n232 1.11056
R4676 VSS.n1555 VSS 1.10328
R4677 VSS.n1553 VSS 1.07702
R4678 VSS.n2529 VSS.n2528 1.07463
R4679 VSS.n2991 VSS.n2990 1.05425
R4680 VSS.n3372 VSS 1.00137
R4681 VSS.n1881 VSS.n1880 0.993972
R4682 VSS.n726 VSS.n718 0.985115
R4683 VSS.n2283 VSS.n876 0.953691
R4684 VSS.n2499 VSS.n2490 0.952566
R4685 VSS.n1295 VSS.n1294 0.952566
R4686 VSS.n1309 VSS.n1308 0.952566
R4687 VSS.n1328 VSS.n1324 0.952566
R4688 VSS.n1964 VSS.n1917 0.952566
R4689 VSS.n472 VSS.n0 0.927421
R4690 VSS.n2498 VSS.n2493 0.899674
R4691 VSS.n2092 VSS.n2037 0.895605
R4692 VSS.n2097 VSS.n909 0.895605
R4693 VSS.n1117 VSS.n1080 0.892621
R4694 VSS.n2715 VSS.n588 0.892621
R4695 VSS.n621 VSS.n620 0.892621
R4696 VSS.n1875 VSS.n1703 0.853
R4697 VSS.n1879 VSS.n1878 0.842928
R4698 VSS.n1978 VSS.n1911 0.833377
R4699 VSS.n1823 VSS.n1714 0.833377
R4700 VSS.n2964 VSS.n2963 0.833377
R4701 VSS.n2783 VSS.n2782 0.830425
R4702 VSS.n3431 VSS.n3430 0.828306
R4703 VSS.n2777 VSS.n561 0.798505
R4704 VSS.n1888 VSS.n1887 0.777453
R4705 VSS.n3373 VSS.n3372 0.761313
R4706 VSS.n3104 VSS.n3103 0.761313
R4707 VSS.n3319 VSS.n79 0.761313
R4708 VSS.n3095 VSS.n3094 0.753441
R4709 VSS.n3089 VSS.n188 0.753441
R4710 VSS.n3123 VSS.n3122 0.753441
R4711 VSS.n3117 VSS.n3116 0.753441
R4712 VSS.n3068 VSS.n3067 0.753441
R4713 VSS.n3061 VSS.n3060 0.753441
R4714 VSS.n3054 VSS.n3053 0.753441
R4715 VSS.n1510 VSS.n1509 0.753441
R4716 VSS.n2352 VSS.n815 0.753441
R4717 VSS.n2480 VSS.n2479 0.753441
R4718 VSS.n1451 VSS.n1450 0.716584
R4719 VSS.n2778 VSS.n559 0.606984
R4720 VSS.n468 VSS.n426 0.577852
R4721 VSS.t419 VSS.t519 0.577852
R4722 VSS.n460 VSS.n438 0.577852
R4723 VSS.n2872 VSS.n518 0.537563
R4724 VSS.n1034 VSS.n986 0.537563
R4725 VSS.n1044 VSS.n979 0.537563
R4726 VSS.n1035 VSS.n985 0.537563
R4727 VSS.n2532 VSS.n705 0.537563
R4728 VSS.n694 VSS.n685 0.537563
R4729 VSS.n2536 VSS.n2535 0.537563
R4730 VSS.n1437 VSS.n1434 0.537563
R4731 VSS.n1436 VSS.n1435 0.537563
R4732 VSS.n1523 VSS.n1461 0.537563
R4733 VSS.n2113 VSS.n2112 0.537563
R4734 VSS.n1838 VSS.n1837 0.537563
R4735 VSS.n1859 VSS.n1850 0.537563
R4736 VSS.n1776 VSS.n1760 0.537563
R4737 VSS.n2923 VSS.n495 0.537563
R4738 VSS.n1755 VSS.n1754 0.537563
R4739 VSS.n1778 VSS.n1777 0.537563
R4740 VSS.n271 VSS.n264 0.537563
R4741 VSS.n2928 VSS.n277 0.537563
R4742 VSS.n1 VSS 0.531208
R4743 VSS.n3072 VSS 0.531208
R4744 VSS.n2313 VSS.n836 0.526527
R4745 VSS.n2317 VSS.n2316 0.526527
R4746 VSS.n1979 VSS.n1899 0.526527
R4747 VSS.n1824 VSS.n1822 0.526527
R4748 VSS.n261 VSS.n259 0.526527
R4749 VSS.n3431 VSS.n3407 0.509828
R4750 VSS.n3321 VSS.n3320 0.482665
R4751 VSS.n2988 VSS.n0 0.473674
R4752 VSS.n329 VSS.n328 0.467019
R4753 VSS.n350 VSS.n228 0.467019
R4754 VSS.n3159 VSS.n3140 0.467019
R4755 VSS.n3212 VSS.n78 0.467019
R4756 VSS.n3233 VSS 0.448179
R4757 VSS.n1660 VSS.n1659 0.448052
R4758 VSS.n1426 VSS.n1375 0.448052
R4759 VSS.n1447 VSS.n1367 0.448052
R4760 VSS.n232 VSS.n210 0.426643
R4761 VSS.n2359 VSS.n2358 0.417891
R4762 VSS.n2366 VSS.n812 0.417891
R4763 VSS.n2233 VSS.n2124 0.417891
R4764 VSS.n2228 VSS.n2227 0.417891
R4765 VSS.n2202 VSS.n2201 0.417891
R4766 VSS.n2200 VSS.n2199 0.417891
R4767 VSS.n2197 VSS.n2196 0.417891
R4768 VSS.n1252 VSS.n1230 0.417891
R4769 VSS.n1937 VSS.n1930 0.417891
R4770 VSS.n1858 VSS.n1851 0.417891
R4771 VSS.n1739 VSS.n278 0.417891
R4772 VSS.n1740 VSS.n1735 0.417891
R4773 VSS.n2979 VSS.n2978 0.417891
R4774 VSS.n2975 VSS.n2974 0.417891
R4775 VSS.n255 VSS.n240 0.417891
R4776 VSS.n1887 VSS.n1546 0.410656
R4777 VSS.n3369 VSS.n58 0.409011
R4778 VSS.n3383 VSS.n40 0.409011
R4779 VSS.n33 VSS.n32 0.409011
R4780 VSS.n3403 VSS.n3 0.409011
R4781 VSS.n7 VSS.n6 0.409011
R4782 VSS.n8 VSS.n4 0.409011
R4783 VSS.n3316 VSS.n81 0.409011
R4784 VSS.n97 VSS.n92 0.409011
R4785 VSS.n3255 VSS.n115 0.409011
R4786 VSS.n3259 VSS.n3258 0.409011
R4787 VSS.n3263 VSS.n3262 0.409011
R4788 VSS.n3291 VSS.n3280 0.409011
R4789 VSS.n1606 VSS.n1605 0.409011
R4790 VSS.n1599 VSS.n1594 0.409011
R4791 VSS.n681 VSS.n678 0.409011
R4792 VSS.n2303 VSS.n2302 0.409011
R4793 VSS.n2312 VSS.n2311 0.409011
R4794 VSS.n2511 VSS.n2486 0.409011
R4795 VSS.n2287 VSS.n868 0.409011
R4796 VSS.n2280 VSS.n878 0.409011
R4797 VSS.n1263 VSS.n1224 0.409011
R4798 VSS.n1270 VSS.n1269 0.409011
R4799 VSS.n1292 VSS.n1291 0.409011
R4800 VSS.n1356 VSS.n1306 0.409011
R4801 VSS.n1323 VSS.n1321 0.409011
R4802 VSS.n2013 VSS.n2012 0.409011
R4803 VSS.n2007 VSS.n926 0.409011
R4804 VSS.n2000 VSS.n1897 0.409011
R4805 VSS.n1916 VSS.n1914 0.409011
R4806 VSS.n1723 VSS.n1719 0.409011
R4807 VSS.n258 VSS.n256 0.409011
R4808 VSS.n2779 VSS.n2777 0.383542
R4809 VSS.n2514 VSS.n2513 0.376971
R4810 VSS.n3408 uio_oe[7] 0.371345
R4811 VSS VSS.n3234 0.366908
R4812 VSS.n2988 VSS.n2987 0.364419
R4813 VSS.n3236 VSS.n116 0.358995
R4814 VSS.n985 VSS.n984 0.358542
R4815 VSS.n2568 VSS.n2567 0.358542
R4816 VSS.n2543 VSS.n2542 0.358542
R4817 VSS.n2084 VSS.n2041 0.358542
R4818 VSS.n2576 VSS.n2575 0.340926
R4819 VSS.n2987 VSS.n2986 0.335802
R4820 VSS.n3430 uo_out[0] 0.3295
R4821 VSS.n3429 uo_out[1] 0.3295
R4822 VSS.n3428 uo_out[2] 0.3295
R4823 VSS.n3427 uo_out[3] 0.3295
R4824 VSS.n3426 uo_out[4] 0.3295
R4825 VSS.n3425 uo_out[5] 0.3295
R4826 VSS.n3424 uo_out[6] 0.3295
R4827 VSS.n3423 uo_out[7] 0.3295
R4828 VSS.n3422 uio_out[0] 0.3295
R4829 VSS.n3421 uio_out[1] 0.3295
R4830 VSS.n3420 uio_out[2] 0.3295
R4831 VSS.n3419 uio_out[3] 0.3295
R4832 VSS.n3418 uio_out[4] 0.3295
R4833 VSS.n3417 uio_out[5] 0.3295
R4834 VSS.n3416 uio_out[6] 0.3295
R4835 VSS.n3415 uio_out[7] 0.3295
R4836 VSS.n3414 uio_oe[0] 0.3295
R4837 VSS.n3413 uio_oe[1] 0.3295
R4838 VSS.n3412 uio_oe[2] 0.3295
R4839 VSS.n3411 uio_oe[3] 0.3295
R4840 VSS.n3410 uio_oe[4] 0.3295
R4841 VSS.n3409 uio_oe[5] 0.3295
R4842 VSS.n3408 uio_oe[6] 0.3295
R4843 VSS.n2318 VSS.n2317 0.307349
R4844 VSS.n1119 VSS.n1078 0.305262
R4845 VSS.n1137 VSS.n1072 0.305262
R4846 VSS.n1138 VSS.n1071 0.305262
R4847 VSS.n1151 VSS.n1150 0.305262
R4848 VSS.n1192 VSS.n1191 0.305262
R4849 VSS.n1177 VSS.n1176 0.305262
R4850 VSS.n2900 VSS.n2899 0.305262
R4851 VSS.n2876 VSS.n516 0.305262
R4852 VSS.n2871 VSS.n519 0.305262
R4853 VSS.n1656 VSS.n1633 0.305262
R4854 VSS.n2721 VSS.n2720 0.305262
R4855 VSS.n2737 VSS.n577 0.305262
R4856 VSS.n2738 VSS.n576 0.305262
R4857 VSS.n2751 VSS.n2750 0.305262
R4858 VSS.n2788 VSS.n2787 0.305262
R4859 VSS.n2798 VSS.n553 0.305262
R4860 VSS.n2800 VSS.n2799 0.305262
R4861 VSS.n2810 VSS.n546 0.305262
R4862 VSS.n2823 VSS.n2822 0.305262
R4863 VSS.n2834 VSS.n542 0.305262
R4864 VSS.n2671 VSS.n2670 0.305262
R4865 VSS.n635 VSS.n634 0.305262
R4866 VSS.n2657 VSS.n2656 0.305262
R4867 VSS.n2645 VSS.n639 0.305262
R4868 VSS.n2628 VSS.n2627 0.305262
R4869 VSS.n2613 VSS.n2612 0.305262
R4870 VSS.n941 VSS.n940 0.305262
R4871 VSS.n961 VSS.n930 0.305262
R4872 VSS.n1880 VSS.n1879 0.298799
R4873 VSS.n1116 VSS.n1115 0.298074
R4874 VSS.n2718 VSS.n2717 0.298074
R4875 VSS.n2674 VSS.n2673 0.298074
R4876 VSS.n471 VSS 0.286698
R4877 VSS.n2293 VSS.n861 0.282581
R4878 VSS.n1394 VSS.n1392 0.281546
R4879 VSS.n1092 VSS.n233 0.281132
R4880 VSS.n2322 VSS.n2321 0.263514
R4881 VSS.n1977 VSS.n1976 0.263514
R4882 VSS.n1831 VSS.n1712 0.263514
R4883 VSS.n2960 VSS.n2959 0.263514
R4884 VSS.n3235 VSS 0.260439
R4885 VSS.n1109 VSS.n1082 0.259086
R4886 VSS.n1684 VSS.n1683 0.259086
R4887 VSS.n1678 VSS.n1673 0.259086
R4888 VSS.n2709 VSS.n590 0.259086
R4889 VSS.n2838 VSS.n2837 0.259086
R4890 VSS.n2845 VSS.n2844 0.259086
R4891 VSS.n2756 VSS.n570 0.259086
R4892 VSS.n2761 VSS.n2760 0.259086
R4893 VSS.n996 VSS.n988 0.259086
R4894 VSS.n1011 VSS.n1010 0.259086
R4895 VSS.n2680 VSS.n617 0.259086
R4896 VSS.n743 VSS.n729 0.259086
R4897 VSS.n737 VSS.n736 0.259086
R4898 VSS.n1410 VSS.n1381 0.259086
R4899 VSS.n1418 VSS.n1379 0.259086
R4900 VSS.n1545 VSS.n1535 0.2565
R4901 VSS.n3406 VSS.n1 0.249698
R4902 VSS.n1298 VSS.n1297 0.239381
R4903 VSS.n1326 VSS.n1322 0.239381
R4904 VSS.n2440 VSS 0.237784
R4905 VSS.n1879 VSS.n116 0.23574
R4906 VSS.n2171 VSS.n2170 0.225061
R4907 VSS.n2179 VSS.n2178 0.225061
R4908 VSS.n1880 VSS.n1876 0.224703
R4909 VSS.n1800 VSS.n237 0.218753
R4910 VSS.n1603 VSS.n1602 0.204755
R4911 VSS.n2162 VSS.n2161 0.204755
R4912 VSS.n2163 VSS.n2162 0.204755
R4913 VSS VSS.n2440 0.200023
R4914 VSS.n1116 VSS 0.199635
R4915 VSS VSS.n2718 0.199635
R4916 VSS.n2673 VSS 0.199635
R4917 VSS.n231 VSS.n181 0.198729
R4918 VSS.n1801 VSS.n1800 0.196532
R4919 VSS.n1729 VSS.n234 0.196532
R4920 VSS.n2993 VSS.n2992 0.194976
R4921 VSS.n560 VSS.n557 0.192021
R4922 VSS.n2986 VSS.n234 0.18942
R4923 VSS.n1876 VSS.n1549 0.184476
R4924 VSS.n330 VSS.n230 0.1838
R4925 VSS.n3322 VSS.n3321 0.1838
R4926 VSS.n1919 VSS.n1915 0.180304
R4927 VSS.n2496 VSS 0.17983
R4928 VSS.n2176 VSS 0.17983
R4929 VSS.n1667 VSS.n1666 0.179521
R4930 VSS.n2568 VSS.n683 0.179521
R4931 VSS.n2085 VSS.n2084 0.179521
R4932 VSS.n1676 VSS 0.179485
R4933 VSS.n1596 VSS 0.179485
R4934 VSS.n1007 VSS 0.179485
R4935 VSS VSS.n734 0.179485
R4936 VSS.n1805 VSS.n1804 0.175416
R4937 VSS.n1555 VSS.n1554 0.175147
R4938 VSS.n1887 VSS.n1886 0.173577
R4939 VSS.n1554 VSS.n503 0.171842
R4940 VSS.n2860 VSS.n526 0.1603
R4941 VSS.n2860 VSS.n2859 0.1603
R4942 VSS.n2859 VSS.n529 0.1603
R4943 VSS.n689 VSS.n529 0.1603
R4944 VSS.n2459 VSS.n689 0.1603
R4945 VSS.n2459 VSS.n770 0.1603
R4946 VSS.n1988 VSS.n770 0.1603
R4947 VSS.n2907 VSS.n2906 0.1603
R4948 VSS.n2906 VSS.n506 0.1603
R4949 VSS.n2605 VSS.n506 0.1603
R4950 VSS.n2605 VSS.n2604 0.1603
R4951 VSS.n2604 VSS.n667 0.1603
R4952 VSS.n2105 VSS.n667 0.1603
R4953 VSS.n2105 VSS.n2028 0.1603
R4954 VSS.n1797 VSS.n565 0.1603
R4955 VSS.n2772 VSS.n565 0.1603
R4956 VSS.n2772 VSS.n566 0.1603
R4957 VSS.n801 VSS.n566 0.1603
R4958 VSS.n2385 VSS.n801 0.1603
R4959 VSS.n2385 VSS.n802 0.1603
R4960 VSS.n1345 VSS.n802 0.1603
R4961 VSS.n581 VSS.n267 0.1603
R4962 VSS.n2732 VSS.n581 0.1603
R4963 VSS.n2732 VSS.n582 0.1603
R4964 VSS.n826 VSS.n582 0.1603
R4965 VSS.n2338 VSS.n826 0.1603
R4966 VSS.n2338 VSS.n827 0.1603
R4967 VSS.n1286 VSS.n827 0.1603
R4968 VSS.n597 VSS.n237 0.1603
R4969 VSS.n2702 VSS.n597 0.1603
R4970 VSS.n2702 VSS.n2688 0.1603
R4971 VSS.n2688 VSS.n599 0.1603
R4972 VSS.n2296 VSS.n599 0.1603
R4973 VSS.n2296 VSS.n2295 0.1603
R4974 VSS.n2295 VSS.n859 0.1603
R4975 VSS.n1703 VSS.n1702 0.158327
R4976 VSS.n1702 VSS.n1623 0.158327
R4977 VSS.n1623 VSS.n713 0.158327
R4978 VSS.n2521 VSS.n713 0.158327
R4979 VSS.n2521 VSS.n2520 0.158327
R4980 VSS.n2520 VSS.n751 0.158327
R4981 VSS.n1173 VSS 0.158169
R4982 VSS.n2609 VSS 0.158169
R4983 VSS.n967 VSS 0.158169
R4984 VSS VSS.n2491 0.156867
R4985 VSS.n1954 VSS.n751 0.152235
R4986 VSS.n1949 VSS.n1919 0.151658
R4987 VSS.n861 VSS 0.146218
R4988 VSS.n1106 VSS.n1105 0.143027
R4989 VSS.n2706 VSS.n2705 0.143027
R4990 VSS.n615 VSS.n614 0.143027
R4991 VSS.n1106 VSS 0.14207
R4992 VSS.n1676 VSS 0.14207
R4993 VSS.n2706 VSS 0.14207
R4994 VSS.n1596 VSS 0.14207
R4995 VSS VSS.n615 0.14207
R4996 VSS.n1007 VSS 0.14207
R4997 VSS.n734 VSS 0.14207
R4998 VSS VSS.n1298 0.14207
R4999 VSS.n1326 VSS 0.14207
R5000 VSS.n2496 VSS 0.141725
R5001 VSS.n2176 VSS 0.141725
R5002 VSS.n1392 VSS.n233 0.141676
R5003 VSS.n3050 VSS.n3044 0.141672
R5004 VSS.n3082 VSS.n211 0.141672
R5005 VSS.n2502 VSS.n2501 0.13667
R5006 VSS.n2755 VSS.n571 0.126617
R5007 VSS.n3386 VSS.n37 0.1255
R5008 VSS.n3113 VSS.n3112 0.1255
R5009 VSS.n3295 VSS.n106 0.1255
R5010 VSS.n3236 VSS.n3235 0.122556
R5011 VSS.n3044 VSS 0.121778
R5012 VSS.n3107 VSS 0.121778
R5013 VSS.n2836 VSS.n2835 0.120632
R5014 VSS.n2308 VSS 0.120408
R5015 VSS.n54 VSS.n53 0.120292
R5016 VSS.n54 VSS.n41 0.120292
R5017 VSS.n3366 VSS.n59 0.120292
R5018 VSS.n3366 VSS.n3365 0.120292
R5019 VSS.n3364 VSS.n61 0.120292
R5020 VSS.n62 VSS.n61 0.120292
R5021 VSS.n3357 VSS.n3349 0.120292
R5022 VSS.n3357 VSS.n3356 0.120292
R5023 VSS.n3355 VSS.n3352 0.120292
R5024 VSS.n3352 VSS.n3351 0.120292
R5025 VSS.n3382 VSS.n3381 0.120292
R5026 VSS.n3378 VSS.n3377 0.120292
R5027 VSS.n51 VSS.n43 0.120292
R5028 VSS.n46 VSS.n43 0.120292
R5029 VSS.n46 VSS.n45 0.120292
R5030 VSS.n12 VSS.n11 0.120292
R5031 VSS.n3395 VSS.n18 0.120292
R5032 VSS.n19 VSS.n18 0.120292
R5033 VSS.n3389 VSS.n20 0.120292
R5034 VSS.n34 VSS.n23 0.120292
R5035 VSS.n28 VSS.n23 0.120292
R5036 VSS.n28 VSS.n27 0.120292
R5037 VSS.n3080 VSS.n213 0.120292
R5038 VSS.n3075 VSS.n213 0.120292
R5039 VSS.n3075 VSS.n3074 0.120292
R5040 VSS.n3031 VSS.n3030 0.120292
R5041 VSS.n3065 VSS.n3038 0.120292
R5042 VSS.n3059 VSS.n3038 0.120292
R5043 VSS.n3058 VSS.n3041 0.120292
R5044 VSS.n3051 VSS.n3050 0.120292
R5045 VSS.n3098 VSS.n3097 0.120292
R5046 VSS.n3097 VSS.n3086 0.120292
R5047 VSS.n3092 VSS.n3091 0.120292
R5048 VSS.n3091 VSS.n3088 0.120292
R5049 VSS.n3126 VSS.n3125 0.120292
R5050 VSS.n3125 VSS.n190 0.120292
R5051 VSS.n3120 VSS.n3119 0.120292
R5052 VSS.n3119 VSS.n193 0.120292
R5053 VSS.n3111 VSS.n3110 0.120292
R5054 VSS.n3245 VSS.n3240 0.120292
R5055 VSS.n3240 VSS.n80 0.120292
R5056 VSS.n3313 VSS.n82 0.120292
R5057 VSS.n3313 VSS.n3312 0.120292
R5058 VSS.n3311 VSS.n84 0.120292
R5059 VSS.n85 VSS.n84 0.120292
R5060 VSS.n3304 VSS.n88 0.120292
R5061 VSS.n3304 VSS.n3303 0.120292
R5062 VSS.n3302 VSS.n90 0.120292
R5063 VSS.n91 VSS.n90 0.120292
R5064 VSS.n105 VSS.n104 0.120292
R5065 VSS.n101 VSS.n100 0.120292
R5066 VSS.n3251 VSS.n3239 0.120292
R5067 VSS.n3252 VSS.n3251 0.120292
R5068 VSS.n3253 VSS.n3252 0.120292
R5069 VSS.n3264 VSS.n114 0.120292
R5070 VSS.n3272 VSS.n109 0.120292
R5071 VSS.n3276 VSS.n109 0.120292
R5072 VSS.n3278 VSS.n3277 0.120292
R5073 VSS.n3290 VSS.n3289 0.120292
R5074 VSS.n3289 VSS.n3281 0.120292
R5075 VSS.n3283 VSS.n3281 0.120292
R5076 VSS.n1111 VSS.n1110 0.120292
R5077 VSS.n1111 VSS.n1081 0.120292
R5078 VSS.n1115 VSS.n1081 0.120292
R5079 VSS.n1140 VSS.n1139 0.120292
R5080 VSS.n1140 VSS.n1070 0.120292
R5081 VSS.n1145 VSS.n1070 0.120292
R5082 VSS.n1146 VSS.n1145 0.120292
R5083 VSS.n1147 VSS.n1146 0.120292
R5084 VSS.n1147 VSS.n1068 0.120292
R5085 VSS.n1152 VSS.n1068 0.120292
R5086 VSS.n1193 VSS.n1162 0.120292
R5087 VSS.n1188 VSS.n1162 0.120292
R5088 VSS.n1188 VSS.n1187 0.120292
R5089 VSS.n1187 VSS.n1186 0.120292
R5090 VSS.n1186 VSS.n1169 0.120292
R5091 VSS.n1181 VSS.n1169 0.120292
R5092 VSS.n1181 VSS.n1180 0.120292
R5093 VSS.n1180 VSS.n1179 0.120292
R5094 VSS.n1179 VSS.n1171 0.120292
R5095 VSS.n2889 VSS.n2888 0.120292
R5096 VSS.n2888 VSS.n513 0.120292
R5097 VSS.n2884 VSS.n513 0.120292
R5098 VSS.n2884 VSS.n2883 0.120292
R5099 VSS.n2883 VSS.n515 0.120292
R5100 VSS.n2878 VSS.n515 0.120292
R5101 VSS.n2878 VSS.n2877 0.120292
R5102 VSS.n2870 VSS.n2869 0.120292
R5103 VSS.n1645 VSS.n1636 0.120292
R5104 VSS.n1649 VSS.n1636 0.120292
R5105 VSS.n1650 VSS.n1649 0.120292
R5106 VSS.n1650 VSS.n1634 0.120292
R5107 VSS.n1654 VSS.n1634 0.120292
R5108 VSS.n1655 VSS.n1654 0.120292
R5109 VSS.n1662 VSS.n1631 0.120292
R5110 VSS.n1663 VSS.n1662 0.120292
R5111 VSS.n1664 VSS.n1663 0.120292
R5112 VSS.n1685 VSS.n1670 0.120292
R5113 VSS.n1680 VSS.n1670 0.120292
R5114 VSS.n1680 VSS.n1679 0.120292
R5115 VSS.n2711 VSS.n2710 0.120292
R5116 VSS.n2711 VSS.n589 0.120292
R5117 VSS.n2717 VSS.n589 0.120292
R5118 VSS.n2740 VSS.n2739 0.120292
R5119 VSS.n2740 VSS.n575 0.120292
R5120 VSS.n2745 VSS.n575 0.120292
R5121 VSS.n2746 VSS.n2745 0.120292
R5122 VSS.n2747 VSS.n2746 0.120292
R5123 VSS.n2747 VSS.n573 0.120292
R5124 VSS.n2752 VSS.n573 0.120292
R5125 VSS.n2758 VSS.n2757 0.120292
R5126 VSS.n2784 VSS.n558 0.120292
R5127 VSS.n2785 VSS.n2784 0.120292
R5128 VSS.n2786 VSS.n556 0.120292
R5129 VSS.n2791 VSS.n556 0.120292
R5130 VSS.n2792 VSS.n2791 0.120292
R5131 VSS.n2792 VSS.n554 0.120292
R5132 VSS.n2796 VSS.n554 0.120292
R5133 VSS.n2797 VSS.n2796 0.120292
R5134 VSS.n2807 VSS.n2801 0.120292
R5135 VSS.n2821 VSS.n545 0.120292
R5136 VSS.n2826 VSS.n545 0.120292
R5137 VSS.n2827 VSS.n2826 0.120292
R5138 VSS.n2827 VSS.n543 0.120292
R5139 VSS.n2831 VSS.n543 0.120292
R5140 VSS.n2833 VSS.n2831 0.120292
R5141 VSS.n2840 VSS.n2839 0.120292
R5142 VSS.n2841 VSS.n2840 0.120292
R5143 VSS.n1573 VSS.n1572 0.120292
R5144 VSS.n1576 VSS.n1573 0.120292
R5145 VSS.n1577 VSS.n1576 0.120292
R5146 VSS.n1578 VSS.n1577 0.120292
R5147 VSS.n1578 VSS.n1569 0.120292
R5148 VSS.n1569 VSS.n1567 0.120292
R5149 VSS.n1583 VSS.n1567 0.120292
R5150 VSS.n1584 VSS.n1583 0.120292
R5151 VSS.n1585 VSS.n1584 0.120292
R5152 VSS.n1585 VSS.n1565 0.120292
R5153 VSS.n1607 VSS.n1592 0.120292
R5154 VSS.n1601 VSS.n1592 0.120292
R5155 VSS.n2679 VSS.n2678 0.120292
R5156 VSS.n2678 VSS.n618 0.120292
R5157 VSS.n2674 VSS.n618 0.120292
R5158 VSS.n2658 VSS.n633 0.120292
R5159 VSS.n2653 VSS.n633 0.120292
R5160 VSS.n2653 VSS.n2652 0.120292
R5161 VSS.n2652 VSS.n2651 0.120292
R5162 VSS.n2651 VSS.n637 0.120292
R5163 VSS.n2647 VSS.n637 0.120292
R5164 VSS.n2647 VSS.n2646 0.120292
R5165 VSS.n2629 VSS.n651 0.120292
R5166 VSS.n2624 VSS.n651 0.120292
R5167 VSS.n2624 VSS.n2623 0.120292
R5168 VSS.n2623 VSS.n2622 0.120292
R5169 VSS.n2622 VSS.n658 0.120292
R5170 VSS.n2617 VSS.n658 0.120292
R5171 VSS.n2617 VSS.n2616 0.120292
R5172 VSS.n2616 VSS.n2615 0.120292
R5173 VSS.n2615 VSS.n660 0.120292
R5174 VSS.n952 VSS.n951 0.120292
R5175 VSS.n952 VSS.n934 0.120292
R5176 VSS.n956 VSS.n934 0.120292
R5177 VSS.n957 VSS.n956 0.120292
R5178 VSS.n957 VSS.n932 0.120292
R5179 VSS.n963 VSS.n932 0.120292
R5180 VSS.n964 VSS.n963 0.120292
R5181 VSS.n1043 VSS.n1042 0.120292
R5182 VSS.n1042 VSS.n980 0.120292
R5183 VSS VSS.n980 0.120292
R5184 VSS.n1037 VSS.n1036 0.120292
R5185 VSS.n1033 VSS.n1032 0.120292
R5186 VSS.n1032 VSS.n987 0.120292
R5187 VSS.n1019 VSS.n995 0.120292
R5188 VSS.n1014 VSS.n995 0.120292
R5189 VSS.n1014 VSS.n1013 0.120292
R5190 VSS.n1013 VSS.n1005 0.120292
R5191 VSS.n1412 VSS.n1411 0.120292
R5192 VSS.n1412 VSS.n1380 0.120292
R5193 VSS.n1416 VSS.n1380 0.120292
R5194 VSS.n1417 VSS.n1416 0.120292
R5195 VSS.n1422 VSS.n1421 0.120292
R5196 VSS.n1427 VSS.n1376 0.120292
R5197 VSS.n1452 VSS.n1366 0.120292
R5198 VSS.n1453 VSS.n1452 0.120292
R5199 VSS.n1454 VSS.n1453 0.120292
R5200 VSS.n1454 VSS.n1364 0.120292
R5201 VSS.n1459 VSS.n1364 0.120292
R5202 VSS.n1460 VSS.n1459 0.120292
R5203 VSS.n1525 VSS.n1524 0.120292
R5204 VSS.n1508 VSS.n1507 0.120292
R5205 VSS.n1507 VSS.n1506 0.120292
R5206 VSS.n1506 VSS.n1479 0.120292
R5207 VSS.n1500 VSS.n1479 0.120292
R5208 VSS.n1500 VSS.n1499 0.120292
R5209 VSS.n1499 VSS.n1498 0.120292
R5210 VSS.n1498 VSS.n1484 0.120292
R5211 VSS.n1491 VSS.n1484 0.120292
R5212 VSS.n1491 VSS.n1490 0.120292
R5213 VSS.n1490 VSS.n1489 0.120292
R5214 VSS.n2588 VSS.n2587 0.120292
R5215 VSS.n2582 VSS.n2581 0.120292
R5216 VSS.n2581 VSS.n680 0.120292
R5217 VSS.n2574 VSS.n680 0.120292
R5218 VSS.n2547 VSS.n2546 0.120292
R5219 VSS.n2546 VSS.n697 0.120292
R5220 VSS.n2540 VSS.n697 0.120292
R5221 VSS.n2540 VSS.n2539 0.120292
R5222 VSS.n2539 VSS.n2538 0.120292
R5223 VSS.n2538 VSS.n702 0.120292
R5224 VSS.n2531 VSS.n2530 0.120292
R5225 VSS.n2530 VSS.n706 0.120292
R5226 VSS.n2525 VSS.n706 0.120292
R5227 VSS.n742 VSS.n741 0.120292
R5228 VSS.n741 VSS.n730 0.120292
R5229 VSS.n735 VSS.n730 0.120292
R5230 VSS.n2307 VSS.n841 0.120292
R5231 VSS.n2309 VSS.n837 0.120292
R5232 VSS.n2314 VSS.n837 0.120292
R5233 VSS.n2315 VSS.n2314 0.120292
R5234 VSS.n2315 VSS.n833 0.120292
R5235 VSS.n2323 VSS.n833 0.120292
R5236 VSS.n2325 VSS.n2324 0.120292
R5237 VSS.n2347 VSS.n2346 0.120292
R5238 VSS.n2347 VSS.n816 0.120292
R5239 VSS.n2353 VSS.n816 0.120292
R5240 VSS.n2354 VSS.n2353 0.120292
R5241 VSS.n2364 VSS.n813 0.120292
R5242 VSS.n2365 VSS.n2364 0.120292
R5243 VSS.n2372 VSS.n2371 0.120292
R5244 VSS.n2395 VSS.n793 0.120292
R5245 VSS.n2401 VSS.n793 0.120292
R5246 VSS.n2402 VSS.n2401 0.120292
R5247 VSS.n2403 VSS.n2402 0.120292
R5248 VSS.n2403 VSS.n791 0.120292
R5249 VSS.n2408 VSS.n791 0.120292
R5250 VSS.n2434 VSS.n2433 0.120292
R5251 VSS.n2435 VSS.n2434 0.120292
R5252 VSS.n2446 VSS.n2445 0.120292
R5253 VSS.n2447 VSS.n2446 0.120292
R5254 VSS.n2467 VSS.n765 0.120292
R5255 VSS.n2468 VSS.n2467 0.120292
R5256 VSS.n2468 VSS.n761 0.120292
R5257 VSS.n2472 VSS.n761 0.120292
R5258 VSS.n2473 VSS.n2472 0.120292
R5259 VSS.n2474 VSS.n2473 0.120292
R5260 VSS.n2474 VSS.n758 0.120292
R5261 VSS.n2481 VSS.n758 0.120292
R5262 VSS.n2482 VSS.n2481 0.120292
R5263 VSS.n2503 VSS.n2488 0.120292
R5264 VSS.n2286 VSS.n2285 0.120292
R5265 VSS.n2277 VSS.n879 0.120292
R5266 VSS.n2277 VSS.n2276 0.120292
R5267 VSS.n2276 VSS.n883 0.120292
R5268 VSS.n884 VSS.n883 0.120292
R5269 VSS.n2270 VSS.n2269 0.120292
R5270 VSS.n2247 VSS.n2246 0.120292
R5271 VSS.n2246 VSS.n2245 0.120292
R5272 VSS.n2242 VSS.n2241 0.120292
R5273 VSS.n2241 VSS.n899 0.120292
R5274 VSS.n2074 VSS.n2044 0.120292
R5275 VSS.n2078 VSS.n2044 0.120292
R5276 VSS.n2080 VSS.n2079 0.120292
R5277 VSS.n2087 VSS.n2040 0.120292
R5278 VSS.n2089 VSS.n2038 0.120292
R5279 VSS.n2093 VSS.n2038 0.120292
R5280 VSS.n2094 VSS.n2093 0.120292
R5281 VSS.n2109 VSS.n908 0.120292
R5282 VSS.n2114 VSS.n908 0.120292
R5283 VSS.n2116 VSS.n2115 0.120292
R5284 VSS.n2116 VSS.n904 0.120292
R5285 VSS.n2121 VSS.n904 0.120292
R5286 VSS.n2122 VSS.n2121 0.120292
R5287 VSS.n2217 VSS.n2131 0.120292
R5288 VSS.n2212 VSS.n2131 0.120292
R5289 VSS.n2212 VSS.n2211 0.120292
R5290 VSS.n2211 VSS.n2210 0.120292
R5291 VSS.n2210 VSS.n2146 0.120292
R5292 VSS.n2205 VSS.n2146 0.120292
R5293 VSS.n2205 VSS.n2204 0.120292
R5294 VSS.n2203 VSS.n2150 0.120292
R5295 VSS.n2195 VSS.n2150 0.120292
R5296 VSS.n2186 VSS.n2158 0.120292
R5297 VSS.n2182 VSS.n2158 0.120292
R5298 VSS.n2182 VSS.n2181 0.120292
R5299 VSS.n2181 VSS.n2173 0.120292
R5300 VSS.n1256 VSS.n1255 0.120292
R5301 VSS.n1260 VSS.n1259 0.120292
R5302 VSS.n1261 VSS.n1260 0.120292
R5303 VSS.n1265 VSS.n1264 0.120292
R5304 VSS.n1265 VSS.n1223 0.120292
R5305 VSS.n1271 VSS.n1223 0.120292
R5306 VSS.n1297 VSS.n1214 0.120292
R5307 VSS.n1304 VSS.n1303 0.120292
R5308 VSS.n1355 VSS.n1354 0.120292
R5309 VSS.n1337 VSS.n1336 0.120292
R5310 VSS.n1332 VSS.n1331 0.120292
R5311 VSS.n1331 VSS.n1322 0.120292
R5312 VSS.n2014 VSS.n924 0.120292
R5313 VSS.n2009 VSS.n924 0.120292
R5314 VSS.n2009 VSS.n2008 0.120292
R5315 VSS.n2004 VSS.n2003 0.120292
R5316 VSS.n1999 VSS.n1998 0.120292
R5317 VSS.n1998 VSS.n1898 0.120292
R5318 VSS.n1984 VSS.n1910 0.120292
R5319 VSS.n1973 VSS.n1972 0.120292
R5320 VSS.n1968 VSS.n1967 0.120292
R5321 VSS.n1967 VSS.n1915 0.120292
R5322 VSS.n1940 VSS.n1928 0.120292
R5323 VSS.n1936 VSS.n1935 0.120292
R5324 VSS.n1935 VSS.n1931 0.120292
R5325 VSS.n2980 VSS.n239 0.120292
R5326 VSS.n2973 VSS.n239 0.120292
R5327 VSS.n2972 VSS.n2971 0.120292
R5328 VSS.n2971 VSS.n257 0.120292
R5329 VSS.n2967 VSS.n257 0.120292
R5330 VSS.n2967 VSS.n2966 0.120292
R5331 VSS.n2966 VSS.n2965 0.120292
R5332 VSS.n2965 VSS.n260 0.120292
R5333 VSS.n2958 VSS.n260 0.120292
R5334 VSS.n2940 VSS.n2939 0.120292
R5335 VSS.n2939 VSS.n274 0.120292
R5336 VSS.n2935 VSS.n274 0.120292
R5337 VSS.n2935 VSS.n2934 0.120292
R5338 VSS.n2934 VSS.n276 0.120292
R5339 VSS.n2930 VSS.n276 0.120292
R5340 VSS.n2930 VSS.n2929 0.120292
R5341 VSS.n1743 VSS.n1738 0.120292
R5342 VSS.n1793 VSS.n1734 0.120292
R5343 VSS.n1789 VSS.n1734 0.120292
R5344 VSS.n1789 VSS.n1788 0.120292
R5345 VSS.n1788 VSS.n1787 0.120292
R5346 VSS.n1787 VSS.n1758 0.120292
R5347 VSS.n1782 VSS.n1758 0.120292
R5348 VSS.n1782 VSS.n1781 0.120292
R5349 VSS.n1781 VSS.n1780 0.120292
R5350 VSS.n1780 VSS 0.120292
R5351 VSS.n1775 VSS.n1774 0.120292
R5352 VSS.n2912 VSS.n2911 0.120292
R5353 VSS.n2912 VSS.n498 0.120292
R5354 VSS.n2916 VSS.n498 0.120292
R5355 VSS.n2917 VSS.n2916 0.120292
R5356 VSS.n2917 VSS.n496 0.120292
R5357 VSS.n2921 VSS.n496 0.120292
R5358 VSS.n2922 VSS.n2921 0.120292
R5359 VSS.n1721 VSS.n1720 0.120292
R5360 VSS.n1821 VSS.n1713 0.120292
R5361 VSS.n1829 VSS.n1713 0.120292
R5362 VSS.n1830 VSS.n1829 0.120292
R5363 VSS.n1835 VSS.n1834 0.120292
R5364 VSS.n1840 VSS.n1709 0.120292
R5365 VSS.n1841 VSS.n1840 0.120292
R5366 VSS.n1842 VSS.n1841 0.120292
R5367 VSS.n1866 VSS.n1865 0.120292
R5368 VSS.n1865 VSS.n1848 0.120292
R5369 VSS.n1861 VSS.n1848 0.120292
R5370 VSS.n1861 VSS.n1860 0.120292
R5371 VSS.n1857 VSS.n1856 0.120292
R5372 VSS.n1856 VSS.n1852 0.120292
R5373 VSS.n116 VSS 0.114397
R5374 VSS.n330 VSS.n329 0.113648
R5375 VSS.n3322 VSS.n78 0.113648
R5376 VSS.n229 VSS 0.11275
R5377 VSS.n130 VSS.n129 0.111077
R5378 VSS.n135 VSS.n134 0.111077
R5379 VSS.n140 VSS.n139 0.111077
R5380 VSS.n145 VSS.n144 0.111077
R5381 VSS.n150 VSS.n149 0.111077
R5382 VSS.n155 VSS.n154 0.111077
R5383 VSS.n160 VSS.n159 0.111077
R5384 VSS.n165 VSS.n164 0.111077
R5385 VSS.n170 VSS.n169 0.111077
R5386 VSS.n968 VSS.n967 0.109992
R5387 VSS.n1802 VSS.n503 0.10744
R5388 VSS.n1804 VSS.n1803 0.10744
R5389 VSS.n1446 VSS.n1445 0.102062
R5390 VSS.n2346 VSS.n820 0.102062
R5391 VSS.n2252 VSS.n2251 0.102062
R5392 VSS.n1289 VSS.n1214 0.102062
R5393 VSS.n2945 VSS.n2940 0.102062
R5394 VSS.n1392 VSS.n861 0.0991735
R5395 VSS.n11 VSS 0.0981562
R5396 VSS.n3030 VSS 0.0981562
R5397 VSS VSS.n114 0.0981562
R5398 VSS.n1139 VSS 0.0981562
R5399 VSS.n1206 VSS 0.0981562
R5400 VSS.n2874 VSS 0.0981562
R5401 VSS VSS.n1631 0.0981562
R5402 VSS.n2739 VSS 0.0981562
R5403 VSS.n2753 VSS 0.0981562
R5404 VSS.n2801 VSS 0.0981562
R5405 VSS.n2821 VSS 0.0981562
R5406 VSS VSS.n2832 0.0981562
R5407 VSS VSS.n2658 0.0981562
R5408 VSS.n2642 VSS 0.0981562
R5409 VSS.n1063 VSS 0.0981562
R5410 VSS.n1033 VSS 0.0981562
R5411 VSS.n1421 VSS 0.0981562
R5412 VSS.n1508 VSS 0.0981562
R5413 VSS.n2565 VSS 0.0981562
R5414 VSS.n2531 VSS 0.0981562
R5415 VSS.n2410 VSS 0.0981562
R5416 VSS VSS.n2281 0.0981562
R5417 VSS.n2247 VSS 0.0981562
R5418 VSS.n2089 VSS 0.0981562
R5419 VSS.n2226 VSS 0.0981562
R5420 VSS.n279 VSS 0.0981562
R5421 VSS.n1775 VSS 0.0981562
R5422 VSS VSS.n494 0.0981562
R5423 VSS.n1857 VSS 0.0981562
R5424 VSS.n1645 VSS.n1644 0.0968542
R5425 VSS.n1572 VSS.n536 0.0968542
R5426 VSS.n1048 VSS.n1047 0.0968542
R5427 VSS.n2552 VSS.n2547 0.0968542
R5428 VSS.n2395 VSS 0.0968542
R5429 VSS VSS.n2270 0.0968542
R5430 VSS.n1985 VSS.n1984 0.0968542
R5431 VSS.n1821 VSS.n1820 0.0968542
R5432 VSS.n1255 VSS 0.0955521
R5433 VSS.n1273 VSS 0.0955521
R5434 VSS.n1303 VSS 0.0955521
R5435 VSS VSS.n1337 0.0955521
R5436 VSS VSS.n2004 0.0955521
R5437 VSS VSS.n1973 0.0955521
R5438 VSS VSS.n1940 0.0955521
R5439 VSS.n1834 VSS 0.0955521
R5440 VSS.n1811 VSS.n1726 0.0950946
R5441 VSS.n1819 VSS.n1818 0.0950946
R5442 VSS.n249 VSS.n243 0.0950946
R5443 VSS.n2982 VSS.n238 0.0950946
R5444 VSS.n1747 VSS.n1737 0.0950946
R5445 VSS.n1795 VSS.n1732 0.0950946
R5446 VSS.n1766 VSS.n1765 0.0950946
R5447 VSS.n2909 VSS.n501 0.0950946
R5448 VSS.n1395 VSS.n1391 0.0950946
R5449 VSS.n1404 VSS.n1383 0.0950946
R5450 VSS.n2523 VSS.n711 0.0950946
R5451 VSS.n748 VSS.n715 0.0950946
R5452 VSS.n2904 VSS.n2903 0.0950946
R5453 VSS.n2895 VSS.n2894 0.0950946
R5454 VSS.n1200 VSS.n1158 0.0950946
R5455 VSS.n1194 VSS.n1161 0.0950946
R5456 VSS.n1123 VSS.n1121 0.0950946
R5457 VSS.n1134 VSS.n1074 0.0950946
R5458 VSS.n1094 VSS.n1093 0.0950946
R5459 VSS.n1104 VSS.n1087 0.0950946
R5460 VSS.n1700 VSS.n1699 0.0950946
R5461 VSS.n1691 VSS.n1690 0.0950946
R5462 VSS.n2864 VSS.n523 0.0950946
R5463 VSS.n1643 VSS.n1642 0.0950946
R5464 VSS.n2730 VSS.n2729 0.0950946
R5465 VSS.n2734 VSS.n579 0.0950946
R5466 VSS.n2700 VSS.n2699 0.0950946
R5467 VSS.n2704 VSS.n595 0.0950946
R5468 VSS.n1621 VSS.n1620 0.0950946
R5469 VSS.n1613 VSS.n1612 0.0950946
R5470 VSS.n2805 VSS.n2803 0.0950946
R5471 VSS.n2818 VSS.n548 0.0950946
R5472 VSS.n2770 VSS.n2769 0.0950946
R5473 VSS.n2774 VSS.n563 0.0950946
R5474 VSS.n2857 VSS.n2856 0.0950946
R5475 VSS.n2850 VSS.n535 0.0950946
R5476 VSS.n2666 VSS.n626 0.0950946
R5477 VSS.n2660 VSS.n629 0.0950946
R5478 VSS.n2686 VSS.n2685 0.0950946
R5479 VSS.n613 VSS.n612 0.0950946
R5480 VSS.n1026 VSS.n990 0.0950946
R5481 VSS.n1021 VSS.n993 0.0950946
R5482 VSS.n2607 VSS.n663 0.0950946
R5483 VSS.n949 VSS.n948 0.0950946
R5484 VSS.n2636 VSS.n647 0.0950946
R5485 VSS.n2630 VSS.n650 0.0950946
R5486 VSS.n1055 VSS.n969 0.0950946
R5487 VSS.n1049 VSS.n972 0.0950946
R5488 VSS.n2457 VSS.n2456 0.0950946
R5489 VSS.n2461 VSS.n768 0.0950946
R5490 VSS.n2224 VSS.n2126 0.0950946
R5491 VSS.n2219 VSS.n2129 0.0950946
R5492 VSS.n1992 VSS.n1902 0.0950946
R5493 VSS.n1986 VSS.n1906 0.0950946
R5494 VSS.n2563 VSS.n688 0.0950946
R5495 VSS.n2551 VSS.n2548 0.0950946
R5496 VSS.n1472 VSS.n1471 0.0950946
R5497 VSS.n1514 VSS.n1469 0.0950946
R5498 VSS.n1430 VSS.n1428 0.0950946
R5499 VSS.n1444 VSS.n1369 0.0950946
R5500 VSS.n2602 VSS.n2601 0.0950946
R5501 VSS.n2594 VSS.n2593 0.0950946
R5502 VSS.n2103 VSS.n2102 0.0950946
R5503 VSS.n2107 VSS.n911 0.0950946
R5504 VSS.n2026 VSS.n2025 0.0950946
R5505 VSS.n2018 VSS.n2017 0.0950946
R5506 VSS.n2418 VSS.n787 0.0950946
R5507 VSS.n2426 VSS.n2425 0.0950946
R5508 VSS.n2336 VSS.n2335 0.0950946
R5509 VSS.n2341 VSS.n2340 0.0950946
R5510 VSS.n2298 VSS.n846 0.0950946
R5511 VSS.n856 VSS.n853 0.0950946
R5512 VSS.n2518 VSS.n2517 0.0950946
R5513 VSS.n2508 VSS.n2507 0.0950946
R5514 VSS.n2383 VSS.n2382 0.0950946
R5515 VSS.n2388 VSS.n2387 0.0950946
R5516 VSS.n1349 VSS.n1311 0.0950946
R5517 VSS.n1343 VSS.n1315 0.0950946
R5518 VSS.n2060 VSS.n2057 0.0950946
R5519 VSS.n2072 VSS.n2049 0.0950946
R5520 VSS.n2292 VSS.n2291 0.0950946
R5521 VSS.n874 VSS.n873 0.0950946
R5522 VSS.n2193 VSS.n2153 0.0950946
R5523 VSS.n2188 VSS.n2156 0.0950946
R5524 VSS.n2257 VSS.n2256 0.0950946
R5525 VSS.n2263 VSS.n2262 0.0950946
R5526 VSS.n1284 VSS.n1283 0.0950946
R5527 VSS.n1288 VSS.n1216 0.0950946
R5528 VSS.n1241 VSS.n1234 0.0950946
R5529 VSS.n1249 VSS.n1248 0.0950946
R5530 VSS.n1952 VSS.n1951 0.0950946
R5531 VSS.n1947 VSS.n1923 0.0950946
R5532 VSS.n1874 VSS.n1873 0.0950946
R5533 VSS.n1846 VSS.n1552 0.0950946
R5534 VSS.n2955 VSS.n266 0.0950946
R5535 VSS.n2944 VSS.n2941 0.0950946
R5536 VSS.n52 VSS 0.09425
R5537 VSS.n3081 VSS 0.09425
R5538 VSS VSS.n3246 0.09425
R5539 VSS.n3107 VSS.n3105 0.0934947
R5540 VSS.n1664 VSS.n1625 0.0916458
R5541 VSS.n1565 VSS.n1559 0.0916458
R5542 VSS.n2525 VSS.n2524 0.0916458
R5543 VSS.n2483 VSS.n753 0.0916458
R5544 VSS.n1842 VSS.n1704 0.0916458
R5545 VSS.n1878 VSS 0.0907344
R5546 VSS.n129 VSS 0.0906442
R5547 VSS.n134 VSS 0.0906442
R5548 VSS.n139 VSS 0.0906442
R5549 VSS.n144 VSS 0.0906442
R5550 VSS.n149 VSS 0.0906442
R5551 VSS.n154 VSS 0.0906442
R5552 VSS.n159 VSS 0.0906442
R5553 VSS.n164 VSS 0.0906442
R5554 VSS.n169 VSS 0.0906442
R5555 VSS.n1659 VSS.n1658 0.0900105
R5556 VSS.n1046 VSS.n1045 0.0900105
R5557 VSS.n1802 VSS.n1801 0.0898892
R5558 VSS.n1803 VSS.n1729 0.0898892
R5559 VSS.n3373 VSS 0.0881354
R5560 VSS.n3104 VSS 0.0881354
R5561 VSS.n79 VSS 0.0881354
R5562 VSS.n1204 VSS.n1153 0.0864375
R5563 VSS.n2758 VSS.n568 0.0864375
R5564 VSS.n2640 VSS.n642 0.0864375
R5565 VSS.n2372 VSS.n804 0.0864375
R5566 VSS.n1354 VSS.n1307 0.0864375
R5567 VSS.n1744 VSS.n1743 0.0864375
R5568 VSS.n3407 VSS.n0 0.0853293
R5569 VSS.n1129 VSS.n1077 0.0838333
R5570 VSS.n1164 VSS.n1163 0.0838333
R5571 VSS.n2896 VSS.n2890 0.0838333
R5572 VSS.n2865 VSS.n522 0.0838333
R5573 VSS.n1669 VSS.n1628 0.0838333
R5574 VSS.n2728 VSS.n2727 0.0838333
R5575 VSS.n2765 VSS.n562 0.0838333
R5576 VSS.n2806 VSS.n2802 0.0838333
R5577 VSS.n2819 VSS.n547 0.0838333
R5578 VSS.n1591 VSS.n1562 0.0838333
R5579 VSS.n2667 VSS.n625 0.0838333
R5580 VSS.n653 VSS.n652 0.0838333
R5581 VSS.n950 VSS.n936 0.0838333
R5582 VSS.n1000 VSS.n998 0.0838333
R5583 VSS.n1439 VSS.n1372 0.0838333
R5584 VSS.n1519 VSS.n1467 0.0838333
R5585 VSS.n2600 VSS.n669 0.0838333
R5586 VSS.n2595 VSS.n2589 0.0838333
R5587 VSS.n2558 VSS.n692 0.0838333
R5588 VSS.n724 VSS.n720 0.0838333
R5589 VSS.n2334 VSS.n2333 0.0838333
R5590 VSS.n2389 VSS.n798 0.0838333
R5591 VSS.n2417 VSS.n2415 0.0838333
R5592 VSS.n2427 VSS.n782 0.0838333
R5593 VSS.n2455 VSS.n2454 0.0838333
R5594 VSS.n2255 VSS.n891 0.0838333
R5595 VSS.n2067 VSS.n2066 0.0838333
R5596 VSS.n2108 VSS.n910 0.0838333
R5597 VSS.n2138 VSS.n2136 0.0838333
R5598 VSS.n1317 VSS.n1316 0.0838333
R5599 VSS.n1993 VSS.n1901 0.0838333
R5600 VSS.n2950 VSS.n269 0.0838333
R5601 VSS.n1752 VSS.n1736 0.0838333
R5602 VSS.n1763 VSS.n1761 0.0838333
R5603 VSS.n2910 VSS.n500 0.0838333
R5604 VSS.n1812 VSS.n1718 0.0838333
R5605 VSS.n1847 VSS.n1707 0.0838333
R5606 VSS VSS.n2491 0.082648
R5607 VSS VSS.n2308 0.082648
R5608 VSS.n1925 VSS 0.0773229
R5609 VSS.n2993 VSS.n228 0.0766574
R5610 VSS.n3140 VSS.n181 0.0766574
R5611 VSS.n1125 VSS.n1124 0.0760208
R5612 VSS.n586 VSS.n584 0.0760208
R5613 VSS.n2668 VSS.n622 0.0760208
R5614 VSS.n1432 VSS.n1431 0.0760208
R5615 VSS.n2331 VSS.n829 0.0760208
R5616 VSS.n889 VSS.n887 0.0760208
R5617 VSS.n1276 VSS.n1219 0.0760208
R5618 VSS.n2956 VSS.n265 0.0760208
R5619 VSS.n1877 VSS.n1546 0.0747188
R5620 VSS.n3378 VSS.n3374 0.0721146
R5621 VSS.n101 VSS.n96 0.0721146
R5622 VSS.n3103 VSS.n210 0.0708554
R5623 VSS.n3397 VSS.n17 0.0708125
R5624 VSS.n3071 VSS.n3070 0.0708125
R5625 VSS.n3270 VSS.n111 0.0708125
R5626 VSS.n1099 VSS.n1098 0.0708125
R5627 VSS.n1201 VSS.n1157 0.0708125
R5628 VSS.n2866 VSS.n520 0.0708125
R5629 VSS.n2696 VSS.n2693 0.0708125
R5630 VSS.n2768 VSS.n2767 0.0708125
R5631 VSS.n533 VSS.n531 0.0708125
R5632 VSS.n605 VSS.n603 0.0708125
R5633 VSS.n2637 VSS.n646 0.0708125
R5634 VSS.n1057 VSS.n968 0.0708125
R5635 VSS.n1399 VSS.n1398 0.0708125
R5636 VSS.n1520 VSS.n1466 0.0708125
R5637 VSS.n2564 VSS.n687 0.0708125
R5638 VSS.n850 VSS.n843 0.0708125
R5639 VSS.n2381 VSS.n2380 0.0708125
R5640 VSS.n2450 VSS.n772 0.0708125
R5641 VSS.n866 VSS.n864 0.0708125
R5642 VSS.n2065 VSS.n2052 0.0708125
R5643 VSS.n1251 VSS.n1231 0.0708125
R5644 VSS.n1350 VSS.n1310 0.0708125
R5645 VSS.n1994 VSS.n1900 0.0708125
R5646 VSS.n254 VSS.n252 0.0708125
R5647 VSS.n1813 VSS.n1725 0.0708125
R5648 VSS.n2902 VSS 0.0695104
R5649 VSS.n938 VSS 0.0695104
R5650 VSS.n2577 VSS.n2576 0.0685851
R5651 VSS.n1173 VSS.n508 0.068325
R5652 VSS.n2609 VSS.n2608 0.068325
R5653 VSS.n1810 VSS.n1727 0.0680676
R5654 VSS.n1727 VSS.n1717 0.0680676
R5655 VSS.n251 VSS.n250 0.0680676
R5656 VSS.n251 VSS.n236 0.0680676
R5657 VSS.n1751 VSS.n1749 0.0680676
R5658 VSS.n1751 VSS.n1750 0.0680676
R5659 VSS.n1769 VSS.n1767 0.0680676
R5660 VSS.n1769 VSS.n1768 0.0680676
R5661 VSS.n1400 VSS.n1385 0.0680676
R5662 VSS.n1401 VSS.n1400 0.0680676
R5663 VSS.n723 VSS.n721 0.0680676
R5664 VSS.n723 VSS.n722 0.0680676
R5665 VSS.n2891 VSS.n509 0.0680676
R5666 VSS.n2893 VSS.n2891 0.0680676
R5667 VSS.n1199 VSS.n1159 0.0680676
R5668 VSS.n1160 VSS.n1159 0.0680676
R5669 VSS.n1130 VSS.n1076 0.0680676
R5670 VSS.n1131 VSS.n1130 0.0680676
R5671 VSS.n1100 VSS.n1089 0.0680676
R5672 VSS.n1101 VSS.n1100 0.0680676
R5673 VSS.n1687 VSS.n1626 0.0680676
R5674 VSS.n1689 VSS.n1687 0.0680676
R5675 VSS.n2863 VSS.n524 0.0680676
R5676 VSS.n1639 VSS.n524 0.0680676
R5677 VSS.n2726 VSS.n585 0.0680676
R5678 VSS.n2726 VSS.n2725 0.0680676
R5679 VSS.n2695 VSS.n2691 0.0680676
R5680 VSS.n2695 VSS.n2694 0.0680676
R5681 VSS.n1609 VSS.n1560 0.0680676
R5682 VSS.n1611 VSS.n1609 0.0680676
R5683 VSS.n2814 VSS.n550 0.0680676
R5684 VSS.n2815 VSS.n2814 0.0680676
R5685 VSS.n2764 VSS.n569 0.0680676
R5686 VSS.n2764 VSS.n2763 0.0680676
R5687 VSS.n2853 VSS.n532 0.0680676
R5688 VSS.n2853 VSS.n2852 0.0680676
R5689 VSS.n2665 VSS.n627 0.0680676
R5690 VSS.n628 VSS.n627 0.0680676
R5691 VSS.n608 VSS.n602 0.0680676
R5692 VSS.n610 VSS.n608 0.0680676
R5693 VSS.n999 VSS.n991 0.0680676
R5694 VSS.n999 VSS.n992 0.0680676
R5695 VSS.n945 VSS.n937 0.0680676
R5696 VSS.n947 VSS.n945 0.0680676
R5697 VSS.n2635 VSS.n648 0.0680676
R5698 VSS.n649 VSS.n648 0.0680676
R5699 VSS.n1054 VSS.n970 0.0680676
R5700 VSS.n971 VSS.n970 0.0680676
R5701 VSS.n2453 VSS.n773 0.0680676
R5702 VSS.n2453 VSS.n2452 0.0680676
R5703 VSS.n2137 VSS.n2127 0.0680676
R5704 VSS.n2137 VSS.n2128 0.0680676
R5705 VSS.n1991 VSS.n1903 0.0680676
R5706 VSS.n1905 VSS.n1903 0.0680676
R5707 VSS.n2560 VSS.n2559 0.0680676
R5708 VSS.n2559 VSS.n691 0.0680676
R5709 VSS.n1518 VSS.n1468 0.0680676
R5710 VSS.n1518 VSS.n1517 0.0680676
R5711 VSS.n1440 VSS.n1371 0.0680676
R5712 VSS.n1441 VSS.n1440 0.0680676
R5713 VSS.n2590 VSS.n670 0.0680676
R5714 VSS.n2592 VSS.n2590 0.0680676
R5715 VSS.n2034 VSS.n2031 0.0680676
R5716 VSS.n2034 VSS.n2033 0.0680676
R5717 VSS.n921 VSS.n916 0.0680676
R5718 VSS.n923 VSS.n921 0.0680676
R5719 VSS.n2420 VSS.n2419 0.0680676
R5720 VSS.n2419 VSS.n785 0.0680676
R5721 VSS.n2332 VSS.n830 0.0680676
R5722 VSS.n2332 VSS.n824 0.0680676
R5723 VSS.n851 VSS.n849 0.0680676
R5724 VSS.n852 VSS.n851 0.0680676
R5725 VSS.n2504 VSS.n754 0.0680676
R5726 VSS.n2506 VSS.n2504 0.0680676
R5727 VSS.n806 VSS.n805 0.0680676
R5728 VSS.n805 VSS.n799 0.0680676
R5729 VSS.n1348 VSS.n1312 0.0680676
R5730 VSS.n1314 VSS.n1312 0.0680676
R5731 VSS.n2068 VSS.n2051 0.0680676
R5732 VSS.n2069 VSS.n2068 0.0680676
R5733 VSS.n869 VSS.n863 0.0680676
R5734 VSS.n871 VSS.n869 0.0680676
R5735 VSS.n2166 VSS.n2154 0.0680676
R5736 VSS.n2166 VSS.n2155 0.0680676
R5737 VSS.n2254 VSS.n2253 0.0680676
R5738 VSS.n2253 VSS.n893 0.0680676
R5739 VSS.n1280 VSS.n1220 0.0680676
R5740 VSS.n1280 VSS.n1279 0.0680676
R5741 VSS.n1243 VSS.n1242 0.0680676
R5742 VSS.n1242 VSS.n1232 0.0680676
R5743 VSS.n1959 VSS.n1922 0.0680676
R5744 VSS.n1959 VSS.n1958 0.0680676
R5745 VSS.n1706 VSS.n1551 0.0680676
R5746 VSS.n1706 VSS.n1550 0.0680676
R5747 VSS.n2952 VSS.n2951 0.0680676
R5748 VSS.n2951 VSS.n268 0.0680676
R5749 VSS.n2024 VSS 0.0669062
R5750 VSS.n1136 VSS.n1073 0.0656042
R5751 VSS.n2897 VSS.n510 0.0656042
R5752 VSS.n1698 VSS.n1697 0.0656042
R5753 VSS.n2736 VSS.n578 0.0656042
R5754 VSS.n2813 VSS.n2812 0.0656042
R5755 VSS.n1619 VSS.n1618 0.0656042
R5756 VSS.n632 VSS.n631 0.0656042
R5757 VSS.n944 VSS.n943 0.0656042
R5758 VSS.n1001 VSS.n997 0.0656042
R5759 VSS.n1020 VSS.n994 0.0656042
R5760 VSS.n1373 VSS.n1368 0.0656042
R5761 VSS.n2596 VSS.n671 0.0656042
R5762 VSS.n725 VSS.n719 0.0656042
R5763 VSS.n747 VSS.n716 0.0656042
R5764 VSS.n2343 VSS.n2342 0.0656042
R5765 VSS.n2428 VSS.n784 0.0656042
R5766 VSS.n2516 VSS.n2515 0.0656042
R5767 VSS.n2510 VSS.n2509 0.0656042
R5768 VSS.n2264 VSS.n892 0.0656042
R5769 VSS.n2035 VSS.n2032 0.0656042
R5770 VSS.n2168 VSS.n2164 0.0656042
R5771 VSS.n2187 VSS.n2157 0.0656042
R5772 VSS.n2020 VSS.n917 0.0656042
R5773 VSS.n1946 VSS.n1926 0.0656042
R5774 VSS.n2946 VSS.n270 0.0656042
R5775 VSS.n1770 VSS.n1764 0.0656042
R5776 VSS.n1872 VSS.n1871 0.0656042
R5777 VSS.n1868 VSS.n1867 0.0656042
R5778 VSS.n227 VSS 0.064875
R5779 VSS.n288 VSS 0.064875
R5780 VSS.n287 VSS 0.064875
R5781 VSS.n327 VSS 0.064875
R5782 VSS.n331 VSS 0.064875
R5783 VSS.n374 VSS 0.064875
R5784 VSS.n351 VSS 0.064875
R5785 VSS.n349 VSS 0.064875
R5786 VSS.n3179 VSS 0.064875
R5787 VSS.n3211 VSS 0.064875
R5788 VSS.n3160 VSS 0.064875
R5789 VSS.n3158 VSS 0.064875
R5790 VSS.n200 VSS 0.064875
R5791 VSS.n3139 VSS 0.064875
R5792 VSS.n3323 VSS 0.064875
R5793 VSS.n3213 VSS 0.064875
R5794 VSS.n1095 VSS 0.0643021
R5795 VSS.n2698 VSS 0.0643021
R5796 VSS.n2684 VSS 0.0643021
R5797 VSS.n1390 VSS 0.0643021
R5798 VSS.n845 VSS 0.0643021
R5799 VSS.n2290 VSS 0.0643021
R5800 VSS.n2061 VSS 0.0643021
R5801 VSS.n1240 VSS 0.0643021
R5802 VSS.n248 VSS 0.0643021
R5803 VSS.n2992 VSS.n2991 0.063797
R5804 VSS.n3007 VSS 0.063625
R5805 VSS.n2987 VSS.n233 0.0635047
R5806 VSS.n3005 VSS 0.063
R5807 VSS.n3371 VSS.n41 0.0616979
R5808 VSS.n3102 VSS.n211 0.0616979
R5809 VSS.n3318 VSS.n80 0.0616979
R5810 VSS.n59 VSS 0.0603958
R5811 VSS VSS.n3364 0.0603958
R5812 VSS.n3348 VSS 0.0603958
R5813 VSS.n3349 VSS 0.0603958
R5814 VSS VSS.n3355 0.0603958
R5815 VSS VSS.n36 0.0603958
R5816 VSS.n3382 VSS 0.0603958
R5817 VSS.n45 VSS 0.0603958
R5818 VSS.n5 VSS 0.0603958
R5819 VSS.n13 VSS 0.0603958
R5820 VSS.n14 VSS 0.0603958
R5821 VSS.n3397 VSS 0.0603958
R5822 VSS VSS.n3396 0.0603958
R5823 VSS VSS.n3395 0.0603958
R5824 VSS.n20 VSS 0.0603958
R5825 VSS.n3389 VSS 0.0603958
R5826 VSS VSS.n34 0.0603958
R5827 VSS.n3074 VSS 0.0603958
R5828 VSS.n3025 VSS 0.0603958
R5829 VSS.n3032 VSS 0.0603958
R5830 VSS VSS.n217 0.0603958
R5831 VSS.n3070 VSS 0.0603958
R5832 VSS.n3066 VSS 0.0603958
R5833 VSS VSS.n3065 0.0603958
R5834 VSS VSS.n3058 0.0603958
R5835 VSS VSS.n3041 0.0603958
R5836 VSS VSS.n3051 0.0603958
R5837 VSS.n3098 VSS 0.0603958
R5838 VSS.n3092 VSS 0.0603958
R5839 VSS.n3127 VSS 0.0603958
R5840 VSS VSS.n3126 0.0603958
R5841 VSS.n3120 VSS 0.0603958
R5842 VSS.n194 VSS 0.0603958
R5843 VSS VSS.n3111 0.0603958
R5844 VSS.n82 VSS 0.0603958
R5845 VSS VSS.n3311 0.0603958
R5846 VSS.n87 VSS 0.0603958
R5847 VSS.n88 VSS 0.0603958
R5848 VSS VSS.n3302 0.0603958
R5849 VSS.n3297 VSS 0.0603958
R5850 VSS VSS.n105 0.0603958
R5851 VSS.n3253 VSS 0.0603958
R5852 VSS.n3257 VSS 0.0603958
R5853 VSS.n3265 VSS 0.0603958
R5854 VSS.n3266 VSS 0.0603958
R5855 VSS VSS.n3270 0.0603958
R5856 VSS.n3271 VSS 0.0603958
R5857 VSS.n3272 VSS 0.0603958
R5858 VSS.n3277 VSS 0.0603958
R5859 VSS.n3278 VSS 0.0603958
R5860 VSS.n3290 VSS 0.0603958
R5861 VSS.n1110 VSS 0.0603958
R5862 VSS.n1120 VSS 0.0603958
R5863 VSS VSS.n1205 0.0603958
R5864 VSS VSS.n1204 0.0603958
R5865 VSS VSS.n1193 0.0603958
R5866 VSS VSS.n2873 0.0603958
R5867 VSS.n2870 VSS 0.0603958
R5868 VSS.n1641 VSS.n1640 0.0603958
R5869 VSS.n1641 VSS.n1638 0.0603958
R5870 VSS VSS.n1685 0.0603958
R5871 VSS.n2710 VSS 0.0603958
R5872 VSS.n2719 VSS 0.0603958
R5873 VSS.n2757 VSS 0.0603958
R5874 VSS.n2776 VSS.n2775 0.0603958
R5875 VSS.n2775 VSS.n558 0.0603958
R5876 VSS.n2786 VSS 0.0603958
R5877 VSS.n2839 VSS 0.0603958
R5878 VSS.n2849 VSS.n2848 0.0603958
R5879 VSS.n1615 VSS 0.0603958
R5880 VSS VSS.n1607 0.0603958
R5881 VSS.n1601 VSS 0.0603958
R5882 VSS VSS.n1600 0.0603958
R5883 VSS.n2679 VSS 0.0603958
R5884 VSS VSS.n2672 0.0603958
R5885 VSS VSS.n2641 0.0603958
R5886 VSS VSS.n2640 0.0603958
R5887 VSS VSS.n2629 0.0603958
R5888 VSS VSS.n1062 0.0603958
R5889 VSS.n976 VSS.n975 0.0603958
R5890 VSS.n975 VSS.n973 0.0603958
R5891 VSS.n1043 VSS 0.0603958
R5892 VSS VSS.n1037 0.0603958
R5893 VSS.n1028 VSS 0.0603958
R5894 VSS.n1407 VSS 0.0603958
R5895 VSS.n1411 VSS 0.0603958
R5896 VSS.n1420 VSS 0.0603958
R5897 VSS.n1422 VSS 0.0603958
R5898 VSS VSS.n1376 0.0603958
R5899 VSS VSS.n1366 0.0603958
R5900 VSS.n1526 VSS 0.0603958
R5901 VSS VSS.n1525 0.0603958
R5902 VSS VSS.n1475 0.0603958
R5903 VSS VSS.n1513 0.0603958
R5904 VSS.n2587 VSS 0.0603958
R5905 VSS.n677 VSS 0.0603958
R5906 VSS VSS.n677 0.0603958
R5907 VSS.n2583 VSS 0.0603958
R5908 VSS VSS.n2582 0.0603958
R5909 VSS VSS.n2573 0.0603958
R5910 VSS VSS.n2572 0.0603958
R5911 VSS.n686 VSS 0.0603958
R5912 VSS.n2557 VSS.n693 0.0603958
R5913 VSS.n2553 VSS.n693 0.0603958
R5914 VSS.n746 VSS 0.0603958
R5915 VSS.n742 VSS 0.0603958
R5916 VSS.n2309 VSS 0.0603958
R5917 VSS.n2324 VSS 0.0603958
R5918 VSS VSS.n813 0.0603958
R5919 VSS.n2370 VSS 0.0603958
R5920 VSS.n2371 VSS 0.0603958
R5921 VSS.n2390 VSS.n796 0.0603958
R5922 VSS.n2393 VSS.n796 0.0603958
R5923 VSS.n2394 VSS 0.0603958
R5924 VSS VSS.n2408 0.0603958
R5925 VSS.n2409 VSS 0.0603958
R5926 VSS.n2414 VSS 0.0603958
R5927 VSS.n2435 VSS 0.0603958
R5928 VSS.n2439 VSS 0.0603958
R5929 VSS.n2441 VSS 0.0603958
R5930 VSS.n2445 VSS 0.0603958
R5931 VSS.n2451 VSS.n767 0.0603958
R5932 VSS.n2463 VSS.n767 0.0603958
R5933 VSS VSS.n765 0.0603958
R5934 VSS.n2483 VSS 0.0603958
R5935 VSS.n2492 VSS 0.0603958
R5936 VSS.n2282 VSS 0.0603958
R5937 VSS.n879 VSS 0.0603958
R5938 VSS VSS.n884 0.0603958
R5939 VSS.n2271 VSS 0.0603958
R5940 VSS.n2251 VSS 0.0603958
R5941 VSS.n894 VSS 0.0603958
R5942 VSS.n2242 VSS 0.0603958
R5943 VSS VSS.n899 0.0603958
R5944 VSS.n901 VSS 0.0603958
R5945 VSS.n2055 VSS 0.0603958
R5946 VSS.n2056 VSS 0.0603958
R5947 VSS.n2073 VSS.n2048 0.0603958
R5948 VSS.n2074 VSS.n2073 0.0603958
R5949 VSS VSS.n2078 0.0603958
R5950 VSS.n2079 VSS 0.0603958
R5951 VSS VSS.n2040 0.0603958
R5952 VSS.n2088 VSS 0.0603958
R5953 VSS.n2115 VSS 0.0603958
R5954 VSS.n2123 VSS 0.0603958
R5955 VSS.n2232 VSS 0.0603958
R5956 VSS VSS.n2231 0.0603958
R5957 VSS.n2135 VSS 0.0603958
R5958 VSS.n2140 VSS.n2139 0.0603958
R5959 VSS.n2139 VSS.n2130 0.0603958
R5960 VSS VSS.n2217 0.0603958
R5961 VSS VSS.n2203 0.0603958
R5962 VSS.n1256 VSS 0.0603958
R5963 VSS.n1259 VSS 0.0603958
R5964 VSS.n1264 VSS 0.0603958
R5965 VSS.n1272 VSS 0.0603958
R5966 VSS.n1290 VSS 0.0603958
R5967 VSS.n1299 VSS 0.0603958
R5968 VSS VSS.n1304 0.0603958
R5969 VSS.n1305 VSS 0.0603958
R5970 VSS.n1355 VSS 0.0603958
R5971 VSS.n1342 VSS.n1318 0.0603958
R5972 VSS.n1342 VSS.n1341 0.0603958
R5973 VSS.n1338 VSS 0.0603958
R5974 VSS.n1336 VSS 0.0603958
R5975 VSS.n1333 VSS 0.0603958
R5976 VSS VSS.n1332 0.0603958
R5977 VSS VSS.n1325 0.0603958
R5978 VSS VSS.n2014 0.0603958
R5979 VSS.n2005 VSS 0.0603958
R5980 VSS.n2003 VSS 0.0603958
R5981 VSS.n1896 VSS 0.0603958
R5982 VSS.n1999 VSS 0.0603958
R5983 VSS.n1908 VSS.n1907 0.0603958
R5984 VSS.n1909 VSS.n1908 0.0603958
R5985 VSS.n1974 VSS 0.0603958
R5986 VSS.n1972 VSS 0.0603958
R5987 VSS.n1969 VSS 0.0603958
R5988 VSS VSS.n1968 0.0603958
R5989 VSS.n1961 VSS 0.0603958
R5990 VSS.n1945 VSS 0.0603958
R5991 VSS.n1942 VSS 0.0603958
R5992 VSS VSS.n1941 0.0603958
R5993 VSS VSS.n1928 0.0603958
R5994 VSS.n1936 VSS 0.0603958
R5995 VSS VSS.n2972 0.0603958
R5996 VSS VSS.n2957 0.0603958
R5997 VSS.n1738 VSS 0.0603958
R5998 VSS.n1753 VSS 0.0603958
R5999 VSS.n1794 VSS.n1733 0.0603958
R6000 VSS.n1794 VSS.n1793 0.0603958
R6001 VSS.n1720 VSS 0.0603958
R6002 VSS.n1724 VSS 0.0603958
R6003 VSS.n1817 VSS.n1816 0.0603958
R6004 VSS.n1817 VSS.n1716 0.0603958
R6005 VSS.n1833 VSS 0.0603958
R6006 VSS.n1835 VSS 0.0603958
R6007 VSS VSS.n1709 0.0603958
R6008 VSS.n3371 VSS.n3370 0.0590938
R6009 VSS VSS.n3388 0.0590938
R6010 VSS.n3043 VSS 0.0590938
R6011 VSS.n3102 VSS.n3101 0.0590938
R6012 VSS.n3318 VSS.n3317 0.0590938
R6013 VSS.n3294 VSS 0.0590938
R6014 VSS.n714 VSS.n712 0.0574697
R6015 VSS.n2892 VSS.n507 0.0574697
R6016 VSS.n1198 VSS.n1196 0.0574697
R6017 VSS.n1132 VSS.n1075 0.0574697
R6018 VSS.n1688 VSS.n1624 0.0574697
R6019 VSS.n2862 VSS.n525 0.0574697
R6020 VSS.n583 VSS.n580 0.0574697
R6021 VSS.n2689 VSS.n596 0.0574697
R6022 VSS.n1610 VSS.n1558 0.0574697
R6023 VSS.n2816 VSS.n549 0.0574697
R6024 VSS.n567 VSS.n564 0.0574697
R6025 VSS.n2851 VSS.n530 0.0574697
R6026 VSS.n2664 VSS.n2662 0.0574697
R6027 VSS.n609 VSS.n600 0.0574697
R6028 VSS.n1024 VSS.n1023 0.0574697
R6029 VSS.n946 VSS.n664 0.0574697
R6030 VSS.n2634 VSS.n2632 0.0574697
R6031 VSS.n1053 VSS.n1051 0.0574697
R6032 VSS.n771 VSS.n769 0.0574697
R6033 VSS.n2222 VSS.n2221 0.0574697
R6034 VSS.n1990 VSS.n1904 0.0574697
R6035 VSS.n2562 VSS.n2561 0.0574697
R6036 VSS.n2550 VSS.n2549 0.0574697
R6037 VSS.n1516 VSS.n1474 0.0574697
R6038 VSS.n1442 VSS.n1370 0.0574697
R6039 VSS.n2591 VSS.n668 0.0574697
R6040 VSS.n2029 VSS.n912 0.0574697
R6041 VSS.n922 VSS.n914 0.0574697
R6042 VSS.n2421 VSS.n786 0.0574697
R6043 VSS.n2424 VSS.n2423 0.0574697
R6044 VSS.n828 VSS.n825 0.0574697
R6045 VSS.n848 VSS.n847 0.0574697
R6046 VSS.n2505 VSS.n752 0.0574697
R6047 VSS.n803 VSS.n800 0.0574697
R6048 VSS.n1347 VSS.n1313 0.0574697
R6049 VSS.n2059 VSS.n2058 0.0574697
R6050 VSS.n2071 VSS.n2070 0.0574697
R6051 VSS.n2191 VSS.n2190 0.0574697
R6052 VSS.n2260 VSS.n2259 0.0574697
R6053 VSS.n1218 VSS.n1217 0.0574697
R6054 VSS.n1244 VSS.n1233 0.0574697
R6055 VSS.n1247 VSS.n1246 0.0574697
R6056 VSS.n1957 VSS.n1924 0.0574697
R6057 VSS.n1957 VSS.n1948 0.0574697
R6058 VSS.n232 VSS.n231 0.0574529
R6059 VSS VSS.n3338 0.0557885
R6060 VSS VSS.n3337 0.0557885
R6061 VSS VSS.n3336 0.0557885
R6062 VSS.n126 VSS 0.0557885
R6063 VSS.n128 VSS 0.0557885
R6064 VSS.n133 VSS 0.0557885
R6065 VSS.n138 VSS 0.0557885
R6066 VSS.n143 VSS 0.0557885
R6067 VSS.n148 VSS 0.0557885
R6068 VSS.n153 VSS 0.0557885
R6069 VSS.n158 VSS 0.0557885
R6070 VSS.n163 VSS 0.0557885
R6071 VSS.n168 VSS 0.0557885
R6072 VSS.n3232 VSS 0.0557885
R6073 VSS.n1128 VSS.n1073 0.0551875
R6074 VSS.n2901 VSS.n510 0.0551875
R6075 VSS.n1698 VSS.n1627 0.0551875
R6076 VSS.n1692 VSS.n1686 0.0551875
R6077 VSS.n2724 VSS.n578 0.0551875
R6078 VSS.n2813 VSS.n551 0.0551875
R6079 VSS.n1619 VSS.n1561 0.0551875
R6080 VSS.n1614 VSS.n1608 0.0551875
R6081 VSS.n631 VSS.n630 0.0551875
R6082 VSS.n944 VSS.n939 0.0551875
R6083 VSS.n997 VSS.n989 0.0551875
R6084 VSS.n1020 VSS.n1019 0.0551875
R6085 VSS.n2599 VSS.n671 0.0551875
R6086 VSS.n719 VSS.n710 0.0551875
R6087 VSS.n747 VSS.n746 0.0551875
R6088 VSS.n2342 VSS.n823 0.0551875
R6089 VSS.n2416 VSS.n784 0.0551875
R6090 VSS.n2516 VSS.n755 0.0551875
R6091 VSS.n2509 VSS.n2503 0.0551875
R6092 VSS.n2265 VSS.n2264 0.0551875
R6093 VSS.n2100 VSS.n2035 0.0551875
R6094 VSS.n2164 VSS.n2152 0.0551875
R6095 VSS.n2187 VSS.n2186 0.0551875
R6096 VSS.n2023 VSS.n917 0.0551875
R6097 VSS.n1946 VSS.n1945 0.0551875
R6098 VSS.n2949 VSS.n270 0.0551875
R6099 VSS.n1771 VSS.n1770 0.0551875
R6100 VSS.n1872 VSS.n1705 0.0551875
R6101 VSS.n1867 VSS.n1866 0.0551875
R6102 VSS.n3320 VSS 0.0527529
R6103 VSS VSS.n2030 0.0525833
R6104 VSS.n1282 VSS 0.0525833
R6105 VSS.n3320 VSS.n3319 0.0519696
R6106 VSS.n3234 VSS 0.0518289
R6107 VSS.n17 VSS.n14 0.0499792
R6108 VSS.n3071 VSS.n217 0.0499792
R6109 VSS.n3266 VSS.n111 0.0499792
R6110 VSS.n1099 VSS.n1096 0.0499792
R6111 VSS.n2869 VSS.n520 0.0499792
R6112 VSS.n2697 VSS.n2696 0.0499792
R6113 VSS.n2841 VSS.n531 0.0499792
R6114 VSS.n2683 VSS.n603 0.0499792
R6115 VSS.n1399 VSS.n1386 0.0499792
R6116 VSS.n2565 VSS.n2564 0.0499792
R6117 VSS.n850 VSS.n844 0.0499792
R6118 VSS.n2381 VSS.n807 0.0499792
R6119 VSS.n2447 VSS.n772 0.0499792
R6120 VSS.n2289 VSS.n864 0.0499792
R6121 VSS.n2062 VSS.n2052 0.0499792
R6122 VSS.n1239 VSS.n1231 0.0499792
R6123 VSS.n1351 VSS.n1350 0.0499792
R6124 VSS.n1900 VSS.n1898 0.0499792
R6125 VSS.n252 VSS.n241 0.0499792
R6126 VSS.n1725 VSS.n1724 0.0499792
R6127 VSS.n3381 VSS.n3374 0.0486771
R6128 VSS.n3110 VSS.n3105 0.0486771
R6129 VSS.n104 VSS.n96 0.0486771
R6130 VSS.n1097 VSS 0.047375
R6131 VSS.n2692 VSS 0.047375
R6132 VSS.n611 VSS 0.047375
R6133 VSS.n1387 VSS 0.047375
R6134 VSS VSS.n854 0.047375
R6135 VSS.n872 VSS 0.047375
R6136 VSS.n1250 VSS 0.047375
R6137 VSS.n253 VSS 0.047375
R6138 VSS.n3405 VSS 0.0460729
R6139 VSS VSS.n3073 0.0460729
R6140 VSS VSS.n3237 0.0460729
R6141 VSS.n1124 VSS.n1120 0.0447708
R6142 VSS.n2719 VSS.n584 0.0447708
R6143 VSS.n2672 VSS.n622 0.0447708
R6144 VSS.n1431 VSS.n1427 0.0447708
R6145 VSS.n2325 VSS.n829 0.0447708
R6146 VSS.n2269 VSS.n887 0.0447708
R6147 VSS.n1273 VSS.n1219 0.0447708
R6148 VSS.n2957 VSS.n2956 0.0447708
R6149 VSS.n3430 VSS.n3429 0.0423452
R6150 VSS.n3429 VSS.n3428 0.0423452
R6151 VSS.n3428 VSS.n3427 0.0423452
R6152 VSS.n3427 VSS.n3426 0.0423452
R6153 VSS.n3426 VSS.n3425 0.0423452
R6154 VSS.n3425 VSS.n3424 0.0423452
R6155 VSS.n3424 VSS.n3423 0.0423452
R6156 VSS.n3423 VSS.n3422 0.0423452
R6157 VSS.n3422 VSS.n3421 0.0423452
R6158 VSS.n3421 VSS.n3420 0.0423452
R6159 VSS.n3420 VSS.n3419 0.0423452
R6160 VSS.n3419 VSS.n3418 0.0423452
R6161 VSS.n3418 VSS.n3417 0.0423452
R6162 VSS.n3417 VSS.n3416 0.0423452
R6163 VSS.n3416 VSS.n3415 0.0423452
R6164 VSS.n3415 VSS.n3414 0.0423452
R6165 VSS.n3414 VSS.n3413 0.0423452
R6166 VSS.n3413 VSS.n3412 0.0423452
R6167 VSS.n3412 VSS.n3411 0.0423452
R6168 VSS.n3411 VSS.n3410 0.0423452
R6169 VSS.n3410 VSS.n3409 0.0423452
R6170 VSS.n3409 VSS.n3408 0.0423452
R6171 VSS.n1956 VSS.n1955 0.0422778
R6172 VSS.n2487 VSS 0.0421667
R6173 VSS VSS.n2165 0.0421667
R6174 VSS.n2019 VSS 0.0421667
R6175 VSS.n2016 VSS 0.0421667
R6176 VSS.n2990 VSS.n230 0.0416941
R6177 VSS.n1885 VSS.n1883 0.0414836
R6178 VSS.n1811 VSS.n1810 0.0410405
R6179 VSS.n1818 VSS.n1717 0.0410405
R6180 VSS.n250 VSS.n249 0.0410405
R6181 VSS.n238 VSS.n236 0.0410405
R6182 VSS.n1749 VSS.n1747 0.0410405
R6183 VSS.n1750 VSS.n1732 0.0410405
R6184 VSS.n1767 VSS.n1766 0.0410405
R6185 VSS.n1768 VSS.n501 0.0410405
R6186 VSS.n1391 VSS.n1385 0.0410405
R6187 VSS.n1401 VSS.n1383 0.0410405
R6188 VSS.n721 VSS.n711 0.0410405
R6189 VSS.n722 VSS.n715 0.0410405
R6190 VSS.n2903 VSS.n509 0.0410405
R6191 VSS.n2895 VSS.n2893 0.0410405
R6192 VSS.n1200 VSS.n1199 0.0410405
R6193 VSS.n1161 VSS.n1160 0.0410405
R6194 VSS.n1121 VSS.n1076 0.0410405
R6195 VSS.n1131 VSS.n1074 0.0410405
R6196 VSS.n1094 VSS.n1089 0.0410405
R6197 VSS.n1101 VSS.n1087 0.0410405
R6198 VSS.n1699 VSS.n1626 0.0410405
R6199 VSS.n1690 VSS.n1689 0.0410405
R6200 VSS.n2864 VSS.n2863 0.0410405
R6201 VSS.n1642 VSS.n1639 0.0410405
R6202 VSS.n2729 VSS.n585 0.0410405
R6203 VSS.n2725 VSS.n579 0.0410405
R6204 VSS.n2699 VSS.n2691 0.0410405
R6205 VSS.n2694 VSS.n595 0.0410405
R6206 VSS.n1620 VSS.n1560 0.0410405
R6207 VSS.n1612 VSS.n1611 0.0410405
R6208 VSS.n2803 VSS.n550 0.0410405
R6209 VSS.n2815 VSS.n548 0.0410405
R6210 VSS.n2769 VSS.n569 0.0410405
R6211 VSS.n2763 VSS.n563 0.0410405
R6212 VSS.n2856 VSS.n532 0.0410405
R6213 VSS.n2852 VSS.n2850 0.0410405
R6214 VSS.n2666 VSS.n2665 0.0410405
R6215 VSS.n629 VSS.n628 0.0410405
R6216 VSS.n2685 VSS.n602 0.0410405
R6217 VSS.n612 VSS.n610 0.0410405
R6218 VSS.n991 VSS.n990 0.0410405
R6219 VSS.n993 VSS.n992 0.0410405
R6220 VSS.n937 VSS.n663 0.0410405
R6221 VSS.n948 VSS.n947 0.0410405
R6222 VSS.n2636 VSS.n2635 0.0410405
R6223 VSS.n650 VSS.n649 0.0410405
R6224 VSS.n1055 VSS.n1054 0.0410405
R6225 VSS.n972 VSS.n971 0.0410405
R6226 VSS.n2456 VSS.n773 0.0410405
R6227 VSS.n2452 VSS.n768 0.0410405
R6228 VSS.n2127 VSS.n2126 0.0410405
R6229 VSS.n2129 VSS.n2128 0.0410405
R6230 VSS.n1992 VSS.n1991 0.0410405
R6231 VSS.n1906 VSS.n1905 0.0410405
R6232 VSS.n2560 VSS.n688 0.0410405
R6233 VSS.n2548 VSS.n691 0.0410405
R6234 VSS.n1471 VSS.n1468 0.0410405
R6235 VSS.n1517 VSS.n1469 0.0410405
R6236 VSS.n1428 VSS.n1371 0.0410405
R6237 VSS.n1441 VSS.n1369 0.0410405
R6238 VSS.n2601 VSS.n670 0.0410405
R6239 VSS.n2594 VSS.n2592 0.0410405
R6240 VSS.n2102 VSS.n2031 0.0410405
R6241 VSS.n2033 VSS.n911 0.0410405
R6242 VSS.n2025 VSS.n916 0.0410405
R6243 VSS.n2018 VSS.n923 0.0410405
R6244 VSS.n2420 VSS.n2418 0.0410405
R6245 VSS.n2426 VSS.n785 0.0410405
R6246 VSS.n2335 VSS.n830 0.0410405
R6247 VSS.n2341 VSS.n824 0.0410405
R6248 VSS.n849 VSS.n846 0.0410405
R6249 VSS.n853 VSS.n852 0.0410405
R6250 VSS.n2517 VSS.n754 0.0410405
R6251 VSS.n2507 VSS.n2506 0.0410405
R6252 VSS.n2382 VSS.n806 0.0410405
R6253 VSS.n2388 VSS.n799 0.0410405
R6254 VSS.n1349 VSS.n1348 0.0410405
R6255 VSS.n1315 VSS.n1314 0.0410405
R6256 VSS.n2057 VSS.n2051 0.0410405
R6257 VSS.n2069 VSS.n2049 0.0410405
R6258 VSS.n2291 VSS.n863 0.0410405
R6259 VSS.n873 VSS.n871 0.0410405
R6260 VSS.n2154 VSS.n2153 0.0410405
R6261 VSS.n2156 VSS.n2155 0.0410405
R6262 VSS.n2256 VSS.n2254 0.0410405
R6263 VSS.n2263 VSS.n893 0.0410405
R6264 VSS.n1283 VSS.n1220 0.0410405
R6265 VSS.n1279 VSS.n1216 0.0410405
R6266 VSS.n1243 VSS.n1241 0.0410405
R6267 VSS.n1249 VSS.n1232 0.0410405
R6268 VSS.n1951 VSS.n1922 0.0410405
R6269 VSS.n1958 VSS.n1923 0.0410405
R6270 VSS.n1873 VSS.n1551 0.0410405
R6271 VSS.n1846 VSS.n1550 0.0410405
R6272 VSS.n2952 VSS.n266 0.0410405
R6273 VSS.n2941 VSS.n268 0.0410405
R6274 VSS.n1554 VSS.n1553 0.0393869
R6275 VSS.n2849 VSS 0.0382604
R6276 VSS.n1105 VSS 0.0369583
R6277 VSS.n2705 VSS 0.0369583
R6278 VSS VSS.n2854 0.0369583
R6279 VSS.n614 VSS 0.0369583
R6280 VSS.n974 VSS 0.0369583
R6281 VSS.n1405 VSS 0.0369583
R6282 VSS.n855 VSS 0.0369583
R6283 VSS.n2462 VSS 0.0369583
R6284 VSS.n875 VSS 0.0369583
R6285 VSS.n2218 VSS 0.0369583
R6286 VSS VSS.n1229 0.0369583
R6287 VSS.n2981 VSS 0.0369583
R6288 VSS.n1878 VSS.n1877 0.0352656
R6289 VSS.n210 VSS 0.0346243
R6290 VSS.n3404 VSS 0.0343542
R6291 VSS VSS.n216 0.0343542
R6292 VSS VSS.n3256 0.0343542
R6293 VSS.n1096 VSS.n1095 0.0343542
R6294 VSS.n1202 VSS.n1153 0.0343542
R6295 VSS.n2698 VSS.n2697 0.0343542
R6296 VSS.n2762 VSS.n568 0.0343542
R6297 VSS.n2684 VSS.n2683 0.0343542
R6298 VSS.n2638 VSS.n642 0.0343542
R6299 VSS.n1390 VSS.n1386 0.0343542
R6300 VSS.n1407 VSS 0.0343542
R6301 VSS.n1470 VSS.n1462 0.0343542
R6302 VSS.n845 VSS.n844 0.0343542
R6303 VSS VSS.n2307 0.0343542
R6304 VSS.n807 VSS.n804 0.0343542
R6305 VSS.n2290 VSS.n2289 0.0343542
R6306 VSS.n2285 VSS 0.0343542
R6307 VSS.n2062 VSS.n2061 0.0343542
R6308 VSS.n2080 VSS 0.0343542
R6309 VSS.n2232 VSS 0.0343542
R6310 VSS.n1240 VSS.n1239 0.0343542
R6311 VSS.n1351 VSS.n1307 0.0343542
R6312 VSS.n248 VSS.n241 0.0343542
R6313 VSS.n1745 VSS.n1744 0.0343542
R6314 VSS.n1721 VSS 0.0343542
R6315 VSS VSS.n3348 0.0330521
R6316 VSS VSS.n13 0.0330521
R6317 VSS.n3032 VSS 0.0330521
R6318 VSS.n3127 VSS 0.0330521
R6319 VSS VSS.n87 0.0330521
R6320 VSS VSS.n3265 0.0330521
R6321 VSS.n1206 VSS 0.0330521
R6322 VSS.n2874 VSS 0.0330521
R6323 VSS.n2753 VSS 0.0330521
R6324 VSS.n2832 VSS 0.0330521
R6325 VSS.n2642 VSS 0.0330521
R6326 VSS.n1063 VSS 0.0330521
R6327 VSS VSS.n1373 0.0330521
R6328 VSS.n1526 VSS 0.0330521
R6329 VSS.n2573 VSS 0.0330521
R6330 VSS VSS.n2370 0.0330521
R6331 VSS VSS.n901 0.0330521
R6332 VSS VSS.n2123 0.0330521
R6333 VSS VSS.n1305 0.0330521
R6334 VSS VSS.n1896 0.0330521
R6335 VSS.n1950 VSS 0.0330521
R6336 VSS VSS.n279 0.0330521
R6337 VSS VSS.n494 0.0330521
R6338 VSS VSS.n37 0.03175
R6339 VSS.n3112 VSS 0.03175
R6340 VSS.n106 VSS 0.03175
R6341 VSS.n1205 VSS 0.03175
R6342 VSS.n1686 VSS 0.03175
R6343 VSS.n2641 VSS 0.03175
R6344 VSS.n1028 VSS 0.03175
R6345 VSS VSS.n1027 0.03175
R6346 VSS VSS.n1406 0.03175
R6347 VSS.n2583 VSS 0.03175
R6348 VSS.n2572 VSS 0.03175
R6349 VSS VSS.n2055 0.03175
R6350 VSS.n2101 VSS 0.03175
R6351 VSS VSS.n2194 0.03175
R6352 VSS VSS.n1281 0.03175
R6353 VSS.n1278 VSS 0.03175
R6354 VSS.n1333 VSS 0.03175
R6355 VSS.n2015 VSS 0.03175
R6356 VSS.n1969 VSS 0.03175
R6357 VSS.n1942 VSS 0.03175
R6358 VSS.n1881 VSS.n1548 0.0308279
R6359 VSS.n3338 VSS 0.0305481
R6360 VSS.n3337 VSS 0.0305481
R6361 VSS.n3336 VSS 0.0305481
R6362 VSS VSS.n126 0.0305481
R6363 VSS VSS.n3232 0.0305481
R6364 VSS.n1990 VSS.n1989 0.0292489
R6365 VSS.n1987 VSS.n1904 0.0292489
R6366 VSS.n2223 VSS.n2222 0.0292489
R6367 VSS.n2221 VSS.n2220 0.0292489
R6368 VSS.n2458 VSS.n771 0.0292489
R6369 VSS.n2460 VSS.n769 0.0292489
R6370 VSS.n1053 VSS.n1052 0.0292489
R6371 VSS.n1051 VSS.n1050 0.0292489
R6372 VSS.n2858 VSS.n530 0.0292489
R6373 VSS.n2851 VSS.n528 0.0292489
R6374 VSS.n2862 VSS.n2861 0.0292489
R6375 VSS.n527 VSS.n525 0.0292489
R6376 VSS.n2549 VSS.n690 0.0292489
R6377 VSS.n2561 VSS.n690 0.0292489
R6378 VSS.n2027 VSS.n914 0.0292489
R6379 VSS.n922 VSS.n913 0.0292489
R6380 VSS.n2104 VSS.n2029 0.0292489
R6381 VSS.n2106 VSS.n912 0.0292489
R6382 VSS.n2603 VSS.n668 0.0292489
R6383 VSS.n2591 VSS.n666 0.0292489
R6384 VSS.n2606 VSS.n664 0.0292489
R6385 VSS.n946 VSS.n665 0.0292489
R6386 VSS.n2804 VSS.n549 0.0292489
R6387 VSS.n2817 VSS.n2816 0.0292489
R6388 VSS.n2905 VSS.n507 0.0292489
R6389 VSS.n2892 VSS.n505 0.0292489
R6390 VSS.n2423 VSS.n2422 0.0292489
R6391 VSS.n2422 VSS.n2421 0.0292489
R6392 VSS.n1347 VSS.n1346 0.0292489
R6393 VSS.n1344 VSS.n1313 0.0292489
R6394 VSS.n2384 VSS.n803 0.0292489
R6395 VSS.n2386 VSS.n800 0.0292489
R6396 VSS.n1474 VSS.n1473 0.0292489
R6397 VSS.n1516 VSS.n1515 0.0292489
R6398 VSS.n2634 VSS.n2633 0.0292489
R6399 VSS.n2632 VSS.n2631 0.0292489
R6400 VSS.n2771 VSS.n567 0.0292489
R6401 VSS.n2773 VSS.n564 0.0292489
R6402 VSS.n1198 VSS.n1197 0.0292489
R6403 VSS.n1196 VSS.n1195 0.0292489
R6404 VSS.n2070 VSS.n2050 0.0292489
R6405 VSS.n2058 VSS.n2050 0.0292489
R6406 VSS.n1285 VSS.n1218 0.0292489
R6407 VSS.n1287 VSS.n1217 0.0292489
R6408 VSS.n2259 VSS.n2258 0.0292489
R6409 VSS.n2261 VSS.n2260 0.0292489
R6410 VSS.n2337 VSS.n828 0.0292489
R6411 VSS.n2339 VSS.n825 0.0292489
R6412 VSS.n1429 VSS.n1370 0.0292489
R6413 VSS.n1443 VSS.n1442 0.0292489
R6414 VSS.n2664 VSS.n2663 0.0292489
R6415 VSS.n2662 VSS.n2661 0.0292489
R6416 VSS.n2731 VSS.n583 0.0292489
R6417 VSS.n2733 VSS.n580 0.0292489
R6418 VSS.n1122 VSS.n1075 0.0292489
R6419 VSS.n1133 VSS.n1132 0.0292489
R6420 VSS.n2297 VSS.n847 0.0292489
R6421 VSS.n857 VSS.n848 0.0292489
R6422 VSS.n2687 VSS.n600 0.0292489
R6423 VSS.n609 VSS.n598 0.0292489
R6424 VSS.n2701 VSS.n2689 0.0292489
R6425 VSS.n2703 VSS.n596 0.0292489
R6426 VSS.n1246 VSS.n1245 0.0292489
R6427 VSS.n1245 VSS.n1244 0.0292489
R6428 VSS.n2192 VSS.n2191 0.0292489
R6429 VSS.n2190 VSS.n2189 0.0292489
R6430 VSS.n2519 VSS.n752 0.0292489
R6431 VSS.n2505 VSS.n750 0.0292489
R6432 VSS.n2522 VSS.n712 0.0292489
R6433 VSS.n749 VSS.n714 0.0292489
R6434 VSS.n1025 VSS.n1024 0.0292489
R6435 VSS.n1023 VSS.n1022 0.0292489
R6436 VSS.n1622 VSS.n1558 0.0292489
R6437 VSS.n1610 VSS.n1557 0.0292489
R6438 VSS.n1701 VSS.n1624 0.0292489
R6439 VSS.n1688 VSS.n1556 0.0292489
R6440 VSS.n1129 VSS.n1128 0.0291458
R6441 VSS.n2902 VSS.n2901 0.0291458
R6442 VSS.n1627 VSS.n1625 0.0291458
R6443 VSS.n2727 VSS.n2724 0.0291458
R6444 VSS.n2802 VSS.n551 0.0291458
R6445 VSS.n1561 VSS.n1559 0.0291458
R6446 VSS.n630 VSS.n625 0.0291458
R6447 VSS.n939 VSS.n938 0.0291458
R6448 VSS.n1027 VSS.n989 0.0291458
R6449 VSS.n1439 VSS.n1438 0.0291458
R6450 VSS.n2600 VSS.n2599 0.0291458
R6451 VSS.n2524 VSS.n710 0.0291458
R6452 VSS.n2333 VSS.n823 0.0291458
R6453 VSS.n2417 VSS.n2416 0.0291458
R6454 VSS.n755 VSS.n753 0.0291458
R6455 VSS.n2265 VSS.n891 0.0291458
R6456 VSS.n2101 VSS.n2100 0.0291458
R6457 VSS.n2194 VSS.n2152 0.0291458
R6458 VSS.n1281 VSS.n1278 0.0291458
R6459 VSS.n2024 VSS.n2023 0.0291458
R6460 VSS.n1949 VSS.n1918 0.0291458
R6461 VSS.n2950 VSS.n2949 0.0291458
R6462 VSS.n1771 VSS.n1763 0.0291458
R6463 VSS.n1705 VSS.n1704 0.0291458
R6464 VSS.n1953 VSS.n1924 0.0290783
R6465 VSS VSS.n1201 0.0278438
R6466 VSS.n2768 VSS 0.0278438
R6467 VSS VSS.n2637 0.0278438
R6468 VSS.n1466 VSS 0.0278438
R6469 VSS VSS.n2225 0.0278438
R6470 VSS.n1746 VSS 0.0278438
R6471 VSS.n1470 VSS 0.0265417
R6472 VSS VSS.n1254 0.0252396
R6473 VSS VSS.n1272 0.0252396
R6474 VSS.n1299 VSS 0.0252396
R6475 VSS.n1338 VSS 0.0252396
R6476 VSS.n2005 VSS 0.0252396
R6477 VSS.n1974 VSS 0.0252396
R6478 VSS.n1941 VSS 0.0252396
R6479 VSS VSS.n1833 0.0252396
R6480 VSS.n2907 VSS.n503 0.0250071
R6481 VSS.n1876 VSS.n1875 0.024993
R6482 VSS.n1165 VSS.n1164 0.0239375
R6483 VSS.n1640 VSS.n522 0.0239375
R6484 VSS.n1644 VSS.n1638 0.0239375
R6485 VSS.n2776 VSS.n562 0.0239375
R6486 VSS.n2854 VSS.n534 0.0239375
R6487 VSS.n2848 VSS.n536 0.0239375
R6488 VSS.n654 VSS.n653 0.0239375
R6489 VSS.n976 VSS.n974 0.0239375
R6490 VSS.n1048 VSS.n973 0.0239375
R6491 VSS.n1406 VSS.n1405 0.0239375
R6492 VSS.n1475 VSS.n1467 0.0239375
R6493 VSS.n2558 VSS.n2557 0.0239375
R6494 VSS.n2553 VSS.n2552 0.0239375
R6495 VSS.n855 VSS.n841 0.0239375
R6496 VSS.n2390 VSS.n2389 0.0239375
R6497 VSS VSS.n2394 0.0239375
R6498 VSS.n2454 VSS.n2451 0.0239375
R6499 VSS.n2463 VSS.n2462 0.0239375
R6500 VSS.n2492 VSS 0.0239375
R6501 VSS.n2286 VSS.n875 0.0239375
R6502 VSS.n2271 VSS 0.0239375
R6503 VSS.n2066 VSS.n2048 0.0239375
R6504 VSS.n2140 VSS.n2138 0.0239375
R6505 VSS.n2218 VSS.n2130 0.0239375
R6506 VSS.n1254 VSS.n1229 0.0239375
R6507 VSS VSS.n1277 0.0239375
R6508 VSS.n1318 VSS.n1317 0.0239375
R6509 VSS.n1907 VSS.n1901 0.0239375
R6510 VSS.n1985 VSS.n1909 0.0239375
R6511 VSS.n2981 VSS.n2980 0.0239375
R6512 VSS.n1736 VSS.n1733 0.0239375
R6513 VSS.n1816 VSS.n1718 0.0239375
R6514 VSS.n1820 VSS.n1716 0.0239375
R6515 VSS.n3370 VSS 0.0226354
R6516 VSS.n3365 VSS 0.0226354
R6517 VSS VSS.n62 0.0226354
R6518 VSS.n3356 VSS 0.0226354
R6519 VSS.n3351 VSS 0.0226354
R6520 VSS.n3377 VSS 0.0226354
R6521 VSS.n5 VSS 0.0226354
R6522 VSS VSS.n12 0.0226354
R6523 VSS.n3396 VSS 0.0226354
R6524 VSS VSS.n19 0.0226354
R6525 VSS.n35 VSS 0.0226354
R6526 VSS.n27 VSS 0.0226354
R6527 VSS.n3025 VSS 0.0226354
R6528 VSS VSS.n3031 0.0226354
R6529 VSS.n3066 VSS 0.0226354
R6530 VSS.n3059 VSS 0.0226354
R6531 VSS.n3052 VSS 0.0226354
R6532 VSS.n3101 VSS 0.0226354
R6533 VSS VSS.n3086 0.0226354
R6534 VSS.n3088 VSS 0.0226354
R6535 VSS VSS.n190 0.0226354
R6536 VSS VSS.n193 0.0226354
R6537 VSS.n3317 VSS 0.0226354
R6538 VSS.n3312 VSS 0.0226354
R6539 VSS VSS.n85 0.0226354
R6540 VSS.n3303 VSS 0.0226354
R6541 VSS VSS.n91 0.0226354
R6542 VSS.n100 VSS 0.0226354
R6543 VSS.n3257 VSS 0.0226354
R6544 VSS VSS.n3264 0.0226354
R6545 VSS VSS.n3271 0.0226354
R6546 VSS VSS.n3276 0.0226354
R6547 VSS.n3293 VSS 0.0226354
R6548 VSS.n3283 VSS 0.0226354
R6549 VSS VSS.n1152 0.0226354
R6550 VSS.n1202 VSS 0.0226354
R6551 VSS.n1165 VSS 0.0226354
R6552 VSS VSS.n1171 0.0226354
R6553 VSS.n2877 VSS 0.0226354
R6554 VSS.n2873 VSS 0.0226354
R6555 VSS.n1655 VSS 0.0226354
R6556 VSS.n1693 VSS 0.0226354
R6557 VSS.n1679 VSS 0.0226354
R6558 VSS VSS.n2752 0.0226354
R6559 VSS VSS.n2762 0.0226354
R6560 VSS VSS.n2785 0.0226354
R6561 VSS.n2797 VSS 0.0226354
R6562 VSS VSS.n2820 0.0226354
R6563 VSS.n2833 VSS 0.0226354
R6564 VSS VSS.n534 0.0226354
R6565 VSS.n1608 VSS 0.0226354
R6566 VSS.n1600 VSS 0.0226354
R6567 VSS.n2646 VSS 0.0226354
R6568 VSS.n2638 VSS 0.0226354
R6569 VSS.n654 VSS 0.0226354
R6570 VSS VSS.n660 0.0226354
R6571 VSS VSS.n964 0.0226354
R6572 VSS.n1062 VSS 0.0226354
R6573 VSS.n1036 VSS 0.0226354
R6574 VSS VSS.n987 0.0226354
R6575 VSS VSS.n1005 0.0226354
R6576 VSS.n1417 VSS 0.0226354
R6577 VSS VSS.n1420 0.0226354
R6578 VSS.n1438 VSS 0.0226354
R6579 VSS.n1446 VSS 0.0226354
R6580 VSS VSS.n1460 0.0226354
R6581 VSS.n1524 VSS 0.0226354
R6582 VSS VSS.n1462 0.0226354
R6583 VSS.n1513 VSS 0.0226354
R6584 VSS.n2574 VSS 0.0226354
R6585 VSS VSS.n686 0.0226354
R6586 VSS VSS.n702 0.0226354
R6587 VSS.n735 VSS 0.0226354
R6588 VSS VSS.n2323 0.0226354
R6589 VSS.n2354 VSS 0.0226354
R6590 VSS.n2365 VSS 0.0226354
R6591 VSS VSS.n2393 0.0226354
R6592 VSS VSS.n2409 0.0226354
R6593 VSS.n2410 VSS 0.0226354
R6594 VSS.n2441 VSS 0.0226354
R6595 VSS VSS.n2482 0.0226354
R6596 VSS VSS.n2488 0.0226354
R6597 VSS.n2282 VSS 0.0226354
R6598 VSS.n2281 VSS 0.0226354
R6599 VSS VSS.n894 0.0226354
R6600 VSS.n2245 VSS 0.0226354
R6601 VSS VSS.n2056 0.0226354
R6602 VSS VSS.n2087 0.0226354
R6603 VSS VSS.n2088 0.0226354
R6604 VSS VSS.n2114 0.0226354
R6605 VSS VSS.n2122 0.0226354
R6606 VSS.n2231 VSS 0.0226354
R6607 VSS.n2226 VSS 0.0226354
R6608 VSS.n2204 VSS 0.0226354
R6609 VSS.n2195 VSS 0.0226354
R6610 VSS VSS.n2173 0.0226354
R6611 VSS VSS.n1271 0.0226354
R6612 VSS.n1341 VSS 0.0226354
R6613 VSS.n2008 VSS 0.0226354
R6614 VSS VSS.n1910 0.0226354
R6615 VSS VSS.n1918 0.0226354
R6616 VSS.n1931 VSS 0.0226354
R6617 VSS.n2973 VSS 0.0226354
R6618 VSS.n2958 VSS 0.0226354
R6619 VSS.n2929 VSS 0.0226354
R6620 VSS VSS.n1745 0.0226354
R6621 VSS.n2922 VSS 0.0226354
R6622 VSS.n1830 VSS 0.0226354
R6623 VSS.n1860 VSS 0.0226354
R6624 VSS.n1852 VSS 0.0226354
R6625 VSS.n3233 VSS 0.0219286
R6626 VSS.n1803 VSS.n1802 0.0218125
R6627 VSS.n1956 VSS.n1954 0.0213889
R6628 VSS.n1955 VSS 0.0213889
R6629 VSS.n1047 VSS 0.0213333
R6630 VSS VSS.n2439 0.0213333
R6631 VSS VSS.n128 0.0209327
R6632 VSS.n130 VSS 0.0209327
R6633 VSS VSS.n133 0.0209327
R6634 VSS.n135 VSS 0.0209327
R6635 VSS VSS.n138 0.0209327
R6636 VSS.n140 VSS 0.0209327
R6637 VSS VSS.n143 0.0209327
R6638 VSS.n145 VSS 0.0209327
R6639 VSS VSS.n148 0.0209327
R6640 VSS.n150 VSS 0.0209327
R6641 VSS VSS.n153 0.0209327
R6642 VSS.n155 VSS 0.0209327
R6643 VSS VSS.n158 0.0209327
R6644 VSS.n160 VSS 0.0209327
R6645 VSS VSS.n163 0.0209327
R6646 VSS.n165 VSS 0.0209327
R6647 VSS VSS.n168 0.0209327
R6648 VSS.n170 VSS 0.0209327
R6649 VSS.n1090 VSS 0.0200312
R6650 VSS VSS.n2690 0.0200312
R6651 VSS VSS.n601 0.0200312
R6652 VSS.n1396 VSS 0.0200312
R6653 VSS.n2299 VSS 0.0200312
R6654 VSS VSS.n862 0.0200312
R6655 VSS.n1235 VSS 0.0200312
R6656 VSS.n1261 VSS 0.0200312
R6657 VSS VSS.n247 0.0200312
R6658 VSS.n1136 VSS.n1135 0.0187292
R6659 VSS.n2897 VSS.n2896 0.0187292
R6660 VSS.n2890 VSS.n2889 0.0187292
R6661 VSS.n1697 VSS.n1628 0.0187292
R6662 VSS.n1693 VSS.n1669 0.0187292
R6663 VSS.n2736 VSS.n2735 0.0187292
R6664 VSS.n2812 VSS.n547 0.0187292
R6665 VSS.n2820 VSS.n2819 0.0187292
R6666 VSS.n1618 VSS.n1562 0.0187292
R6667 VSS.n1615 VSS.n1591 0.0187292
R6668 VSS.n2659 VSS.n632 0.0187292
R6669 VSS.n943 VSS.n936 0.0187292
R6670 VSS.n951 VSS.n950 0.0187292
R6671 VSS.n1001 VSS.n1000 0.0187292
R6672 VSS.n998 VSS.n994 0.0187292
R6673 VSS.n1445 VSS.n1368 0.0187292
R6674 VSS.n2596 VSS.n2595 0.0187292
R6675 VSS.n2589 VSS.n2588 0.0187292
R6676 VSS.n725 VSS.n724 0.0187292
R6677 VSS.n720 VSS.n716 0.0187292
R6678 VSS.n2343 VSS.n820 0.0187292
R6679 VSS.n2428 VSS.n2427 0.0187292
R6680 VSS.n2433 VSS.n782 0.0187292
R6681 VSS.n2515 VSS.n756 0.0187292
R6682 VSS.n2510 VSS.n2487 0.0187292
R6683 VSS.n2252 VSS.n892 0.0187292
R6684 VSS.n2032 VSS.n910 0.0187292
R6685 VSS.n2109 VSS.n2108 0.0187292
R6686 VSS.n2168 VSS.n2167 0.0187292
R6687 VSS.n2165 VSS.n2157 0.0187292
R6688 VSS.n1290 VSS.n1289 0.0187292
R6689 VSS.n2020 VSS.n2019 0.0187292
R6690 VSS.n2016 VSS.n2015 0.0187292
R6691 VSS.n1961 VSS.n1960 0.0187292
R6692 VSS.n1926 VSS.n1925 0.0187292
R6693 VSS.n2946 VSS.n2945 0.0187292
R6694 VSS.n1764 VSS.n500 0.0187292
R6695 VSS.n2911 VSS.n2910 0.0187292
R6696 VSS.n1871 VSS.n1707 0.0187292
R6697 VSS.n1868 VSS.n1847 0.0187292
R6698 VSS.n1800 VSS.n1799 0.0183038
R6699 VSS.n1801 VSS.n1798 0.0182893
R6700 VSS VSS.n915 0.0174271
R6701 VSS.n472 VSS.n471 0.0158654
R6702 VSS.n3405 VSS.n3404 0.0148229
R6703 VSS.n3073 VSS.n216 0.0148229
R6704 VSS.n3256 VSS.n3237 0.0148229
R6705 VSS VSS.n508 0.0148229
R6706 VSS.n2608 VSS 0.0148229
R6707 VSS.n2986 VSS 0.0140546
R6708 VSS.n1954 VSS 0.0135556
R6709 VSS.n1098 VSS.n1097 0.0135208
R6710 VSS.n1163 VSS.n1157 0.0135208
R6711 VSS.n2866 VSS.n2865 0.0135208
R6712 VSS.n2693 VSS.n2692 0.0135208
R6713 VSS.n2767 VSS.n2765 0.0135208
R6714 VSS.n2855 VSS.n533 0.0135208
R6715 VSS.n611 VSS.n605 0.0135208
R6716 VSS.n652 VSS.n646 0.0135208
R6717 VSS.n1057 VSS.n1056 0.0135208
R6718 VSS.n1398 VSS.n1387 0.0135208
R6719 VSS.n1520 VSS.n1519 0.0135208
R6720 VSS.n692 VSS.n687 0.0135208
R6721 VSS.n854 VSS.n843 0.0135208
R6722 VSS.n2380 VSS.n798 0.0135208
R6723 VSS.n2455 VSS.n2450 0.0135208
R6724 VSS.n872 VSS.n866 0.0135208
R6725 VSS.n2067 VSS.n2065 0.0135208
R6726 VSS.n2136 VSS.n2135 0.0135208
R6727 VSS.n1251 VSS.n1250 0.0135208
R6728 VSS.n1316 VSS.n1310 0.0135208
R6729 VSS.n1994 VSS.n1993 0.0135208
R6730 VSS.n254 VSS.n253 0.0135208
R6731 VSS.n1753 VSS.n1752 0.0135208
R6732 VSS.n1813 VSS.n1812 0.0135208
R6733 VSS.n2225 VSS 0.0109167
R6734 VSS.n1746 VSS 0.0109167
R6735 VSS.n2855 VSS 0.00961458
R6736 VSS.n1056 VSS 0.00961458
R6737 VSS.n1402 VSS.n1384 0.00878194
R6738 VSS.n1102 VSS.n1088 0.00878194
R6739 VSS.n870 VSS.n860 0.00878194
R6740 VSS.n242 VSS.n235 0.00838554
R6741 VSS.n2984 VSS.n2983 0.00838554
R6742 VSS.n1125 VSS.n1077 0.0083125
R6743 VSS.n2728 VSS.n586 0.0083125
R6744 VSS.n2807 VSS.n2806 0.0083125
R6745 VSS.n2668 VSS.n2667 0.0083125
R6746 VSS.n1432 VSS.n1372 0.0083125
R6747 VSS.n1489 VSS.n669 0.0083125
R6748 VSS.n2334 VSS.n2331 0.0083125
R6749 VSS.n2415 VSS.n2414 0.0083125
R6750 VSS.n2255 VSS.n889 0.0083125
R6751 VSS.n2094 VSS.n2030 0.0083125
R6752 VSS.n1282 VSS.n1276 0.0083125
R6753 VSS.n1325 VSS.n915 0.0083125
R6754 VSS.n269 VSS.n265 0.0083125
R6755 VSS.n1774 VSS.n1761 0.0083125
R6756 VSS.n1886 VSS.n1881 0.00808197
R6757 VSS.n2985 VSS.n235 0.00790157
R6758 VSS.n2985 VSS.n2984 0.00790157
R6759 VSS.n1988 VSS 0.00755
R6760 VSS.n2028 VSS 0.00755
R6761 VSS.n1345 VSS 0.00755
R6762 VSS.n1286 VSS 0.00755
R6763 VSS.n859 VSS 0.00755
R6764 VSS.n2986 VSS.n2985 0.0070355
R6765 VSS.n1960 VSS 0.00701042
R6766 VSS.n1731 VSS.n1729 0.00653911
R6767 VSS.n2942 VSS.n234 0.00640857
R6768 VSS.n2954 VSS.n2953 0.00636298
R6769 VSS.n2943 VSS.n2942 0.00636298
R6770 VSS.n1804 VSS.n502 0.00631183
R6771 VSS.n1748 VSS.n1730 0.00624332
R6772 VSS.n1796 VSS.n1731 0.00624332
R6773 VSS.n1728 VSS.n504 0.00604629
R6774 VSS.n2908 VSS.n502 0.00604629
R6775 VSS.n1809 VSS.n1808 0.00579577
R6776 VSS VSS.n1692 0.00570833
R6777 VSS VSS.n1614 0.00570833
R6778 VSS.n1277 VSS 0.00570833
R6779 VSS.n1950 VSS 0.00570833
R6780 VSS.n2953 VSS.n234 0.00533429
R6781 VSS.n1553 VSS.n526 0.0052
R6782 VSS.n1798 VSS.n1797 0.0052
R6783 VSS.n1799 VSS.n267 0.0052
R6784 VSS.n1703 VSS.n1555 0.00514198
R6785 VSS.n1394 VSS.n1393 0.00513595
R6786 VSS.n1092 VSS.n1091 0.00513595
R6787 VSS.n2294 VSS.n2293 0.00513595
R6788 VSS.n2294 VSS.n860 0.00513595
R6789 VSS.n870 VSS.n858 0.00513595
R6790 VSS.n1393 VSS.n1384 0.00513595
R6791 VSS.n1403 VSS.n1402 0.00513595
R6792 VSS.n1091 VSS.n1088 0.00513595
R6793 VSS.n1103 VSS.n1102 0.00513595
R6794 VSS.n1748 VSS.n1729 0.00496369
R6795 VSS.n1804 VSS.n1728 0.0047957
R6796 VSS.n52 VSS.n51 0.00440625
R6797 VSS.n3081 VSS.n3080 0.00440625
R6798 VSS.n3246 VSS.n3239 0.00440625
R6799 VSS.n1135 VSS 0.00440625
R6800 VSS.n2735 VSS 0.00440625
R6801 VSS.n2659 VSS 0.00440625
R6802 VSS.n2167 VSS 0.00440625
R6803 VSS.n1809 VSS.n1806 0.00364583
R6804 VSS.n1807 VSS.n1549 0.00364583
R6805 VSS.n1808 VSS.n1807 0.00364583
R6806 VSS.n1806 VSS.n1805 0.00364583
R6807 VSS VSS.n756 0.00310417
R6808 VSS.n37 VSS.n36 0.00180208
R6809 VSS.n3388 VSS.n35 0.00180208
R6810 VSS.n3052 VSS.n3043 0.00180208
R6811 VSS.n3112 VSS.n194 0.00180208
R6812 VSS.n3297 VSS.n106 0.00180208
R6813 VSS.n3294 VSS.n3293 0.00180208
R6814 VSS.n1886 VSS.n1885 0.00152459
R6815 VDPWR.n710 VDPWR.n706 8629.41
R6816 VDPWR.n710 VDPWR.n707 8629.41
R6817 VDPWR.n712 VDPWR.n706 8629.41
R6818 VDPWR.n712 VDPWR.n707 8629.41
R6819 VDPWR.n695 VDPWR.n691 8629.41
R6820 VDPWR.n695 VDPWR.n692 8629.41
R6821 VDPWR.n697 VDPWR.n691 8629.41
R6822 VDPWR.n697 VDPWR.n692 8629.41
R6823 VDPWR.n679 VDPWR.n675 8629.41
R6824 VDPWR.n679 VDPWR.n676 8629.41
R6825 VDPWR.n681 VDPWR.n675 8629.41
R6826 VDPWR.n681 VDPWR.n676 8629.41
R6827 VDPWR.n665 VDPWR.n659 8629.41
R6828 VDPWR.n663 VDPWR.n659 8629.41
R6829 VDPWR.n665 VDPWR.n661 8629.41
R6830 VDPWR.n663 VDPWR.n661 8629.41
R6831 VDPWR.n521 VDPWR.n517 8629.41
R6832 VDPWR.n521 VDPWR.n518 8629.41
R6833 VDPWR.n523 VDPWR.n517 8629.41
R6834 VDPWR.n523 VDPWR.n518 8629.41
R6835 VDPWR.n506 VDPWR.n502 8629.41
R6836 VDPWR.n506 VDPWR.n503 8629.41
R6837 VDPWR.n508 VDPWR.n502 8629.41
R6838 VDPWR.n508 VDPWR.n503 8629.41
R6839 VDPWR.n490 VDPWR.n486 8629.41
R6840 VDPWR.n490 VDPWR.n487 8629.41
R6841 VDPWR.n492 VDPWR.n486 8629.41
R6842 VDPWR.n492 VDPWR.n487 8629.41
R6843 VDPWR.n473 VDPWR.n469 8629.41
R6844 VDPWR.n473 VDPWR.n470 8629.41
R6845 VDPWR.n475 VDPWR.n469 8629.41
R6846 VDPWR.n475 VDPWR.n470 8629.41
R6847 VDPWR.n411 VDPWR.n405 8629.41
R6848 VDPWR.n411 VDPWR.n406 8629.41
R6849 VDPWR.n409 VDPWR.n406 8629.41
R6850 VDPWR.n409 VDPWR.n405 8629.41
R6851 VDPWR.n384 VDPWR.n378 8629.41
R6852 VDPWR.n381 VDPWR.n380 8629.41
R6853 VDPWR.n396 VDPWR.n390 8629.41
R6854 VDPWR.n393 VDPWR.n392 8629.41
R6855 VDPWR.n452 VDPWR.n448 8629.41
R6856 VDPWR.n452 VDPWR.n449 8629.41
R6857 VDPWR.n454 VDPWR.n448 8629.41
R6858 VDPWR.n454 VDPWR.n449 8629.41
R6859 VDPWR.n436 VDPWR.n432 8629.41
R6860 VDPWR.n436 VDPWR.n433 8629.41
R6861 VDPWR.n438 VDPWR.n432 8629.41
R6862 VDPWR.n438 VDPWR.n433 8629.41
R6863 VDPWR.n422 VDPWR.n416 8629.41
R6864 VDPWR.n420 VDPWR.n416 8629.41
R6865 VDPWR.n422 VDPWR.n418 8629.41
R6866 VDPWR.n420 VDPWR.n418 8629.41
R6867 VDPWR.n765 VDPWR.n761 8629.41
R6868 VDPWR.n765 VDPWR.n762 8629.41
R6869 VDPWR.n767 VDPWR.n761 8629.41
R6870 VDPWR.n767 VDPWR.n762 8629.41
R6871 VDPWR.n3098 VDPWR.n3092 8629.41
R6872 VDPWR.n3098 VDPWR.n3093 8629.41
R6873 VDPWR.n3096 VDPWR.n3093 8629.41
R6874 VDPWR.n3096 VDPWR.n3092 8629.41
R6875 VDPWR.n3082 VDPWR.n3076 8629.41
R6876 VDPWR.n3082 VDPWR.n3077 8629.41
R6877 VDPWR.n3080 VDPWR.n3077 8629.41
R6878 VDPWR.n3080 VDPWR.n3076 8629.41
R6879 VDPWR.n3063 VDPWR.n3059 8629.41
R6880 VDPWR.n3063 VDPWR.n3060 8629.41
R6881 VDPWR.n3065 VDPWR.n3059 8629.41
R6882 VDPWR.n3065 VDPWR.n3060 8629.41
R6883 VDPWR.n733 VDPWR.n730 5460
R6884 VDPWR.n735 VDPWR.n730 5460
R6885 VDPWR.n733 VDPWR.n731 5460
R6886 VDPWR.n735 VDPWR.n731 5460
R6887 VDPWR.n747 VDPWR.n741 4260
R6888 VDPWR.n745 VDPWR.n744 4260
R6889 VDPWR.t536 VDPWR.n710 2459.29
R6890 VDPWR.n712 VDPWR.t535 2459.29
R6891 VDPWR.t111 VDPWR.n695 2459.29
R6892 VDPWR.n697 VDPWR.t94 2459.29
R6893 VDPWR.t75 VDPWR.n679 2459.29
R6894 VDPWR.n681 VDPWR.t76 2459.29
R6895 VDPWR.t5 VDPWR.n659 2459.29
R6896 VDPWR.t4 VDPWR.n661 2459.29
R6897 VDPWR.t660 VDPWR.n521 2459.29
R6898 VDPWR.n523 VDPWR.t659 2459.29
R6899 VDPWR.t246 VDPWR.n506 2459.29
R6900 VDPWR.n508 VDPWR.t49 2459.29
R6901 VDPWR.t713 VDPWR.n490 2459.29
R6902 VDPWR.n492 VDPWR.t712 2459.29
R6903 VDPWR.t464 VDPWR.n473 2459.29
R6904 VDPWR.n475 VDPWR.t465 2459.29
R6905 VDPWR.t662 VDPWR.n409 2459.29
R6906 VDPWR.n411 VDPWR.t661 2459.29
R6907 VDPWR.t247 VDPWR.n452 2459.29
R6908 VDPWR.n454 VDPWR.t248 2459.29
R6909 VDPWR.t711 VDPWR.n436 2459.29
R6910 VDPWR.n438 VDPWR.t714 2459.29
R6911 VDPWR.t466 VDPWR.n416 2459.29
R6912 VDPWR.t467 VDPWR.n418 2459.29
R6913 VDPWR.t602 VDPWR.n765 2459.29
R6914 VDPWR.n767 VDPWR.t176 2459.29
R6915 VDPWR.t470 VDPWR.n3096 2459.29
R6916 VDPWR.n3098 VDPWR.t64 2459.29
R6917 VDPWR.t556 VDPWR.n3080 2459.29
R6918 VDPWR.n3082 VDPWR.t557 2459.29
R6919 VDPWR.t363 VDPWR.n3063 2459.29
R6920 VDPWR.n3065 VDPWR.t463 2459.29
R6921 VDPWR.n711 VDPWR.t536 2298.92
R6922 VDPWR.t535 VDPWR.n711 2298.92
R6923 VDPWR.n696 VDPWR.t111 2298.92
R6924 VDPWR.t94 VDPWR.n696 2298.92
R6925 VDPWR.n680 VDPWR.t75 2298.92
R6926 VDPWR.t76 VDPWR.n680 2298.92
R6927 VDPWR.n664 VDPWR.t5 2298.92
R6928 VDPWR.n664 VDPWR.t4 2298.92
R6929 VDPWR.n522 VDPWR.t660 2298.92
R6930 VDPWR.t659 VDPWR.n522 2298.92
R6931 VDPWR.n507 VDPWR.t246 2298.92
R6932 VDPWR.t49 VDPWR.n507 2298.92
R6933 VDPWR.n491 VDPWR.t713 2298.92
R6934 VDPWR.t712 VDPWR.n491 2298.92
R6935 VDPWR.n474 VDPWR.t464 2298.92
R6936 VDPWR.t465 VDPWR.n474 2298.92
R6937 VDPWR.n410 VDPWR.t662 2298.92
R6938 VDPWR.t661 VDPWR.n410 2298.92
R6939 VDPWR.n453 VDPWR.t247 2298.92
R6940 VDPWR.t248 VDPWR.n453 2298.92
R6941 VDPWR.n437 VDPWR.t711 2298.92
R6942 VDPWR.t714 VDPWR.n437 2298.92
R6943 VDPWR.n421 VDPWR.t466 2298.92
R6944 VDPWR.n421 VDPWR.t467 2298.92
R6945 VDPWR.n766 VDPWR.t602 2298.92
R6946 VDPWR.t176 VDPWR.n766 2298.92
R6947 VDPWR.n3097 VDPWR.t470 2298.92
R6948 VDPWR.t64 VDPWR.n3097 2298.92
R6949 VDPWR.n3081 VDPWR.t556 2298.92
R6950 VDPWR.t557 VDPWR.n3081 2298.92
R6951 VDPWR.n3064 VDPWR.t363 2298.92
R6952 VDPWR.t463 VDPWR.n3064 2298.92
R6953 VDPWR.n1525 VDPWR.n1507 2296.22
R6954 VDPWR.n1300 VDPWR.n1282 2296.22
R6955 VDPWR.n1923 VDPWR.n1922 2296.22
R6956 VDPWR.n2695 VDPWR.n2694 2291.62
R6957 VDPWR.n2694 VDPWR.n2684 1418.92
R6958 VDPWR.n1525 VDPWR.n1524 1408
R6959 VDPWR.n1300 VDPWR.n1299 1408
R6960 VDPWR.n1922 VDPWR.n1921 1408
R6961 VDPWR VDPWR.t970 975.178
R6962 VDPWR VDPWR.t870 975.178
R6963 VDPWR VDPWR.t864 975.178
R6964 VDPWR.n709 VDPWR.n708 920.471
R6965 VDPWR.n694 VDPWR.n693 920.471
R6966 VDPWR.n678 VDPWR.n677 920.471
R6967 VDPWR.n662 VDPWR.n658 920.471
R6968 VDPWR.n520 VDPWR.n519 920.471
R6969 VDPWR.n505 VDPWR.n504 920.471
R6970 VDPWR.n489 VDPWR.n488 920.471
R6971 VDPWR.n472 VDPWR.n471 920.471
R6972 VDPWR.n408 VDPWR.n407 920.471
R6973 VDPWR.n385 VDPWR.n379 920.471
R6974 VDPWR.n397 VDPWR.n391 920.471
R6975 VDPWR.n451 VDPWR.n450 920.471
R6976 VDPWR.n435 VDPWR.n434 920.471
R6977 VDPWR.n419 VDPWR.n415 920.471
R6978 VDPWR.n764 VDPWR.n763 920.471
R6979 VDPWR.n3095 VDPWR.n3094 920.471
R6980 VDPWR.n3079 VDPWR.n3078 920.471
R6981 VDPWR.n3062 VDPWR.n3061 920.471
R6982 VDPWR.n386 VDPWR.n385 917.46
R6983 VDPWR.n398 VDPWR.n397 917.46
R6984 VDPWR.n708 VDPWR.n704 914.447
R6985 VDPWR.n693 VDPWR.n688 914.447
R6986 VDPWR.n677 VDPWR.n672 914.447
R6987 VDPWR.n662 VDPWR.n657 914.447
R6988 VDPWR.n519 VDPWR.n515 914.447
R6989 VDPWR.n504 VDPWR.n499 914.447
R6990 VDPWR.n488 VDPWR.n483 914.447
R6991 VDPWR.n471 VDPWR.n467 914.447
R6992 VDPWR.n407 VDPWR.n403 914.447
R6993 VDPWR.n450 VDPWR.n445 914.447
R6994 VDPWR.n434 VDPWR.n429 914.447
R6995 VDPWR.n419 VDPWR.n414 914.447
R6996 VDPWR.n763 VDPWR.n759 914.447
R6997 VDPWR.n3094 VDPWR.n3089 914.447
R6998 VDPWR.n3078 VDPWR.n3073 914.447
R6999 VDPWR.n3061 VDPWR.n3057 914.447
R7000 VDPWR.t970 VDPWR 877.827
R7001 VDPWR.t870 VDPWR 877.827
R7002 VDPWR.t864 VDPWR 877.827
R7003 VDPWR.n2622 VDPWR.t826 843.261
R7004 VDPWR.n1409 VDPWR.t206 842.073
R7005 VDPWR.n2925 VDPWR.t722 842.073
R7006 VDPWR.n2018 VDPWR.t14 832.876
R7007 VDPWR.n1788 VDPWR.t981 812.014
R7008 VDPWR.n2222 VDPWR.t898 811.918
R7009 VDPWR.n2287 VDPWR.t1111 811.793
R7010 VDPWR.n1098 VDPWR.t570 808.141
R7011 VDPWR.n1354 VDPWR.t1017 807.567
R7012 VDPWR.n2701 VDPWR.t917 807.548
R7013 VDPWR.n1811 VDPWR.t1056 807.481
R7014 VDPWR.n1835 VDPWR.t1158 807.481
R7015 VDPWR.n1841 VDPWR.t957 807.462
R7016 VDPWR.n1383 VDPWR.t859 806.484
R7017 VDPWR.n1485 VDPWR.t1080 806.423
R7018 VDPWR.n1964 VDPWR.t952 806.423
R7019 VDPWR.n803 VDPWR.t280 804.845
R7020 VDPWR.n1710 VDPWR.t1014 804.731
R7021 VDPWR.n1446 VDPWR.t1013 804.731
R7022 VDPWR.n1710 VDPWR.t866 804.731
R7023 VDPWR.n1446 VDPWR.t865 804.731
R7024 VDPWR.n1447 VDPWR.t1060 804.731
R7025 VDPWR.n1458 VDPWR.t1059 804.731
R7026 VDPWR.n1646 VDPWR.t1028 804.731
R7027 VDPWR.n1470 VDPWR.t1027 804.731
R7028 VDPWR.n1646 VDPWR.t872 804.731
R7029 VDPWR.n1470 VDPWR.t871 804.731
R7030 VDPWR.n1471 VDPWR.t1115 804.731
R7031 VDPWR.n1594 VDPWR.t1114 804.731
R7032 VDPWR.n1471 VDPWR.t972 804.731
R7033 VDPWR.n1594 VDPWR.t971 804.731
R7034 VDPWR.n1484 VDPWR.t893 804.731
R7035 VDPWR.n1486 VDPWR.t1026 804.731
R7036 VDPWR.n1563 VDPWR.t1079 804.731
R7037 VDPWR.n1555 VDPWR.t1025 804.731
R7038 VDPWR.n1497 VDPWR.t929 804.731
R7039 VDPWR.n1508 VDPWR.t928 804.731
R7040 VDPWR.n1511 VDPWR.t863 804.731
R7041 VDPWR.n1514 VDPWR.t1052 804.731
R7042 VDPWR.n1518 VDPWR.t836 804.731
R7043 VDPWR.n1523 VDPWR.t1039 804.731
R7044 VDPWR.n1440 VDPWR.t857 804.731
R7045 VDPWR.n1723 VDPWR.t1054 804.731
R7046 VDPWR.n1396 VDPWR.t860 804.731
R7047 VDPWR.t1150 VDPWR.n1378 804.731
R7048 VDPWR.n1355 VDPWR.t980 804.731
R7049 VDPWR.n1376 VDPWR.t1057 804.731
R7050 VDPWR.n1333 VDPWR.t1016 804.731
R7051 VDPWR.n1816 VDPWR.t1159 804.731
R7052 VDPWR.n1840 VDPWR.t1130 804.731
R7053 VDPWR.n1329 VDPWR.t875 804.731
R7054 VDPWR.n1861 VDPWR.t956 804.731
R7055 VDPWR.n1309 VDPWR.t874 804.731
R7056 VDPWR.n1866 VDPWR.t987 804.731
R7057 VDPWR.n1283 VDPWR.t986 804.731
R7058 VDPWR.n1286 VDPWR.t1096 804.731
R7059 VDPWR.n1289 VDPWR.t943 804.731
R7060 VDPWR.n1293 VDPWR.t926 804.731
R7061 VDPWR.n1298 VDPWR.t1108 804.731
R7062 VDPWR.n1416 VDPWR.t1153 804.731
R7063 VDPWR.n1421 VDPWR.t1020 804.731
R7064 VDPWR.n1424 VDPWR.t1148 804.731
R7065 VDPWR.n1429 VDPWR.t1009 804.731
R7066 VDPWR.n1902 VDPWR.t983 804.731
R7067 VDPWR.n1946 VDPWR.t965 804.731
R7068 VDPWR.n1268 VDPWR.t984 804.731
R7069 VDPWR.n2175 VDPWR.t966 804.731
R7070 VDPWR.n1954 VDPWR.t951 804.731
R7071 VDPWR.t853 VDPWR.n2164 804.731
R7072 VDPWR.n2163 VDPWR.t1155 804.731
R7073 VDPWR.n1971 VDPWR.t1070 804.731
R7074 VDPWR.n2143 VDPWR.t1156 804.731
R7075 VDPWR.n1992 VDPWR.t1071 804.731
R7076 VDPWR.n1990 VDPWR.t1049 804.731
R7077 VDPWR.n1993 VDPWR.t1064 804.731
R7078 VDPWR.n2011 VDPWR.t1050 804.731
R7079 VDPWR.n2110 VDPWR.t1065 804.731
R7080 VDPWR.n1906 VDPWR.t1023 804.731
R7081 VDPWR.n1912 VDPWR.t1100 804.731
R7082 VDPWR.n1915 VDPWR.t848 804.731
R7083 VDPWR.n1919 VDPWR.t940 804.731
R7084 VDPWR.t1011 VDPWR.n2039 804.731
R7085 VDPWR.n2054 VDPWR.t920 804.731
R7086 VDPWR.n2057 VDPWR.t998 804.731
R7087 VDPWR.n2213 VDPWR.t932 804.731
R7088 VDPWR.n2216 VDPWR.t1041 804.731
R7089 VDPWR.n2432 VDPWR.t996 804.731
R7090 VDPWR.n1184 VDPWR.t995 804.731
R7091 VDPWR.n1187 VDPWR.t1037 804.731
R7092 VDPWR.n1203 VDPWR.t1036 804.731
R7093 VDPWR.n1204 VDPWR.t1143 804.731
R7094 VDPWR.n2336 VDPWR.t1142 804.731
R7095 VDPWR.n1223 VDPWR.t839 804.731
R7096 VDPWR.n2300 VDPWR.t838 804.731
R7097 VDPWR.n1249 VDPWR.t968 804.731
R7098 VDPWR.n2281 VDPWR.t1047 804.731
R7099 VDPWR.n2256 VDPWR.t1110 804.731
R7100 VDPWR.n2251 VDPWR.t1046 804.731
R7101 VDPWR.n2195 VDPWR.t899 804.731
R7102 VDPWR.n2209 VDPWR.t1084 804.731
R7103 VDPWR.n1176 VDPWR.t990 804.731
R7104 VDPWR.n2445 VDPWR.t1098 804.731
R7105 VDPWR.n964 VDPWR.t1031 804.731
R7106 VDPWR.n967 VDPWR.t1128 804.731
R7107 VDPWR.n2461 VDPWR.t1094 804.731
R7108 VDPWR.n2499 VDPWR.t1093 804.731
R7109 VDPWR.n1151 VDPWR.t1121 804.731
R7110 VDPWR.n1136 VDPWR.t1120 804.731
R7111 VDPWR.t993 VDPWR.n960 804.731
R7112 VDPWR.t977 VDPWR.n961 804.731
R7113 VDPWR.n976 VDPWR.t992 804.731
R7114 VDPWR.n2465 VDPWR.t1082 804.731
R7115 VDPWR.n2468 VDPWR.t851 804.731
R7116 VDPWR.n2597 VDPWR.t1113 804.731
R7117 VDPWR.n2600 VDPWR.t896 804.731
R7118 VDPWR.n2590 VDPWR.t1126 804.731
R7119 VDPWR.n2593 VDPWR.t905 804.731
R7120 VDPWR.n927 VDPWR.t902 804.731
R7121 VDPWR.n2923 VDPWR.t1137 804.731
R7122 VDPWR.n2961 VDPWR.t833 804.731
R7123 VDPWR.n2969 VDPWR.t954 804.731
R7124 VDPWR.n815 VDPWR.t914 804.731
R7125 VDPWR.n2633 VDPWR.t881 804.731
R7126 VDPWR.n2636 VDPWR.t1000 804.731
R7127 VDPWR.n2716 VDPWR.t1139 804.731
R7128 VDPWR.n2692 VDPWR.t916 804.731
R7129 VDPWR.n828 VDPWR.t938 804.731
R7130 VDPWR.n832 VDPWR.t1062 804.731
R7131 VDPWR.n2564 VDPWR.t397 783.403
R7132 VDPWR.n2343 VDPWR.t812 779.372
R7133 VDPWR.n2423 VDPWR.t314 779.372
R7134 VDPWR.t1069 VDPWR.t1154 772.086
R7135 VDPWR.t1063 VDPWR.t1048 772.086
R7136 VDPWR.n1379 VDPWR.t1150 751.692
R7137 VDPWR.t1130 VDPWR.n1839 751.692
R7138 VDPWR.t1153 VDPWR.n1415 751.692
R7139 VDPWR.t1020 VDPWR.n1420 751.692
R7140 VDPWR.n2165 VDPWR.t853 751.692
R7141 VDPWR.n2040 VDPWR.t1011 751.692
R7142 VDPWR.t968 VDPWR.n1248 751.692
R7143 VDPWR.n973 VDPWR.t993 751.692
R7144 VDPWR.n983 VDPWR.t977 751.692
R7145 VDPWR.t992 VDPWR.n975 751.692
R7146 VDPWR.t1126 VDPWR.n2589 751.692
R7147 VDPWR.t905 VDPWR.n2592 751.692
R7148 VDPWR.t1139 VDPWR.n2715 751.692
R7149 VDPWR.t893 VDPWR.n1483 725.173
R7150 VDPWR.t863 VDPWR.n1510 725.173
R7151 VDPWR.t1052 VDPWR.n1513 725.173
R7152 VDPWR.t836 VDPWR.n1517 725.173
R7153 VDPWR.t1039 VDPWR.n1522 725.173
R7154 VDPWR.t857 VDPWR.n1439 725.173
R7155 VDPWR.t1054 VDPWR.n1722 725.173
R7156 VDPWR.t1096 VDPWR.n1285 725.173
R7157 VDPWR.t943 VDPWR.n1288 725.173
R7158 VDPWR.t926 VDPWR.n1292 725.173
R7159 VDPWR.t1108 VDPWR.n1297 725.173
R7160 VDPWR.t1148 VDPWR.n1423 725.173
R7161 VDPWR.t1009 VDPWR.n1428 725.173
R7162 VDPWR.t1023 VDPWR.n1905 725.173
R7163 VDPWR.t1100 VDPWR.n1911 725.173
R7164 VDPWR.t848 VDPWR.n1914 725.173
R7165 VDPWR.t940 VDPWR.n1918 725.173
R7166 VDPWR.t920 VDPWR.n2053 725.173
R7167 VDPWR.t998 VDPWR.n2056 725.173
R7168 VDPWR.t932 VDPWR.n2212 725.173
R7169 VDPWR.t1041 VDPWR.n2215 725.173
R7170 VDPWR.t1084 VDPWR.n2208 725.173
R7171 VDPWR.t990 VDPWR.n1175 725.173
R7172 VDPWR.t1098 VDPWR.n2444 725.173
R7173 VDPWR.t1031 VDPWR.n963 725.173
R7174 VDPWR.t1128 VDPWR.n966 725.173
R7175 VDPWR.t1082 VDPWR.n2464 725.173
R7176 VDPWR.t851 VDPWR.n2467 725.173
R7177 VDPWR.t1113 VDPWR.n2596 725.173
R7178 VDPWR.t896 VDPWR.n2599 725.173
R7179 VDPWR.t902 VDPWR.n926 725.173
R7180 VDPWR.t1137 VDPWR.n2922 725.173
R7181 VDPWR.t833 VDPWR.n2960 725.173
R7182 VDPWR.t954 VDPWR.n2968 725.173
R7183 VDPWR.t914 VDPWR.n814 725.173
R7184 VDPWR.t881 VDPWR.n2632 725.173
R7185 VDPWR.t1000 VDPWR.n2635 725.173
R7186 VDPWR.t938 VDPWR.n827 725.173
R7187 VDPWR.t1062 VDPWR.n831 725.173
R7188 VDPWR.n2892 VDPWR.n900 717.729
R7189 VDPWR.n2887 VDPWR.n903 717.729
R7190 VDPWR.n2034 VDPWR.n2031 713.462
R7191 VDPWR.n570 VDPWR.t265 675.542
R7192 VDPWR.n290 VDPWR.t102 675.542
R7193 VDPWR.n33 VDPWR.t16 675.542
R7194 VDPWR.n2905 VDPWR.t156 671.408
R7195 VDPWR.n785 VDPWR.t636 671.408
R7196 VDPWR.n3031 VDPWR.t634 671.408
R7197 VDPWR.n559 VDPWR.t274 671.376
R7198 VDPWR.n279 VDPWR.t38 671.376
R7199 VDPWR.n22 VDPWR.t684 671.376
R7200 VDPWR.n1085 VDPWR.t734 669.655
R7201 VDPWR.n1759 VDPWR.t3 667.734
R7202 VDPWR.n2081 VDPWR.t186 667.734
R7203 VDPWR.n1032 VDPWR.t225 667.734
R7204 VDPWR.n2810 VDPWR.t123 667.734
R7205 VDPWR.n2810 VDPWR.t828 667.734
R7206 VDPWR.n2931 VDPWR.t115 667.734
R7207 VDPWR.n2938 VDPWR.t194 667.734
R7208 VDPWR.n1065 VDPWR.t771 666.677
R7209 VDPWR.n2868 VDPWR.t544 666.677
R7210 VDPWR.n2824 VDPWR.t152 666.677
R7211 VDPWR.n2824 VDPWR.t257 666.677
R7212 VDPWR.n2994 VDPWR.t682 666.677
R7213 VDPWR.n2989 VDPWR.t587 666.677
R7214 VDPWR.t909 VDPWR 666.343
R7215 VDPWR.t1122 VDPWR 666.343
R7216 VDPWR.t1157 VDPWR 666.343
R7217 VDPWR.t1055 VDPWR 666.343
R7218 VDPWR.t882 VDPWR 666.343
R7219 VDPWR.t961 VDPWR 666.343
R7220 VDPWR VDPWR.t1089 664.664
R7221 VDPWR.n2885 VDPWR.t581 664.37
R7222 VDPWR.n2523 VDPWR.t93 664.279
R7223 VDPWR.n2859 VDPWR.t188 664.279
R7224 VDPWR.n2850 VDPWR.t335 664.279
R7225 VDPWR.n1156 VDPWR.t579 663.024
R7226 VDPWR.n1387 VDPWR.t282 662.571
R7227 VDPWR.n2102 VDPWR.t676 662.571
R7228 VDPWR.n1017 VDPWR.t726 659.593
R7229 VDPWR.n2660 VDPWR.t127 659.593
R7230 VDPWR.n2676 VDPWR.t577 659.593
R7231 VDPWR.n1043 VDPWR.n1042 642.188
R7232 VDPWR.n251 VDPWR.t613 633.369
R7233 VDPWR VDPWR.t921 630.375
R7234 VDPWR VDPWR.t840 630.375
R7235 VDPWR VDPWR.t973 630.375
R7236 VDPWR.t1078 VDPWR.t1024 617.668
R7237 VDPWR.t955 VDPWR.t873 617.668
R7238 VDPWR.t950 VDPWR.t964 617.668
R7239 VDPWR.n810 VDPWR.n809 614.562
R7240 VDPWR.n1093 VDPWR.n1092 613.71
R7241 VDPWR.n2083 VDPWR.n2082 611.178
R7242 VDPWR.n2895 VDPWR.n2894 611.178
R7243 VDPWR.n2885 VDPWR.n907 611.178
R7244 VDPWR.n995 VDPWR.n994 610.861
R7245 VDPWR.n2557 VDPWR.n990 609.847
R7246 VDPWR.n2555 VDPWR.n993 609.717
R7247 VDPWR.n2408 VDPWR.n1186 609.303
R7248 VDPWR.n2329 VDPWR.n2328 606.42
R7249 VDPWR.n2326 VDPWR.n1225 606.42
R7250 VDPWR.n2335 VDPWR.n1222 606.42
R7251 VDPWR.n2416 VDPWR.n2415 606.42
R7252 VDPWR.n2413 VDPWR.n1183 606.42
R7253 VDPWR.n2548 VDPWR.n999 606.42
R7254 VDPWR.n1220 VDPWR.n1219 605.581
R7255 VDPWR.n2421 VDPWR.n1180 605.581
R7256 VDPWR.n2311 VDPWR.n2310 605.186
R7257 VDPWR.n2309 VDPWR.n1239 605.186
R7258 VDPWR.n1241 VDPWR.n1240 605.186
R7259 VDPWR.n2392 VDPWR.n2390 605.186
R7260 VDPWR.n1197 VDPWR.n1196 605.186
R7261 VDPWR.n2384 VDPWR.n1199 605.186
R7262 VDPWR.n1001 VDPWR.n1000 605.186
R7263 VDPWR.n1016 VDPWR.n1009 605.186
R7264 VDPWR.n1020 VDPWR.n1019 605.186
R7265 VDPWR.n2105 VDPWR.n2104 604.394
R7266 VDPWR.n1061 VDPWR.n1060 604.394
R7267 VDPWR.n2886 VDPWR.n904 604.394
R7268 VDPWR.n909 VDPWR.n908 604.394
R7269 VDPWR.n2829 VDPWR.n939 604.394
R7270 VDPWR.n2829 VDPWR.n2828 604.394
R7271 VDPWR.n2946 VDPWR.n2945 604.394
R7272 VDPWR.n2893 VDPWR.n898 603.231
R7273 VDPWR.n2788 VDPWR.n2787 603.231
R7274 VDPWR.n2075 VDPWR.n2042 603.052
R7275 VDPWR.n629 VDPWR.n564 602.456
R7276 VDPWR.n650 VDPWR.n539 602.456
R7277 VDPWR.n349 VDPWR.n284 602.456
R7278 VDPWR.n370 VDPWR.n259 602.456
R7279 VDPWR.n992 VDPWR.n991 602.456
R7280 VDPWR.n92 VDPWR.n27 602.456
R7281 VDPWR.n113 VDPWR.n2 602.456
R7282 VDPWR.n1781 VDPWR.n1384 601.097
R7283 VDPWR.n2497 VDPWR.n1157 601.097
R7284 VDPWR.n2984 VDPWR.n2949 601.097
R7285 VDPWR.n1122 VDPWR.n1120 599.159
R7286 VDPWR.n1011 VDPWR.n1010 596.442
R7287 VDPWR.n2776 VDPWR.n2662 596.442
R7288 VDPWR.n2752 VDPWR.n2678 596.442
R7289 VDPWR.n2560 VDPWR.n2559 589.481
R7290 VDPWR.n1105 VDPWR.n1028 588.318
R7291 VDPWR.n545 VDPWR.n544 585
R7292 VDPWR.n543 VDPWR.n542 585
R7293 VDPWR.n265 VDPWR.n264 585
R7294 VDPWR.n263 VDPWR.n262 585
R7295 VDPWR.n1067 VDPWR.n1066 585
R7296 VDPWR.n1107 VDPWR.n1106 585
R7297 VDPWR.n2558 VDPWR.n988 585
R7298 VDPWR.n8 VDPWR.n7 585
R7299 VDPWR.n6 VDPWR.n5 585
R7300 VDPWR.n736 VDPWR.n729 582.4
R7301 VDPWR.n732 VDPWR.n729 582.4
R7302 VDPWR VDPWR.t1015 568.994
R7303 VDPWR VDPWR.t979 568.994
R7304 VDPWR VDPWR.t852 568.994
R7305 VDPWR.t903 VDPWR.t894 540.46
R7306 VDPWR VDPWR.n250 535.705
R7307 VDPWR.n732 VDPWR.n728 531.923
R7308 VDPWR.n737 VDPWR.n736 531.427
R7309 VDPWR.t1045 VDPWR 511.926
R7310 VDPWR VDPWR.t1075 510.248
R7311 VDPWR.t313 VDPWR.t1101 496.82
R7312 VDPWR VDPWR.n2002 491.784
R7313 VDPWR.n408 VDPWR.n404 480.764
R7314 VDPWR.n3095 VDPWR.n3090 480.764
R7315 VDPWR.n3079 VDPWR.n3074 480.764
R7316 VDPWR.n709 VDPWR.n705 480.764
R7317 VDPWR.n694 VDPWR.n689 480.764
R7318 VDPWR.n678 VDPWR.n673 480.764
R7319 VDPWR.n666 VDPWR.n658 480.764
R7320 VDPWR.n520 VDPWR.n516 480.764
R7321 VDPWR.n505 VDPWR.n500 480.764
R7322 VDPWR.n489 VDPWR.n484 480.764
R7323 VDPWR.n472 VDPWR.n468 480.764
R7324 VDPWR.n379 VDPWR.n377 480.764
R7325 VDPWR.n391 VDPWR.n389 480.764
R7326 VDPWR.n451 VDPWR.n446 480.764
R7327 VDPWR.n435 VDPWR.n430 480.764
R7328 VDPWR.n423 VDPWR.n415 480.764
R7329 VDPWR.n764 VDPWR.n760 480.764
R7330 VDPWR.n3062 VDPWR.n3058 480.764
R7331 VDPWR VDPWR.t172 470.562
R7332 VDPWR VDPWR.t783 470.562
R7333 VDPWR VDPWR.t768 470.562
R7334 VDPWR VDPWR.t321 470.562
R7335 VDPWR VDPWR.t327 470.562
R7336 VDPWR VDPWR.t527 470.562
R7337 VDPWR VDPWR.t548 470.562
R7338 VDPWR VDPWR.t554 470.562
R7339 VDPWR.t834 VDPWR.t861 463.252
R7340 VDPWR.t924 VDPWR.t941 463.252
R7341 VDPWR.t1021 VDPWR.t846 463.252
R7342 VDPWR.t1083 VDPWR.t930 463.252
R7343 VDPWR.t1109 VDPWR.t1045 463.252
R7344 VDPWR.t1092 VDPWR.t867 463.252
R7345 VDPWR VDPWR.t1104 458.724
R7346 VDPWR.t921 VDPWR 458.724
R7347 VDPWR VDPWR.t1001 458.724
R7348 VDPWR.t840 VDPWR 458.724
R7349 VDPWR VDPWR.t1116 458.724
R7350 VDPWR.t973 VDPWR 458.724
R7351 VDPWR.t689 VDPWR.t749 458.216
R7352 VDPWR.n748 VDPWR.n740 454.401
R7353 VDPWR.n742 VDPWR.n740 454.401
R7354 VDPWR.n742 VDPWR.n739 448.736
R7355 VDPWR.n749 VDPWR.n748 448.288
R7356 VDPWR.n178 VDPWR 435.082
R7357 VDPWR.n620 VDPWR.t700 420.25
R7358 VDPWR.n340 VDPWR.t751 420.25
R7359 VDPWR.t179 VDPWR.n176 420.25
R7360 VDPWR.n83 VDPWR.t706 420.25
R7361 VDPWR.t1058 VDPWR 414.577
R7362 VDPWR VDPWR.t897 414.577
R7363 VDPWR VDPWR.t1109 414.577
R7364 VDPWR.t867 VDPWR 414.577
R7365 VDPWR.t1075 VDPWR 414.577
R7366 VDPWR.n854 VDPWR.t878 390.875
R7367 VDPWR.n1837 VDPWR.t1131 389.526
R7368 VDPWR.n2713 VDPWR.t1140 389.361
R7369 VDPWR.n1381 VDPWR.t1151 388.721
R7370 VDPWR.n319 VDPWR.t842 388.656
R7371 VDPWR.n1508 VDPWR.t910 388.656
R7372 VDPWR.n1549 VDPWR.t911 388.656
R7373 VDPWR.n1663 VDPWR.t1090 388.656
R7374 VDPWR.n1673 VDPWR.t1091 388.656
R7375 VDPWR.n1283 VDPWR.t1123 388.656
R7376 VDPWR.n1308 VDPWR.t1124 388.656
R7377 VDPWR.n1970 VDPWR.t854 388.656
R7378 VDPWR.n1902 VDPWR.t883 388.656
R7379 VDPWR.n1940 VDPWR.t884 388.656
R7380 VDPWR.n2205 VDPWR.t962 388.656
R7381 VDPWR.n2197 VDPWR.t963 388.656
R7382 VDPWR.n2294 VDPWR.t969 388.656
R7383 VDPWR.n2900 VDPWR.t889 388.656
R7384 VDPWR.n2904 VDPWR.t890 388.656
R7385 VDPWR.n824 VDPWR.t949 388.656
R7386 VDPWR.n595 VDPWR.t922 388.656
R7387 VDPWR.n599 VDPWR.t923 388.656
R7388 VDPWR.n587 VDPWR.t1105 388.656
R7389 VDPWR.n623 VDPWR.t1106 388.656
R7390 VDPWR.n573 VDPWR.t1073 388.656
R7391 VDPWR.n582 VDPWR.t1074 388.656
R7392 VDPWR.n547 VDPWR.t1087 388.656
R7393 VDPWR.n552 VDPWR.t1088 388.656
R7394 VDPWR.n315 VDPWR.t841 388.656
R7395 VDPWR.n307 VDPWR.t1002 388.656
R7396 VDPWR.n343 VDPWR.t1003 388.656
R7397 VDPWR.n293 VDPWR.t1005 388.656
R7398 VDPWR.n302 VDPWR.t1006 388.656
R7399 VDPWR.n267 VDPWR.t945 388.656
R7400 VDPWR.n272 VDPWR.t946 388.656
R7401 VDPWR.n2013 VDPWR.t1145 388.656
R7402 VDPWR.n2110 VDPWR.t1146 388.656
R7403 VDPWR.n2043 VDPWR.t1012 388.656
R7404 VDPWR.n2349 VDPWR.t1133 388.656
R7405 VDPWR.n1206 VDPWR.t1134 388.656
R7406 VDPWR.n2429 VDPWR.t1102 388.656
R7407 VDPWR.n2432 VDPWR.t1103 388.656
R7408 VDPWR.n1117 VDPWR.t907 388.656
R7409 VDPWR.n1121 VDPWR.t908 388.656
R7410 VDPWR.n986 VDPWR.t978 388.656
R7411 VDPWR.n1162 VDPWR.t868 388.656
R7412 VDPWR.n2461 VDPWR.t869 388.656
R7413 VDPWR.n2947 VDPWR.t959 388.656
R7414 VDPWR.n2957 VDPWR.t960 388.656
R7415 VDPWR.n2659 VDPWR.t1043 388.656
R7416 VDPWR.n2775 VDPWR.t1044 388.656
R7417 VDPWR.n2653 VDPWR.t844 388.656
R7418 VDPWR.n2795 VDPWR.t845 388.656
R7419 VDPWR.n2758 VDPWR.t886 388.656
R7420 VDPWR.n2679 VDPWR.t887 388.656
R7421 VDPWR.n2692 VDPWR.t1076 388.656
R7422 VDPWR.n2727 VDPWR.t1077 388.656
R7423 VDPWR.n788 VDPWR.t1033 388.656
R7424 VDPWR.n794 VDPWR.t1034 388.656
R7425 VDPWR.n861 VDPWR.t877 388.656
R7426 VDPWR.n58 VDPWR.t974 388.656
R7427 VDPWR.n62 VDPWR.t975 388.656
R7428 VDPWR.n50 VDPWR.t1117 388.656
R7429 VDPWR.n86 VDPWR.t1118 388.656
R7430 VDPWR.n36 VDPWR.t934 388.656
R7431 VDPWR.n45 VDPWR.t935 388.656
R7432 VDPWR.n10 VDPWR.t1067 388.656
R7433 VDPWR.n15 VDPWR.t1068 388.656
R7434 VDPWR.n1414 VDPWR.t1152 387.682
R7435 VDPWR.n1419 VDPWR.t1019 387.682
R7436 VDPWR.n2588 VDPWR.t1125 387.682
R7437 VDPWR.n2591 VDPWR.t904 387.682
R7438 VDPWR.n2003 VDPWR.t1144 386.043
R7439 VDPWR.n816 VDPWR.t948 385.026
R7440 VDPWR.n2206 VDPWR.t1085 383.42
R7441 VDPWR VDPWR.t130 381.007
R7442 VDPWR.n1482 VDPWR.t892 380.193
R7443 VDPWR.n1509 VDPWR.t862 380.193
R7444 VDPWR.n1512 VDPWR.t1051 380.193
R7445 VDPWR.n1516 VDPWR.t835 380.193
R7446 VDPWR.n1521 VDPWR.t1038 380.193
R7447 VDPWR.n1438 VDPWR.t856 380.193
R7448 VDPWR.n1721 VDPWR.t1053 380.193
R7449 VDPWR.n1284 VDPWR.t1095 380.193
R7450 VDPWR.n1287 VDPWR.t942 380.193
R7451 VDPWR.n1291 VDPWR.t925 380.193
R7452 VDPWR.n1296 VDPWR.t1107 380.193
R7453 VDPWR.n1422 VDPWR.t1147 380.193
R7454 VDPWR.n1427 VDPWR.t1008 380.193
R7455 VDPWR.n1904 VDPWR.t1022 380.193
R7456 VDPWR.n1910 VDPWR.t1099 380.193
R7457 VDPWR.n1913 VDPWR.t847 380.193
R7458 VDPWR.n1917 VDPWR.t939 380.193
R7459 VDPWR.n2052 VDPWR.t919 380.193
R7460 VDPWR.n2055 VDPWR.t997 380.193
R7461 VDPWR.n2211 VDPWR.t931 380.193
R7462 VDPWR.n2214 VDPWR.t1040 380.193
R7463 VDPWR.n1174 VDPWR.t989 380.193
R7464 VDPWR.n2443 VDPWR.t1097 380.193
R7465 VDPWR.n962 VDPWR.t1030 380.193
R7466 VDPWR.n965 VDPWR.t1127 380.193
R7467 VDPWR.n2463 VDPWR.t1081 380.193
R7468 VDPWR.n2466 VDPWR.t850 380.193
R7469 VDPWR.n2595 VDPWR.t1112 380.193
R7470 VDPWR.n2598 VDPWR.t895 380.193
R7471 VDPWR.n925 VDPWR.t901 380.193
R7472 VDPWR.n2921 VDPWR.t1136 380.193
R7473 VDPWR.n2959 VDPWR.t832 380.193
R7474 VDPWR.n2967 VDPWR.t953 380.193
R7475 VDPWR.n813 VDPWR.t913 380.193
R7476 VDPWR.n2631 VDPWR.t880 380.193
R7477 VDPWR.n2634 VDPWR.t999 380.193
R7478 VDPWR.n826 VDPWR.t937 380.193
R7479 VDPWR.n830 VDPWR.t1061 380.193
R7480 VDPWR.n715 VDPWR.n705 379.2
R7481 VDPWR.n699 VDPWR.n689 379.2
R7482 VDPWR.n683 VDPWR.n673 379.2
R7483 VDPWR.n667 VDPWR.n666 379.2
R7484 VDPWR.n526 VDPWR.n516 379.2
R7485 VDPWR.n510 VDPWR.n500 379.2
R7486 VDPWR.n494 VDPWR.n484 379.2
R7487 VDPWR.n478 VDPWR.n468 379.2
R7488 VDPWR.n462 VDPWR.n404 379.2
R7489 VDPWR.n387 VDPWR.n377 379.2
R7490 VDPWR.n399 VDPWR.n389 379.2
R7491 VDPWR.n456 VDPWR.n446 379.2
R7492 VDPWR.n440 VDPWR.n430 379.2
R7493 VDPWR.n424 VDPWR.n423 379.2
R7494 VDPWR.n3106 VDPWR.n760 379.2
R7495 VDPWR.n3100 VDPWR.n3090 379.2
R7496 VDPWR.n3084 VDPWR.n3074 379.2
R7497 VDPWR.n3068 VDPWR.n3058 379.2
R7498 VDPWR VDPWR.t422 369.938
R7499 VDPWR VDPWR.t50 369.938
R7500 VDPWR VDPWR.t350 369.938
R7501 VDPWR VDPWR.t629 369.938
R7502 VDPWR.t584 VDPWR 369.938
R7503 VDPWR.t137 VDPWR 369.938
R7504 VDPWR.t360 VDPWR 369.938
R7505 VDPWR.t356 VDPWR 369.938
R7506 VDPWR.t519 VDPWR 369.938
R7507 VDPWR.t216 VDPWR 369.938
R7508 VDPWR.t214 VDPWR 369.938
R7509 VDPWR.t619 VDPWR 369.938
R7510 VDPWR VDPWR.t262 369.938
R7511 VDPWR VDPWR.t461 369.938
R7512 VDPWR VDPWR.t1018 360.866
R7513 VDPWR.t1024 VDPWR 357.51
R7514 VDPWR.t873 VDPWR 357.51
R7515 VDPWR.t964 VDPWR 357.51
R7516 VDPWR.t991 VDPWR 355.83
R7517 VDPWR.t565 VDPWR.t92 352.474
R7518 VDPWR.t122 VDPWR.t332 352.474
R7519 VDPWR.n141 VDPWR.t650 348.849
R7520 VDPWR.n1059 VDPWR.t742 340.212
R7521 VDPWR VDPWR.t879 337.368
R7522 VDPWR.n2292 VDPWR.t472 336.524
R7523 VDPWR.n2369 VDPWR.t494 336.524
R7524 VDPWR.n929 VDPWR.n928 334.247
R7525 VDPWR VDPWR.t1029 334.012
R7526 VDPWR.n2037 VDPWR.n2036 333.99
R7527 VDPWR.n1756 VDPWR.n1412 333.348
R7528 VDPWR.n1137 VDPWR.n1135 333.348
R7529 VDPWR.n949 VDPWR.n948 333.348
R7530 VDPWR.n880 VDPWR.n879 333.348
R7531 VDPWR.n1099 VDPWR.n1031 333.346
R7532 VDPWR.n2853 VDPWR.n2852 333.346
R7533 VDPWR.n949 VDPWR.n947 333.346
R7534 VDPWR.n2933 VDPWR.n2932 333.346
R7535 VDPWR.n2646 VDPWR.n2625 328.036
R7536 VDPWR.n1561 VDPWR.t1192 328.005
R7537 VDPWR.n1311 VDPWR.t1286 328.005
R7538 VDPWR.n1952 VDPWR.t1208 328.005
R7539 VDPWR.n2712 VDPWR.n2703 326.202
R7540 VDPWR.n2924 VDPWR.n883 325.639
R7541 VDPWR.n1757 VDPWR.n1411 324.74
R7542 VDPWR.n576 VDPWR.n569 322.329
R7543 VDPWR.n554 VDPWR.n550 322.329
R7544 VDPWR.n296 VDPWR.n289 322.329
R7545 VDPWR.n274 VDPWR.n270 322.329
R7546 VDPWR.n2901 VDPWR.n894 322.329
R7547 VDPWR.n792 VDPWR.n791 322.329
R7548 VDPWR.n39 VDPWR.n32 322.329
R7549 VDPWR.n17 VDPWR.n13 322.329
R7550 VDPWR.t319 VDPWR.t195 322.262
R7551 VDPWR.n2378 VDPWR.t1216 321.911
R7552 VDPWR.n140 VDPWR.n139 320.976
R7553 VDPWR.n1403 VDPWR.n1402 320.976
R7554 VDPWR.n1141 VDPWR.n1140 320.976
R7555 VDPWR.n2860 VDPWR.n922 320.976
R7556 VDPWR.n2817 VDPWR.n944 320.976
R7557 VDPWR.n2940 VDPWR.n876 320.976
R7558 VDPWR.n2033 VDPWR.n2032 320.976
R7559 VDPWR.n1086 VDPWR.n1084 320.976
R7560 VDPWR.n2867 VDPWR.n919 320.976
R7561 VDPWR.n2817 VDPWR.n943 320.976
R7562 VDPWR.n2943 VDPWR.n2942 320.976
R7563 VDPWR.t240 VDPWR.t151 315.548
R7564 VDPWR.t431 VDPWR.t825 315.548
R7565 VDPWR.n1047 VDPWR.n1046 315.089
R7566 VDPWR.n1055 VDPWR.n1054 314.447
R7567 VDPWR.t224 VDPWR.t569 313.87
R7568 VDPWR.n2097 VDPWR.n2096 312.829
R7569 VDPWR.n2790 VDPWR.n2789 312.053
R7570 VDPWR.n2646 VDPWR.n2628 312.053
R7571 VDPWR.n2641 VDPWR.n2630 312.053
R7572 VDPWR.n2746 VDPWR.n2683 312.053
R7573 VDPWR.n1055 VDPWR.n1053 312.051
R7574 VDPWR.n2294 VDPWR.n2293 311.151
R7575 VDPWR.n2374 VDPWR.n1202 311.151
R7576 VDPWR.n2301 VDPWR.n1243 310.904
R7577 VDPWR.n2377 VDPWR.n2376 310.904
R7578 VDPWR.n2747 VDPWR.n2680 310.5
R7579 VDPWR.n850 VDPWR.n849 309.533
R7580 VDPWR.t927 VDPWR.t909 308.834
R7581 VDPWR.n1588 VDPWR.t891 308.834
R7582 VDPWR.t985 VDPWR.t1122 308.834
R7583 VDPWR.t1015 VDPWR.t1157 308.834
R7584 VDPWR.t979 VDPWR.t1055 308.834
R7585 VDPWR.t982 VDPWR.t882 308.834
R7586 VDPWR.t1141 VDPWR.t1132 308.834
R7587 VDPWR.t976 VDPWR.t991 308.834
R7588 VDPWR.n820 VDPWR.n819 308.755
R7589 VDPWR.n796 VDPWR.n795 308.755
R7590 VDPWR.n2705 VDPWR.n2704 308.755
R7591 VDPWR.n2700 VDPWR.n2699 308.755
R7592 VDPWR.n2764 VDPWR.n2671 308.755
R7593 VDPWR.n1683 VDPWR.n1453 308.755
R7594 VDPWR.n2568 VDPWR.n985 308.755
R7595 VDPWR.n2549 VDPWR.n998 307.204
R7596 VDPWR.n2673 VDPWR.n2672 307.204
R7597 VDPWR.n1600 VDPWR.t1252 306.735
R7598 VDPWR.n1600 VDPWR.t1281 306.735
R7599 VDPWR.n1468 VDPWR.t1168 306.735
R7600 VDPWR.n1468 VDPWR.t1191 306.735
R7601 VDPWR.n1501 VDPWR.t1272 306.735
R7602 VDPWR.n1569 VDPWR.t1213 306.735
R7603 VDPWR.n1666 VDPWR.t1222 306.735
R7604 VDPWR.n1444 VDPWR.t1170 306.735
R7605 VDPWR.n1444 VDPWR.t1195 306.735
R7606 VDPWR.n1306 VDPWR.t1246 306.735
R7607 VDPWR.n1320 VDPWR.t1260 306.735
R7608 VDPWR.n1335 VDPWR.t1235 306.735
R7609 VDPWR.n1830 VDPWR.t1175 306.735
R7610 VDPWR.n1357 VDPWR.t1177 306.735
R7611 VDPWR.n1806 VDPWR.t1223 306.735
R7612 VDPWR.n1782 VDPWR.t1219 306.735
R7613 VDPWR.n1995 VDPWR.t1174 306.735
R7614 VDPWR.n1991 VDPWR.t1184 306.735
R7615 VDPWR.n1987 VDPWR.t1172 306.735
R7616 VDPWR.n1969 VDPWR.t1271 306.735
R7617 VDPWR.n1960 VDPWR.t1224 306.735
R7618 VDPWR.n1272 VDPWR.t1210 306.735
R7619 VDPWR.n2232 VDPWR.t1238 306.735
R7620 VDPWR.n2194 VDPWR.t1209 306.735
R7621 VDPWR.n2192 VDPWR.t1279 306.735
R7622 VDPWR.n2307 VDPWR.t1283 306.735
R7623 VDPWR.n2342 VDPWR.t1173 306.735
R7624 VDPWR.n1181 VDPWR.t1230 306.735
R7625 VDPWR.n1138 VDPWR.t1178 306.735
R7626 VDPWR.n1161 VDPWR.t1187 306.735
R7627 VDPWR.n2698 VDPWR.t1264 306.735
R7628 VDPWR.t811 VDPWR 290.372
R7629 VDPWR VDPWR.t855 280.3
R7630 VDPWR VDPWR.t1007 280.3
R7631 VDPWR.t183 VDPWR 280.3
R7632 VDPWR VDPWR.t918 280.3
R7633 VDPWR VDPWR.t988 280.3
R7634 VDPWR VDPWR.t849 280.3
R7635 VDPWR VDPWR.t831 280.3
R7636 VDPWR VDPWR.t936 280.3
R7637 VDPWR.t65 VDPWR.t663 278.623
R7638 VDPWR.n147 VDPWR.n146 272.274
R7639 VDPWR.n147 VDPWR.n134 272.274
R7640 VDPWR.n176 VDPWR.n134 272.274
R7641 VDPWR.t210 VDPWR 261.837
R7642 VDPWR VDPWR.t927 260.159
R7643 VDPWR VDPWR.t1078 260.159
R7644 VDPWR VDPWR.t985 260.159
R7645 VDPWR VDPWR.t955 260.159
R7646 VDPWR VDPWR.t1129 260.159
R7647 VDPWR.t1149 VDPWR 260.159
R7648 VDPWR.t1018 VDPWR 260.159
R7649 VDPWR VDPWR.t982 260.159
R7650 VDPWR VDPWR.t950 260.159
R7651 VDPWR.t1144 VDPWR 260.159
R7652 VDPWR.t1132 VDPWR 260.159
R7653 VDPWR.t1101 VDPWR 260.159
R7654 VDPWR VDPWR.t903 260.159
R7655 VDPWR VDPWR.t843 260.159
R7656 VDPWR.t220 VDPWR 260.159
R7657 VDPWR.t258 VDPWR 260.159
R7658 VDPWR.t329 VDPWR 260.159
R7659 VDPWR.n633 VDPWR.n631 259.697
R7660 VDPWR.n353 VDPWR.n351 259.697
R7661 VDPWR.n96 VDPWR.n94 259.697
R7662 VDPWR.n609 VDPWR.t51 255.905
R7663 VDPWR.n614 VDPWR.t423 255.905
R7664 VDPWR.n590 VDPWR.t701 255.905
R7665 VDPWR.n630 VDPWR.t428 255.905
R7666 VDPWR.n538 VDPWR.t534 255.905
R7667 VDPWR.n329 VDPWR.t630 255.905
R7668 VDPWR.n334 VDPWR.t351 255.905
R7669 VDPWR.n310 VDPWR.t752 255.905
R7670 VDPWR.n350 VDPWR.t757 255.905
R7671 VDPWR.n258 VDPWR.t132 255.905
R7672 VDPWR.n183 VDPWR.t620 255.905
R7673 VDPWR.n188 VDPWR.t215 255.905
R7674 VDPWR.n193 VDPWR.t217 255.905
R7675 VDPWR.n198 VDPWR.t520 255.905
R7676 VDPWR.n129 VDPWR.t357 255.905
R7677 VDPWR.n159 VDPWR.t361 255.905
R7678 VDPWR.n164 VDPWR.t138 255.905
R7679 VDPWR.n169 VDPWR.t585 255.905
R7680 VDPWR.n135 VDPWR.t180 255.905
R7681 VDPWR.n72 VDPWR.t462 255.905
R7682 VDPWR.n77 VDPWR.t263 255.905
R7683 VDPWR.n53 VDPWR.t707 255.905
R7684 VDPWR.n93 VDPWR.t778 255.905
R7685 VDPWR.n1 VDPWR.t591 255.905
R7686 VDPWR.n246 VDPWR.t173 255.904
R7687 VDPWR.n123 VDPWR.t784 255.904
R7688 VDPWR.n124 VDPWR.t769 255.904
R7689 VDPWR.n125 VDPWR.t322 255.904
R7690 VDPWR.n126 VDPWR.t328 255.904
R7691 VDPWR.n204 VDPWR.t528 255.904
R7692 VDPWR.n205 VDPWR.t549 255.904
R7693 VDPWR.n206 VDPWR.t555 255.904
R7694 VDPWR.n119 VDPWR.t614 255.904
R7695 VDPWR.n580 VDPWR.t231 254.475
R7696 VDPWR.n300 VDPWR.t773 254.475
R7697 VDPWR.n43 VDPWR.t148 254.475
R7698 VDPWR.n605 VDPWR.t460 252.95
R7699 VDPWR.n610 VDPWR.t421 252.95
R7700 VDPWR.n615 VDPWR.t710 252.95
R7701 VDPWR.n649 VDPWR.t532 252.95
R7702 VDPWR.n644 VDPWR.t656 252.95
R7703 VDPWR.n325 VDPWR.t626 252.95
R7704 VDPWR.n330 VDPWR.t433 252.95
R7705 VDPWR.n335 VDPWR.t754 252.95
R7706 VDPWR.n369 VDPWR.t134 252.95
R7707 VDPWR.n364 VDPWR.t345 252.95
R7708 VDPWR.n179 VDPWR.t618 252.95
R7709 VDPWR.n184 VDPWR.t213 252.95
R7710 VDPWR.n189 VDPWR.t219 252.95
R7711 VDPWR.n194 VDPWR.t518 252.95
R7712 VDPWR.n199 VDPWR.t355 252.95
R7713 VDPWR.n155 VDPWR.t359 252.95
R7714 VDPWR.n160 VDPWR.t136 252.95
R7715 VDPWR.n165 VDPWR.t583 252.95
R7716 VDPWR.n170 VDPWR.t178 252.95
R7717 VDPWR.n68 VDPWR.t425 252.95
R7718 VDPWR.n73 VDPWR.t18 252.95
R7719 VDPWR.n78 VDPWR.t704 252.95
R7720 VDPWR.n112 VDPWR.t589 252.95
R7721 VDPWR.n107 VDPWR.t610 252.95
R7722 VDPWR.n120 VDPWR.t171 252.948
R7723 VDPWR.n245 VDPWR.t782 252.948
R7724 VDPWR.n240 VDPWR.t767 252.948
R7725 VDPWR.n235 VDPWR.t324 252.948
R7726 VDPWR.n230 VDPWR.t326 252.948
R7727 VDPWR.n225 VDPWR.t530 252.948
R7728 VDPWR.n220 VDPWR.t551 252.948
R7729 VDPWR.n215 VDPWR.t553 252.948
R7730 VDPWR.n210 VDPWR.t616 252.948
R7731 VDPWR.n629 VDPWR.t229 251.516
R7732 VDPWR.n349 VDPWR.t775 251.516
R7733 VDPWR.n92 VDPWR.t146 251.516
R7734 VDPWR.n540 VDPWR.t658 250.724
R7735 VDPWR.n260 VDPWR.t343 250.724
R7736 VDPWR.n3 VDPWR.t612 250.724
R7737 VDPWR.n144 VDPWR.t252 249.363
R7738 VDPWR.t700 VDPWR.t709 248.599
R7739 VDPWR.t422 VDPWR.t420 248.599
R7740 VDPWR.t50 VDPWR.t459 248.599
R7741 VDPWR.t751 VDPWR.t753 248.599
R7742 VDPWR.t350 VDPWR.t432 248.599
R7743 VDPWR.t629 VDPWR.t625 248.599
R7744 VDPWR.t172 VDPWR.t170 248.599
R7745 VDPWR.t783 VDPWR.t781 248.599
R7746 VDPWR.t768 VDPWR.t766 248.599
R7747 VDPWR.t321 VDPWR.t323 248.599
R7748 VDPWR.t327 VDPWR.t325 248.599
R7749 VDPWR.t527 VDPWR.t529 248.599
R7750 VDPWR.t548 VDPWR.t550 248.599
R7751 VDPWR.t554 VDPWR.t552 248.599
R7752 VDPWR.t613 VDPWR.t615 248.599
R7753 VDPWR.t651 VDPWR.t649 248.599
R7754 VDPWR.t253 VDPWR.t651 248.599
R7755 VDPWR.t251 VDPWR.t253 248.599
R7756 VDPWR.t177 VDPWR.t179 248.599
R7757 VDPWR.t582 VDPWR.t584 248.599
R7758 VDPWR.t135 VDPWR.t137 248.599
R7759 VDPWR.t358 VDPWR.t360 248.599
R7760 VDPWR.t354 VDPWR.t356 248.599
R7761 VDPWR.t517 VDPWR.t519 248.599
R7762 VDPWR.t218 VDPWR.t216 248.599
R7763 VDPWR.t212 VDPWR.t214 248.599
R7764 VDPWR.t617 VDPWR.t619 248.599
R7765 VDPWR.t706 VDPWR.t703 248.599
R7766 VDPWR.t262 VDPWR.t17 248.599
R7767 VDPWR.t461 VDPWR.t424 248.599
R7768 VDPWR.n632 VDPWR.t430 248.219
R7769 VDPWR.n352 VDPWR.t759 248.219
R7770 VDPWR.n95 VDPWR.t777 248.219
R7771 VDPWR.n2208 VDPWR.t1188 246.71
R7772 VDPWR.n1483 VDPWR.t1244 245.667
R7773 VDPWR.n1510 VDPWR.t1258 245.667
R7774 VDPWR.n1513 VDPWR.t1225 245.667
R7775 VDPWR.n1517 VDPWR.t1262 245.667
R7776 VDPWR.n1522 VDPWR.t1233 245.667
R7777 VDPWR.n1439 VDPWR.t1257 245.667
R7778 VDPWR.n1722 VDPWR.t1226 245.667
R7779 VDPWR.n1285 VDPWR.t1221 245.667
R7780 VDPWR.n1288 VDPWR.t1266 245.667
R7781 VDPWR.n1292 VDPWR.t1227 245.667
R7782 VDPWR.n1297 VDPWR.t1197 245.667
R7783 VDPWR.n1423 VDPWR.t1220 245.667
R7784 VDPWR.n1428 VDPWR.t1242 245.667
R7785 VDPWR.n1905 VDPWR.t1186 245.667
R7786 VDPWR.n1911 VDPWR.t1169 245.667
R7787 VDPWR.n1914 VDPWR.t1251 245.667
R7788 VDPWR.n1918 VDPWR.t1229 245.667
R7789 VDPWR.n2053 VDPWR.t1232 245.667
R7790 VDPWR.n2056 VDPWR.t1203 245.667
R7791 VDPWR.n2212 VDPWR.t1254 245.667
R7792 VDPWR.n2215 VDPWR.t1183 245.667
R7793 VDPWR.n1175 VDPWR.t1234 245.667
R7794 VDPWR.n2444 VDPWR.t1167 245.667
R7795 VDPWR.n963 VDPWR.t1218 245.667
R7796 VDPWR.n966 VDPWR.t1277 245.667
R7797 VDPWR.n2464 VDPWR.t1190 245.667
R7798 VDPWR.n2467 VDPWR.t1253 245.667
R7799 VDPWR.n2596 VDPWR.t1179 245.667
R7800 VDPWR.n2599 VDPWR.t1278 245.667
R7801 VDPWR.n926 VDPWR.t1267 245.667
R7802 VDPWR.n2922 VDPWR.t1180 245.667
R7803 VDPWR.n2960 VDPWR.t1285 245.667
R7804 VDPWR.n2968 VDPWR.t1256 245.667
R7805 VDPWR.n814 VDPWR.t1265 245.667
R7806 VDPWR.n2632 VDPWR.t1274 245.667
R7807 VDPWR.n2635 VDPWR.t1211 245.667
R7808 VDPWR.n827 VDPWR.t1248 245.667
R7809 VDPWR.n831 VDPWR.t1185 245.667
R7810 VDPWR.n1029 VDPWR.t78 245.064
R7811 VDPWR.n2016 VDPWR.t506 243.512
R7812 VDPWR.n793 VDPWR.t750 241.767
R7813 VDPWR.n1160 VDPWR.t638 240.215
R7814 VDPWR.n2957 VDPWR.t642 240.214
R7815 VDPWR.n1379 VDPWR.t1181 235.319
R7816 VDPWR.n2674 VDPWR.t621 234.982
R7817 VDPWR VDPWR.t637 233.304
R7818 VDPWR.t1138 VDPWR.t762 231.625
R7819 VDPWR.t77 VDPWR.t199 229.947
R7820 VDPWR.n146 VDPWR 224.923
R7821 VDPWR.n2656 VDPWR.n2655 223.868
R7822 VDPWR.t124 VDPWR 223.233
R7823 VDPWR.t336 VDPWR 223.233
R7824 VDPWR.n620 VDPWR 221.964
R7825 VDPWR.n340 VDPWR 221.964
R7826 VDPWR.n83 VDPWR 221.964
R7827 VDPWR.t755 VDPWR.t371 221.555
R7828 VDPWR.t69 VDPWR.t71 221.555
R7829 VDPWR.t191 VDPWR.t270 221.555
R7830 VDPWR.n2895 VDPWR.n897 221.314
R7831 VDPWR.n1839 VDPWR.t1189 215.827
R7832 VDPWR.n2715 VDPWR.t1280 215.827
R7833 VDPWR VDPWR.t561 213.163
R7834 VDPWR VDPWR.t1163 213.163
R7835 VDPWR.n1415 VDPWR.t1166 213.148
R7836 VDPWR.n1420 VDPWR.t1237 213.148
R7837 VDPWR.n2589 VDPWR.t1176 213.148
R7838 VDPWR.n2592 VDPWR.t1276 213.148
R7839 VDPWR.n580 VDPWR.n577 213.119
R7840 VDPWR.n300 VDPWR.n297 213.119
R7841 VDPWR.n43 VDPWR.n40 213.119
R7842 VDPWR.n621 VDPWR.n620 213.119
R7843 VDPWR.n640 VDPWR.n639 213.119
R7844 VDPWR.n341 VDPWR.n340 213.119
R7845 VDPWR.n360 VDPWR.n359 213.119
R7846 VDPWR.n176 VDPWR.n175 213.119
R7847 VDPWR.n136 VDPWR.n134 213.119
R7848 VDPWR.n148 VDPWR.n147 213.119
R7849 VDPWR.n146 VDPWR.n145 213.119
R7850 VDPWR.n2531 VDPWR.n2530 213.119
R7851 VDPWR.n2847 VDPWR.n882 213.119
R7852 VDPWR.n3036 VDPWR.n787 213.119
R7853 VDPWR.n84 VDPWR.n83 213.119
R7854 VDPWR.n103 VDPWR.n102 213.119
R7855 VDPWR.n532 VDPWR.t699 212.081
R7856 VDPWR.n533 VDPWR.t708 212.081
R7857 VDPWR.n3111 VDPWR.t705 212.081
R7858 VDPWR.n3112 VDPWR.t702 212.081
R7859 VDPWR.n1247 VDPWR.t1240 211.263
R7860 VDPWR.n597 VDPWR.t1205 210.964
R7861 VDPWR.n588 VDPWR.t1261 210.964
R7862 VDPWR.n574 VDPWR.t1214 210.964
R7863 VDPWR.n549 VDPWR.t1207 210.964
R7864 VDPWR.n317 VDPWR.t1263 210.964
R7865 VDPWR.n308 VDPWR.t1201 210.964
R7866 VDPWR.n294 VDPWR.t1200 210.964
R7867 VDPWR.n269 VDPWR.t1228 210.964
R7868 VDPWR.n2015 VDPWR.t1275 210.964
R7869 VDPWR.n2350 VDPWR.t1273 210.964
R7870 VDPWR.n2430 VDPWR.t1284 210.964
R7871 VDPWR.n1118 VDPWR.t1236 210.964
R7872 VDPWR.n2902 VDPWR.t1270 210.964
R7873 VDPWR.n2654 VDPWR.t1269 210.964
R7874 VDPWR.n60 VDPWR.t1215 210.964
R7875 VDPWR.n51 VDPWR.t1282 210.964
R7876 VDPWR.n37 VDPWR.t1268 210.964
R7877 VDPWR.n12 VDPWR.t1217 210.964
R7878 VDPWR.n1589 VDPWR.n1588 209.368
R7879 VDPWR.n1789 VDPWR.n1367 209.368
R7880 VDPWR.n1846 VDPWR.n1330 209.368
R7881 VDPWR.n2116 VDPWR.n2003 209.368
R7882 VDPWR.n2002 VDPWR.n1963 209.368
R7883 VDPWR.n2365 VDPWR.n1205 209.368
R7884 VDPWR.n1251 VDPWR.n1250 209.368
R7885 VDPWR.n2533 VDPWR.n2532 209.368
R7886 VDPWR.n2849 VDPWR.n2848 209.368
R7887 VDPWR.t6 VDPWR 206.45
R7888 VDPWR VDPWR.t1149 203.093
R7889 VDPWR.t852 VDPWR 203.093
R7890 VDPWR.t1154 VDPWR 203.093
R7891 VDPWR.t1048 VDPWR 203.093
R7892 VDPWR VDPWR.t876 203.093
R7893 VDPWR VDPWR.t675 201.413
R7894 VDPWR VDPWR.t181 199.736
R7895 VDPWR VDPWR.t693 199.736
R7896 VDPWR.t709 VDPWR 198.287
R7897 VDPWR.t420 VDPWR 198.287
R7898 VDPWR.t459 VDPWR 198.287
R7899 VDPWR.t753 VDPWR 198.287
R7900 VDPWR.t432 VDPWR 198.287
R7901 VDPWR.t625 VDPWR 198.287
R7902 VDPWR VDPWR.t177 198.287
R7903 VDPWR VDPWR.t582 198.287
R7904 VDPWR VDPWR.t135 198.287
R7905 VDPWR VDPWR.t358 198.287
R7906 VDPWR VDPWR.t354 198.287
R7907 VDPWR VDPWR.t517 198.287
R7908 VDPWR VDPWR.t218 198.287
R7909 VDPWR VDPWR.t212 198.287
R7910 VDPWR VDPWR.t617 198.287
R7911 VDPWR.t703 VDPWR 198.287
R7912 VDPWR.t17 VDPWR 198.287
R7913 VDPWR.t424 VDPWR 198.287
R7914 VDPWR.t721 VDPWR.t112 198.058
R7915 VDPWR.n2167 VDPWR.n2166 197.508
R7916 VDPWR.t370 VDPWR.t2 191.344
R7917 VDPWR.t92 VDPWR.t513 191.344
R7918 VDPWR.t159 VDPWR.t122 191.344
R7919 VDPWR.t717 VDPWR.t679 189.665
R7920 VDPWR VDPWR.t251 189.409
R7921 VDPWR.n2531 VDPWR 184.63
R7922 VDPWR.n787 VDPWR 184.63
R7923 VDPWR.n642 VDPWR.n641 183.673
R7924 VDPWR.n362 VDPWR.n361 183.673
R7925 VDPWR.n105 VDPWR.n104 183.673
R7926 VDPWR.n534 VDPWR.n533 183.441
R7927 VDPWR.n3113 VDPWR.n3112 183.441
R7928 VDPWR VDPWR.t35 182.952
R7929 VDPWR VDPWR.n640 182.952
R7930 VDPWR.t515 VDPWR 182.952
R7931 VDPWR VDPWR.t623 182.952
R7932 VDPWR VDPWR.n360 182.952
R7933 VDPWR.t118 VDPWR 182.952
R7934 VDPWR VDPWR.t834 182.952
R7935 VDPWR.t891 VDPWR 182.952
R7936 VDPWR.t855 VDPWR 182.952
R7937 VDPWR VDPWR.t924 182.952
R7938 VDPWR.n1367 VDPWR 182.952
R7939 VDPWR.t1007 VDPWR 182.952
R7940 VDPWR VDPWR.t1021 182.952
R7941 VDPWR.t918 VDPWR 182.952
R7942 VDPWR.t988 VDPWR 182.952
R7943 VDPWR.t849 VDPWR 182.952
R7944 VDPWR.t831 VDPWR 182.952
R7945 VDPWR.t912 VDPWR 182.952
R7946 VDPWR.t936 VDPWR 182.952
R7947 VDPWR VDPWR.t143 182.952
R7948 VDPWR VDPWR.n103 182.952
R7949 VDPWR.t450 VDPWR 182.952
R7950 VDPWR.t255 VDPWR.t27 181.273
R7951 VDPWR.n1587 VDPWR 179.595
R7952 VDPWR VDPWR.n1330 179.595
R7953 VDPWR.n1250 VDPWR 179.595
R7954 VDPWR.n1205 VDPWR 179.595
R7955 VDPWR.n2674 VDPWR 179.595
R7956 VDPWR.t29 VDPWR.t486 174.559
R7957 VDPWR.t670 VDPWR.t81 174.559
R7958 VDPWR.t525 VDPWR.t755 172.881
R7959 VDPWR.t71 VDPWR.t563 172.881
R7960 VDPWR.t242 VDPWR.t191 172.881
R7961 VDPWR.t232 VDPWR.t412 172.881
R7962 VDPWR.t155 VDPWR 169.524
R7963 VDPWR.t486 VDPWR.t126 167.845
R7964 VDPWR.t523 VDPWR.t858 164.488
R7965 VDPWR.t600 VDPWR.t719 162.81
R7966 VDPWR.t97 VDPWR.t120 162.81
R7967 VDPWR.t681 VDPWR.t1162 161.131
R7968 VDPWR.t153 VDPWR.t25 161.131
R7969 VDPWR.n544 VDPWR.n543 159.476
R7970 VDPWR.n264 VDPWR.n263 159.476
R7971 VDPWR.n1106 VDPWR.n1105 159.476
R7972 VDPWR.n2559 VDPWR.n2558 159.476
R7973 VDPWR.n7 VDPWR.n6 159.476
R7974 VDPWR.t369 VDPWR.t525 159.452
R7975 VDPWR.t605 VDPWR.t234 159.452
R7976 VDPWR.t779 VDPWR.t237 159.452
R7977 VDPWR.t563 VDPWR.t514 159.452
R7978 VDPWR.t270 VDPWR.t243 159.452
R7979 VDPWR.t160 VDPWR.t242 159.452
R7980 VDPWR.t558 VDPWR.t348 159.452
R7981 VDPWR.t1160 VDPWR.t947 157.774
R7982 VDPWR.n631 VDPWR.t267 157.014
R7983 VDPWR.n351 VDPWR.t435 157.014
R7984 VDPWR.n94 VDPWR.t20 157.014
R7985 VDPWR.t657 VDPWR.t56 154.417
R7986 VDPWR.t342 VDPWR.t107 154.417
R7987 VDPWR.t1089 VDPWR.t1058 154.417
R7988 VDPWR.t11 VDPWR.t283 154.417
R7989 VDPWR.t897 VDPWR.t961 154.417
R7990 VDPWR.t1162 VDPWR.t508 154.417
R7991 VDPWR.t611 VDPWR.t457 154.417
R7992 VDPWR VDPWR.t747 152.739
R7993 VDPWR.t858 VDPWR.t281 151.06
R7994 VDPWR.t906 VDPWR.t819 151.06
R7995 VDPWR.t576 VDPWR.t885 151.06
R7996 VDPWR.t653 VDPWR.t73 149.382
R7997 VDPWR.t436 VDPWR.t210 149.382
R7998 VDPWR.t226 VDPWR.t266 147.703
R7999 VDPWR.t238 VDPWR.t434 147.703
R8000 VDPWR.t67 VDPWR.t203 147.703
R8001 VDPWR.t598 VDPWR.t8 147.703
R8002 VDPWR.t693 VDPWR.t95 147.703
R8003 VDPWR.t621 VDPWR.t83 147.703
R8004 VDPWR.t666 VDPWR.t220 147.703
R8005 VDPWR.t249 VDPWR.t258 147.703
R8006 VDPWR.t477 VDPWR.t1160 147.703
R8007 VDPWR.t442 VDPWR.t260 147.703
R8008 VDPWR.t631 VDPWR.t19 147.703
R8009 VDPWR.t479 VDPWR.t436 144.346
R8010 VDPWR.t471 VDPWR.t62 144.346
R8011 VDPWR.t475 VDPWR.t473 144.346
R8012 VDPWR.t473 VDPWR.t809 144.346
R8013 VDPWR.t809 VDPWR.t803 144.346
R8014 VDPWR.t803 VDPWR.t813 144.346
R8015 VDPWR.t813 VDPWR.t817 144.346
R8016 VDPWR.t817 VDPWR.t789 144.346
R8017 VDPWR.t793 VDPWR.t815 144.346
R8018 VDPWR.t815 VDPWR.t787 144.346
R8019 VDPWR.t791 VDPWR.t795 144.346
R8020 VDPWR.t795 VDPWR.t805 144.346
R8021 VDPWR.t799 VDPWR.t801 144.346
R8022 VDPWR.t801 VDPWR.t797 144.346
R8023 VDPWR.t797 VDPWR.t807 144.346
R8024 VDPWR.t807 VDPWR.t811 144.346
R8025 VDPWR.t493 VDPWR.t499 144.346
R8026 VDPWR.t499 VDPWR.t497 144.346
R8027 VDPWR.t497 VDPWR.t491 144.346
R8028 VDPWR.t491 VDPWR.t293 144.346
R8029 VDPWR.t293 VDPWR.t299 144.346
R8030 VDPWR.t303 VDPWR.t307 144.346
R8031 VDPWR.t307 VDPWR.t297 144.346
R8032 VDPWR.t297 VDPWR.t301 144.346
R8033 VDPWR.t301 VDPWR.t305 144.346
R8034 VDPWR.t305 VDPWR.t295 144.346
R8035 VDPWR.t311 VDPWR.t317 144.346
R8036 VDPWR.t317 VDPWR.t289 144.346
R8037 VDPWR.t289 VDPWR.t291 144.346
R8038 VDPWR.t291 VDPWR.t315 144.346
R8039 VDPWR.t315 VDPWR.t287 144.346
R8040 VDPWR.t287 VDPWR.t309 144.346
R8041 VDPWR.t390 VDPWR.t396 144.346
R8042 VDPWR.t400 VDPWR.t408 144.346
R8043 VDPWR.t394 VDPWR.t404 144.346
R8044 VDPWR.t384 VDPWR.t386 144.346
R8045 VDPWR.t743 VDPWR.t741 144.346
R8046 VDPWR.t81 VDPWR.t163 144.346
R8047 VDPWR.t281 VDPWR.t369 142.668
R8048 VDPWR.t787 VDPWR.t791 142.668
R8049 VDPWR.t402 VDPWR.t398 142.668
R8050 VDPWR.t514 VDPWR.t578 142.668
R8051 VDPWR.t151 VDPWR.t160 142.668
R8052 VDPWR.t543 VDPWR.t232 142.668
R8053 VDPWR.t426 VDPWR.t264 140.989
R8054 VDPWR.t266 VDPWR.t429 140.989
R8055 VDPWR.t531 VDPWR.t533 140.989
R8056 VDPWR.t655 VDPWR.t657 140.989
R8057 VDPWR.t273 VDPWR.t116 140.989
R8058 VDPWR.t109 VDPWR.t101 140.989
R8059 VDPWR.t434 VDPWR.t758 140.989
R8060 VDPWR.t133 VDPWR.t131 140.989
R8061 VDPWR.t344 VDPWR.t342 140.989
R8062 VDPWR.t37 VDPWR.t346 140.989
R8063 VDPWR.t244 VDPWR.t523 140.989
R8064 VDPWR.t205 VDPWR.t440 140.989
R8065 VDPWR.t181 VDPWR.t183 140.989
R8066 VDPWR.t90 VDPWR.t565 140.989
R8067 VDPWR.t513 VDPWR.t564 140.989
R8068 VDPWR.t561 VDPWR.t58 140.989
R8069 VDPWR.t332 VDPWR.t124 140.989
R8070 VDPWR.t243 VDPWR.t159 140.989
R8071 VDPWR.t539 VDPWR.t240 140.989
R8072 VDPWR.t412 VDPWR.t643 140.989
R8073 VDPWR.t574 VDPWR.t664 140.989
R8074 VDPWR.t85 VDPWR.t448 140.989
R8075 VDPWR.t511 VDPWR.t510 140.989
R8076 VDPWR.t1163 VDPWR.t60 140.989
R8077 VDPWR.t168 VDPWR.t824 140.989
R8078 VDPWR.t373 VDPWR.t168 140.989
R8079 VDPWR.t633 VDPWR.t645 140.989
R8080 VDPWR.t54 VDPWR.t15 140.989
R8081 VDPWR.t19 VDPWR.t776 140.989
R8082 VDPWR.t588 VDPWR.t590 140.989
R8083 VDPWR.t609 VDPWR.t611 140.989
R8084 VDPWR.t683 VDPWR.t41 140.989
R8085 VDPWR.n532 VDPWR.t1193 139.78
R8086 VDPWR.n533 VDPWR.t1202 139.78
R8087 VDPWR.n3111 VDPWR.t1206 139.78
R8088 VDPWR.n3112 VDPWR.t1212 139.78
R8089 VDPWR.t719 VDPWR.t770 139.311
R8090 VDPWR.t440 VDPWR.t607 137.633
R8091 VDPWR.t444 VDPWR.t0 137.633
R8092 VDPWR.n631 VDPWR.t724 137.079
R8093 VDPWR.n351 VDPWR.t568 137.079
R8094 VDPWR.n94 VDPWR.t698 137.079
R8095 VDPWR.t13 VDPWR.t736 135.954
R8096 VDPWR.t739 VDPWR.t268 135.954
R8097 VDPWR.t364 VDPWR.t446 135.954
R8098 VDPWR.t413 VDPWR.t79 135.954
R8099 VDPWR.t121 VDPWR.t88 135.954
R8100 VDPWR.t641 VDPWR 135.954
R8101 VDPWR.n1066 VDPWR.t365 135.268
R8102 VDPWR.t166 VDPWR.t594 134.276
R8103 VDPWR.t510 VDPWR.t193 130.919
R8104 VDPWR.t512 VDPWR.t545 130.919
R8105 VDPWR.n2487 VDPWR.t1247 129.344
R8106 VDPWR.n2985 VDPWR.t1250 129.344
R8107 VDPWR.n860 VDPWR.t1259 129.344
R8108 VDPWR.n2757 VDPWR.t1255 129.344
R8109 VDPWR.n2782 VDPWR.t1194 129.344
R8110 VDPWR VDPWR.t526 129.24
R8111 VDPWR.n2695 VDPWR.t1182 127.695
R8112 VDPWR.t521 VDPWR.t392 127.562
R8113 VDPWR.n2848 VDPWR.t334 127.562
R8114 VDPWR.t23 VDPWR.t31 127.562
R8115 VDPWR VDPWR.t255 127.562
R8116 VDPWR.n577 VDPWR 125.883
R8117 VDPWR.n641 VDPWR 125.883
R8118 VDPWR.n297 VDPWR 125.883
R8119 VDPWR.n361 VDPWR 125.883
R8120 VDPWR.t861 VDPWR 125.883
R8121 VDPWR.n1588 VDPWR 125.883
R8122 VDPWR VDPWR.n1587 125.883
R8123 VDPWR.t941 VDPWR 125.883
R8124 VDPWR.n1330 VDPWR 125.883
R8125 VDPWR.n1367 VDPWR 125.883
R8126 VDPWR.t846 VDPWR 125.883
R8127 VDPWR.n2002 VDPWR 125.883
R8128 VDPWR.n2003 VDPWR 125.883
R8129 VDPWR.t930 VDPWR 125.883
R8130 VDPWR.n1250 VDPWR 125.883
R8131 VDPWR VDPWR.n1205 125.883
R8132 VDPWR.t1029 VDPWR 125.883
R8133 VDPWR.t606 VDPWR.t731 125.883
R8134 VDPWR VDPWR.n2531 125.883
R8135 VDPWR.t894 VDPWR 125.883
R8136 VDPWR.n2848 VDPWR 125.883
R8137 VDPWR.t348 VDPWR.t187 125.883
R8138 VDPWR.t149 VDPWR.t501 125.883
R8139 VDPWR VDPWR.n2847 125.883
R8140 VDPWR.t879 VDPWR 125.883
R8141 VDPWR VDPWR.n787 125.883
R8142 VDPWR.n40 VDPWR 125.883
R8143 VDPWR.n104 VDPWR 125.883
R8144 VDPWR.n974 VDPWR.t1231 124.953
R8145 VDPWR.t677 VDPWR.t390 124.206
R8146 VDPWR.t334 VDPWR.t189 124.206
R8147 VDPWR.t157 VDPWR.t727 124.206
R8148 VDPWR.t209 VDPWR 122.526
R8149 VDPWR.t406 VDPWR.t33 122.526
R8150 VDPWR.t380 VDPWR.t488 122.526
R8151 VDPWR.n2532 VDPWR.t384 122.526
R8152 VDPWR.t603 VDPWR.t821 122.526
R8153 VDPWR.t994 VDPWR.t313 120.849
R8154 VDPWR.t165 VDPWR.t733 120.849
R8155 VDPWR.t637 VDPWR.t490 120.849
R8156 VDPWR.t692 VDPWR.t641 120.849
R8157 VDPWR.n817 VDPWR.t1245 120.76
R8158 VDPWR.n983 VDPWR.t1204 119.007
R8159 VDPWR.n2040 VDPWR.t1196 118.853
R8160 VDPWR.n1066 VDPWR.t593 118.549
R8161 VDPWR.t112 VDPWR.t674 117.492
R8162 VDPWR.n998 VDPWR.t34 117.451
R8163 VDPWR.n2672 VDPWR.t597 117.451
R8164 VDPWR.n2680 VDPWR.t164 117.451
R8165 VDPWR.n1665 VDPWR.t1171 117.294
R8166 VDPWR.n2231 VDPWR.t1243 117.294
R8167 VDPWR.n3030 VDPWR.t1198 117.294
R8168 VDPWR.n2703 VDPWR.t748 116.343
R8169 VDPWR.n569 VDPWR.t427 116.341
R8170 VDPWR.n550 VDPWR.t117 116.341
R8171 VDPWR.n289 VDPWR.t110 116.341
R8172 VDPWR.n270 VDPWR.t347 116.341
R8173 VDPWR.n894 VDPWR.t28 116.341
R8174 VDPWR.n791 VDPWR.t646 116.341
R8175 VDPWR.n32 VDPWR.t55 116.341
R8176 VDPWR.n13 VDPWR.t42 116.341
R8177 VDPWR.t729 VDPWR 115.814
R8178 VDPWR.n1092 VDPWR.t732 114.918
R8179 VDPWR.n809 VDPWR.t718 114.918
R8180 VDPWR.n1507 VDPWR.t1239 114.546
R8181 VDPWR.n1282 VDPWR.t1199 114.546
R8182 VDPWR.n1923 VDPWR.t1241 114.546
R8183 VDPWR.t505 VDPWR.t285 114.135
R8184 VDPWR.t398 VDPWR.t764 114.135
R8185 VDPWR.n1402 VDPWR.t756 113.98
R8186 VDPWR.n2032 VDPWR.t654 113.98
R8187 VDPWR.n1084 VDPWR.t447 113.98
R8188 VDPWR.n1140 VDPWR.t72 113.98
R8189 VDPWR.n919 VDPWR.t233 113.98
R8190 VDPWR.n922 VDPWR.t339 113.98
R8191 VDPWR.n944 VDPWR.t272 113.98
R8192 VDPWR.n943 VDPWR.t192 113.98
R8193 VDPWR.n2942 VDPWR.t546 113.98
R8194 VDPWR.n876 VDPWR.t100 113.98
R8195 VDPWR.t264 VDPWR 112.457
R8196 VDPWR.t429 VDPWR 112.457
R8197 VDPWR VDPWR.t273 112.457
R8198 VDPWR.t101 VDPWR 112.457
R8199 VDPWR.t758 VDPWR 112.457
R8200 VDPWR VDPWR.t37 112.457
R8201 VDPWR VDPWR.t633 112.457
R8202 VDPWR.t15 VDPWR 112.457
R8203 VDPWR.t776 VDPWR 112.457
R8204 VDPWR VDPWR.t683 112.457
R8205 VDPWR.t687 VDPWR 110.778
R8206 VDPWR.t62 VDPWR 110.778
R8207 VDPWR.t114 VDPWR.t277 110.778
R8208 VDPWR VDPWR.t737 109.1
R8209 VDPWR VDPWR.t340 109.1
R8210 VDPWR.t203 VDPWR 109.1
R8211 VDPWR VDPWR.t598 109.1
R8212 VDPWR VDPWR.t822 109.1
R8213 VDPWR.t819 VDPWR 109.1
R8214 VDPWR.t503 VDPWR 109.1
R8215 VDPWR.t695 VDPWR 109.1
R8216 VDPWR VDPWR.t352 109.1
R8217 VDPWR VDPWR.t375 109.1
R8218 VDPWR.t21 VDPWR 109.1
R8219 VDPWR.t679 VDPWR 109.1
R8220 VDPWR.t260 VDPWR 109.1
R8221 VDPWR VDPWR.t197 109.1
R8222 VDPWR.t760 VDPWR 107.421
R8223 VDPWR.t438 VDPWR.t185 107.421
R8224 VDPWR.t490 VDPWR 107.421
R8225 VDPWR.t958 VDPWR 107.421
R8226 VDPWR.n1587 VDPWR.n1459 106.561
R8227 VDPWR.n2675 VDPWR.n2674 106.559
R8228 VDPWR.n716 VDPWR.n704 105.788
R8229 VDPWR.n700 VDPWR.n688 105.788
R8230 VDPWR.n684 VDPWR.n672 105.788
R8231 VDPWR.n668 VDPWR.n657 105.788
R8232 VDPWR.n527 VDPWR.n515 105.788
R8233 VDPWR.n511 VDPWR.n499 105.788
R8234 VDPWR.n495 VDPWR.n483 105.788
R8235 VDPWR.n479 VDPWR.n467 105.788
R8236 VDPWR.n463 VDPWR.n403 105.788
R8237 VDPWR.n457 VDPWR.n445 105.788
R8238 VDPWR.n441 VDPWR.n429 105.788
R8239 VDPWR.n425 VDPWR.n414 105.788
R8240 VDPWR.n3107 VDPWR.n759 105.788
R8241 VDPWR.n3101 VDPWR.n3089 105.788
R8242 VDPWR.n3085 VDPWR.n3073 105.788
R8243 VDPWR.n3069 VDPWR.n3057 105.788
R8244 VDPWR VDPWR.t1069 105.743
R8245 VDPWR VDPWR.t1063 105.743
R8246 VDPWR VDPWR.t976 105.743
R8247 VDPWR.t915 VDPWR 105.743
R8248 VDPWR.t279 VDPWR.t329 105.743
R8249 VDPWR.t1072 VDPWR.t426 104.064
R8250 VDPWR.t116 VDPWR.t1086 104.064
R8251 VDPWR.t1004 VDPWR.t109 104.064
R8252 VDPWR.t346 VDPWR.t944 104.064
R8253 VDPWR.t382 VDPWR 104.064
R8254 VDPWR.t537 VDPWR 104.064
R8255 VDPWR VDPWR.t128 104.064
R8256 VDPWR.t645 VDPWR.t1032 104.064
R8257 VDPWR.t933 VDPWR.t54 104.064
R8258 VDPWR.t41 VDPWR.t1066 104.064
R8259 VDPWR.t52 VDPWR 102.385
R8260 VDPWR.t627 VDPWR 102.385
R8261 VDPWR.t222 VDPWR.t77 102.385
R8262 VDPWR.t578 VDPWR 102.385
R8263 VDPWR.t580 VDPWR 102.385
R8264 VDPWR.t947 VDPWR 102.385
R8265 VDPWR.t647 VDPWR 102.385
R8266 VDPWR.n2166 VDPWR.n2165 101.591
R8267 VDPWR VDPWR.t452 100.707
R8268 VDPWR.t230 VDPWR 99.0288
R8269 VDPWR.t772 VDPWR 99.0288
R8270 VDPWR.t1035 VDPWR.t303 99.0288
R8271 VDPWR.t199 VDPWR 99.0288
R8272 VDPWR VDPWR.t141 99.0288
R8273 VDPWR.t147 VDPWR 99.0288
R8274 VDPWR.t170 VDPWR 97.6641
R8275 VDPWR.t781 VDPWR 97.6641
R8276 VDPWR.t766 VDPWR 97.6641
R8277 VDPWR.t323 VDPWR 97.6641
R8278 VDPWR.t325 VDPWR 97.6641
R8279 VDPWR.t529 VDPWR 97.6641
R8280 VDPWR.t550 VDPWR 97.6641
R8281 VDPWR.t552 VDPWR 97.6641
R8282 VDPWR.t615 VDPWR 97.6641
R8283 VDPWR.t592 VDPWR.t605 97.3503
R8284 VDPWR.n564 VDPWR.t227 96.1553
R8285 VDPWR.n539 VDPWR.t106 96.1553
R8286 VDPWR.n284 VDPWR.t239 96.1553
R8287 VDPWR.n259 VDPWR.t686 96.1553
R8288 VDPWR.n1042 VDPWR.t720 96.1553
R8289 VDPWR.n1120 VDPWR.t96 96.1553
R8290 VDPWR.n991 VDPWR.t522 96.1553
R8291 VDPWR.n27 VDPWR.t632 96.1553
R8292 VDPWR.n2 VDPWR.t40 96.1553
R8293 VDPWR.t187 VDPWR.t338 95.6719
R8294 VDPWR.t338 VDPWR.t830 95.6719
R8295 VDPWR.t415 VDPWR.t139 95.6719
R8296 VDPWR.n2031 VDPWR.t208 93.81
R8297 VDPWR.n900 VDPWR.t150 93.81
R8298 VDPWR.n903 VDPWR.t80 93.81
R8299 VDPWR.n745 VDPWR.n740 92.5005
R8300 VDPWR.n741 VDPWR.n739 92.5005
R8301 VDPWR VDPWR.t105 92.315
R8302 VDPWR VDPWR.t685 92.315
R8303 VDPWR.t378 VDPWR.t668 92.315
R8304 VDPWR VDPWR.t39 92.315
R8305 VDPWR.t526 VDPWR.t10 90.6365
R8306 VDPWR.t888 VDPWR.t155 90.6365
R8307 VDPWR.t1165 VDPWR.t507 90.6365
R8308 VDPWR.t275 VDPWR.t512 90.6365
R8309 VDPWR.n743 VDPWR.n741 89.0328
R8310 VDPWR.n746 VDPWR.n745 89.0328
R8311 VDPWR.t805 VDPWR 88.9581
R8312 VDPWR.t367 VDPWR.t207 87.2797
R8313 VDPWR.t745 VDPWR.t635 87.2797
R8314 VDPWR VDPWR.t691 87.2797
R8315 VDPWR.n543 VDPWR.t57 86.7743
R8316 VDPWR.n263 VDPWR.t108 86.7743
R8317 VDPWR.n1105 VDPWR.t694 86.7743
R8318 VDPWR.n2559 VDPWR.t678 86.7743
R8319 VDPWR.n1010 VDPWR.t489 86.7743
R8320 VDPWR.n1010 VDPWR.t669 86.7743
R8321 VDPWR.n2662 VDPWR.t487 86.7743
R8322 VDPWR.n2662 VDPWR.t30 86.7743
R8323 VDPWR.n2678 VDPWR.t671 86.7743
R8324 VDPWR.n2678 VDPWR.t82 86.7743
R8325 VDPWR.n6 VDPWR.t458 86.7743
R8326 VDPWR VDPWR.t311 85.6012
R8327 VDPWR.t130 VDPWR 85.6012
R8328 VDPWR.n577 VDPWR.t230 83.9228
R8329 VDPWR.n297 VDPWR.t772 83.9228
R8330 VDPWR.t284 VDPWR.t454 83.9228
R8331 VDPWR.t735 VDPWR.t438 83.9228
R8332 VDPWR.t141 VDPWR.t900 83.9228
R8333 VDPWR.n40 VDPWR.t147 83.9228
R8334 VDPWR.t741 VDPWR 82.2443
R8335 VDPWR.t99 VDPWR.t1165 82.2443
R8336 VDPWR.n640 VDPWR.t723 80.5659
R8337 VDPWR.n360 VDPWR.t567 80.5659
R8338 VDPWR.t495 VDPWR 80.5659
R8339 VDPWR.t564 VDPWR.t1119 80.5659
R8340 VDPWR.t58 VDPWR 80.5659
R8341 VDPWR VDPWR.t539 80.5659
R8342 VDPWR.t541 VDPWR 80.5659
R8343 VDPWR.t277 VDPWR.t511 80.5659
R8344 VDPWR.t60 VDPWR 80.5659
R8345 VDPWR.n103 VDPWR.t697 80.5659
R8346 VDPWR.t733 VDPWR.t779 78.8874
R8347 VDPWR.t1119 VDPWR.t69 78.8874
R8348 VDPWR.t572 VDPWR.t543 78.8874
R8349 VDPWR VDPWR.t596 78.8874
R8350 VDPWR.t163 VDPWR 78.8874
R8351 VDPWR.t35 VDPWR.t1072 77.209
R8352 VDPWR.t1086 VDPWR.t515 77.209
R8353 VDPWR.t623 VDPWR.t1004 77.209
R8354 VDPWR.t944 VDPWR.t118 77.209
R8355 VDPWR.t830 VDPWR.t559 77.209
R8356 VDPWR.t1032 VDPWR.t689 77.209
R8357 VDPWR.t876 VDPWR.t912 77.209
R8358 VDPWR.t143 VDPWR.t933 77.209
R8359 VDPWR.t1066 VDPWR.t450 77.209
R8360 VDPWR.t789 VDPWR.t837 75.5305
R8361 VDPWR.t725 VDPWR.t378 75.5305
R8362 VDPWR VDPWR.t153 75.5305
R8363 VDPWR.t596 VDPWR 75.5305
R8364 VDPWR.t43 VDPWR.n733 75.1466
R8365 VDPWR.n735 VDPWR.t47 75.1466
R8366 VDPWR.t2 VDPWR.t205 73.8521
R8367 VDPWR.t140 VDPWR.t785 73.8521
R8368 VDPWR.t448 VDPWR.t1135 73.8521
R8369 VDPWR.t586 VDPWR 73.8521
R8370 VDPWR.t73 VDPWR.t367 72.1736
R8371 VDPWR.t207 VDPWR.t284 72.1736
R8372 VDPWR.t386 VDPWR 72.1736
R8373 VDPWR VDPWR.t495 72.1736
R8374 VDPWR.n744 VDPWR.n743 70.6952
R8375 VDPWR.n747 VDPWR.n746 70.6952
R8376 VDPWR.t837 VDPWR.t793 68.8168
R8377 VDPWR.t388 VDPWR.t725 68.8168
R8378 VDPWR.t507 VDPWR.t275 68.8168
R8379 VDPWR VDPWR.t29 68.8168
R8380 VDPWR VDPWR.t90 67.1383
R8381 VDPWR.t189 VDPWR.t140 67.1383
R8382 VDPWR.t785 VDPWR.t558 67.1383
R8383 VDPWR.t1135 VDPWR.t729 67.1383
R8384 VDPWR.t691 VDPWR 67.1383
R8385 VDPWR.n544 VDPWR.t738 66.8398
R8386 VDPWR.n264 VDPWR.t341 66.8398
R8387 VDPWR.n1106 VDPWR.t200 66.8398
R8388 VDPWR.n2558 VDPWR.t7 66.8398
R8389 VDPWR.n7 VDPWR.t198 66.8398
R8390 VDPWR.t731 VDPWR.t224 65.4599
R8391 VDPWR VDPWR.t85 65.4599
R8392 VDPWR.t824 VDPWR 65.4599
R8393 VDPWR.n386 VDPWR.n378 64.4072
R8394 VDPWR.n398 VDPWR.n390 64.4072
R8395 VDPWR.t410 VDPWR.t606 63.7814
R8396 VDPWR.t559 VDPWR.t415 63.7814
R8397 VDPWR.t139 VDPWR.t572 63.7814
R8398 VDPWR.n699 VDPWR.n698 63.3551
R8399 VDPWR.n683 VDPWR.n682 63.3551
R8400 VDPWR.n510 VDPWR.n509 63.3551
R8401 VDPWR.n494 VDPWR.n493 63.3551
R8402 VDPWR.n456 VDPWR.n455 63.3551
R8403 VDPWR.n440 VDPWR.n439 63.3551
R8404 VDPWR.n3100 VDPWR.n3099 63.3551
R8405 VDPWR.n3084 VDPWR.n3083 63.3551
R8406 VDPWR.n564 VDPWR.t53 63.3219
R8407 VDPWR.n539 VDPWR.t417 63.3219
R8408 VDPWR.n284 VDPWR.t628 63.3219
R8409 VDPWR.n259 VDPWR.t104 63.3219
R8410 VDPWR.n2082 VDPWR.t455 63.3219
R8411 VDPWR.n2082 VDPWR.t439 63.3219
R8412 VDPWR.n1120 VDPWR.t820 63.3219
R8413 VDPWR.n991 VDPWR.t823 63.3219
R8414 VDPWR.n2894 VDPWR.t24 63.3219
R8415 VDPWR.n2894 VDPWR.t504 63.3219
R8416 VDPWR.n907 VDPWR.t575 63.3219
R8417 VDPWR.n907 VDPWR.t665 63.3219
R8418 VDPWR.n27 VDPWR.t648 63.3219
R8419 VDPWR.n2 VDPWR.t419 63.3219
R8420 VDPWR.n715 VDPWR.n714 62.2257
R8421 VDPWR.n526 VDPWR.n525 62.2257
R8422 VDPWR.n462 VDPWR.n461 62.2257
R8423 VDPWR.n3106 VDPWR.n3105 62.2257
R8424 VDPWR VDPWR.t226 62.103
R8425 VDPWR VDPWR.t238 62.103
R8426 VDPWR.t829 VDPWR 62.103
R8427 VDPWR VDPWR.t631 62.103
R8428 VDPWR.n710 VDPWR.n709 61.6672
R8429 VDPWR.n713 VDPWR.n712 61.6672
R8430 VDPWR.n695 VDPWR.n694 61.6672
R8431 VDPWR.n698 VDPWR.n697 61.6672
R8432 VDPWR.n679 VDPWR.n678 61.6672
R8433 VDPWR.n682 VDPWR.n681 61.6672
R8434 VDPWR.n659 VDPWR.n658 61.6672
R8435 VDPWR.n661 VDPWR.n660 61.6672
R8436 VDPWR.n521 VDPWR.n520 61.6672
R8437 VDPWR.n524 VDPWR.n523 61.6672
R8438 VDPWR.n506 VDPWR.n505 61.6672
R8439 VDPWR.n509 VDPWR.n508 61.6672
R8440 VDPWR.n490 VDPWR.n489 61.6672
R8441 VDPWR.n493 VDPWR.n492 61.6672
R8442 VDPWR.n473 VDPWR.n472 61.6672
R8443 VDPWR.n476 VDPWR.n475 61.6672
R8444 VDPWR.n409 VDPWR.n408 61.6672
R8445 VDPWR.n412 VDPWR.n411 61.6672
R8446 VDPWR.n380 VDPWR.n379 61.6672
R8447 VDPWR.n392 VDPWR.n391 61.6672
R8448 VDPWR.n452 VDPWR.n451 61.6672
R8449 VDPWR.n455 VDPWR.n454 61.6672
R8450 VDPWR.n436 VDPWR.n435 61.6672
R8451 VDPWR.n439 VDPWR.n438 61.6672
R8452 VDPWR.n416 VDPWR.n415 61.6672
R8453 VDPWR.n418 VDPWR.n417 61.6672
R8454 VDPWR.n765 VDPWR.n764 61.6672
R8455 VDPWR.n768 VDPWR.n767 61.6672
R8456 VDPWR.n3096 VDPWR.n3095 61.6672
R8457 VDPWR.n3099 VDPWR.n3098 61.6672
R8458 VDPWR.n3080 VDPWR.n3079 61.6672
R8459 VDPWR.n3083 VDPWR.n3082 61.6672
R8460 VDPWR.n3063 VDPWR.n3062 61.6672
R8461 VDPWR.n3066 VDPWR.n3065 61.6672
R8462 VDPWR.n667 VDPWR.n656 61.4728
R8463 VDPWR.n478 VDPWR.n477 61.4728
R8464 VDPWR.n424 VDPWR.n413 61.4728
R8465 VDPWR.n3068 VDPWR.n3067 61.4728
R8466 VDPWR.n533 VDPWR.n532 61.346
R8467 VDPWR.n3112 VDPWR.n3111 61.346
R8468 VDPWR.n382 VDPWR.n378 60.9564
R8469 VDPWR.n383 VDPWR.n380 60.9564
R8470 VDPWR.n394 VDPWR.n390 60.9564
R8471 VDPWR.n395 VDPWR.n392 60.9564
R8472 VDPWR.t635 VDPWR.t21 60.4245
R8473 VDPWR.t120 VDPWR.t99 58.7461
R8474 VDPWR VDPWR.t653 57.0676
R8475 VDPWR.t454 VDPWR.t735 57.0676
R8476 VDPWR.t295 VDPWR 57.0676
R8477 VDPWR.t900 VDPWR.t336 57.0676
R8478 VDPWR.t56 VDPWR 55.3892
R8479 VDPWR.t107 VDPWR 55.3892
R8480 VDPWR VDPWR.t799 55.3892
R8481 VDPWR.t457 VDPWR 55.3892
R8482 VDPWR VDPWR.t493 53.7107
R8483 VDPWR.t416 VDPWR 52.0323
R8484 VDPWR.t103 VDPWR 52.0323
R8485 VDPWR VDPWR.t67 52.0323
R8486 VDPWR VDPWR.t244 52.0323
R8487 VDPWR VDPWR.t86 52.0323
R8488 VDPWR VDPWR.t1141 52.0323
R8489 VDPWR.t8 VDPWR 52.0323
R8490 VDPWR.t668 VDPWR.t380 52.0323
R8491 VDPWR VDPWR.t201 52.0323
R8492 VDPWR VDPWR.t537 52.0323
R8493 VDPWR VDPWR.t410 52.0323
R8494 VDPWR VDPWR.t580 52.0323
R8495 VDPWR VDPWR.t574 52.0323
R8496 VDPWR.t128 VDPWR 52.0323
R8497 VDPWR.t452 VDPWR 52.0323
R8498 VDPWR.t161 VDPWR 52.0323
R8499 VDPWR.t83 VDPWR 52.0323
R8500 VDPWR VDPWR.t576 52.0323
R8501 VDPWR VDPWR.t249 52.0323
R8502 VDPWR VDPWR.t745 52.0323
R8503 VDPWR VDPWR.t639 52.0323
R8504 VDPWR VDPWR.t477 52.0323
R8505 VDPWR VDPWR.t442 52.0323
R8506 VDPWR.t418 VDPWR 52.0323
R8507 VDPWR.n2166 VDPWR.t1249 50.5057
R8508 VDPWR.t10 VDPWR.t370 50.3539
R8509 VDPWR VDPWR.t1092 50.3539
R8510 VDPWR.t27 VDPWR.t888 50.3539
R8511 VDPWR VDPWR.t692 50.3539
R8512 VDPWR.t1129 VDPWR 48.6754
R8513 VDPWR VDPWR.t1010 48.6754
R8514 VDPWR VDPWR.t967 48.6754
R8515 VDPWR VDPWR.t958 48.6754
R8516 VDPWR.t1042 VDPWR 48.6754
R8517 VDPWR VDPWR.t915 48.6754
R8518 VDPWR VDPWR.t1138 48.6754
R8519 VDPWR.n2167 VDPWR.n1967 46.0805
R8520 VDPWR VDPWR.t723 45.3185
R8521 VDPWR VDPWR.t567 45.3185
R8522 VDPWR.t299 VDPWR.t1035 45.3185
R8523 VDPWR.t770 VDPWR.t592 45.3185
R8524 VDPWR VDPWR.t65 45.3185
R8525 VDPWR VDPWR.t672 45.3185
R8526 VDPWR VDPWR.t697 45.3185
R8527 VDPWR VDPWR.t695 43.6401
R8528 VDPWR.t352 VDPWR 43.6401
R8529 VDPWR.n998 VDPWR.t765 42.3555
R8530 VDPWR.n2672 VDPWR.t622 42.3555
R8531 VDPWR.n2680 VDPWR.t673 42.3555
R8532 VDPWR VDPWR.t228 41.9616
R8533 VDPWR VDPWR.t774 41.9616
R8534 VDPWR.t639 VDPWR.t279 41.9616
R8535 VDPWR VDPWR.t145 41.9616
R8536 VDPWR.n1384 VDPWR.t245 41.5552
R8537 VDPWR.n1384 VDPWR.t524 41.5552
R8538 VDPWR.n2104 VDPWR.t87 41.5552
R8539 VDPWR.n2104 VDPWR.t286 41.5552
R8540 VDPWR.n1060 VDPWR.t538 41.5552
R8541 VDPWR.n1060 VDPWR.t236 41.5552
R8542 VDPWR.n1157 VDPWR.t562 41.5552
R8543 VDPWR.n1157 VDPWR.t59 41.5552
R8544 VDPWR.n904 VDPWR.t414 41.5552
R8545 VDPWR.n904 VDPWR.t542 41.5552
R8546 VDPWR.n908 VDPWR.t560 41.5552
R8547 VDPWR.n908 VDPWR.t644 41.5552
R8548 VDPWR.n939 VDPWR.t331 41.5552
R8549 VDPWR.n939 VDPWR.t571 41.5552
R8550 VDPWR.n2828 VDPWR.t241 41.5552
R8551 VDPWR.n2828 VDPWR.t540 41.5552
R8552 VDPWR.n2945 VDPWR.t509 41.5552
R8553 VDPWR.n2945 VDPWR.t89 41.5552
R8554 VDPWR.n2949 VDPWR.t1164 41.5552
R8555 VDPWR.n2949 VDPWR.t61 41.5552
R8556 VDPWR.t482 VDPWR.t43 40.7512
R8557 VDPWR.t715 VDPWR.t482 40.7512
R8558 VDPWR.t468 VDPWR.t715 40.7512
R8559 VDPWR.t484 VDPWR.t45 40.7512
R8560 VDPWR.t480 VDPWR.t484 40.7512
R8561 VDPWR.t47 VDPWR.t480 40.7512
R8562 VDPWR VDPWR.t388 40.2832
R8563 VDPWR.t569 VDPWR.t603 38.6047
R8564 VDPWR.n384 VDPWR.n383 38.5759
R8565 VDPWR.n382 VDPWR.n381 38.5759
R8566 VDPWR.n396 VDPWR.n395 38.5759
R8567 VDPWR.n394 VDPWR.n393 38.5759
R8568 VDPWR VDPWR.t235 36.9263
R8569 VDPWR.t234 VDPWR.t364 36.9263
R8570 VDPWR.t663 VDPWR.t157 36.9263
R8571 VDPWR.n2096 VDPWR.t12 36.4455
R8572 VDPWR.n1453 VDPWR.t68 36.1587
R8573 VDPWR.n1453 VDPWR.t204 36.1587
R8574 VDPWR.n985 VDPWR.t9 36.1587
R8575 VDPWR.n985 VDPWR.t599 36.1587
R8576 VDPWR.n1053 VDPWR.t202 36.1587
R8577 VDPWR.n1053 VDPWR.t269 36.1587
R8578 VDPWR.n819 VDPWR.t443 36.1587
R8579 VDPWR.n819 VDPWR.t261 36.1587
R8580 VDPWR.n795 VDPWR.t640 36.1587
R8581 VDPWR.n795 VDPWR.t330 36.1587
R8582 VDPWR.n2704 VDPWR.t746 36.1587
R8583 VDPWR.n2704 VDPWR.t22 36.1587
R8584 VDPWR.n2699 VDPWR.t250 36.1587
R8585 VDPWR.n2699 VDPWR.t259 36.1587
R8586 VDPWR.n2671 VDPWR.t84 36.1587
R8587 VDPWR.n2671 VDPWR.t761 36.1587
R8588 VDPWR.n2789 VDPWR.t162 36.1587
R8589 VDPWR.n2789 VDPWR.t167 36.1587
R8590 VDPWR.n2628 VDPWR.t169 36.1587
R8591 VDPWR.n2628 VDPWR.t376 36.1587
R8592 VDPWR.n2630 VDPWR.t129 36.1587
R8593 VDPWR.n2630 VDPWR.t353 36.1587
R8594 VDPWR.n2683 VDPWR.t667 36.1587
R8595 VDPWR.n2683 VDPWR.t221 36.1587
R8596 VDPWR.n849 VDPWR.t478 36.1587
R8597 VDPWR.n849 VDPWR.t1161 36.1587
R8598 VDPWR.n1402 VDPWR.t372 35.4605
R8599 VDPWR.n2032 VDPWR.t368 35.4605
R8600 VDPWR.n1084 VDPWR.t780 35.4605
R8601 VDPWR.n1140 VDPWR.t70 35.4605
R8602 VDPWR.n919 VDPWR.t573 35.4605
R8603 VDPWR.n922 VDPWR.t349 35.4605
R8604 VDPWR.n944 VDPWR.t271 35.4605
R8605 VDPWR.n943 VDPWR.t456 35.4605
R8606 VDPWR.n2942 VDPWR.t276 35.4605
R8607 VDPWR.n876 VDPWR.t98 35.4605
R8608 VDPWR.t727 VDPWR.t149 35.2479
R8609 VDPWR.n2084 VDPWR.n2035 34.6358
R8610 VDPWR.n2764 VDPWR.n2763 34.6358
R8611 VDPWR.n2711 VDPWR.n2705 34.6358
R8612 VDPWR.n3019 VDPWR.n796 34.6358
R8613 VDPWR.n1764 VDPWR.n1763 34.6358
R8614 VDPWR.n1763 VDPWR.n1762 34.6358
R8615 VDPWR.n1755 VDPWR.n1413 34.6358
R8616 VDPWR.n1751 VDPWR.n1413 34.6358
R8617 VDPWR.n2084 VDPWR.n2083 34.6358
R8618 VDPWR.n2095 VDPWR.n2020 34.6358
R8619 VDPWR.n1087 VDPWR.n1083 34.6358
R8620 VDPWR.n1091 VDPWR.n1034 34.6358
R8621 VDPWR.n1101 VDPWR.n1100 34.6358
R8622 VDPWR.n2891 VDPWR.n901 34.6358
R8623 VDPWR.n2858 VDPWR.n923 34.6358
R8624 VDPWR.n2862 VDPWR.n2861 34.6358
R8625 VDPWR.n2862 VDPWR.n920 34.6358
R8626 VDPWR.n2866 VDPWR.n920 34.6358
R8627 VDPWR.n2854 VDPWR.n2851 34.6358
R8628 VDPWR.n2606 VDPWR.n2605 34.6358
R8629 VDPWR.n2811 VDPWR.n945 34.6358
R8630 VDPWR.n2815 VDPWR.n945 34.6358
R8631 VDPWR.n2816 VDPWR.n2815 34.6358
R8632 VDPWR.n2818 VDPWR.n941 34.6358
R8633 VDPWR.n2822 VDPWR.n941 34.6358
R8634 VDPWR.n2823 VDPWR.n2822 34.6358
R8635 VDPWR.n2927 VDPWR.n2926 34.6358
R8636 VDPWR.n2999 VDPWR.n2941 34.6358
R8637 VDPWR.n2999 VDPWR.n2998 34.6358
R8638 VDPWR.n2645 VDPWR.n2629 34.6358
R8639 VDPWR.n2745 VDPWR.n2684 34.6358
R8640 VDPWR.n808 VDPWR.n804 34.6358
R8641 VDPWR.n897 VDPWR.t32 34.4755
R8642 VDPWR.n2655 VDPWR.t595 34.4755
R8643 VDPWR.n2547 VDPWR.n2546 33.6462
R8644 VDPWR.n1015 VDPWR.n1014 33.6462
R8645 VDPWR.n2534 VDPWR.n2533 33.6462
R8646 VDPWR VDPWR.t475 33.5694
R8647 VDPWR.t749 VDPWR 33.5694
R8648 VDPWR.n1092 VDPWR.t411 33.4905
R8649 VDPWR.n897 VDPWR.t696 33.4905
R8650 VDPWR.n2655 VDPWR.t453 33.4905
R8651 VDPWR.n809 VDPWR.t680 33.4905
R8652 VDPWR.n1042 VDPWR.t601 32.7439
R8653 VDPWR.n387 VDPWR.n386 32.5881
R8654 VDPWR.n399 VDPWR.n398 32.5881
R8655 VDPWR.n898 VDPWR.t728 32.5055
R8656 VDPWR.n898 VDPWR.t502 32.5055
R8657 VDPWR.n2787 VDPWR.t26 32.5055
R8658 VDPWR.n2787 VDPWR.t154 32.5055
R8659 VDPWR.n2098 VDPWR.n2018 32.377
R8660 VDPWR.n1083 VDPWR.n1036 32.2581
R8661 VDPWR.n2103 VDPWR.n2102 32.0005
R8662 VDPWR.t404 VDPWR 31.891
R8663 VDPWR.n751 VDPWR.t175 31.6605
R8664 VDPWR.n2853 VDPWR.n923 31.624
R8665 VDPWR.n2809 VDPWR.n949 31.624
R8666 VDPWR.n2930 VDPWR.n880 31.624
R8667 VDPWR.n2933 VDPWR.n877 31.624
R8668 VDPWR.n143 VDPWR.n140 30.8711
R8669 VDPWR.n1757 VDPWR.n1756 30.8711
R8670 VDPWR.n1099 VDPWR.n1098 30.8711
R8671 VDPWR.n1048 VDPWR.n1047 30.7205
R8672 VDPWR.n2042 VDPWR.t211 30.5355
R8673 VDPWR.n1759 VDPWR.n1758 30.4946
R8674 VDPWR.n2810 VDPWR.n2809 30.4946
R8675 VDPWR.n2931 VDPWR.n2930 30.4946
R8676 VDPWR.n2938 VDPWR.n877 30.4946
R8677 VDPWR.t371 VDPWR 30.2125
R8678 VDPWR VDPWR.t1083 30.2125
R8679 VDPWR.t396 VDPWR.t6 30.2125
R8680 VDPWR.t764 VDPWR.t394 30.2125
R8681 VDPWR.t501 VDPWR.t23 30.2125
R8682 VDPWR.t195 VDPWR.t114 30.2125
R8683 VDPWR.n2673 VDPWR.n2663 29.3652
R8684 VDPWR.n2550 VDPWR.n995 29.2576
R8685 VDPWR.n1108 VDPWR.n1104 29.1064
R8686 VDPWR.n722 VDPWR.t44 28.6596
R8687 VDPWR.n724 VDPWR.t48 28.6583
R8688 VDPWR.n641 VDPWR 28.5341
R8689 VDPWR.n361 VDPWR 28.5341
R8690 VDPWR.n2847 VDPWR 28.5341
R8691 VDPWR.t193 VDPWR.t97 28.5341
R8692 VDPWR.t762 VDPWR 28.5341
R8693 VDPWR.n104 VDPWR 28.5341
R8694 VDPWR.n894 VDPWR.t256 28.4453
R8695 VDPWR.n569 VDPWR.t36 28.4453
R8696 VDPWR.n550 VDPWR.t516 28.4453
R8697 VDPWR.n289 VDPWR.t624 28.4453
R8698 VDPWR.n270 VDPWR.t119 28.4453
R8699 VDPWR.n791 VDPWR.t690 28.4453
R8700 VDPWR.n32 VDPWR.t144 28.4453
R8701 VDPWR.n13 VDPWR.t451 28.4453
R8702 VDPWR.n2703 VDPWR.t763 28.4433
R8703 VDPWR.n2096 VDPWR.t688 27.5805
R8704 VDPWR.n2042 VDPWR.t437 27.5805
R8705 VDPWR.n1186 VDPWR.t296 27.5805
R8706 VDPWR.n2293 VDPWR.t63 27.5805
R8707 VDPWR.n2293 VDPWR.t476 27.5805
R8708 VDPWR.n2328 VDPWR.t796 27.5805
R8709 VDPWR.n2328 VDPWR.t806 27.5805
R8710 VDPWR.n1225 VDPWR.t788 27.5805
R8711 VDPWR.n2310 VDPWR.t794 27.5805
R8712 VDPWR.n2310 VDPWR.t816 27.5805
R8713 VDPWR.n1239 VDPWR.t818 27.5805
R8714 VDPWR.n1239 VDPWR.t790 27.5805
R8715 VDPWR.n1240 VDPWR.t804 27.5805
R8716 VDPWR.n1240 VDPWR.t814 27.5805
R8717 VDPWR.n1243 VDPWR.t474 27.5805
R8718 VDPWR.n1243 VDPWR.t810 27.5805
R8719 VDPWR.n1219 VDPWR.t798 27.5805
R8720 VDPWR.n1219 VDPWR.t808 27.5805
R8721 VDPWR.n1222 VDPWR.t800 27.5805
R8722 VDPWR.n1222 VDPWR.t802 27.5805
R8723 VDPWR.n1202 VDPWR.t500 27.5805
R8724 VDPWR.n1202 VDPWR.t498 27.5805
R8725 VDPWR.n2390 VDPWR.t302 27.5805
R8726 VDPWR.n2390 VDPWR.t306 27.5805
R8727 VDPWR.n1196 VDPWR.t308 27.5805
R8728 VDPWR.n1196 VDPWR.t298 27.5805
R8729 VDPWR.n1199 VDPWR.t300 27.5805
R8730 VDPWR.n1199 VDPWR.t304 27.5805
R8731 VDPWR.n2376 VDPWR.t492 27.5805
R8732 VDPWR.n2376 VDPWR.t294 27.5805
R8733 VDPWR.n1180 VDPWR.t288 27.5805
R8734 VDPWR.n1180 VDPWR.t310 27.5805
R8735 VDPWR.n2415 VDPWR.t292 27.5805
R8736 VDPWR.n2415 VDPWR.t316 27.5805
R8737 VDPWR.n1183 VDPWR.t318 27.5805
R8738 VDPWR.n1183 VDPWR.t290 27.5805
R8739 VDPWR.n1054 VDPWR.t740 27.5805
R8740 VDPWR.n1054 VDPWR.t744 27.5805
R8741 VDPWR.n1046 VDPWR.t387 27.5805
R8742 VDPWR.n1046 VDPWR.t496 27.5805
R8743 VDPWR.n990 VDPWR.t391 27.5805
R8744 VDPWR.n990 VDPWR.t393 27.5805
R8745 VDPWR.n993 VDPWR.t409 27.5805
R8746 VDPWR.n993 VDPWR.t401 27.5805
R8747 VDPWR.n994 VDPWR.t405 27.5805
R8748 VDPWR.n994 VDPWR.t395 27.5805
R8749 VDPWR.n999 VDPWR.t403 27.5805
R8750 VDPWR.n1000 VDPWR.t407 27.5805
R8751 VDPWR.n1000 VDPWR.t381 27.5805
R8752 VDPWR.n1009 VDPWR.t379 27.5805
R8753 VDPWR.n1009 VDPWR.t389 27.5805
R8754 VDPWR.n1019 VDPWR.t383 27.5805
R8755 VDPWR.n1019 VDPWR.t385 27.5805
R8756 VDPWR.n1068 VDPWR.n1065 27.4829
R8757 VDPWR.n1093 VDPWR.n1091 27.4829
R8758 VDPWR.n2895 VDPWR.n2893 27.4829
R8759 VDPWR.n2824 VDPWR.n2823 27.4829
R8760 VDPWR.n2995 VDPWR.n2994 27.4829
R8761 VDPWR.n1659 VDPWR.n1658 27.0566
R8762 VDPWR.n2529 VDPWR.n1133 27.0566
R8763 VDPWR.n2031 VDPWR.t74 26.9729
R8764 VDPWR.n900 VDPWR.t158 26.9729
R8765 VDPWR.n903 VDPWR.t66 26.9729
R8766 VDPWR.t86 VDPWR.t505 26.8556
R8767 VDPWR.n1764 VDPWR.n1408 26.7859
R8768 VDPWR.n644 VDPWR.n643 26.7299
R8769 VDPWR.n364 VDPWR.n363 26.7299
R8770 VDPWR.n107 VDPWR.n106 26.7299
R8771 VDPWR.n2851 VDPWR.n2850 26.7299
R8772 VDPWR.n139 VDPWR.t652 26.5955
R8773 VDPWR.n139 VDPWR.t254 26.5955
R8774 VDPWR.n1411 VDPWR.t441 26.5955
R8775 VDPWR.n1411 VDPWR.t445 26.5955
R8776 VDPWR.n1412 VDPWR.t608 26.5955
R8777 VDPWR.n1412 VDPWR.t1 26.5955
R8778 VDPWR.n2036 VDPWR.t182 26.5955
R8779 VDPWR.n2036 VDPWR.t184 26.5955
R8780 VDPWR.n1186 VDPWR.t312 26.5955
R8781 VDPWR.n1225 VDPWR.t792 26.5955
R8782 VDPWR.n1031 VDPWR.t604 26.5955
R8783 VDPWR.n1031 VDPWR.t223 26.5955
R8784 VDPWR.n999 VDPWR.t399 26.5955
R8785 VDPWR.n1135 VDPWR.t91 26.5955
R8786 VDPWR.n1135 VDPWR.t566 26.5955
R8787 VDPWR.n2852 VDPWR.t190 26.5955
R8788 VDPWR.n2852 VDPWR.t786 26.5955
R8789 VDPWR.n948 VDPWR.t827 26.5955
R8790 VDPWR.n948 VDPWR.t366 26.5955
R8791 VDPWR.n947 VDPWR.t125 26.5955
R8792 VDPWR.n947 VDPWR.t333 26.5955
R8793 VDPWR.n928 VDPWR.t337 26.5955
R8794 VDPWR.n928 VDPWR.t142 26.5955
R8795 VDPWR.n883 VDPWR.t449 26.5955
R8796 VDPWR.n883 VDPWR.t730 26.5955
R8797 VDPWR.n879 VDPWR.t113 26.5955
R8798 VDPWR.n879 VDPWR.t320 26.5955
R8799 VDPWR.n2932 VDPWR.t196 26.5955
R8800 VDPWR.n2932 VDPWR.t278 26.5955
R8801 VDPWR.n2625 VDPWR.t377 26.5955
R8802 VDPWR.n2625 VDPWR.t374 26.5955
R8803 VDPWR.n853 VDPWR.n816 26.3341
R8804 VDPWR.n144 VDPWR.n143 25.977
R8805 VDPWR.n643 VDPWR.n642 25.6953
R8806 VDPWR.n363 VDPWR.n362 25.6953
R8807 VDPWR.n106 VDPWR.n105 25.6953
R8808 VDPWR.n609 VDPWR.n593 25.224
R8809 VDPWR.n605 VDPWR.n593 25.224
R8810 VDPWR.n614 VDPWR.n592 25.224
R8811 VDPWR.n610 VDPWR.n592 25.224
R8812 VDPWR.n616 VDPWR.n590 25.224
R8813 VDPWR.n616 VDPWR.n615 25.224
R8814 VDPWR.n634 VDPWR.n630 25.224
R8815 VDPWR.n329 VDPWR.n313 25.224
R8816 VDPWR.n325 VDPWR.n313 25.224
R8817 VDPWR.n334 VDPWR.n312 25.224
R8818 VDPWR.n330 VDPWR.n312 25.224
R8819 VDPWR.n336 VDPWR.n310 25.224
R8820 VDPWR.n336 VDPWR.n335 25.224
R8821 VDPWR.n354 VDPWR.n350 25.224
R8822 VDPWR.n247 VDPWR.n120 25.224
R8823 VDPWR.n247 VDPWR.n246 25.224
R8824 VDPWR.n245 VDPWR.n244 25.224
R8825 VDPWR.n244 VDPWR.n123 25.224
R8826 VDPWR.n240 VDPWR.n239 25.224
R8827 VDPWR.n239 VDPWR.n124 25.224
R8828 VDPWR.n235 VDPWR.n234 25.224
R8829 VDPWR.n234 VDPWR.n125 25.224
R8830 VDPWR.n230 VDPWR.n229 25.224
R8831 VDPWR.n229 VDPWR.n126 25.224
R8832 VDPWR.n225 VDPWR.n224 25.224
R8833 VDPWR.n224 VDPWR.n204 25.224
R8834 VDPWR.n220 VDPWR.n219 25.224
R8835 VDPWR.n219 VDPWR.n205 25.224
R8836 VDPWR.n215 VDPWR.n214 25.224
R8837 VDPWR.n214 VDPWR.n206 25.224
R8838 VDPWR.n210 VDPWR.n209 25.224
R8839 VDPWR.n209 VDPWR.n119 25.224
R8840 VDPWR.n183 VDPWR.n133 25.224
R8841 VDPWR.n179 VDPWR.n133 25.224
R8842 VDPWR.n188 VDPWR.n132 25.224
R8843 VDPWR.n184 VDPWR.n132 25.224
R8844 VDPWR.n193 VDPWR.n131 25.224
R8845 VDPWR.n189 VDPWR.n131 25.224
R8846 VDPWR.n198 VDPWR.n130 25.224
R8847 VDPWR.n194 VDPWR.n130 25.224
R8848 VDPWR.n200 VDPWR.n129 25.224
R8849 VDPWR.n200 VDPWR.n199 25.224
R8850 VDPWR.n159 VDPWR.n154 25.224
R8851 VDPWR.n155 VDPWR.n154 25.224
R8852 VDPWR.n164 VDPWR.n153 25.224
R8853 VDPWR.n160 VDPWR.n153 25.224
R8854 VDPWR.n169 VDPWR.n152 25.224
R8855 VDPWR.n165 VDPWR.n152 25.224
R8856 VDPWR.n171 VDPWR.n135 25.224
R8857 VDPWR.n171 VDPWR.n170 25.224
R8858 VDPWR.n72 VDPWR.n56 25.224
R8859 VDPWR.n68 VDPWR.n56 25.224
R8860 VDPWR.n77 VDPWR.n55 25.224
R8861 VDPWR.n73 VDPWR.n55 25.224
R8862 VDPWR.n79 VDPWR.n53 25.224
R8863 VDPWR.n79 VDPWR.n78 25.224
R8864 VDPWR.n97 VDPWR.n93 25.224
R8865 VDPWR.n2899 VDPWR.n895 25.1912
R8866 VDPWR.n2774 VDPWR.n2663 25.1912
R8867 VDPWR.n2786 VDPWR.n2658 25.1912
R8868 VDPWR.n3020 VDPWR.n3019 25.1912
R8869 VDPWR.t237 VDPWR 25.1772
R8870 VDPWR VDPWR.t721 25.1772
R8871 VDPWR.t825 VDPWR 25.1772
R8872 VDPWR.n724 VDPWR.n723 25.0224
R8873 VDPWR.n726 VDPWR.n725 25.0224
R8874 VDPWR.n722 VDPWR.n721 25.0224
R8875 VDPWR.n2647 VDPWR.n2622 24.0841
R8876 VDPWR.n1248 VDPWR.n1247 24.0557
R8877 VDPWR.n2849 VDPWR.n929 23.7181
R8878 VDPWR.n580 VDPWR.n563 23.7181
R8879 VDPWR.n639 VDPWR.n561 23.7181
R8880 VDPWR.n300 VDPWR.n283 23.7181
R8881 VDPWR.n359 VDPWR.n281 23.7181
R8882 VDPWR.n1658 VDPWR.n1459 23.7181
R8883 VDPWR.n1751 VDPWR.n1750 23.7181
R8884 VDPWR.n971 VDPWR.n968 23.7181
R8885 VDPWR.n977 VDPWR.n971 23.7181
R8886 VDPWR.n2530 VDPWR.n2529 23.7181
R8887 VDPWR.n2895 VDPWR.n895 23.7181
R8888 VDPWR.n2885 VDPWR.n2884 23.7181
R8889 VDPWR.n2605 VDPWR.n2594 23.7181
R8890 VDPWR.n2830 VDPWR.n929 23.7181
R8891 VDPWR.n2763 VDPWR.n2675 23.7181
R8892 VDPWR.n2640 VDPWR.n2637 23.7181
R8893 VDPWR.n3037 VDPWR.n3036 23.7181
R8894 VDPWR.n43 VDPWR.n26 23.7181
R8895 VDPWR.n102 VDPWR.n24 23.7181
R8896 VDPWR.t309 VDPWR.t994 23.4987
R8897 VDPWR.t674 VDPWR.t319 23.4987
R8898 VDPWR.t25 VDPWR.t166 23.4987
R8899 VDPWR.n804 VDPWR.n803 22.9652
R8900 VDPWR.n2105 VDPWR.n2103 22.9652
R8901 VDPWR.n2886 VDPWR.n2885 22.9652
R8902 VDPWR.n2869 VDPWR.n909 22.9652
R8903 VDPWR.n2829 VDPWR.n938 22.9652
R8904 VDPWR.n2993 VDPWR.n2946 22.9652
R8905 VDPWR.n1048 VDPWR.n1020 22.6748
R8906 VDPWR.n1059 VDPWR.n1044 22.5887
R8907 VDPWR.n2887 VDPWR.n901 22.5887
R8908 VDPWR.n2892 VDPWR.n2891 22.5887
R8909 VDPWR.n2556 VDPWR.n2555 22.3091
R8910 VDPWR.n2097 VDPWR.n2095 22.2123
R8911 VDPWR.n2098 VDPWR.n2097 22.2123
R8912 VDPWR.n1055 VDPWR.n1052 22.2123
R8913 VDPWR.n1055 VDPWR.n1044 22.2123
R8914 VDPWR.n2647 VDPWR.n2646 22.2123
R8915 VDPWR.n2641 VDPWR.n2629 22.2123
R8916 VDPWR.n2646 VDPWR.n2645 22.2123
R8917 VDPWR.n2641 VDPWR.n2640 22.2123
R8918 VDPWR.n2746 VDPWR.n2745 22.2123
R8919 VDPWR.n2869 VDPWR.n2868 21.8358
R8920 VDPWR.n2824 VDPWR.n938 21.8358
R8921 VDPWR.n2994 VDPWR.n2993 21.8358
R8922 VDPWR.t33 VDPWR.t402 21.8203
R8923 VDPWR.t488 VDPWR.t406 21.8203
R8924 VDPWR.n2532 VDPWR.t382 21.8203
R8925 VDPWR.t446 VDPWR.t165 21.8203
R8926 VDPWR.n629 VDPWR.n563 21.4593
R8927 VDPWR.n349 VDPWR.n283 21.4593
R8928 VDPWR.n2884 VDPWR.n909 21.4593
R8929 VDPWR.n2830 VDPWR.n2829 21.4593
R8930 VDPWR.n92 VDPWR.n26 21.4593
R8931 VDPWR.n2565 VDPWR.n2564 21.05
R8932 VDPWR.n2221 VDPWR.n2206 20.912
R8933 VDPWR.n2555 VDPWR.n2554 20.8462
R8934 VDPWR.n854 VDPWR.n853 20.4852
R8935 VDPWR.n2557 VDPWR.n2556 20.4805
R8936 VDPWR.n734 VDPWR.t468 20.3758
R8937 VDPWR.t45 VDPWR.n734 20.3758
R8938 VDPWR.n610 VDPWR.n609 20.3299
R8939 VDPWR.n615 VDPWR.n614 20.3299
R8940 VDPWR.n330 VDPWR.n329 20.3299
R8941 VDPWR.n335 VDPWR.n334 20.3299
R8942 VDPWR.n246 VDPWR.n245 20.3299
R8943 VDPWR.n240 VDPWR.n123 20.3299
R8944 VDPWR.n235 VDPWR.n124 20.3299
R8945 VDPWR.n230 VDPWR.n125 20.3299
R8946 VDPWR.n225 VDPWR.n126 20.3299
R8947 VDPWR.n220 VDPWR.n204 20.3299
R8948 VDPWR.n215 VDPWR.n205 20.3299
R8949 VDPWR.n210 VDPWR.n206 20.3299
R8950 VDPWR.n184 VDPWR.n183 20.3299
R8951 VDPWR.n189 VDPWR.n188 20.3299
R8952 VDPWR.n194 VDPWR.n193 20.3299
R8953 VDPWR.n199 VDPWR.n198 20.3299
R8954 VDPWR.n155 VDPWR.n129 20.3299
R8955 VDPWR.n160 VDPWR.n159 20.3299
R8956 VDPWR.n165 VDPWR.n164 20.3299
R8957 VDPWR.n170 VDPWR.n169 20.3299
R8958 VDPWR.n73 VDPWR.n72 20.3299
R8959 VDPWR.n78 VDPWR.n77 20.3299
R8960 VDPWR.t105 VDPWR.t531 20.1418
R8961 VDPWR.t685 VDPWR.t133 20.1418
R8962 VDPWR.t392 VDPWR.t677 20.1418
R8963 VDPWR.t664 VDPWR.t413 20.1418
R8964 VDPWR.t39 VDPWR.t588 20.1418
R8965 VDPWR.n2554 VDPWR.n995 20.1148
R8966 VDPWR.n2169 VDPWR.n1967 20.0749
R8967 VDPWR.n2705 VDPWR.n785 19.9534
R8968 VDPWR.n975 VDPWR.n974 19.9237
R8969 VDPWR.n649 VDPWR.n648 19.8181
R8970 VDPWR.n369 VDPWR.n368 19.8181
R8971 VDPWR.n112 VDPWR.n111 19.8181
R8972 VDPWR.n2549 VDPWR.n2548 19.7491
R8973 VDPWR.n2546 VDPWR.n1001 19.7491
R8974 VDPWR.n645 VDPWR.n644 19.6946
R8975 VDPWR.n365 VDPWR.n364 19.6946
R8976 VDPWR.n108 VDPWR.n107 19.6946
R8977 VDPWR.n2081 VDPWR.n2037 19.577
R8978 VDPWR.n2370 VDPWR.n2368 19.2067
R8979 VDPWR.n2334 VDPWR.n2333 18.7808
R8980 VDPWR.n1380 VDPWR.n1378 18.7591
R8981 VDPWR.t821 VDPWR.t222 18.4634
R8982 VDPWR.t643 VDPWR.t829 18.4634
R8983 VDPWR.n2033 VDPWR.n2020 18.4476
R8984 VDPWR.n1087 VDPWR.n1086 18.4476
R8985 VDPWR.n2861 VDPWR.n2860 18.4476
R8986 VDPWR.n2818 VDPWR.n2817 18.4476
R8987 VDPWR.n2941 VDPWR.n2940 18.4476
R8988 VDPWR.n2995 VDPWR.n2943 18.4476
R8989 VDPWR.n1052 VDPWR.n1045 18.0711
R8990 VDPWR.n2794 VDPWR.n2656 18.0382
R8991 VDPWR.n1694 VDPWR.n1693 17.9678
R8992 VDPWR.n2299 VDPWR.n1244 17.612
R8993 VDPWR.n621 VDPWR.n590 17.3181
R8994 VDPWR.n633 VDPWR.n632 17.3181
R8995 VDPWR.n639 VDPWR.n538 17.3181
R8996 VDPWR.n341 VDPWR.n310 17.3181
R8997 VDPWR.n353 VDPWR.n352 17.3181
R8998 VDPWR.n359 VDPWR.n258 17.3181
R8999 VDPWR.n251 VDPWR.n119 17.3181
R9000 VDPWR.n175 VDPWR.n135 17.3181
R9001 VDPWR.n84 VDPWR.n53 17.3181
R9002 VDPWR.n96 VDPWR.n95 17.3181
R9003 VDPWR.n102 VDPWR.n1 17.3181
R9004 VDPWR.n605 VDPWR.n604 17.2853
R9005 VDPWR.n325 VDPWR.n324 17.2853
R9006 VDPWR.n68 VDPWR.n67 17.2853
R9007 VDPWR.n2925 VDPWR.n2924 16.9417
R9008 VDPWR.n2788 VDPWR.n2786 16.9417
R9009 VDPWR.t408 VDPWR.t521 16.785
R9010 VDPWR.t843 VDPWR.t431 16.785
R9011 VDPWR.t885 VDPWR.t670 16.785
R9012 VDPWR.n1787 VDPWR.n1378 16.7729
R9013 VDPWR.n2288 VDPWR.n1249 16.7729
R9014 VDPWR.n1624 VDPWR.n1623 16.6847
R9015 VDPWR.n2500 VDPWR.n1156 16.5825
R9016 VDPWR.n630 VDPWR.n629 16.5652
R9017 VDPWR.n634 VDPWR.n633 16.5652
R9018 VDPWR.n350 VDPWR.n349 16.5652
R9019 VDPWR.n354 VDPWR.n353 16.5652
R9020 VDPWR.n93 VDPWR.n92 16.5652
R9021 VDPWR.n97 VDPWR.n96 16.5652
R9022 VDPWR.n1017 VDPWR.n1016 16.4576
R9023 VDPWR.n2867 VDPWR.n2866 16.1887
R9024 VDPWR.n2817 VDPWR.n2816 16.1887
R9025 VDPWR.n2940 VDPWR.n2939 16.1887
R9026 VDPWR.n2998 VDPWR.n2943 16.1887
R9027 VDPWR.n250 VDPWR.n120 15.8123
R9028 VDPWR.n179 VDPWR.n178 15.8123
R9029 VDPWR.n731 VDPWR.n729 15.4172
R9030 VDPWR.n734 VDPWR.n731 15.4172
R9031 VDPWR.n730 VDPWR.n728 15.4172
R9032 VDPWR.n734 VDPWR.n730 15.4172
R9033 VDPWR.n1016 VDPWR.n1015 15.3605
R9034 VDPWR.n1248 VDPWR.n1246 15.2281
R9035 VDPWR.n1381 VDPWR.n1380 15.101
R9036 VDPWR.n1094 VDPWR.n1032 15.0593
R9037 VDPWR.n2811 VDPWR.n2810 15.0593
R9038 VDPWR.n2934 VDPWR.n2931 15.0593
R9039 VDPWR.n2939 VDPWR.n2938 15.0593
R9040 VDPWR.n2790 VDPWR.n2788 15.0593
R9041 VDPWR.n2747 VDPWR.n2746 15.0593
R9042 VDPWR.n1593 VDPWR.n1592 14.9
R9043 VDPWR.n3037 VDPWR.n785 14.6829
R9044 VDPWR.n2109 VDPWR.n2016 14.6484
R9045 VDPWR.n643 VDPWR.n559 14.6078
R9046 VDPWR.n363 VDPWR.n279 14.6078
R9047 VDPWR.n106 VDPWR.n22 14.6078
R9048 VDPWR.n1645 VDPWR.n1459 14.5851
R9049 VDPWR.n1724 VDPWR.n1437 14.5851
R9050 VDPWR.n1086 VDPWR.n1085 14.3064
R9051 VDPWR.n2887 VDPWR.n2886 14.3064
R9052 VDPWR.n2989 VDPWR.n2946 14.3064
R9053 VDPWR.n622 VDPWR.n621 14.2735
R9054 VDPWR.n581 VDPWR.n580 14.2735
R9055 VDPWR.n342 VDPWR.n341 14.2735
R9056 VDPWR.n301 VDPWR.n300 14.2735
R9057 VDPWR.n2063 VDPWR.n2051 14.2735
R9058 VDPWR.n2530 VDPWR.n1021 14.2735
R9059 VDPWR.n2903 VDPWR.n882 14.2735
R9060 VDPWR.n2970 VDPWR.n2958 14.2735
R9061 VDPWR.n2759 VDPWR.n2675 14.2735
R9062 VDPWR.n3036 VDPWR.n3035 14.2735
R9063 VDPWR.n837 VDPWR.n825 14.2735
R9064 VDPWR.n85 VDPWR.n84 14.2735
R9065 VDPWR.n44 VDPWR.n43 14.2735
R9066 VDPWR.n2034 VDPWR.n2033 13.9299
R9067 VDPWR.n2446 VDPWR.n1173 13.8955
R9068 VDPWR.n2474 VDPWR.n2462 13.8955
R9069 VDPWR.n650 VDPWR.n649 13.5534
R9070 VDPWR.n370 VDPWR.n369 13.5534
R9071 VDPWR.n113 VDPWR.n112 13.5534
R9072 VDPWR VDPWR.n570 13.4732
R9073 VDPWR VDPWR.n290 13.4732
R9074 VDPWR VDPWR.n33 13.4732
R9075 VDPWR.t235 VDPWR.t600 13.4281
R9076 VDPWR.t95 VDPWR.t906 13.4281
R9077 VDPWR.t31 VDPWR.t503 13.4281
R9078 VDPWR.t594 VDPWR.t161 13.4281
R9079 VDPWR VDPWR.t717 13.4281
R9080 VDPWR.n2564 VDPWR.n2563 12.9181
R9081 VDPWR.n175 VDPWR.n136 12.8005
R9082 VDPWR.n148 VDPWR.n136 12.8005
R9083 VDPWR.n148 VDPWR.n145 12.8005
R9084 VDPWR.n145 VDPWR.n144 12.8005
R9085 VDPWR.n1524 VDPWR.n1515 12.8005
R9086 VDPWR.n1299 VDPWR.n1290 12.8005
R9087 VDPWR.n1750 VDPWR.n1749 12.8005
R9088 VDPWR.n1921 VDPWR.n1920 12.8005
R9089 VDPWR.n2217 VDPWR.n2210 12.8005
R9090 VDPWR.n2601 VDPWR.n2594 12.8005
R9091 VDPWR.n2924 VDPWR.n882 12.8005
R9092 VDPWR.n1068 VDPWR.n1067 12.3976
R9093 VDPWR.n2989 VDPWR.n2988 12.3912
R9094 VDPWR.n650 VDPWR.n538 12.0476
R9095 VDPWR.n370 VDPWR.n258 12.0476
R9096 VDPWR.n113 VDPWR.n1 12.0476
R9097 VDPWR.t201 VDPWR.t739 11.7496
R9098 VDPWR.t545 VDPWR.t681 11.7496
R9099 VDPWR.n810 VDPWR.n808 11.6993
R9100 VDPWR.n803 VDPWR.n796 11.6711
R9101 VDPWR.n586 VDPWR.n585 11.4366
R9102 VDPWR.n306 VDPWR.n305 11.4366
R9103 VDPWR.n49 VDPWR.n48 11.4366
R9104 VDPWR VDPWR.n534 11.4331
R9105 VDPWR VDPWR.n3113 11.4331
R9106 VDPWR.n388 VDPWR.n387 11.3235
R9107 VDPWR.n400 VDPWR.n399 11.3235
R9108 VDPWR.n1061 VDPWR.n1059 11.2946
R9109 VDPWR.n2868 VDPWR.n2867 11.2946
R9110 VDPWR.n642 VDPWR.n560 11.2937
R9111 VDPWR.n362 VDPWR.n280 11.2937
R9112 VDPWR.n105 VDPWR.n23 11.2937
R9113 VDPWR.n627 VDPWR.n626 11.2737
R9114 VDPWR.n347 VDPWR.n346 11.2737
R9115 VDPWR.n90 VDPWR.n89 11.2737
R9116 VDPWR.n2533 VDPWR.n1020 10.9719
R9117 VDPWR.n141 VDPWR.n140 10.9345
R9118 VDPWR.n1094 VDPWR.n1093 10.9181
R9119 VDPWR.n2168 VDPWR.n2167 10.912
R9120 VDPWR.n977 VDPWR.n976 10.5744
R9121 VDPWR.n2790 VDPWR.n2656 10.5417
R9122 VDPWR.n559 VDPWR.n558 10.1786
R9123 VDPWR.n279 VDPWR.n278 10.1786
R9124 VDPWR.n22 VDPWR.n21 10.1786
R9125 VDPWR.n1065 VDPWR.n1043 10.1652
R9126 VDPWR.t228 VDPWR.t52 10.0712
R9127 VDPWR.t774 VDPWR.t627 10.0712
R9128 VDPWR.t1010 VDPWR.t479 10.0712
R9129 VDPWR.t145 VDPWR.t647 10.0712
R9130 VDPWR.n2222 VDPWR.n2221 9.8812
R9131 VDPWR.n1061 VDPWR.n1043 9.78874
R9132 VDPWR.n2893 VDPWR.n2892 9.78874
R9133 VDPWR.n1683 VDPWR.n1682 9.73273
R9134 VDPWR.n1846 VDPWR.n1331 9.73273
R9135 VDPWR.n1780 VDPWR.n1385 9.73273
R9136 VDPWR.n1776 VDPWR.n1775 9.73273
R9137 VDPWR.n1775 VDPWR.n1774 9.73273
R9138 VDPWR.n1774 VDPWR.n1388 9.73273
R9139 VDPWR.n1404 VDPWR.n1388 9.73273
R9140 VDPWR.n2286 VDPWR.n1251 9.73273
R9141 VDPWR.n2344 VDPWR.n1217 9.73273
R9142 VDPWR.n2379 VDPWR.n2375 9.73273
R9143 VDPWR.n2525 VDPWR.n2524 9.73273
R9144 VDPWR.n2519 VDPWR.n2518 9.73273
R9145 VDPWR.n2518 VDPWR.n2517 9.73273
R9146 VDPWR.n2514 VDPWR.n2513 9.73273
R9147 VDPWR.n2513 VDPWR.n2512 9.73273
R9148 VDPWR.n2512 VDPWR.n1143 9.73273
R9149 VDPWR.n2496 VDPWR.n1158 9.73273
R9150 VDPWR.n2492 VDPWR.n2491 9.73273
R9151 VDPWR.n2725 VDPWR.n2700 9.73273
R9152 VDPWR.n2721 VDPWR.n2700 9.73273
R9153 VDPWR.n2721 VDPWR.n2720 9.73273
R9154 VDPWR.n2341 VDPWR.n2340 9.71972
R9155 VDPWR.n2424 VDPWR.n2422 9.71972
R9156 VDPWR.n2288 VDPWR.n2287 9.71084
R9157 VDPWR.n2303 VDPWR.n2302 9.65296
R9158 VDPWR.n2313 VDPWR.n2312 9.65296
R9159 VDPWR.n2325 VDPWR.n1226 9.65296
R9160 VDPWR.n2330 VDPWR.n2327 9.65296
R9161 VDPWR.n2383 VDPWR.n1200 9.65296
R9162 VDPWR.n2386 VDPWR.n2385 9.65296
R9163 VDPWR.n2393 VDPWR.n2389 9.65296
R9164 VDPWR.n2417 VDPWR.n2414 9.65296
R9165 VDPWR.n599 VDPWR.n598 9.60526
R9166 VDPWR.n587 VDPWR.n586 9.60526
R9167 VDPWR.n552 VDPWR.n551 9.60526
R9168 VDPWR.n319 VDPWR.n318 9.60526
R9169 VDPWR.n307 VDPWR.n306 9.60526
R9170 VDPWR.n272 VDPWR.n271 9.60526
R9171 VDPWR.n62 VDPWR.n61 9.60526
R9172 VDPWR.n50 VDPWR.n49 9.60526
R9173 VDPWR.n15 VDPWR.n14 9.60526
R9174 VDPWR.n975 VDPWR.n972 9.6005
R9175 VDPWR.n2552 VDPWR.n995 9.56172
R9176 VDPWR.n2497 VDPWR.n2496 9.52116
R9177 VDPWR.n1788 VDPWR.n1787 9.49016
R9178 VDPWR.n2409 VDPWR.n2408 9.35121
R9179 VDPWR.n250 VDPWR 9.30627
R9180 VDPWR.n589 VDPWR.n565 9.3005
R9181 VDPWR.n625 VDPWR.n624 9.3005
R9182 VDPWR.n622 VDPWR.n566 9.3005
R9183 VDPWR.n621 VDPWR.n619 9.3005
R9184 VDPWR.n618 VDPWR.n590 9.3005
R9185 VDPWR.n617 VDPWR.n616 9.3005
R9186 VDPWR.n615 VDPWR.n591 9.3005
R9187 VDPWR.n614 VDPWR.n613 9.3005
R9188 VDPWR.n612 VDPWR.n592 9.3005
R9189 VDPWR.n611 VDPWR.n610 9.3005
R9190 VDPWR.n609 VDPWR.n608 9.3005
R9191 VDPWR.n607 VDPWR.n593 9.3005
R9192 VDPWR.n606 VDPWR.n605 9.3005
R9193 VDPWR.n604 VDPWR.n603 9.3005
R9194 VDPWR.n602 VDPWR.n601 9.3005
R9195 VDPWR.n600 VDPWR.n596 9.3005
R9196 VDPWR.n572 VDPWR.n571 9.3005
R9197 VDPWR.n575 VDPWR.n567 9.3005
R9198 VDPWR.n584 VDPWR.n583 9.3005
R9199 VDPWR.n581 VDPWR.n568 9.3005
R9200 VDPWR.n580 VDPWR.n579 9.3005
R9201 VDPWR.n578 VDPWR.n563 9.3005
R9202 VDPWR.n629 VDPWR.n628 9.3005
R9203 VDPWR.n630 VDPWR.n562 9.3005
R9204 VDPWR.n635 VDPWR.n634 9.3005
R9205 VDPWR.n636 VDPWR.n561 9.3005
R9206 VDPWR.n639 VDPWR.n638 9.3005
R9207 VDPWR.n637 VDPWR.n538 9.3005
R9208 VDPWR.n651 VDPWR.n650 9.3005
R9209 VDPWR.n649 VDPWR.n537 9.3005
R9210 VDPWR.n648 VDPWR.n647 9.3005
R9211 VDPWR.n646 VDPWR.n645 9.3005
R9212 VDPWR.n644 VDPWR.n541 9.3005
R9213 VDPWR.n643 VDPWR.n546 9.3005
R9214 VDPWR.n558 VDPWR.n557 9.3005
R9215 VDPWR.n556 VDPWR.n555 9.3005
R9216 VDPWR.n553 VDPWR.n548 9.3005
R9217 VDPWR.n309 VDPWR.n285 9.3005
R9218 VDPWR.n345 VDPWR.n344 9.3005
R9219 VDPWR.n342 VDPWR.n286 9.3005
R9220 VDPWR.n341 VDPWR.n339 9.3005
R9221 VDPWR.n338 VDPWR.n310 9.3005
R9222 VDPWR.n337 VDPWR.n336 9.3005
R9223 VDPWR.n335 VDPWR.n311 9.3005
R9224 VDPWR.n334 VDPWR.n333 9.3005
R9225 VDPWR.n332 VDPWR.n312 9.3005
R9226 VDPWR.n331 VDPWR.n330 9.3005
R9227 VDPWR.n329 VDPWR.n328 9.3005
R9228 VDPWR.n327 VDPWR.n313 9.3005
R9229 VDPWR.n326 VDPWR.n325 9.3005
R9230 VDPWR.n324 VDPWR.n323 9.3005
R9231 VDPWR.n322 VDPWR.n321 9.3005
R9232 VDPWR.n320 VDPWR.n316 9.3005
R9233 VDPWR.n292 VDPWR.n291 9.3005
R9234 VDPWR.n295 VDPWR.n287 9.3005
R9235 VDPWR.n304 VDPWR.n303 9.3005
R9236 VDPWR.n301 VDPWR.n288 9.3005
R9237 VDPWR.n300 VDPWR.n299 9.3005
R9238 VDPWR.n298 VDPWR.n283 9.3005
R9239 VDPWR.n349 VDPWR.n348 9.3005
R9240 VDPWR.n350 VDPWR.n282 9.3005
R9241 VDPWR.n355 VDPWR.n354 9.3005
R9242 VDPWR.n356 VDPWR.n281 9.3005
R9243 VDPWR.n359 VDPWR.n358 9.3005
R9244 VDPWR.n357 VDPWR.n258 9.3005
R9245 VDPWR.n371 VDPWR.n370 9.3005
R9246 VDPWR.n369 VDPWR.n257 9.3005
R9247 VDPWR.n368 VDPWR.n367 9.3005
R9248 VDPWR.n366 VDPWR.n365 9.3005
R9249 VDPWR.n364 VDPWR.n261 9.3005
R9250 VDPWR.n363 VDPWR.n266 9.3005
R9251 VDPWR.n278 VDPWR.n277 9.3005
R9252 VDPWR.n276 VDPWR.n275 9.3005
R9253 VDPWR.n273 VDPWR.n268 9.3005
R9254 VDPWR.n143 VDPWR.n142 9.3005
R9255 VDPWR.n144 VDPWR.n138 9.3005
R9256 VDPWR.n145 VDPWR.n137 9.3005
R9257 VDPWR.n149 VDPWR.n148 9.3005
R9258 VDPWR.n150 VDPWR.n136 9.3005
R9259 VDPWR.n175 VDPWR.n174 9.3005
R9260 VDPWR.n173 VDPWR.n135 9.3005
R9261 VDPWR.n172 VDPWR.n171 9.3005
R9262 VDPWR.n170 VDPWR.n151 9.3005
R9263 VDPWR.n169 VDPWR.n168 9.3005
R9264 VDPWR.n167 VDPWR.n152 9.3005
R9265 VDPWR.n166 VDPWR.n165 9.3005
R9266 VDPWR.n164 VDPWR.n163 9.3005
R9267 VDPWR.n162 VDPWR.n153 9.3005
R9268 VDPWR.n161 VDPWR.n160 9.3005
R9269 VDPWR.n159 VDPWR.n158 9.3005
R9270 VDPWR.n157 VDPWR.n154 9.3005
R9271 VDPWR.n156 VDPWR.n155 9.3005
R9272 VDPWR.n129 VDPWR.n127 9.3005
R9273 VDPWR.n201 VDPWR.n200 9.3005
R9274 VDPWR.n199 VDPWR.n128 9.3005
R9275 VDPWR.n198 VDPWR.n197 9.3005
R9276 VDPWR.n196 VDPWR.n130 9.3005
R9277 VDPWR.n195 VDPWR.n194 9.3005
R9278 VDPWR.n193 VDPWR.n192 9.3005
R9279 VDPWR.n191 VDPWR.n131 9.3005
R9280 VDPWR.n190 VDPWR.n189 9.3005
R9281 VDPWR.n188 VDPWR.n187 9.3005
R9282 VDPWR.n186 VDPWR.n132 9.3005
R9283 VDPWR.n185 VDPWR.n184 9.3005
R9284 VDPWR.n183 VDPWR.n182 9.3005
R9285 VDPWR.n181 VDPWR.n133 9.3005
R9286 VDPWR.n180 VDPWR.n179 9.3005
R9287 VDPWR.n178 VDPWR.n177 9.3005
R9288 VDPWR.n252 VDPWR.n251 9.3005
R9289 VDPWR.n249 VDPWR.n120 9.3005
R9290 VDPWR.n248 VDPWR.n247 9.3005
R9291 VDPWR.n246 VDPWR.n121 9.3005
R9292 VDPWR.n245 VDPWR.n122 9.3005
R9293 VDPWR.n244 VDPWR.n243 9.3005
R9294 VDPWR.n242 VDPWR.n123 9.3005
R9295 VDPWR.n241 VDPWR.n240 9.3005
R9296 VDPWR.n239 VDPWR.n238 9.3005
R9297 VDPWR.n237 VDPWR.n124 9.3005
R9298 VDPWR.n236 VDPWR.n235 9.3005
R9299 VDPWR.n234 VDPWR.n233 9.3005
R9300 VDPWR.n232 VDPWR.n125 9.3005
R9301 VDPWR.n231 VDPWR.n230 9.3005
R9302 VDPWR.n229 VDPWR.n228 9.3005
R9303 VDPWR.n227 VDPWR.n126 9.3005
R9304 VDPWR.n226 VDPWR.n225 9.3005
R9305 VDPWR.n224 VDPWR.n223 9.3005
R9306 VDPWR.n222 VDPWR.n204 9.3005
R9307 VDPWR.n221 VDPWR.n220 9.3005
R9308 VDPWR.n219 VDPWR.n218 9.3005
R9309 VDPWR.n217 VDPWR.n205 9.3005
R9310 VDPWR.n216 VDPWR.n215 9.3005
R9311 VDPWR.n214 VDPWR.n213 9.3005
R9312 VDPWR.n212 VDPWR.n206 9.3005
R9313 VDPWR.n211 VDPWR.n210 9.3005
R9314 VDPWR.n209 VDPWR.n208 9.3005
R9315 VDPWR.n207 VDPWR.n119 9.3005
R9316 VDPWR.n1725 VDPWR.n1724 9.3005
R9317 VDPWR.n1724 VDPWR.n1436 9.3005
R9318 VDPWR.n1724 VDPWR.n1720 9.3005
R9319 VDPWR.n1527 VDPWR.n1526 9.3005
R9320 VDPWR.n1534 VDPWR.n1533 9.3005
R9321 VDPWR.n1536 VDPWR.n1506 9.3005
R9322 VDPWR.n1538 VDPWR.n1537 9.3005
R9323 VDPWR.n1547 VDPWR.n1546 9.3005
R9324 VDPWR.n1548 VDPWR.n1500 9.3005
R9325 VDPWR.n1551 VDPWR.n1550 9.3005
R9326 VDPWR.n1552 VDPWR.n1499 9.3005
R9327 VDPWR.n1554 VDPWR.n1553 9.3005
R9328 VDPWR.n1556 VDPWR.n1498 9.3005
R9329 VDPWR.n1558 VDPWR.n1557 9.3005
R9330 VDPWR.n1560 VDPWR.n1559 9.3005
R9331 VDPWR.n1562 VDPWR.n1496 9.3005
R9332 VDPWR.n1565 VDPWR.n1564 9.3005
R9333 VDPWR.n1566 VDPWR.n1495 9.3005
R9334 VDPWR.n1568 VDPWR.n1567 9.3005
R9335 VDPWR.n1570 VDPWR.n1493 9.3005
R9336 VDPWR.n1573 VDPWR.n1572 9.3005
R9337 VDPWR.n1571 VDPWR.n1487 9.3005
R9338 VDPWR.n1586 VDPWR.n1585 9.3005
R9339 VDPWR.n1590 VDPWR.n1589 9.3005
R9340 VDPWR.n1593 VDPWR.n1481 9.3005
R9341 VDPWR.n1596 VDPWR.n1595 9.3005
R9342 VDPWR.n1597 VDPWR.n1480 9.3005
R9343 VDPWR.n1599 VDPWR.n1598 9.3005
R9344 VDPWR.n1601 VDPWR.n1479 9.3005
R9345 VDPWR.n1604 VDPWR.n1603 9.3005
R9346 VDPWR.n1602 VDPWR.n1478 9.3005
R9347 VDPWR.n1610 VDPWR.n1473 9.3005
R9348 VDPWR.n1619 VDPWR.n1618 9.3005
R9349 VDPWR.n1620 VDPWR.n1472 9.3005
R9350 VDPWR.n1622 VDPWR.n1621 9.3005
R9351 VDPWR.n1623 VDPWR 9.3005
R9352 VDPWR.n1625 VDPWR.n1624 9.3005
R9353 VDPWR.n1627 VDPWR.n1626 9.3005
R9354 VDPWR.n1628 VDPWR.n1469 9.3005
R9355 VDPWR.n1630 VDPWR.n1629 9.3005
R9356 VDPWR.n1632 VDPWR.n1631 9.3005
R9357 VDPWR.n1633 VDPWR.n1467 9.3005
R9358 VDPWR.n1635 VDPWR.n1634 9.3005
R9359 VDPWR.n1636 VDPWR.n1466 9.3005
R9360 VDPWR.n1643 VDPWR.n1642 9.3005
R9361 VDPWR.n1644 VDPWR.n1464 9.3005
R9362 VDPWR.n1648 VDPWR.n1647 9.3005
R9363 VDPWR.n1645 VDPWR.n1460 9.3005
R9364 VDPWR.n1656 VDPWR.n1459 9.3005
R9365 VDPWR.n1658 VDPWR.n1657 9.3005
R9366 VDPWR.n1660 VDPWR.n1659 9.3005
R9367 VDPWR.n1662 VDPWR.n1661 9.3005
R9368 VDPWR.n1664 VDPWR.n1457 9.3005
R9369 VDPWR.n1668 VDPWR.n1667 9.3005
R9370 VDPWR.n1669 VDPWR.n1456 9.3005
R9371 VDPWR.n1671 VDPWR.n1670 9.3005
R9372 VDPWR.n1672 VDPWR.n1455 9.3005
R9373 VDPWR.n1675 VDPWR.n1674 9.3005
R9374 VDPWR.n1676 VDPWR.n1454 9.3005
R9375 VDPWR.n1682 VDPWR.n1681 9.3005
R9376 VDPWR.n1684 VDPWR.n1683 9.3005
R9377 VDPWR.n1693 VDPWR.n1692 9.3005
R9378 VDPWR.n1695 VDPWR.n1694 9.3005
R9379 VDPWR.n1697 VDPWR.n1696 9.3005
R9380 VDPWR.n1698 VDPWR.n1445 9.3005
R9381 VDPWR.n1700 VDPWR.n1699 9.3005
R9382 VDPWR.n1702 VDPWR.n1701 9.3005
R9383 VDPWR.n1703 VDPWR.n1443 9.3005
R9384 VDPWR.n1705 VDPWR.n1704 9.3005
R9385 VDPWR.n1706 VDPWR.n1442 9.3005
R9386 VDPWR.n1708 VDPWR.n1707 9.3005
R9387 VDPWR.n1709 VDPWR.n1441 9.3005
R9388 VDPWR.n1712 VDPWR.n1711 9.3005
R9389 VDPWR.n1713 VDPWR.n1437 9.3005
R9390 VDPWR.n1749 VDPWR.n1748 9.3005
R9391 VDPWR.n1749 VDPWR.n1426 9.3005
R9392 VDPWR.n1749 VDPWR.n1425 9.3005
R9393 VDPWR.n1302 VDPWR.n1301 9.3005
R9394 VDPWR.n1304 VDPWR.n1303 9.3005
R9395 VDPWR.n1889 VDPWR.n1888 9.3005
R9396 VDPWR.n1887 VDPWR.n1886 9.3005
R9397 VDPWR.n1878 VDPWR.n1877 9.3005
R9398 VDPWR.n1876 VDPWR.n1307 9.3005
R9399 VDPWR.n1875 VDPWR.n1874 9.3005
R9400 VDPWR.n1873 VDPWR.n1872 9.3005
R9401 VDPWR.n1871 VDPWR.n1870 9.3005
R9402 VDPWR.n1869 VDPWR.n1868 9.3005
R9403 VDPWR.n1867 VDPWR.n1310 9.3005
R9404 VDPWR.n1865 VDPWR.n1864 9.3005
R9405 VDPWR.n1863 VDPWR.n1862 9.3005
R9406 VDPWR.n1860 VDPWR.n1312 9.3005
R9407 VDPWR.n1859 VDPWR.n1858 9.3005
R9408 VDPWR.n1857 VDPWR.n1313 9.3005
R9409 VDPWR.n1321 VDPWR.n1314 9.3005
R9410 VDPWR.n1327 VDPWR.n1326 9.3005
R9411 VDPWR.n1328 VDPWR.n1319 9.3005
R9412 VDPWR.n1848 VDPWR.n1847 9.3005
R9413 VDPWR.n1846 VDPWR.n1845 9.3005
R9414 VDPWR.n1844 VDPWR.n1331 9.3005
R9415 VDPWR.n1834 VDPWR.n1833 9.3005
R9416 VDPWR.n1832 VDPWR.n1831 9.3005
R9417 VDPWR.n1829 VDPWR.n1334 9.3005
R9418 VDPWR.n1828 VDPWR.n1827 9.3005
R9419 VDPWR.n1344 VDPWR.n1336 9.3005
R9420 VDPWR.n1352 VDPWR.n1351 9.3005
R9421 VDPWR.n1353 VDPWR.n1342 9.3005
R9422 VDPWR.n1819 VDPWR.n1818 9.3005
R9423 VDPWR.n1817 VDPWR.n1343 9.3005
R9424 VDPWR.n1815 VDPWR.n1814 9.3005
R9425 VDPWR.n1810 VDPWR.n1809 9.3005
R9426 VDPWR.n1808 VDPWR.n1807 9.3005
R9427 VDPWR.n1805 VDPWR.n1356 9.3005
R9428 VDPWR.n1804 VDPWR.n1803 9.3005
R9429 VDPWR.n1802 VDPWR.n1801 9.3005
R9430 VDPWR.n1800 VDPWR.n1358 9.3005
R9431 VDPWR.n1799 VDPWR.n1798 9.3005
R9432 VDPWR.n1368 VDPWR.n1359 9.3005
R9433 VDPWR.n1375 VDPWR.n1374 9.3005
R9434 VDPWR.n1377 VDPWR.n1366 9.3005
R9435 VDPWR.n1790 VDPWR.n1789 9.3005
R9436 VDPWR.n1787 VDPWR.n1786 9.3005
R9437 VDPWR.n1784 VDPWR.n1783 9.3005
R9438 VDPWR.n1780 VDPWR.n1779 9.3005
R9439 VDPWR.n1778 VDPWR.n1385 9.3005
R9440 VDPWR.n1777 VDPWR.n1776 9.3005
R9441 VDPWR.n1775 VDPWR.n1386 9.3005
R9442 VDPWR.n1774 VDPWR.n1773 9.3005
R9443 VDPWR.n1389 VDPWR.n1388 9.3005
R9444 VDPWR.n1405 VDPWR.n1404 9.3005
R9445 VDPWR.n1408 VDPWR.n1407 9.3005
R9446 VDPWR.n1765 VDPWR.n1764 9.3005
R9447 VDPWR.n1763 VDPWR.n1395 9.3005
R9448 VDPWR.n1762 VDPWR.n1761 9.3005
R9449 VDPWR.n1760 VDPWR.n1759 9.3005
R9450 VDPWR.n1758 VDPWR.n1410 9.3005
R9451 VDPWR.n1755 VDPWR.n1754 9.3005
R9452 VDPWR.n1753 VDPWR.n1413 9.3005
R9453 VDPWR.n1752 VDPWR.n1751 9.3005
R9454 VDPWR.n1750 VDPWR.n1417 9.3005
R9455 VDPWR.n2063 VDPWR.n2062 9.3005
R9456 VDPWR.n2064 VDPWR.n2063 9.3005
R9457 VDPWR.n2063 VDPWR.n2049 9.3005
R9458 VDPWR.n1908 VDPWR.n1903 9.3005
R9459 VDPWR.n1907 VDPWR.n1901 9.3005
R9460 VDPWR.n1928 VDPWR.n1927 9.3005
R9461 VDPWR.n1926 VDPWR.n1925 9.3005
R9462 VDPWR.n1938 VDPWR.n1937 9.3005
R9463 VDPWR.n1939 VDPWR.n1271 9.3005
R9464 VDPWR.n1942 VDPWR.n1941 9.3005
R9465 VDPWR.n1943 VDPWR.n1270 9.3005
R9466 VDPWR.n1945 VDPWR.n1944 9.3005
R9467 VDPWR.n1947 VDPWR.n1269 9.3005
R9468 VDPWR.n1949 VDPWR.n1948 9.3005
R9469 VDPWR.n1951 VDPWR.n1950 9.3005
R9470 VDPWR.n1953 VDPWR.n1267 9.3005
R9471 VDPWR.n1956 VDPWR.n1955 9.3005
R9472 VDPWR.n1957 VDPWR.n1266 9.3005
R9473 VDPWR.n1959 VDPWR.n1958 9.3005
R9474 VDPWR.n1961 VDPWR.n1262 9.3005
R9475 VDPWR.n1962 VDPWR.n1263 9.3005
R9476 VDPWR.n2177 VDPWR.n2176 9.3005
R9477 VDPWR.n2174 VDPWR.n2173 9.3005
R9478 VDPWR.n2172 VDPWR.n1963 9.3005
R9479 VDPWR.n2170 VDPWR.n2169 9.3005
R9480 VDPWR.n2162 VDPWR.n1966 9.3005
R9481 VDPWR.n2161 VDPWR.n2160 9.3005
R9482 VDPWR.n2159 VDPWR.n1968 9.3005
R9483 VDPWR.n2158 VDPWR.n2157 9.3005
R9484 VDPWR.n2156 VDPWR.n2155 9.3005
R9485 VDPWR.n1979 VDPWR.n1972 9.3005
R9486 VDPWR.n1985 VDPWR.n1984 9.3005
R9487 VDPWR.n1986 VDPWR.n1977 9.3005
R9488 VDPWR.n2146 VDPWR.n2145 9.3005
R9489 VDPWR.n2144 VDPWR.n1978 9.3005
R9490 VDPWR.n2142 VDPWR.n2141 9.3005
R9491 VDPWR.n2140 VDPWR.n1988 9.3005
R9492 VDPWR.n2139 VDPWR.n2138 9.3005
R9493 VDPWR.n2137 VDPWR.n1989 9.3005
R9494 VDPWR.n2136 VDPWR.n2135 9.3005
R9495 VDPWR.n2134 VDPWR.n2133 9.3005
R9496 VDPWR.n2132 VDPWR.n2131 9.3005
R9497 VDPWR.n2130 VDPWR.n2129 9.3005
R9498 VDPWR.n2128 VDPWR.n1994 9.3005
R9499 VDPWR.n2127 VDPWR.n2126 9.3005
R9500 VDPWR.n2005 VDPWR.n2004 9.3005
R9501 VDPWR.n2010 VDPWR.n2009 9.3005
R9502 VDPWR.n2012 VDPWR.n2001 9.3005
R9503 VDPWR.n2117 VDPWR.n2116 9.3005
R9504 VDPWR.n2115 VDPWR.n2114 9.3005
R9505 VDPWR.n2113 VDPWR.n2112 9.3005
R9506 VDPWR.n2111 VDPWR.n2014 9.3005
R9507 VDPWR.n2109 VDPWR.n2108 9.3005
R9508 VDPWR.n2107 VDPWR.n2016 9.3005
R9509 VDPWR.n2106 VDPWR.n2105 9.3005
R9510 VDPWR.n2103 VDPWR.n2017 9.3005
R9511 VDPWR.n2101 VDPWR.n2100 9.3005
R9512 VDPWR.n2099 VDPWR.n2098 9.3005
R9513 VDPWR.n2097 VDPWR.n2019 9.3005
R9514 VDPWR.n2095 VDPWR 9.3005
R9515 VDPWR.n2027 VDPWR.n2020 9.3005
R9516 VDPWR.n2035 VDPWR.n2029 9.3005
R9517 VDPWR.n2085 VDPWR.n2084 9.3005
R9518 VDPWR.n2081 VDPWR.n2080 9.3005
R9519 VDPWR.n2078 VDPWR.n2037 9.3005
R9520 VDPWR.n2077 VDPWR.n2076 9.3005
R9521 VDPWR.n2074 VDPWR.n2038 9.3005
R9522 VDPWR.n2073 VDPWR.n2072 9.3005
R9523 VDPWR.n2051 VDPWR.n2044 9.3005
R9524 VDPWR.n2447 VDPWR.n2446 9.3005
R9525 VDPWR.n2446 VDPWR.n1172 9.3005
R9526 VDPWR.n2446 VDPWR.n2442 9.3005
R9527 VDPWR.n2221 VDPWR.n2220 9.3005
R9528 VDPWR.n2224 VDPWR.n2223 9.3005
R9529 VDPWR.n2230 VDPWR.n2229 9.3005
R9530 VDPWR.n2234 VDPWR.n2233 9.3005
R9531 VDPWR.n2235 VDPWR.n2199 9.3005
R9532 VDPWR.n2244 VDPWR.n2243 9.3005
R9533 VDPWR.n2245 VDPWR.n2198 9.3005
R9534 VDPWR.n2247 VDPWR.n2246 9.3005
R9535 VDPWR.n2249 VDPWR.n2248 9.3005
R9536 VDPWR.n2250 VDPWR.n2196 9.3005
R9537 VDPWR.n2253 VDPWR.n2252 9.3005
R9538 VDPWR.n2255 VDPWR.n2254 9.3005
R9539 VDPWR.n2258 VDPWR.n2257 9.3005
R9540 VDPWR.n2260 VDPWR.n2259 9.3005
R9541 VDPWR.n2261 VDPWR.n2193 9.3005
R9542 VDPWR.n2263 VDPWR.n2262 9.3005
R9543 VDPWR.n2265 VDPWR.n2264 9.3005
R9544 VDPWR.n2267 VDPWR.n2266 9.3005
R9545 VDPWR.n1254 VDPWR.n1253 9.3005
R9546 VDPWR.n2280 VDPWR.n2279 9.3005
R9547 VDPWR.n2283 VDPWR.n2282 9.3005
R9548 VDPWR.n2284 VDPWR.n1251 9.3005
R9549 VDPWR.n2286 VDPWR.n2285 9.3005
R9550 VDPWR.n2289 VDPWR.n2288 9.3005
R9551 VDPWR.n2291 VDPWR.n2290 9.3005
R9552 VDPWR.n2296 VDPWR.n2295 9.3005
R9553 VDPWR.n2297 VDPWR.n1244 9.3005
R9554 VDPWR.n2299 VDPWR.n2298 9.3005
R9555 VDPWR.n2302 VDPWR.n1242 9.3005
R9556 VDPWR.n2304 VDPWR.n2303 9.3005
R9557 VDPWR.n2306 VDPWR.n2305 9.3005
R9558 VDPWR.n2308 VDPWR.n1234 9.3005
R9559 VDPWR.n2314 VDPWR.n2313 9.3005
R9560 VDPWR.n2312 VDPWR.n1227 9.3005
R9561 VDPWR.n2323 VDPWR.n1226 9.3005
R9562 VDPWR.n2325 VDPWR.n2324 9.3005
R9563 VDPWR.n2327 VDPWR.n1224 9.3005
R9564 VDPWR.n2331 VDPWR.n2330 9.3005
R9565 VDPWR.n2333 VDPWR.n2332 9.3005
R9566 VDPWR.n2334 VDPWR.n1221 9.3005
R9567 VDPWR.n2338 VDPWR.n2337 9.3005
R9568 VDPWR.n2340 VDPWR.n2339 9.3005
R9569 VDPWR.n2341 VDPWR.n1218 9.3005
R9570 VDPWR.n2345 VDPWR.n2344 9.3005
R9571 VDPWR.n2346 VDPWR.n1217 9.3005
R9572 VDPWR.n2348 VDPWR.n2347 9.3005
R9573 VDPWR.n2354 VDPWR.n2353 9.3005
R9574 VDPWR.n2352 VDPWR.n2351 9.3005
R9575 VDPWR.n2364 VDPWR.n2363 9.3005
R9576 VDPWR.n2366 VDPWR.n2365 9.3005
R9577 VDPWR.n2368 VDPWR.n2367 9.3005
R9578 VDPWR.n2371 VDPWR.n2370 9.3005
R9579 VDPWR.n2373 VDPWR.n2372 9.3005
R9580 VDPWR.n2375 VDPWR.n1201 9.3005
R9581 VDPWR.n2380 VDPWR.n2379 9.3005
R9582 VDPWR.n2381 VDPWR.n1200 9.3005
R9583 VDPWR.n2383 VDPWR.n2382 9.3005
R9584 VDPWR.n2385 VDPWR.n1198 9.3005
R9585 VDPWR.n2387 VDPWR.n2386 9.3005
R9586 VDPWR.n2389 VDPWR.n2388 9.3005
R9587 VDPWR.n2394 VDPWR.n2393 9.3005
R9588 VDPWR.n2391 VDPWR.n1188 9.3005
R9589 VDPWR.n2407 VDPWR.n2406 9.3005
R9590 VDPWR.n2410 VDPWR.n2409 9.3005
R9591 VDPWR.n2412 VDPWR.n2411 9.3005
R9592 VDPWR.n2414 VDPWR.n1182 9.3005
R9593 VDPWR.n2418 VDPWR.n2417 9.3005
R9594 VDPWR.n2420 VDPWR.n2419 9.3005
R9595 VDPWR.n2422 VDPWR.n1179 9.3005
R9596 VDPWR.n2425 VDPWR.n2424 9.3005
R9597 VDPWR.n2426 VDPWR.n1178 9.3005
R9598 VDPWR.n2428 VDPWR.n2427 9.3005
R9599 VDPWR.n2431 VDPWR.n1177 9.3005
R9600 VDPWR.n2434 VDPWR.n2433 9.3005
R9601 VDPWR.n2435 VDPWR.n1173 9.3005
R9602 VDPWR.n2474 VDPWR.n2473 9.3005
R9603 VDPWR.n2475 VDPWR.n2474 9.3005
R9604 VDPWR.n2474 VDPWR.n2459 9.3005
R9605 VDPWR.n971 VDPWR.n970 9.3005
R9606 VDPWR.n978 VDPWR.n977 9.3005
R9607 VDPWR.n2577 VDPWR.n2576 9.3005
R9608 VDPWR.n2576 VDPWR.n2575 9.3005
R9609 VDPWR.n2570 VDPWR.n2569 9.3005
R9610 VDPWR.n2568 VDPWR.n2567 9.3005
R9611 VDPWR.n2566 VDPWR.n2565 9.3005
R9612 VDPWR.n2564 VDPWR.n987 9.3005
R9613 VDPWR.n2563 VDPWR.n2562 9.3005
R9614 VDPWR.n2561 VDPWR.n2560 9.3005
R9615 VDPWR.n2556 VDPWR.n989 9.3005
R9616 VDPWR.n996 VDPWR.n992 9.3005
R9617 VDPWR.n2554 VDPWR.n2553 9.3005
R9618 VDPWR.n2551 VDPWR.n2550 9.3005
R9619 VDPWR.n2547 VDPWR.n997 9.3005
R9620 VDPWR.n2546 VDPWR.n2545 9.3005
R9621 VDPWR.n1014 VDPWR.n1013 9.3005
R9622 VDPWR.n1015 VDPWR.n1008 9.3005
R9623 VDPWR.n2535 VDPWR.n2534 9.3005
R9624 VDPWR.n2533 VDPWR.n1018 9.3005
R9625 VDPWR.n1049 VDPWR.n1048 9.3005
R9626 VDPWR.n1050 VDPWR.n1045 9.3005
R9627 VDPWR.n1052 VDPWR.n1051 9.3005
R9628 VDPWR.n1056 VDPWR.n1055 9.3005
R9629 VDPWR.n1057 VDPWR.n1044 9.3005
R9630 VDPWR.n1059 VDPWR.n1058 9.3005
R9631 VDPWR.n1062 VDPWR.n1061 9.3005
R9632 VDPWR.n1063 VDPWR.n1043 9.3005
R9633 VDPWR.n1065 VDPWR.n1064 9.3005
R9634 VDPWR.n1069 VDPWR.n1068 9.3005
R9635 VDPWR.n1070 VDPWR.n1036 9.3005
R9636 VDPWR.n1083 VDPWR.n1082 9.3005
R9637 VDPWR.n1088 VDPWR.n1087 9.3005
R9638 VDPWR.n1089 VDPWR.n1034 9.3005
R9639 VDPWR.n1091 VDPWR.n1090 9.3005
R9640 VDPWR.n1093 VDPWR.n1033 9.3005
R9641 VDPWR.n1095 VDPWR.n1094 9.3005
R9642 VDPWR.n1096 VDPWR.n1032 9.3005
R9643 VDPWR.n1098 VDPWR.n1097 9.3005
R9644 VDPWR.n1100 VDPWR.n1030 9.3005
R9645 VDPWR.n1102 VDPWR.n1101 9.3005
R9646 VDPWR.n1104 VDPWR.n1103 9.3005
R9647 VDPWR.n1109 VDPWR.n1108 9.3005
R9648 VDPWR.n1116 VDPWR.n1115 9.3005
R9649 VDPWR.n1119 VDPWR.n1026 9.3005
R9650 VDPWR.n1124 VDPWR.n1123 9.3005
R9651 VDPWR.n1022 VDPWR.n1021 9.3005
R9652 VDPWR.n2530 VDPWR.n1132 9.3005
R9653 VDPWR.n2529 VDPWR.n2528 9.3005
R9654 VDPWR.n2527 VDPWR.n1133 9.3005
R9655 VDPWR.n2526 VDPWR.n2525 9.3005
R9656 VDPWR.n2524 VDPWR.n1134 9.3005
R9657 VDPWR.n2522 VDPWR.n2521 9.3005
R9658 VDPWR.n2520 VDPWR.n2519 9.3005
R9659 VDPWR.n2518 VDPWR.n1139 9.3005
R9660 VDPWR.n2517 VDPWR.n2516 9.3005
R9661 VDPWR.n2515 VDPWR.n2514 9.3005
R9662 VDPWR.n2513 VDPWR.n1142 9.3005
R9663 VDPWR.n2512 VDPWR.n2511 9.3005
R9664 VDPWR.n1152 VDPWR.n1143 9.3005
R9665 VDPWR.n1155 VDPWR.n1154 9.3005
R9666 VDPWR.n2501 VDPWR.n2500 9.3005
R9667 VDPWR.n2498 VDPWR.n1150 9.3005
R9668 VDPWR.n2496 VDPWR.n2495 9.3005
R9669 VDPWR.n2494 VDPWR.n1158 9.3005
R9670 VDPWR.n2493 VDPWR.n2492 9.3005
R9671 VDPWR.n2491 VDPWR.n1159 9.3005
R9672 VDPWR.n2490 VDPWR.n2489 9.3005
R9673 VDPWR.n2488 VDPWR.n2487 9.3005
R9674 VDPWR.n2486 VDPWR.n1163 9.3005
R9675 VDPWR.n2485 VDPWR.n2484 9.3005
R9676 VDPWR.n2483 VDPWR.n1164 9.3005
R9677 VDPWR.n2462 VDPWR.n1165 9.3005
R9678 VDPWR.n2971 VDPWR.n2970 9.3005
R9679 VDPWR.n2970 VDPWR.n2966 9.3005
R9680 VDPWR.n2970 VDPWR.n2963 9.3005
R9681 VDPWR.n2605 VDPWR.n2604 9.3005
R9682 VDPWR.n2607 VDPWR.n2606 9.3005
R9683 VDPWR.n2809 VDPWR.n2808 9.3005
R9684 VDPWR.n2810 VDPWR.n946 9.3005
R9685 VDPWR.n2812 VDPWR.n2811 9.3005
R9686 VDPWR.n2813 VDPWR.n945 9.3005
R9687 VDPWR.n2815 VDPWR.n2814 9.3005
R9688 VDPWR.n2816 VDPWR.n942 9.3005
R9689 VDPWR.n2819 VDPWR.n2818 9.3005
R9690 VDPWR.n2820 VDPWR.n941 9.3005
R9691 VDPWR.n2822 VDPWR.n2821 9.3005
R9692 VDPWR.n2823 VDPWR.n940 9.3005
R9693 VDPWR.n2825 VDPWR.n2824 9.3005
R9694 VDPWR.n2826 VDPWR.n938 9.3005
R9695 VDPWR.n2829 VDPWR.n2827 9.3005
R9696 VDPWR.n2831 VDPWR.n2830 9.3005
R9697 VDPWR.n2833 VDPWR.n929 9.3005
R9698 VDPWR.n930 VDPWR.n929 9.3005
R9699 VDPWR.n2845 VDPWR.n929 9.3005
R9700 VDPWR.n2849 VDPWR.n2846 9.3005
R9701 VDPWR.n2851 VDPWR.n924 9.3005
R9702 VDPWR.n2855 VDPWR.n2854 9.3005
R9703 VDPWR.n2856 VDPWR.n923 9.3005
R9704 VDPWR.n2858 VDPWR.n2857 9.3005
R9705 VDPWR.n2861 VDPWR.n921 9.3005
R9706 VDPWR.n2863 VDPWR.n2862 9.3005
R9707 VDPWR.n2864 VDPWR.n920 9.3005
R9708 VDPWR.n2866 VDPWR.n2865 9.3005
R9709 VDPWR.n2868 VDPWR.n918 9.3005
R9710 VDPWR.n2870 VDPWR.n2869 9.3005
R9711 VDPWR.n2874 VDPWR.n909 9.3005
R9712 VDPWR.n2884 VDPWR.n2883 9.3005
R9713 VDPWR.n2885 VDPWR.n906 9.3005
R9714 VDPWR.n2885 VDPWR.n905 9.3005
R9715 VDPWR.n2886 VDPWR.n902 9.3005
R9716 VDPWR.n2888 VDPWR.n2887 9.3005
R9717 VDPWR.n2889 VDPWR.n901 9.3005
R9718 VDPWR.n2891 VDPWR.n2890 9.3005
R9719 VDPWR.n2892 VDPWR.n899 9.3005
R9720 VDPWR.n2893 VDPWR.n896 9.3005
R9721 VDPWR.n2897 VDPWR.n895 9.3005
R9722 VDPWR.n2899 VDPWR.n2898 9.3005
R9723 VDPWR.n2910 VDPWR.n2909 9.3005
R9724 VDPWR.n2908 VDPWR.n2907 9.3005
R9725 VDPWR.n2903 VDPWR.n884 9.3005
R9726 VDPWR.n2919 VDPWR.n882 9.3005
R9727 VDPWR.n2926 VDPWR.n881 9.3005
R9728 VDPWR.n2928 VDPWR.n2927 9.3005
R9729 VDPWR.n2930 VDPWR.n2929 9.3005
R9730 VDPWR.n2931 VDPWR.n878 9.3005
R9731 VDPWR.n2935 VDPWR.n2934 9.3005
R9732 VDPWR.n2936 VDPWR.n877 9.3005
R9733 VDPWR.n2938 VDPWR.n2937 9.3005
R9734 VDPWR.n2939 VDPWR.n872 9.3005
R9735 VDPWR.n2941 VDPWR.n873 9.3005
R9736 VDPWR.n3000 VDPWR.n2999 9.3005
R9737 VDPWR.n2998 VDPWR.n2997 9.3005
R9738 VDPWR.n2996 VDPWR.n2995 9.3005
R9739 VDPWR.n2994 VDPWR.n2944 9.3005
R9740 VDPWR.n2993 VDPWR.n2992 9.3005
R9741 VDPWR.n2991 VDPWR.n2946 9.3005
R9742 VDPWR.n2990 VDPWR.n2989 9.3005
R9743 VDPWR.n2988 VDPWR.n2987 9.3005
R9744 VDPWR.n2986 VDPWR.n2985 9.3005
R9745 VDPWR.n2983 VDPWR.n2948 9.3005
R9746 VDPWR.n2982 VDPWR.n2981 9.3005
R9747 VDPWR.n2980 VDPWR.n2950 9.3005
R9748 VDPWR.n2958 VDPWR.n2951 9.3005
R9749 VDPWR.n837 VDPWR.n836 9.3005
R9750 VDPWR.n837 VDPWR.n829 9.3005
R9751 VDPWR.n838 VDPWR.n837 9.3005
R9752 VDPWR.n2640 VDPWR.n2639 9.3005
R9753 VDPWR.n2642 VDPWR.n2641 9.3005
R9754 VDPWR.n2643 VDPWR.n2629 9.3005
R9755 VDPWR.n2645 VDPWR.n2644 9.3005
R9756 VDPWR.n2646 VDPWR.n2627 9.3005
R9757 VDPWR.n2648 VDPWR.n2647 9.3005
R9758 VDPWR.n2652 VDPWR.n2651 9.3005
R9759 VDPWR.n2798 VDPWR.n2797 9.3005
R9760 VDPWR.n2796 VDPWR.n2621 9.3005
R9761 VDPWR.n2794 VDPWR.n2793 9.3005
R9762 VDPWR.n2792 VDPWR.n2656 9.3005
R9763 VDPWR.n2791 VDPWR.n2790 9.3005
R9764 VDPWR.n2788 VDPWR.n2657 9.3005
R9765 VDPWR.n2786 VDPWR.n2785 9.3005
R9766 VDPWR.n2784 VDPWR.n2658 9.3005
R9767 VDPWR.n2783 VDPWR.n2782 9.3005
R9768 VDPWR.n2781 VDPWR.n2780 9.3005
R9769 VDPWR.n2779 VDPWR.n2778 9.3005
R9770 VDPWR.n2777 VDPWR.n2661 9.3005
R9771 VDPWR.n2774 VDPWR.n2773 9.3005
R9772 VDPWR.n2669 VDPWR.n2663 9.3005
R9773 VDPWR.n2765 VDPWR.n2764 9.3005
R9774 VDPWR.n2763 VDPWR.n2762 9.3005
R9775 VDPWR.n2761 VDPWR.n2675 9.3005
R9776 VDPWR.n2760 VDPWR.n2759 9.3005
R9777 VDPWR.n2757 VDPWR.n2756 9.3005
R9778 VDPWR.n2755 VDPWR.n2754 9.3005
R9779 VDPWR.n2753 VDPWR.n2677 9.3005
R9780 VDPWR.n2751 VDPWR.n2750 9.3005
R9781 VDPWR.n2749 VDPWR.n2748 9.3005
R9782 VDPWR.n2747 VDPWR.n2681 9.3005
R9783 VDPWR.n2746 VDPWR.n2682 9.3005
R9784 VDPWR.n2745 VDPWR.n2744 9.3005
R9785 VDPWR.n2685 VDPWR.n2684 9.3005
R9786 VDPWR.n2693 VDPWR.n2690 9.3005
R9787 VDPWR.n2735 VDPWR.n2734 9.3005
R9788 VDPWR.n2732 VDPWR.n2731 9.3005
R9789 VDPWR.n2730 VDPWR.n2696 9.3005
R9790 VDPWR.n2729 VDPWR.n2728 9.3005
R9791 VDPWR.n2726 VDPWR.n2697 9.3005
R9792 VDPWR.n2725 VDPWR.n2724 9.3005
R9793 VDPWR.n2723 VDPWR.n2700 9.3005
R9794 VDPWR.n2722 VDPWR.n2721 9.3005
R9795 VDPWR.n2720 VDPWR.n2719 9.3005
R9796 VDPWR.n2711 VDPWR.n2710 9.3005
R9797 VDPWR.n2705 VDPWR.n783 9.3005
R9798 VDPWR.n3038 VDPWR.n3037 9.3005
R9799 VDPWR.n3036 VDPWR.n786 9.3005
R9800 VDPWR.n3035 VDPWR.n3034 9.3005
R9801 VDPWR.n3033 VDPWR.n3032 9.3005
R9802 VDPWR.n3029 VDPWR.n3028 9.3005
R9803 VDPWR.n3027 VDPWR.n789 9.3005
R9804 VDPWR.n3026 VDPWR.n3025 9.3005
R9805 VDPWR.n3024 VDPWR.n790 9.3005
R9806 VDPWR.n3023 VDPWR.n3022 9.3005
R9807 VDPWR.n3021 VDPWR.n3020 9.3005
R9808 VDPWR.n3019 VDPWR.n3018 9.3005
R9809 VDPWR.n3017 VDPWR.n796 9.3005
R9810 VDPWR.n804 VDPWR.n797 9.3005
R9811 VDPWR.n808 VDPWR.n807 9.3005
R9812 VDPWR.n863 VDPWR.n862 9.3005
R9813 VDPWR.n860 VDPWR.n859 9.3005
R9814 VDPWR.n858 VDPWR.n811 9.3005
R9815 VDPWR.n857 VDPWR.n856 9.3005
R9816 VDPWR.n855 VDPWR.n812 9.3005
R9817 VDPWR.n853 VDPWR.n852 9.3005
R9818 VDPWR.n851 VDPWR.n850 9.3005
R9819 VDPWR.n847 VDPWR.n846 9.3005
R9820 VDPWR.n845 VDPWR.n844 9.3005
R9821 VDPWR.n843 VDPWR.n820 9.3005
R9822 VDPWR.n825 VDPWR.n821 9.3005
R9823 VDPWR.n52 VDPWR.n28 9.3005
R9824 VDPWR.n88 VDPWR.n87 9.3005
R9825 VDPWR.n85 VDPWR.n29 9.3005
R9826 VDPWR.n84 VDPWR.n82 9.3005
R9827 VDPWR.n81 VDPWR.n53 9.3005
R9828 VDPWR.n80 VDPWR.n79 9.3005
R9829 VDPWR.n78 VDPWR.n54 9.3005
R9830 VDPWR.n77 VDPWR.n76 9.3005
R9831 VDPWR.n75 VDPWR.n55 9.3005
R9832 VDPWR.n74 VDPWR.n73 9.3005
R9833 VDPWR.n72 VDPWR.n71 9.3005
R9834 VDPWR.n70 VDPWR.n56 9.3005
R9835 VDPWR.n69 VDPWR.n68 9.3005
R9836 VDPWR.n67 VDPWR.n66 9.3005
R9837 VDPWR.n65 VDPWR.n64 9.3005
R9838 VDPWR.n63 VDPWR.n59 9.3005
R9839 VDPWR.n35 VDPWR.n34 9.3005
R9840 VDPWR.n38 VDPWR.n30 9.3005
R9841 VDPWR.n47 VDPWR.n46 9.3005
R9842 VDPWR.n44 VDPWR.n31 9.3005
R9843 VDPWR.n43 VDPWR.n42 9.3005
R9844 VDPWR.n41 VDPWR.n26 9.3005
R9845 VDPWR.n92 VDPWR.n91 9.3005
R9846 VDPWR.n93 VDPWR.n25 9.3005
R9847 VDPWR.n98 VDPWR.n97 9.3005
R9848 VDPWR.n99 VDPWR.n24 9.3005
R9849 VDPWR.n102 VDPWR.n101 9.3005
R9850 VDPWR.n100 VDPWR.n1 9.3005
R9851 VDPWR.n114 VDPWR.n113 9.3005
R9852 VDPWR.n112 VDPWR.n0 9.3005
R9853 VDPWR.n111 VDPWR.n110 9.3005
R9854 VDPWR.n109 VDPWR.n108 9.3005
R9855 VDPWR.n107 VDPWR.n4 9.3005
R9856 VDPWR.n106 VDPWR.n9 9.3005
R9857 VDPWR.n21 VDPWR.n20 9.3005
R9858 VDPWR.n19 VDPWR.n18 9.3005
R9859 VDPWR.n16 VDPWR.n11 9.3005
R9860 VDPWR.n1683 VDPWR.n1447 9.09802
R9861 VDPWR.n2365 VDPWR.n1204 9.09802
R9862 VDPWR.n2373 VDPWR.n1203 9.09802
R9863 VDPWR.n2374 VDPWR.n2373 9.09802
R9864 VDPWR.n1151 VDPWR.n1143 9.09802
R9865 VDPWR.n2499 VDPWR.n2498 9.09802
R9866 VDPWR.n2337 VDPWR.n2336 9.02345
R9867 VDPWR.n2391 VDPWR.n1187 9.02345
R9868 VDPWR.n2412 VDPWR.n1184 9.02345
R9869 VDPWR.n1387 VDPWR.n1385 8.99224
R9870 VDPWR.n817 VDPWR.n816 8.9761
R9871 VDPWR.n2525 VDPWR.n1137 8.88645
R9872 VDPWR.n2548 VDPWR.n2547 8.77764
R9873 VDPWR.n2337 VDPWR.n1220 8.60378
R9874 VDPWR.n2421 VDPWR.n2420 8.60378
R9875 VDPWR.n1589 VDPWR.n1586 8.44958
R9876 VDPWR.n1847 VDPWR.n1846 8.44958
R9877 VDPWR.n1789 VDPWR.n1377 8.44958
R9878 VDPWR.n2116 VDPWR.n2012 8.44958
R9879 VDPWR.n2174 VDPWR.n1963 8.44958
R9880 VDPWR.n2282 VDPWR.n1251 8.44958
R9881 VDPWR.t268 VDPWR.t743 8.39273
R9882 VDPWR.n2414 VDPWR.n2413 8.28902
R9883 VDPWR.n1759 VDPWR.n1409 8.28285
R9884 VDPWR.n2860 VDPWR.n2859 8.28285
R9885 VDPWR.n670 VDPWR.n656 8.23557
R9886 VDPWR.n427 VDPWR.n413 8.23557
R9887 VDPWR.n1011 VDPWR.n1001 8.04621
R9888 VDPWR.n2424 VDPWR.n2423 8.04017
R9889 VDPWR.n1837 VDPWR.n1836 7.98741
R9890 VDPWR.n2859 VDPWR.n2858 7.90638
R9891 VDPWR.n2850 VDPWR.n2849 7.90638
R9892 VDPWR.n1682 VDPWR.n1454 7.75995
R9893 VDPWR.n2116 VDPWR.n2115 7.75995
R9894 VDPWR.n2348 VDPWR.n1217 7.75995
R9895 VDPWR.n2365 VDPWR.n2364 7.75995
R9896 VDPWR.n2428 VDPWR.n1178 7.75995
R9897 VDPWR.n2491 VDPWR.n2490 7.75995
R9898 VDPWR.n2726 VDPWR.n2725 7.75995
R9899 VDPWR.n2329 VDPWR.n1223 7.65952
R9900 VDPWR.n717 VDPWR.n716 7.54407
R9901 VDPWR.n701 VDPWR.n700 7.54407
R9902 VDPWR.n685 VDPWR.n684 7.54407
R9903 VDPWR.n669 VDPWR.n668 7.54407
R9904 VDPWR.n528 VDPWR.n527 7.54407
R9905 VDPWR.n512 VDPWR.n511 7.54407
R9906 VDPWR.n496 VDPWR.n495 7.54407
R9907 VDPWR.n480 VDPWR.n479 7.54407
R9908 VDPWR.n458 VDPWR.n457 7.54407
R9909 VDPWR.n442 VDPWR.n441 7.54407
R9910 VDPWR.n426 VDPWR.n425 7.54407
R9911 VDPWR.n3108 VDPWR.n3107 7.54407
R9912 VDPWR.n3070 VDPWR.n3069 7.54407
R9913 VDPWR.n464 VDPWR.n463 7.54307
R9914 VDPWR.n3102 VDPWR.n3101 7.54307
R9915 VDPWR.n3086 VDPWR.n3085 7.54307
R9916 VDPWR.n2523 VDPWR.n2522 7.51124
R9917 VDPWR.n2748 VDPWR.n2747 7.49704
R9918 VDPWR.n1249 VDPWR.n1246 7.28326
R9919 VDPWR.n1247 VDPWR.n1245 7.23528
R9920 VDPWR.n2133 VDPWR.n2132 7.21067
R9921 VDPWR.n2142 VDPWR.n1988 7.21067
R9922 VDPWR.n2257 VDPWR.n2255 7.21067
R9923 VDPWR.n2301 VDPWR.n2300 7.17134
R9924 VDPWR.n1662 VDPWR.n1458 7.12524
R9925 VDPWR.n536 VDPWR.n531 7.10511
R9926 VDPWR.n2327 VDPWR.n2326 7.03001
R9927 VDPWR.n545 VDPWR.n542 6.8005
R9928 VDPWR.n265 VDPWR.n262 6.8005
R9929 VDPWR.n8 VDPWR.n5 6.8005
R9930 VDPWR.n1762 VDPWR.n1409 6.77697
R9931 VDPWR.n2105 VDPWR.n2016 6.77697
R9932 VDPWR.n2926 VDPWR.n2925 6.77697
R9933 VDPWR.n855 VDPWR.n854 6.73838
R9934 VDPWR.t285 VDPWR.t760 6.71428
R9935 VDPWR.t675 VDPWR.t13 6.71428
R9936 VDPWR.t88 VDPWR.t586 6.71428
R9937 VDPWR.t375 VDPWR.t373 6.71428
R9938 VDPWR.t672 VDPWR.t666 6.71428
R9939 VDPWR.n1589 VDPWR.n1485 6.66496
R9940 VDPWR.n1841 VDPWR.n1331 6.66496
R9941 VDPWR.n1789 VDPWR.n1788 6.66496
R9942 VDPWR.n1783 VDPWR.n1383 6.66496
R9943 VDPWR.n1964 VDPWR.n1963 6.66496
R9944 VDPWR.n2287 VDPWR.n2286 6.66496
R9945 VDPWR.n2720 VDPWR.n2701 6.66496
R9946 VDPWR.n1554 VDPWR.n1499 6.52104
R9947 VDPWR.n1872 VDPWR.n1871 6.52104
R9948 VDPWR.n2250 VDPWR.n2249 6.52104
R9949 VDPWR.n2157 VDPWR.n2156 6.52104
R9950 VDPWR.n1945 VDPWR.n1270 6.52104
R9951 VDPWR.n2303 VDPWR.n1241 6.50542
R9952 VDPWR.n2384 VDPWR.n2383 6.50542
R9953 VDPWR.n1842 VDPWR.n1840 6.48583
R9954 VDPWR.n2717 VDPWR.n2716 6.48583
R9955 VDPWR.n2713 VDPWR.n2712 6.46951
R9956 VDPWR.n1098 VDPWR.n1032 6.4005
R9957 VDPWR.n2712 VDPWR.n2711 6.4005
R9958 VDPWR.n748 VDPWR.n747 6.37981
R9959 VDPWR.n744 VDPWR.n742 6.37981
R9960 VDPWR.n736 VDPWR.n735 6.37981
R9961 VDPWR.n733 VDPWR.n732 6.37981
R9962 VDPWR.n2560 VDPWR.n988 6.3005
R9963 VDPWR.n719 VDPWR.n655 6.18087
R9964 VDPWR.n3115 VDPWR.n3110 6.12434
R9965 VDPWR.n713 VDPWR.n704 6.02403
R9966 VDPWR.n660 VDPWR.n657 6.02403
R9967 VDPWR.n524 VDPWR.n515 6.02403
R9968 VDPWR.n476 VDPWR.n467 6.02403
R9969 VDPWR.n412 VDPWR.n403 6.02403
R9970 VDPWR.n417 VDPWR.n414 6.02403
R9971 VDPWR.n768 VDPWR.n759 6.02403
R9972 VDPWR.n3066 VDPWR.n3057 6.02403
R9973 VDPWR.n974 VDPWR.n973 5.97436
R9974 VDPWR.n1839 VDPWR.n1838 5.8885
R9975 VDPWR.n2715 VDPWR.n2714 5.8885
R9976 VDPWR.n1014 VDPWR.n1011 5.85193
R9977 VDPWR.n3115 VDPWR.n3114 5.75618
R9978 VDPWR.n2311 VDPWR.n1226 5.66607
R9979 VDPWR.n2392 VDPWR.n2391 5.66607
R9980 VDPWR.n1595 VDPWR.n1480 5.66204
R9981 VDPWR.n1599 VDPWR.n1480 5.66204
R9982 VDPWR.n1603 VDPWR.n1601 5.66204
R9983 VDPWR.n1603 VDPWR.n1602 5.66204
R9984 VDPWR.n1602 VDPWR.n1473 5.66204
R9985 VDPWR.n1619 VDPWR.n1473 5.66204
R9986 VDPWR.n1620 VDPWR.n1619 5.66204
R9987 VDPWR.n1621 VDPWR.n1620 5.66204
R9988 VDPWR.n1628 VDPWR.n1627 5.66204
R9989 VDPWR.n1629 VDPWR.n1628 5.66204
R9990 VDPWR.n1633 VDPWR.n1632 5.66204
R9991 VDPWR.n1634 VDPWR.n1633 5.66204
R9992 VDPWR.n1634 VDPWR.n1466 5.66204
R9993 VDPWR.n1643 VDPWR.n1466 5.66204
R9994 VDPWR.n1644 VDPWR.n1643 5.66204
R9995 VDPWR.n1647 VDPWR.n1644 5.66204
R9996 VDPWR.n1557 VDPWR.n1556 5.66204
R9997 VDPWR.n1564 VDPWR.n1495 5.66204
R9998 VDPWR.n1568 VDPWR.n1495 5.66204
R9999 VDPWR.n1572 VDPWR.n1570 5.66204
R10000 VDPWR.n1572 VDPWR.n1571 5.66204
R10001 VDPWR.n1698 VDPWR.n1697 5.66204
R10002 VDPWR.n1699 VDPWR.n1698 5.66204
R10003 VDPWR.n1703 VDPWR.n1702 5.66204
R10004 VDPWR.n1704 VDPWR.n1703 5.66204
R10005 VDPWR.n1704 VDPWR.n1442 5.66204
R10006 VDPWR.n1708 VDPWR.n1442 5.66204
R10007 VDPWR.n1709 VDPWR.n1708 5.66204
R10008 VDPWR.n1711 VDPWR.n1709 5.66204
R10009 VDPWR.n1868 VDPWR.n1867 5.66204
R10010 VDPWR.n1860 VDPWR.n1859 5.66204
R10011 VDPWR.n1859 VDPWR.n1313 5.66204
R10012 VDPWR.n1327 VDPWR.n1321 5.66204
R10013 VDPWR.n1328 VDPWR.n1327 5.66204
R10014 VDPWR.n1829 VDPWR.n1828 5.66204
R10015 VDPWR.n1352 VDPWR.n1344 5.66204
R10016 VDPWR.n1353 VDPWR.n1352 5.66204
R10017 VDPWR.n1818 VDPWR.n1353 5.66204
R10018 VDPWR.n1818 VDPWR.n1817 5.66204
R10019 VDPWR.n1805 VDPWR.n1804 5.66204
R10020 VDPWR.n1801 VDPWR.n1800 5.66204
R10021 VDPWR.n1800 VDPWR.n1799 5.66204
R10022 VDPWR.n1799 VDPWR.n1359 5.66204
R10023 VDPWR.n1375 VDPWR.n1359 5.66204
R10024 VDPWR.n2129 VDPWR.n2128 5.66204
R10025 VDPWR.n2128 VDPWR.n2127 5.66204
R10026 VDPWR.n2010 VDPWR.n2004 5.66204
R10027 VDPWR.n2138 VDPWR.n2137 5.66204
R10028 VDPWR.n2137 VDPWR.n2136 5.66204
R10029 VDPWR.n1985 VDPWR.n1979 5.66204
R10030 VDPWR.n1986 VDPWR.n1985 5.66204
R10031 VDPWR.n2145 VDPWR.n2144 5.66204
R10032 VDPWR.n1955 VDPWR.n1266 5.66204
R10033 VDPWR.n1959 VDPWR.n1266 5.66204
R10034 VDPWR.n1962 VDPWR.n1961 5.66204
R10035 VDPWR.n2176 VDPWR.n1962 5.66204
R10036 VDPWR.n1948 VDPWR.n1947 5.66204
R10037 VDPWR.n2261 VDPWR.n2260 5.66204
R10038 VDPWR.n2262 VDPWR.n2261 5.66204
R10039 VDPWR.n2266 VDPWR.n2265 5.66204
R10040 VDPWR.n2266 VDPWR.n1253 5.66204
R10041 VDPWR.n2280 VDPWR.n1253 5.66204
R10042 VDPWR.n534 VDPWR 5.6325
R10043 VDPWR.n3113 VDPWR 5.6325
R10044 VDPWR.n1815 VDPWR.n1354 5.48759
R10045 VDPWR.n1835 VDPWR.n1834 5.42606
R10046 VDPWR.n1811 VDPWR.n1810 5.42606
R10047 VDPWR.n1382 VDPWR.n1381 5.3712
R10048 VDPWR.n1595 VDPWR.n1594 5.29281
R10049 VDPWR.n1621 VDPWR.n1471 5.29281
R10050 VDPWR.n1627 VDPWR.n1470 5.29281
R10051 VDPWR.n1647 VDPWR.n1646 5.29281
R10052 VDPWR.n1556 VDPWR.n1555 5.29281
R10053 VDPWR.n1557 VDPWR.n1497 5.29281
R10054 VDPWR.n1564 VDPWR.n1563 5.29281
R10055 VDPWR.n1571 VDPWR.n1486 5.29281
R10056 VDPWR.n1697 VDPWR.n1446 5.29281
R10057 VDPWR.n1711 VDPWR.n1710 5.29281
R10058 VDPWR.n1868 VDPWR.n1309 5.29281
R10059 VDPWR.n1867 VDPWR.n1866 5.29281
R10060 VDPWR.n1861 VDPWR.n1860 5.29281
R10061 VDPWR.n1329 VDPWR.n1328 5.29281
R10062 VDPWR.n1831 VDPWR.n1333 5.29281
R10063 VDPWR.n1817 VDPWR.n1816 5.29281
R10064 VDPWR.n1807 VDPWR.n1355 5.29281
R10065 VDPWR.n1376 VDPWR.n1375 5.29281
R10066 VDPWR.n2129 VDPWR.n1993 5.29281
R10067 VDPWR.n2011 VDPWR.n2010 5.29281
R10068 VDPWR.n2138 VDPWR.n1990 5.29281
R10069 VDPWR.n1979 VDPWR.n1971 5.29281
R10070 VDPWR.n2144 VDPWR.n2143 5.29281
R10071 VDPWR.n1955 VDPWR.n1954 5.29281
R10072 VDPWR.n2176 VDPWR.n2175 5.29281
R10073 VDPWR.n1947 VDPWR.n1946 5.29281
R10074 VDPWR.n1948 VDPWR.n1268 5.29281
R10075 VDPWR.n2252 VDPWR.n2251 5.29281
R10076 VDPWR.n2252 VDPWR.n2195 5.29281
R10077 VDPWR.n2281 VDPWR.n2280 5.29281
R10078 VDPWR.n1104 VDPWR.n1029 5.27109
R10079 VDPWR.n2764 VDPWR.n2673 5.27109
R10080 VDPWR.n2210 VDPWR.n2209 5.25888
R10081 VDPWR.n2309 VDPWR.n2308 5.2464
R10082 VDPWR.n2386 VDPWR.n1197 5.2464
R10083 VDPWR.n1783 VDPWR.n1782 5.18397
R10084 VDPWR.n1404 VDPWR.n1403 5.18397
R10085 VDPWR.n2342 VDPWR.n2341 5.18397
R10086 VDPWR.n2522 VDPWR.n1138 5.18397
R10087 VDPWR.n2514 VDPWR.n1141 5.18397
R10088 VDPWR.n716 VDPWR.n715 5.18145
R10089 VDPWR.n700 VDPWR.n699 5.18145
R10090 VDPWR.n684 VDPWR.n683 5.18145
R10091 VDPWR.n668 VDPWR.n667 5.18145
R10092 VDPWR.n527 VDPWR.n526 5.18145
R10093 VDPWR.n511 VDPWR.n510 5.18145
R10094 VDPWR.n495 VDPWR.n494 5.18145
R10095 VDPWR.n479 VDPWR.n478 5.18145
R10096 VDPWR.n463 VDPWR.n462 5.18145
R10097 VDPWR.n457 VDPWR.n456 5.18145
R10098 VDPWR.n441 VDPWR.n440 5.18145
R10099 VDPWR.n425 VDPWR.n424 5.18145
R10100 VDPWR.n3107 VDPWR.n3106 5.18145
R10101 VDPWR.n3101 VDPWR.n3100 5.18145
R10102 VDPWR.n3085 VDPWR.n3084 5.18145
R10103 VDPWR.n3069 VDPWR.n3068 5.18145
R10104 VDPWR.n2307 VDPWR.n2306 5.14148
R10105 VDPWR.n2550 VDPWR.n2549 5.1205
R10106 VDPWR.n2379 VDPWR.n2378 5.103
R10107 VDPWR.n2416 VDPWR.n1181 5.03657
R10108 VDPWR.t736 VDPWR.t11 5.03584
R10109 VDPWR.t283 VDPWR.t687 5.03584
R10110 VDPWR.t967 VDPWR.t471 5.03584
R10111 VDPWR.t79 VDPWR.t541 5.03584
R10112 VDPWR.t508 VDPWR.t121 5.03584
R10113 VDPWR.n850 VDPWR.n818 4.98336
R10114 VDPWR.n1107 VDPWR.n1028 4.9005
R10115 VDPWR.n698 VDPWR.n690 4.89462
R10116 VDPWR.n674 VDPWR.n672 4.89462
R10117 VDPWR.n509 VDPWR.n501 4.89462
R10118 VDPWR.n485 VDPWR.n483 4.89462
R10119 VDPWR.n455 VDPWR.n447 4.89462
R10120 VDPWR.n431 VDPWR.n429 4.89462
R10121 VDPWR.n3099 VDPWR.n3091 4.89462
R10122 VDPWR.n3075 VDPWR.n3073 4.89462
R10123 VDPWR.n3071 VDPWR.n3056 4.72727
R10124 VDPWR.n2223 VDPWR.n2222 4.69218
R10125 VDPWR.n601 VDPWR.n600 4.67352
R10126 VDPWR.n624 VDPWR.n589 4.67352
R10127 VDPWR.n321 VDPWR.n320 4.67352
R10128 VDPWR.n344 VDPWR.n309 4.67352
R10129 VDPWR.n2074 VDPWR.n2073 4.67352
R10130 VDPWR.n1123 VDPWR.n1119 4.67352
R10131 VDPWR.n2569 VDPWR.n2568 4.67352
R10132 VDPWR.n2909 VDPWR.n2908 4.67352
R10133 VDPWR.n2983 VDPWR.n2982 4.67352
R10134 VDPWR.n2982 VDPWR.n2950 4.67352
R10135 VDPWR.n2782 VDPWR.n2781 4.67352
R10136 VDPWR.n2778 VDPWR.n2777 4.67352
R10137 VDPWR.n2797 VDPWR.n2796 4.67352
R10138 VDPWR.n2754 VDPWR.n2753 4.67352
R10139 VDPWR.n3029 VDPWR.n789 4.67352
R10140 VDPWR.n3025 VDPWR.n3024 4.67352
R10141 VDPWR.n3024 VDPWR.n3023 4.67352
R10142 VDPWR.n860 VDPWR.n811 4.67352
R10143 VDPWR.n856 VDPWR.n811 4.67352
R10144 VDPWR.n856 VDPWR.n855 4.67352
R10145 VDPWR.n846 VDPWR.n845 4.67352
R10146 VDPWR.n845 VDPWR.n820 4.67352
R10147 VDPWR.n64 VDPWR.n63 4.67352
R10148 VDPWR.n87 VDPWR.n52 4.67352
R10149 VDPWR.n750 VDPWR.n749 4.6505
R10150 VDPWR.n2083 VDPWR.n2030 4.62124
R10151 VDPWR.n2896 VDPWR.n2895 4.62124
R10152 VDPWR.n1843 VDPWR.n1842 4.62124
R10153 VDPWR.n1836 VDPWR.n1332 4.62124
R10154 VDPWR.n1813 VDPWR.n1812 4.62124
R10155 VDPWR.n2219 VDPWR.n2210 4.62124
R10156 VDPWR.n2718 VDPWR.n2717 4.62124
R10157 VDPWR.n2712 VDPWR.n2702 4.62124
R10158 VDPWR.n850 VDPWR.n848 4.62124
R10159 VDPWR.n976 VDPWR.n972 4.5918
R10160 VDPWR.n2076 VDPWR.n2075 4.57193
R10161 VDPWR.n2984 VDPWR.n2983 4.57193
R10162 VDPWR.n2519 VDPWR.n1138 4.54926
R10163 VDPWR.n2517 VDPWR.n1141 4.54926
R10164 VDPWR.n1161 VDPWR.n1160 4.54926
R10165 VDPWR.n2492 VDPWR.n1161 4.54926
R10166 VDPWR.n2295 VDPWR.n2292 4.52113
R10167 VDPWR.n1101 VDPWR.n1029 4.51815
R10168 VDPWR.n2839 VDPWR.n936 4.51401
R10169 VDPWR.n2844 VDPWR.n2843 4.51401
R10170 VDPWR.n2877 VDPWR.n916 4.51401
R10171 VDPWR.n2882 VDPWR.n2881 4.51401
R10172 VDPWR.n2743 VDPWR.n2742 4.51401
R10173 VDPWR.n2691 VDPWR.n2688 4.51401
R10174 VDPWR.n1641 VDPWR.n1640 4.51401
R10175 VDPWR.n1655 VDPWR.n1654 4.51401
R10176 VDPWR.n1607 VDPWR.n1605 4.51401
R10177 VDPWR.n1617 VDPWR.n1616 4.51401
R10178 VDPWR.n1579 VDPWR.n1491 4.51401
R10179 VDPWR.n1584 VDPWR.n1583 4.51401
R10180 VDPWR.n1532 VDPWR.n1531 4.51401
R10181 VDPWR.n1545 VDPWR.n1544 4.51401
R10182 VDPWR.n1715 VDPWR.n1714 4.51401
R10183 VDPWR.n1726 VDPWR.n1433 4.51401
R10184 VDPWR.n1680 VDPWR.n1679 4.51401
R10185 VDPWR.n1691 VDPWR.n1690 4.51401
R10186 VDPWR.n1797 VDPWR.n1796 4.51401
R10187 VDPWR.n1792 VDPWR.n1791 4.51401
R10188 VDPWR.n1826 VDPWR.n1825 4.51401
R10189 VDPWR.n1821 VDPWR.n1820 4.51401
R10190 VDPWR.n1856 VDPWR.n1855 4.51401
R10191 VDPWR.n1850 VDPWR.n1849 4.51401
R10192 VDPWR.n1892 VDPWR.n1279 4.51401
R10193 VDPWR.n1883 VDPWR.n1879 4.51401
R10194 VDPWR.n1737 VDPWR.n1735 4.51401
R10195 VDPWR.n1747 VDPWR.n1746 4.51401
R10196 VDPWR.n1772 VDPWR.n1771 4.51401
R10197 VDPWR.n1767 VDPWR.n1766 4.51401
R10198 VDPWR.n2125 VDPWR.n2124 4.51401
R10199 VDPWR.n2119 VDPWR.n2118 4.51401
R10200 VDPWR.n2154 VDPWR.n2153 4.51401
R10201 VDPWR.n2148 VDPWR.n2147 4.51401
R10202 VDPWR.n2186 VDPWR.n1260 4.51401
R10203 VDPWR.n1265 VDPWR.n1264 4.51401
R10204 VDPWR.n1931 VDPWR.n1896 4.51401
R10205 VDPWR.n1936 VDPWR.n1935 4.51401
R10206 VDPWR.n2071 VDPWR.n2070 4.51401
R10207 VDPWR.n2061 VDPWR.n2060 4.51401
R10208 VDPWR.n2022 VDPWR.n2021 4.51401
R10209 VDPWR.n2087 VDPWR.n2086 4.51401
R10210 VDPWR.n1146 VDPWR.n1144 4.51401
R10211 VDPWR.n2503 VDPWR.n2502 4.51401
R10212 VDPWR.n3009 VDPWR.n870 4.51401
R10213 VDPWR.n875 VDPWR.n874 4.51401
R10214 VDPWR.n2399 VDPWR.n1194 4.51401
R10215 VDPWR.n2403 VDPWR.n1185 4.51401
R10216 VDPWR.n2317 VDPWR.n1232 4.51401
R10217 VDPWR.n2322 VDPWR.n2321 4.51401
R10218 VDPWR.n2272 VDPWR.n2190 4.51401
R10219 VDPWR.n2276 VDPWR.n1252 4.51401
R10220 VDPWR.n2228 VDPWR.n2227 4.51401
R10221 VDPWR.n2242 VDPWR.n2241 4.51401
R10222 VDPWR.n2437 VDPWR.n2436 4.51401
R10223 VDPWR.n2448 VDPWR.n1169 4.51401
R10224 VDPWR.n2357 VDPWR.n1212 4.51401
R10225 VDPWR.n2362 VDPWR.n2361 4.51401
R10226 VDPWR.n1114 VDPWR.n1113 4.51401
R10227 VDPWR.n1131 VDPWR.n1130 4.51401
R10228 VDPWR.n2913 VDPWR.n889 4.51401
R10229 VDPWR.n2918 VDPWR.n2917 4.51401
R10230 VDPWR.n2706 VDPWR.n781 4.51401
R10231 VDPWR.n784 VDPWR.n780 4.51401
R10232 VDPWR.n1041 VDPWR.n1040 4.51401
R10233 VDPWR.n1079 VDPWR.n1035 4.51401
R10234 VDPWR.n1004 VDPWR.n1002 4.51401
R10235 VDPWR.n2537 VDPWR.n2536 4.51401
R10236 VDPWR.n2482 VDPWR.n2481 4.51401
R10237 VDPWR.n2472 VDPWR.n2471 4.51401
R10238 VDPWR.n2580 VDPWR.n957 4.51401
R10239 VDPWR.n2572 VDPWR.n2571 4.51401
R10240 VDPWR.n2610 VDPWR.n2585 4.51401
R10241 VDPWR.n2805 VDPWR.n951 4.51401
R10242 VDPWR.n2979 VDPWR.n2978 4.51401
R10243 VDPWR.n2973 VDPWR.n2972 4.51401
R10244 VDPWR.n2665 VDPWR.n2664 4.51401
R10245 VDPWR.n2670 VDPWR.n2667 4.51401
R10246 VDPWR.n2626 VDPWR.n2617 4.51401
R10247 VDPWR.n2800 VDPWR.n2799 4.51401
R10248 VDPWR.n842 VDPWR.n841 4.51401
R10249 VDPWR.n835 VDPWR.n771 4.51401
R10250 VDPWR.n3016 VDPWR.n3015 4.51401
R10251 VDPWR.n802 VDPWR.n800 4.51401
R10252 VDPWR.n2308 VDPWR.n2307 4.51198
R10253 VDPWR.n2420 VDPWR.n1181 4.51198
R10254 VDPWR.n536 VDPWR.n535 4.5005
R10255 VDPWR.n1718 VDPWR.n1717 4.5005
R10256 VDPWR.n1719 VDPWR.n1435 4.5005
R10257 VDPWR.n1728 VDPWR.n1727 4.5005
R10258 VDPWR.n1529 VDPWR.n1528 4.5005
R10259 VDPWR.n1540 VDPWR.n1539 4.5005
R10260 VDPWR.n1503 VDPWR.n1502 4.5005
R10261 VDPWR.n1578 VDPWR.n1577 4.5005
R10262 VDPWR.n1576 VDPWR.n1575 4.5005
R10263 VDPWR.n1494 VDPWR.n1488 4.5005
R10264 VDPWR.n1609 VDPWR.n1608 4.5005
R10265 VDPWR.n1612 VDPWR.n1611 4.5005
R10266 VDPWR.n1475 VDPWR.n1474 4.5005
R10267 VDPWR.n1638 VDPWR.n1637 4.5005
R10268 VDPWR.n1650 VDPWR.n1649 4.5005
R10269 VDPWR.n1465 VDPWR.n1461 4.5005
R10270 VDPWR.n1677 VDPWR.n1452 4.5005
R10271 VDPWR.n1686 VDPWR.n1685 4.5005
R10272 VDPWR.n1449 VDPWR.n1448 4.5005
R10273 VDPWR.n1739 VDPWR.n1738 4.5005
R10274 VDPWR.n1742 VDPWR.n1741 4.5005
R10275 VDPWR.n1431 VDPWR.n1430 4.5005
R10276 VDPWR.n1891 VDPWR.n1890 4.5005
R10277 VDPWR.n1880 VDPWR.n1281 4.5005
R10278 VDPWR.n1885 VDPWR.n1884 4.5005
R10279 VDPWR.n1322 VDPWR.n1315 4.5005
R10280 VDPWR.n1324 VDPWR.n1323 4.5005
R10281 VDPWR.n1325 VDPWR.n1318 4.5005
R10282 VDPWR.n1345 VDPWR.n1337 4.5005
R10283 VDPWR.n1350 VDPWR.n1349 4.5005
R10284 VDPWR.n1346 VDPWR.n1341 4.5005
R10285 VDPWR.n1361 VDPWR.n1360 4.5005
R10286 VDPWR.n1372 VDPWR.n1371 4.5005
R10287 VDPWR.n1373 VDPWR.n1365 4.5005
R10288 VDPWR.n1397 VDPWR.n1390 4.5005
R10289 VDPWR.n1401 VDPWR.n1400 4.5005
R10290 VDPWR.n1406 VDPWR.n1394 4.5005
R10291 VDPWR.n2048 VDPWR.n2045 4.5005
R10292 VDPWR.n2066 VDPWR.n2065 4.5005
R10293 VDPWR.n2058 VDPWR.n2050 4.5005
R10294 VDPWR.n1930 VDPWR.n1929 4.5005
R10295 VDPWR.n1900 VDPWR.n1899 4.5005
R10296 VDPWR.n1274 VDPWR.n1273 4.5005
R10297 VDPWR.n2185 VDPWR.n2184 4.5005
R10298 VDPWR.n2183 VDPWR.n2182 4.5005
R10299 VDPWR.n2179 VDPWR.n2178 4.5005
R10300 VDPWR.n1980 VDPWR.n1973 4.5005
R10301 VDPWR.n1983 VDPWR.n1982 4.5005
R10302 VDPWR.n1981 VDPWR.n1976 4.5005
R10303 VDPWR.n1997 VDPWR.n1996 4.5005
R10304 VDPWR.n2007 VDPWR.n2006 4.5005
R10305 VDPWR.n2008 VDPWR.n2000 4.5005
R10306 VDPWR.n2094 VDPWR.n2093 4.5005
R10307 VDPWR.n2026 VDPWR.n2023 4.5005
R10308 VDPWR.n2028 VDPWR.n2025 4.5005
R10309 VDPWR.n2440 VDPWR.n2439 4.5005
R10310 VDPWR.n2441 VDPWR.n1171 4.5005
R10311 VDPWR.n2450 VDPWR.n2449 4.5005
R10312 VDPWR.n2225 VDPWR.n2204 4.5005
R10313 VDPWR.n2237 VDPWR.n2236 4.5005
R10314 VDPWR.n2201 VDPWR.n2200 4.5005
R10315 VDPWR.n2271 VDPWR.n2270 4.5005
R10316 VDPWR.n2269 VDPWR.n2268 4.5005
R10317 VDPWR.n2278 VDPWR.n2277 4.5005
R10318 VDPWR.n2316 VDPWR.n2315 4.5005
R10319 VDPWR.n1238 VDPWR.n1237 4.5005
R10320 VDPWR.n1235 VDPWR.n1228 4.5005
R10321 VDPWR.n2398 VDPWR.n2397 4.5005
R10322 VDPWR.n2396 VDPWR.n2395 4.5005
R10323 VDPWR.n2405 VDPWR.n2404 4.5005
R10324 VDPWR.n2356 VDPWR.n2355 4.5005
R10325 VDPWR.n1216 VDPWR.n1215 4.5005
R10326 VDPWR.n1208 VDPWR.n1207 4.5005
R10327 VDPWR.n2458 VDPWR.n1166 4.5005
R10328 VDPWR.n2477 VDPWR.n2476 4.5005
R10329 VDPWR.n2469 VDPWR.n2460 4.5005
R10330 VDPWR.n2544 VDPWR.n2543 4.5005
R10331 VDPWR.n1005 VDPWR.n1003 4.5005
R10332 VDPWR.n1012 VDPWR.n1007 4.5005
R10333 VDPWR.n1072 VDPWR.n1071 4.5005
R10334 VDPWR.n1073 VDPWR.n1037 4.5005
R10335 VDPWR.n1081 VDPWR.n1080 4.5005
R10336 VDPWR.n1111 VDPWR.n1110 4.5005
R10337 VDPWR.n1126 VDPWR.n1125 4.5005
R10338 VDPWR.n1027 VDPWR.n1023 4.5005
R10339 VDPWR.n2510 VDPWR.n2509 4.5005
R10340 VDPWR.n1147 VDPWR.n1145 4.5005
R10341 VDPWR.n1153 VDPWR.n1149 4.5005
R10342 VDPWR.n2579 VDPWR.n2578 4.5005
R10343 VDPWR.n980 VDPWR.n959 4.5005
R10344 VDPWR.n2574 VDPWR.n2573 4.5005
R10345 VDPWR.n2609 VDPWR.n2608 4.5005
R10346 VDPWR.n2586 VDPWR.n950 4.5005
R10347 VDPWR.n2807 VDPWR.n2806 4.5005
R10348 VDPWR.n2838 VDPWR.n2837 4.5005
R10349 VDPWR.n2836 VDPWR.n2835 4.5005
R10350 VDPWR.n2832 VDPWR.n931 4.5005
R10351 VDPWR.n2876 VDPWR.n2875 4.5005
R10352 VDPWR.n2873 VDPWR.n2872 4.5005
R10353 VDPWR.n911 VDPWR.n910 4.5005
R10354 VDPWR.n2912 VDPWR.n2911 4.5005
R10355 VDPWR.n893 VDPWR.n892 4.5005
R10356 VDPWR.n2906 VDPWR.n885 4.5005
R10357 VDPWR.n3008 VDPWR.n3007 4.5005
R10358 VDPWR.n3006 VDPWR.n3005 4.5005
R10359 VDPWR.n3002 VDPWR.n3001 4.5005
R10360 VDPWR.n2962 VDPWR.n2952 4.5005
R10361 VDPWR.n2965 VDPWR.n2964 4.5005
R10362 VDPWR.n2956 VDPWR.n2955 4.5005
R10363 VDPWR.n840 VDPWR.n839 4.5005
R10364 VDPWR.n823 VDPWR.n822 4.5005
R10365 VDPWR.n834 VDPWR.n833 4.5005
R10366 VDPWR.n2624 VDPWR.n2623 4.5005
R10367 VDPWR.n2650 VDPWR.n2649 4.5005
R10368 VDPWR.n2620 VDPWR.n2619 4.5005
R10369 VDPWR.n2772 VDPWR.n2771 4.5005
R10370 VDPWR.n2668 VDPWR.n2666 4.5005
R10371 VDPWR.n2767 VDPWR.n2766 4.5005
R10372 VDPWR.n2689 VDPWR.n2686 4.5005
R10373 VDPWR.n2739 VDPWR.n2738 4.5005
R10374 VDPWR.n2737 VDPWR.n2736 4.5005
R10375 VDPWR.n2708 VDPWR.n2707 4.5005
R10376 VDPWR.n2709 VDPWR.n782 4.5005
R10377 VDPWR.n3040 VDPWR.n3039 4.5005
R10378 VDPWR.n805 VDPWR.n798 4.5005
R10379 VDPWR.n806 VDPWR.n801 4.5005
R10380 VDPWR.n865 VDPWR.n864 4.5005
R10381 VDPWR.n2164 VDPWR.n1967 4.49637
R10382 VDPWR.n2313 VDPWR.n2309 4.40706
R10383 VDPWR.n2389 VDPWR.n1197 4.40706
R10384 VDPWR.n758 VDPWR.n757 4.38372
R10385 VDPWR.n600 VDPWR.n599 4.36875
R10386 VDPWR.n624 VDPWR.n623 4.36875
R10387 VDPWR.n583 VDPWR.n582 4.36875
R10388 VDPWR.n553 VDPWR.n552 4.36875
R10389 VDPWR.n320 VDPWR.n319 4.36875
R10390 VDPWR.n344 VDPWR.n343 4.36875
R10391 VDPWR.n303 VDPWR.n302 4.36875
R10392 VDPWR.n273 VDPWR.n272 4.36875
R10393 VDPWR.n2073 VDPWR.n2043 4.36875
R10394 VDPWR.n2295 VDPWR.n2294 4.36875
R10395 VDPWR.n2568 VDPWR.n986 4.36875
R10396 VDPWR.n2985 VDPWR.n2947 4.36875
R10397 VDPWR.n2957 VDPWR.n2950 4.36875
R10398 VDPWR.n2782 VDPWR.n2659 4.36875
R10399 VDPWR.n2778 VDPWR.n2660 4.36875
R10400 VDPWR.n2796 VDPWR.n2795 4.36875
R10401 VDPWR.n2758 VDPWR.n2757 4.36875
R10402 VDPWR.n2754 VDPWR.n2676 4.36875
R10403 VDPWR.n2751 VDPWR.n2679 4.36875
R10404 VDPWR.n3032 VDPWR.n788 4.36875
R10405 VDPWR.n861 VDPWR.n860 4.36875
R10406 VDPWR.n824 VDPWR.n820 4.36875
R10407 VDPWR.n63 VDPWR.n62 4.36875
R10408 VDPWR.n87 VDPWR.n86 4.36875
R10409 VDPWR.n46 VDPWR.n45 4.36875
R10410 VDPWR.n16 VDPWR.n15 4.36875
R10411 VDPWR.n1782 VDPWR.n1781 4.33769
R10412 VDPWR.n2208 VDPWR.n2207 4.29023
R10413 VDPWR.n1122 VDPWR.n1121 4.26717
R10414 VDPWR.n2083 VDPWR.n2081 4.14168
R10415 VDPWR.n3110 VDPWR.n3109 4.06613
R10416 VDPWR.n719 VDPWR.n718 4.05291
R10417 VDPWR.n1592 VDPWR.n1484 4.02033
R10418 VDPWR.n1515 VDPWR.n1511 4.02033
R10419 VDPWR.n1515 VDPWR.n1514 4.02033
R10420 VDPWR.n1524 VDPWR.n1518 4.02033
R10421 VDPWR.n1524 VDPWR.n1523 4.02033
R10422 VDPWR.n1724 VDPWR.n1440 4.02033
R10423 VDPWR.n1724 VDPWR.n1723 4.02033
R10424 VDPWR.n1290 VDPWR.n1286 4.02033
R10425 VDPWR.n1290 VDPWR.n1289 4.02033
R10426 VDPWR.n1299 VDPWR.n1293 4.02033
R10427 VDPWR.n1299 VDPWR.n1298 4.02033
R10428 VDPWR.n1749 VDPWR.n1424 4.02033
R10429 VDPWR.n1749 VDPWR.n1429 4.02033
R10430 VDPWR.n2164 VDPWR.n1965 4.02033
R10431 VDPWR.n1921 VDPWR.n1906 4.02033
R10432 VDPWR.n1921 VDPWR.n1912 4.02033
R10433 VDPWR.n1920 VDPWR.n1915 4.02033
R10434 VDPWR.n1920 VDPWR.n1919 4.02033
R10435 VDPWR.n2063 VDPWR.n2054 4.02033
R10436 VDPWR.n2063 VDPWR.n2057 4.02033
R10437 VDPWR.n2217 VDPWR.n2213 4.02033
R10438 VDPWR.n2217 VDPWR.n2216 4.02033
R10439 VDPWR.n2446 VDPWR.n1176 4.02033
R10440 VDPWR.n2446 VDPWR.n2445 4.02033
R10441 VDPWR.n968 VDPWR.n964 4.02033
R10442 VDPWR.n968 VDPWR.n967 4.02033
R10443 VDPWR.n2474 VDPWR.n2465 4.02033
R10444 VDPWR.n2474 VDPWR.n2468 4.02033
R10445 VDPWR.n2601 VDPWR.n2597 4.02033
R10446 VDPWR.n2601 VDPWR.n2600 4.02033
R10447 VDPWR.n929 VDPWR.n927 4.02033
R10448 VDPWR.n2924 VDPWR.n2923 4.02033
R10449 VDPWR.n2970 VDPWR.n2961 4.02033
R10450 VDPWR.n2970 VDPWR.n2969 4.02033
R10451 VDPWR.n2637 VDPWR.n2633 4.02033
R10452 VDPWR.n2637 VDPWR.n2636 4.02033
R10453 VDPWR.n837 VDPWR.n828 4.02033
R10454 VDPWR.n837 VDPWR.n832 4.02033
R10455 VDPWR.n2312 VDPWR.n2311 3.98739
R10456 VDPWR.n2393 VDPWR.n2392 3.98739
R10457 VDPWR.n1403 VDPWR.n1396 3.91455
R10458 VDPWR.n2752 VDPWR.n2751 3.86082
R10459 VDPWR.n1836 VDPWR.n1835 3.78037
R10460 VDPWR.n1812 VDPWR.n1811 3.78037
R10461 VDPWR.n1842 VDPWR.n1841 3.75517
R10462 VDPWR.n1380 VDPWR.n1379 3.75222
R10463 VDPWR.n1812 VDPWR.n1354 3.69446
R10464 VDPWR.n2717 VDPWR.n2701 3.66983
R10465 VDPWR.n723 VDPWR.t485 3.61217
R10466 VDPWR.n723 VDPWR.t481 3.61217
R10467 VDPWR.n725 VDPWR.t469 3.61217
R10468 VDPWR.n725 VDPWR.t46 3.61217
R10469 VDPWR.n721 VDPWR.t483 3.61217
R10470 VDPWR.n721 VDPWR.t716 3.61217
R10471 VDPWR.n2776 VDPWR.n2775 3.55606
R10472 VDPWR.n2207 VDPWR.n2206 3.53179
R10473 VDPWR.n1067 VDPWR.n1036 3.4812
R10474 VDPWR.n1537 VDPWR.n1536 3.47425
R10475 VDPWR.n1548 VDPWR.n1547 3.47425
R10476 VDPWR.n1550 VDPWR.n1548 3.47425
R10477 VDPWR.n1671 VDPWR.n1456 3.47425
R10478 VDPWR.n1672 VDPWR.n1671 3.47425
R10479 VDPWR.n1674 VDPWR.n1672 3.47425
R10480 VDPWR.n1888 VDPWR.n1887 3.47425
R10481 VDPWR.n1877 VDPWR.n1876 3.47425
R10482 VDPWR.n1876 VDPWR.n1875 3.47425
R10483 VDPWR.n2112 VDPWR.n2111 3.47425
R10484 VDPWR.n2162 VDPWR.n2161 3.47425
R10485 VDPWR.n2161 VDPWR.n1968 3.47425
R10486 VDPWR.n1927 VDPWR.n1926 3.47425
R10487 VDPWR.n1939 VDPWR.n1938 3.47425
R10488 VDPWR.n1941 VDPWR.n1939 3.47425
R10489 VDPWR.n2244 VDPWR.n2199 3.47425
R10490 VDPWR.n2245 VDPWR.n2244 3.47425
R10491 VDPWR.n2246 VDPWR.n2245 3.47425
R10492 VDPWR.n2353 VDPWR.n2352 3.47425
R10493 VDPWR.n2433 VDPWR.n2431 3.47425
R10494 VDPWR.n2487 VDPWR.n2486 3.47425
R10495 VDPWR.n2486 VDPWR.n2485 3.47425
R10496 VDPWR.n2485 VDPWR.n1164 3.47425
R10497 VDPWR.n2732 VDPWR.n2696 3.47425
R10498 VDPWR.n3116 VDPWR.n3115 3.44037
R10499 VDPWR.n2843 VDPWR.n2842 3.43925
R10500 VDPWR.n2840 VDPWR.n2839 3.43925
R10501 VDPWR.n2881 VDPWR.n2880 3.43925
R10502 VDPWR.n2878 VDPWR.n2877 3.43925
R10503 VDPWR.n1654 VDPWR.n1653 3.43925
R10504 VDPWR.n1640 VDPWR.n1639 3.43925
R10505 VDPWR.n1616 VDPWR.n1615 3.43925
R10506 VDPWR.n1607 VDPWR.n1606 3.43925
R10507 VDPWR.n1583 VDPWR.n1582 3.43925
R10508 VDPWR.n1580 VDPWR.n1579 3.43925
R10509 VDPWR.n1544 VDPWR.n1543 3.43925
R10510 VDPWR.n1531 VDPWR.n1530 3.43925
R10511 VDPWR.n1731 VDPWR.n1433 3.43925
R10512 VDPWR.n1715 VDPWR.n1432 3.43925
R10513 VDPWR.n1690 VDPWR.n1689 3.43925
R10514 VDPWR.n1679 VDPWR.n1678 3.43925
R10515 VDPWR.n1793 VDPWR.n1792 3.43925
R10516 VDPWR.n1796 VDPWR.n1795 3.43925
R10517 VDPWR.n1822 VDPWR.n1821 3.43925
R10518 VDPWR.n1825 VDPWR.n1824 3.43925
R10519 VDPWR.n1851 VDPWR.n1850 3.43925
R10520 VDPWR.n1855 VDPWR.n1854 3.43925
R10521 VDPWR.n1883 VDPWR.n1277 3.43925
R10522 VDPWR.n1893 VDPWR.n1892 3.43925
R10523 VDPWR.n1746 VDPWR.n1745 3.43925
R10524 VDPWR.n1737 VDPWR.n1736 3.43925
R10525 VDPWR.n1768 VDPWR.n1767 3.43925
R10526 VDPWR.n1771 VDPWR.n1770 3.43925
R10527 VDPWR.n2120 VDPWR.n2119 3.43925
R10528 VDPWR.n2124 VDPWR.n2123 3.43925
R10529 VDPWR.n2149 VDPWR.n2148 3.43925
R10530 VDPWR.n2153 VDPWR.n2152 3.43925
R10531 VDPWR.n1264 VDPWR.n1258 3.43925
R10532 VDPWR.n2187 VDPWR.n2186 3.43925
R10533 VDPWR.n1935 VDPWR.n1934 3.43925
R10534 VDPWR.n1932 VDPWR.n1931 3.43925
R10535 VDPWR.n2060 VDPWR.n2059 3.43925
R10536 VDPWR.n2070 VDPWR.n2069 3.43925
R10537 VDPWR.n2088 VDPWR.n2087 3.43925
R10538 VDPWR.n2090 VDPWR.n2022 3.43925
R10539 VDPWR.n2504 VDPWR.n2503 3.43925
R10540 VDPWR.n2506 VDPWR.n1146 3.43925
R10541 VDPWR.n874 VDPWR.n868 3.43925
R10542 VDPWR.n3010 VDPWR.n3009 3.43925
R10543 VDPWR.n2321 VDPWR.n2320 3.43925
R10544 VDPWR.n2318 VDPWR.n2317 3.43925
R10545 VDPWR.n2276 VDPWR.n2275 3.43925
R10546 VDPWR.n2273 VDPWR.n2272 3.43925
R10547 VDPWR.n2241 VDPWR.n2240 3.43925
R10548 VDPWR.n2227 VDPWR.n2226 3.43925
R10549 VDPWR.n2453 VDPWR.n1169 3.43925
R10550 VDPWR.n2437 VDPWR.n1168 3.43925
R10551 VDPWR.n2361 VDPWR.n2360 3.43925
R10552 VDPWR.n2358 VDPWR.n2357 3.43925
R10553 VDPWR.n1130 VDPWR.n1129 3.43925
R10554 VDPWR.n1113 VDPWR.n1112 3.43925
R10555 VDPWR.n2917 VDPWR.n2916 3.43925
R10556 VDPWR.n2914 VDPWR.n2913 3.43925
R10557 VDPWR.n2538 VDPWR.n2537 3.43925
R10558 VDPWR.n2540 VDPWR.n1004 3.43925
R10559 VDPWR.n2471 VDPWR.n2470 3.43925
R10560 VDPWR.n2481 VDPWR.n2480 3.43925
R10561 VDPWR.n2572 VDPWR.n955 3.43925
R10562 VDPWR.n2581 VDPWR.n2580 3.43925
R10563 VDPWR.n2974 VDPWR.n2973 3.43925
R10564 VDPWR.n2978 VDPWR.n2977 3.43925
R10565 VDPWR.n2733 VDPWR.n2732 3.43649
R10566 VDPWR.n655 VDPWR.n654 3.4105
R10567 VDPWR.n937 VDPWR.n935 3.4105
R10568 VDPWR.n2834 VDPWR.n932 3.4105
R10569 VDPWR.n917 VDPWR.n915 3.4105
R10570 VDPWR.n2871 VDPWR.n912 3.4105
R10571 VDPWR.n1463 VDPWR.n1462 3.4105
R10572 VDPWR.n1652 VDPWR.n1651 3.4105
R10573 VDPWR.n1477 VDPWR.n1476 3.4105
R10574 VDPWR.n1614 VDPWR.n1613 3.4105
R10575 VDPWR.n1492 VDPWR.n1490 3.4105
R10576 VDPWR.n1574 VDPWR.n1489 3.4105
R10577 VDPWR.n1505 VDPWR.n1504 3.4105
R10578 VDPWR.n1542 VDPWR.n1541 3.4105
R10579 VDPWR.n1716 VDPWR.n1434 3.4105
R10580 VDPWR.n1730 VDPWR.n1729 3.4105
R10581 VDPWR.n1451 VDPWR.n1450 3.4105
R10582 VDPWR.n1688 VDPWR.n1687 3.4105
R10583 VDPWR.n1369 VDPWR.n1362 3.4105
R10584 VDPWR.n1370 VDPWR.n1364 3.4105
R10585 VDPWR.n1347 VDPWR.n1338 3.4105
R10586 VDPWR.n1348 VDPWR.n1340 3.4105
R10587 VDPWR.n1853 VDPWR.n1316 3.4105
R10588 VDPWR.n1852 VDPWR.n1317 3.4105
R10589 VDPWR.n1280 VDPWR.n1278 3.4105
R10590 VDPWR.n1882 VDPWR.n1881 3.4105
R10591 VDPWR.n1740 VDPWR.n1734 3.4105
R10592 VDPWR.n1744 VDPWR.n1743 3.4105
R10593 VDPWR.n1398 VDPWR.n1391 3.4105
R10594 VDPWR.n1399 VDPWR.n1393 3.4105
R10595 VDPWR.n2122 VDPWR.n1998 3.4105
R10596 VDPWR.n2121 VDPWR.n1999 3.4105
R10597 VDPWR.n2151 VDPWR.n1974 3.4105
R10598 VDPWR.n2150 VDPWR.n1975 3.4105
R10599 VDPWR.n1261 VDPWR.n1259 3.4105
R10600 VDPWR.n2181 VDPWR.n2180 3.4105
R10601 VDPWR.n1897 VDPWR.n1895 3.4105
R10602 VDPWR.n1898 VDPWR.n1275 3.4105
R10603 VDPWR.n2068 VDPWR.n2067 3.4105
R10604 VDPWR.n2047 VDPWR.n2046 3.4105
R10605 VDPWR.n2092 VDPWR.n2091 3.4105
R10606 VDPWR.n2089 VDPWR.n2024 3.4105
R10607 VDPWR.n2508 VDPWR.n2507 3.4105
R10608 VDPWR.n2505 VDPWR.n1148 3.4105
R10609 VDPWR.n871 VDPWR.n869 3.4105
R10610 VDPWR.n3004 VDPWR.n3003 3.4105
R10611 VDPWR.n2402 VDPWR.n2401 3.4105
R10612 VDPWR.n2401 VDPWR.n2400 3.4105
R10613 VDPWR.n2403 VDPWR.n2402 3.4105
R10614 VDPWR.n2400 VDPWR.n2399 3.4105
R10615 VDPWR.n1195 VDPWR.n1193 3.4105
R10616 VDPWR.n1190 VDPWR.n1189 3.4105
R10617 VDPWR.n1233 VDPWR.n1231 3.4105
R10618 VDPWR.n1236 VDPWR.n1229 3.4105
R10619 VDPWR.n2191 VDPWR.n2189 3.4105
R10620 VDPWR.n1256 VDPWR.n1255 3.4105
R10621 VDPWR.n2203 VDPWR.n2202 3.4105
R10622 VDPWR.n2239 VDPWR.n2238 3.4105
R10623 VDPWR.n2438 VDPWR.n1170 3.4105
R10624 VDPWR.n2452 VDPWR.n2451 3.4105
R10625 VDPWR.n1213 VDPWR.n1211 3.4105
R10626 VDPWR.n1214 VDPWR.n1209 3.4105
R10627 VDPWR.n1025 VDPWR.n1024 3.4105
R10628 VDPWR.n1128 VDPWR.n1127 3.4105
R10629 VDPWR.n890 VDPWR.n888 3.4105
R10630 VDPWR.n891 VDPWR.n886 3.4105
R10631 VDPWR.n3042 VDPWR.n780 3.4105
R10632 VDPWR.n3042 VDPWR.n781 3.4105
R10633 VDPWR.n3042 VDPWR.n779 3.4105
R10634 VDPWR.n3042 VDPWR.n3041 3.4105
R10635 VDPWR.n2741 VDPWR.n2688 3.4105
R10636 VDPWR.n2742 VDPWR.n2741 3.4105
R10637 VDPWR.n2741 VDPWR.n2740 3.4105
R10638 VDPWR.n2741 VDPWR.n2687 3.4105
R10639 VDPWR.n1078 VDPWR.n913 3.4105
R10640 VDPWR.n1039 VDPWR.n913 3.4105
R10641 VDPWR.n1079 VDPWR.n1078 3.4105
R10642 VDPWR.n1040 VDPWR.n1039 3.4105
R10643 VDPWR.n1075 VDPWR.n1074 3.4105
R10644 VDPWR.n1077 VDPWR.n1038 3.4105
R10645 VDPWR.n2542 VDPWR.n2541 3.4105
R10646 VDPWR.n2539 VDPWR.n1006 3.4105
R10647 VDPWR.n2479 VDPWR.n2478 3.4105
R10648 VDPWR.n2457 VDPWR.n2456 3.4105
R10649 VDPWR.n958 VDPWR.n956 3.4105
R10650 VDPWR.n982 VDPWR.n981 3.4105
R10651 VDPWR.n2804 VDPWR.n2803 3.4105
R10652 VDPWR.n2803 VDPWR.n2611 3.4105
R10653 VDPWR.n2805 VDPWR.n2804 3.4105
R10654 VDPWR.n2611 VDPWR.n2610 3.4105
R10655 VDPWR.n2587 VDPWR.n2584 3.4105
R10656 VDPWR.n953 VDPWR.n952 3.4105
R10657 VDPWR.n2976 VDPWR.n2953 3.4105
R10658 VDPWR.n2975 VDPWR.n2954 3.4105
R10659 VDPWR.n2769 VDPWR.n2667 3.4105
R10660 VDPWR.n2769 VDPWR.n2665 3.4105
R10661 VDPWR.n2770 VDPWR.n2769 3.4105
R10662 VDPWR.n2769 VDPWR.n2768 3.4105
R10663 VDPWR.n2801 VDPWR.n2800 3.4105
R10664 VDPWR.n2801 VDPWR.n2617 3.4105
R10665 VDPWR.n2801 VDPWR.n2616 3.4105
R10666 VDPWR.n2801 VDPWR.n2615 3.4105
R10667 VDPWR.n3014 VDPWR.n800 3.4105
R10668 VDPWR.n3015 VDPWR.n3014 3.4105
R10669 VDPWR.n3014 VDPWR.n799 3.4105
R10670 VDPWR.n3014 VDPWR.n866 3.4105
R10671 VDPWR.n3050 VDPWR.n770 3.4105
R10672 VDPWR.n841 VDPWR.n770 3.4105
R10673 VDPWR.n3051 VDPWR.n772 3.4105
R10674 VDPWR.n3051 VDPWR.n773 3.4105
R10675 VDPWR.n3051 VDPWR.n771 3.4105
R10676 VDPWR.t533 VDPWR.t416 3.35739
R10677 VDPWR.t737 VDPWR.t655 3.35739
R10678 VDPWR.t131 VDPWR.t103 3.35739
R10679 VDPWR.t340 VDPWR.t344 3.35739
R10680 VDPWR.t607 VDPWR.t444 3.35739
R10681 VDPWR.t0 VDPWR.t209 3.35739
R10682 VDPWR.t822 VDPWR.t400 3.35739
R10683 VDPWR.t126 VDPWR.t1042 3.35739
R10684 VDPWR.t590 VDPWR.t418 3.35739
R10685 VDPWR.t197 VDPWR.t609 3.35739
R10686 VDPWR.n1534 VDPWR.n1508 3.2477
R10687 VDPWR.n1550 VDPWR.n1549 3.2477
R10688 VDPWR.n1664 VDPWR.n1663 3.2477
R10689 VDPWR.n1674 VDPWR.n1673 3.2477
R10690 VDPWR.n1304 VDPWR.n1283 3.2477
R10691 VDPWR.n1875 VDPWR.n1308 3.2477
R10692 VDPWR.n2111 VDPWR.n2110 3.2477
R10693 VDPWR.n2163 VDPWR.n2162 3.2477
R10694 VDPWR.n1902 VDPWR.n1901 3.2477
R10695 VDPWR.n1941 VDPWR.n1940 3.2477
R10696 VDPWR.n2230 VDPWR.n2205 3.2477
R10697 VDPWR.n2246 VDPWR.n2197 3.2477
R10698 VDPWR.n2352 VDPWR.n1206 3.2477
R10699 VDPWR.n2433 VDPWR.n2432 3.2477
R10700 VDPWR.n2487 VDPWR.n1162 3.2477
R10701 VDPWR.n2461 VDPWR.n1164 3.2477
R10702 VDPWR.n2734 VDPWR.n2692 3.2477
R10703 VDPWR.n2728 VDPWR.n2727 3.2477
R10704 VDPWR.n477 VDPWR.n466 3.24308
R10705 VDPWR.n3067 VDPWR.n3056 3.24308
R10706 VDPWR.n690 VDPWR.n687 3.23917
R10707 VDPWR.n501 VDPWR.n498 3.23917
R10708 VDPWR.n447 VDPWR.n444 3.23917
R10709 VDPWR.n3091 VDPWR.n3088 3.23917
R10710 VDPWR.n674 VDPWR.n671 3.23136
R10711 VDPWR.n485 VDPWR.n482 3.23136
R10712 VDPWR.n431 VDPWR.n428 3.23136
R10713 VDPWR.n3075 VDPWR.n3072 3.23136
R10714 VDPWR.n461 VDPWR.n460 3.22655
R10715 VDPWR.n714 VDPWR.n703 3.22655
R10716 VDPWR.n525 VDPWR.n514 3.22655
R10717 VDPWR.n3105 VDPWR.n3104 3.22655
R10718 VDPWR.n2569 VDPWR.n984 3.2005
R10719 VDPWR.n1838 VDPWR.n1837 3.151
R10720 VDPWR.n2306 VDPWR.n1241 3.14804
R10721 VDPWR.n2385 VDPWR.n2384 3.14804
R10722 VDPWR.n856 VDPWR.n815 3.12116
R10723 VDPWR.n1519 VDPWR.n1515 3.05586
R10724 VDPWR.n1294 VDPWR.n1290 3.05586
R10725 VDPWR.n1920 VDPWR.n1916 3.05586
R10726 VDPWR.n2218 VDPWR.n2217 3.05586
R10727 VDPWR.n969 VDPWR.n968 3.05586
R10728 VDPWR.n2602 VDPWR.n2601 3.05586
R10729 VDPWR.n2638 VDPWR.n2637 3.05586
R10730 VDPWR.n1524 VDPWR.n1520 3.04861
R10731 VDPWR.n1299 VDPWR.n1295 3.04861
R10732 VDPWR.n1750 VDPWR.n1418 3.04861
R10733 VDPWR.n1921 VDPWR.n1909 3.04861
R10734 VDPWR.n2924 VDPWR.n2920 3.04861
R10735 VDPWR.n1592 VDPWR.n1591 3.04861
R10736 VDPWR.n1785 VDPWR.n1382 3.04861
R10737 VDPWR.n2171 VDPWR.n1965 3.04861
R10738 VDPWR.n2079 VDPWR.n2037 3.04861
R10739 VDPWR.n2576 VDPWR.n979 3.04861
R10740 VDPWR.n1600 VDPWR.n1599 3.01588
R10741 VDPWR.n1629 VDPWR.n1468 3.01588
R10742 VDPWR.n1569 VDPWR.n1568 3.01588
R10743 VDPWR.n1699 VDPWR.n1444 3.01588
R10744 VDPWR.n1320 VDPWR.n1313 3.01588
R10745 VDPWR.n1831 VDPWR.n1830 3.01588
R10746 VDPWR.n1828 VDPWR.n1335 3.01588
R10747 VDPWR.n1807 VDPWR.n1806 3.01588
R10748 VDPWR.n1804 VDPWR.n1357 3.01588
R10749 VDPWR.n2127 VDPWR.n1995 3.01588
R10750 VDPWR.n2136 VDPWR.n1991 3.01588
R10751 VDPWR.n1987 VDPWR.n1986 3.01588
R10752 VDPWR.n1960 VDPWR.n1959 3.01588
R10753 VDPWR.n2262 VDPWR.n2192 3.01588
R10754 VDPWR.n1756 VDPWR.n1755 3.01226
R10755 VDPWR.n1100 VDPWR.n1099 3.01226
R10756 VDPWR.n2854 VDPWR.n2853 3.01226
R10757 VDPWR.n2606 VDPWR.n949 3.01226
R10758 VDPWR.n2927 VDPWR.n880 3.01226
R10759 VDPWR.n2934 VDPWR.n2933 3.01226
R10760 VDPWR.n2076 VDPWR.n2041 2.99733
R10761 VDPWR.n846 VDPWR.n818 2.99733
R10762 VDPWR.n1750 VDPWR.n1416 2.91308
R10763 VDPWR.n1750 VDPWR.n1421 2.91308
R10764 VDPWR.n2594 VDPWR.n2590 2.91308
R10765 VDPWR.n2594 VDPWR.n2593 2.91308
R10766 VDPWR.n2039 VDPWR.n2037 2.87861
R10767 VDPWR.n2343 VDPWR.n2342 2.8567
R10768 VDPWR.n708 VDPWR.n707 2.84665
R10769 VDPWR.n711 VDPWR.n707 2.84665
R10770 VDPWR.n706 VDPWR.n705 2.84665
R10771 VDPWR.n711 VDPWR.n706 2.84665
R10772 VDPWR.n693 VDPWR.n692 2.84665
R10773 VDPWR.n696 VDPWR.n692 2.84665
R10774 VDPWR.n691 VDPWR.n689 2.84665
R10775 VDPWR.n696 VDPWR.n691 2.84665
R10776 VDPWR.n677 VDPWR.n676 2.84665
R10777 VDPWR.n680 VDPWR.n676 2.84665
R10778 VDPWR.n675 VDPWR.n673 2.84665
R10779 VDPWR.n680 VDPWR.n675 2.84665
R10780 VDPWR.n663 VDPWR.n662 2.84665
R10781 VDPWR.n664 VDPWR.n663 2.84665
R10782 VDPWR.n666 VDPWR.n665 2.84665
R10783 VDPWR.n665 VDPWR.n664 2.84665
R10784 VDPWR.n519 VDPWR.n518 2.84665
R10785 VDPWR.n522 VDPWR.n518 2.84665
R10786 VDPWR.n517 VDPWR.n516 2.84665
R10787 VDPWR.n522 VDPWR.n517 2.84665
R10788 VDPWR.n504 VDPWR.n503 2.84665
R10789 VDPWR.n507 VDPWR.n503 2.84665
R10790 VDPWR.n502 VDPWR.n500 2.84665
R10791 VDPWR.n507 VDPWR.n502 2.84665
R10792 VDPWR.n488 VDPWR.n487 2.84665
R10793 VDPWR.n491 VDPWR.n487 2.84665
R10794 VDPWR.n486 VDPWR.n484 2.84665
R10795 VDPWR.n491 VDPWR.n486 2.84665
R10796 VDPWR.n471 VDPWR.n470 2.84665
R10797 VDPWR.n474 VDPWR.n470 2.84665
R10798 VDPWR.n469 VDPWR.n468 2.84665
R10799 VDPWR.n474 VDPWR.n469 2.84665
R10800 VDPWR.n405 VDPWR.n404 2.84665
R10801 VDPWR.n410 VDPWR.n405 2.84665
R10802 VDPWR.n407 VDPWR.n406 2.84665
R10803 VDPWR.n410 VDPWR.n406 2.84665
R10804 VDPWR.n385 VDPWR.n384 2.84665
R10805 VDPWR.n381 VDPWR.n377 2.84665
R10806 VDPWR.n397 VDPWR.n396 2.84665
R10807 VDPWR.n393 VDPWR.n389 2.84665
R10808 VDPWR.n450 VDPWR.n449 2.84665
R10809 VDPWR.n453 VDPWR.n449 2.84665
R10810 VDPWR.n448 VDPWR.n446 2.84665
R10811 VDPWR.n453 VDPWR.n448 2.84665
R10812 VDPWR.n434 VDPWR.n433 2.84665
R10813 VDPWR.n437 VDPWR.n433 2.84665
R10814 VDPWR.n432 VDPWR.n430 2.84665
R10815 VDPWR.n437 VDPWR.n432 2.84665
R10816 VDPWR.n420 VDPWR.n419 2.84665
R10817 VDPWR.n421 VDPWR.n420 2.84665
R10818 VDPWR.n423 VDPWR.n422 2.84665
R10819 VDPWR.n422 VDPWR.n421 2.84665
R10820 VDPWR.n763 VDPWR.n762 2.84665
R10821 VDPWR.n766 VDPWR.n762 2.84665
R10822 VDPWR.n761 VDPWR.n760 2.84665
R10823 VDPWR.n766 VDPWR.n761 2.84665
R10824 VDPWR.n3092 VDPWR.n3090 2.84665
R10825 VDPWR.n3097 VDPWR.n3092 2.84665
R10826 VDPWR.n3094 VDPWR.n3093 2.84665
R10827 VDPWR.n3097 VDPWR.n3093 2.84665
R10828 VDPWR.n3076 VDPWR.n3074 2.84665
R10829 VDPWR.n3081 VDPWR.n3076 2.84665
R10830 VDPWR.n3078 VDPWR.n3077 2.84665
R10831 VDPWR.n3081 VDPWR.n3077 2.84665
R10832 VDPWR.n3061 VDPWR.n3060 2.84665
R10833 VDPWR.n3064 VDPWR.n3060 2.84665
R10834 VDPWR.n3059 VDPWR.n3058 2.84665
R10835 VDPWR.n3064 VDPWR.n3059 2.84665
R10836 VDPWR.n1840 VDPWR.n1838 2.8165
R10837 VDPWR.n2716 VDPWR.n2714 2.8165
R10838 VDPWR.n1535 VDPWR.n1507 2.6965
R10839 VDPWR.n1305 VDPWR.n1282 2.6965
R10840 VDPWR.n1924 VDPWR.n1923 2.6965
R10841 VDPWR.n2908 VDPWR.n2905 2.69256
R10842 VDPWR.n1601 VDPWR.n1600 2.64665
R10843 VDPWR.n1632 VDPWR.n1468 2.64665
R10844 VDPWR.n1570 VDPWR.n1569 2.64665
R10845 VDPWR.n1702 VDPWR.n1444 2.64665
R10846 VDPWR.n1321 VDPWR.n1320 2.64665
R10847 VDPWR.n1830 VDPWR.n1829 2.64665
R10848 VDPWR.n1344 VDPWR.n1335 2.64665
R10849 VDPWR.n1806 VDPWR.n1805 2.64665
R10850 VDPWR.n1801 VDPWR.n1357 2.64665
R10851 VDPWR.n2004 VDPWR.n1995 2.64665
R10852 VDPWR.n2145 VDPWR.n1987 2.64665
R10853 VDPWR.n1961 VDPWR.n1960 2.64665
R10854 VDPWR.n2256 VDPWR.n2194 2.64665
R10855 VDPWR.n2260 VDPWR.n2194 2.64665
R10856 VDPWR.n2265 VDPWR.n2192 2.64665
R10857 VDPWR.n2102 VDPWR.n2101 2.63579
R10858 VDPWR.n1484 VDPWR.n1482 2.63539
R10859 VDPWR.n1511 VDPWR.n1509 2.63539
R10860 VDPWR.n1514 VDPWR.n1512 2.63539
R10861 VDPWR.n1518 VDPWR.n1516 2.63539
R10862 VDPWR.n1523 VDPWR.n1521 2.63539
R10863 VDPWR.n1440 VDPWR.n1438 2.63539
R10864 VDPWR.n1723 VDPWR.n1721 2.63539
R10865 VDPWR.n1286 VDPWR.n1284 2.63539
R10866 VDPWR.n1289 VDPWR.n1287 2.63539
R10867 VDPWR.n1293 VDPWR.n1291 2.63539
R10868 VDPWR.n1298 VDPWR.n1296 2.63539
R10869 VDPWR.n1424 VDPWR.n1422 2.63539
R10870 VDPWR.n1429 VDPWR.n1427 2.63539
R10871 VDPWR.n1906 VDPWR.n1904 2.63539
R10872 VDPWR.n1912 VDPWR.n1910 2.63539
R10873 VDPWR.n1915 VDPWR.n1913 2.63539
R10874 VDPWR.n1919 VDPWR.n1917 2.63539
R10875 VDPWR.n2054 VDPWR.n2052 2.63539
R10876 VDPWR.n2057 VDPWR.n2055 2.63539
R10877 VDPWR.n2213 VDPWR.n2211 2.63539
R10878 VDPWR.n2216 VDPWR.n2214 2.63539
R10879 VDPWR.n1176 VDPWR.n1174 2.63539
R10880 VDPWR.n2445 VDPWR.n2443 2.63539
R10881 VDPWR.n964 VDPWR.n962 2.63539
R10882 VDPWR.n967 VDPWR.n965 2.63539
R10883 VDPWR.n2465 VDPWR.n2463 2.63539
R10884 VDPWR.n2468 VDPWR.n2466 2.63539
R10885 VDPWR.n2597 VDPWR.n2595 2.63539
R10886 VDPWR.n2600 VDPWR.n2598 2.63539
R10887 VDPWR.n927 VDPWR.n925 2.63539
R10888 VDPWR.n2923 VDPWR.n2921 2.63539
R10889 VDPWR.n2961 VDPWR.n2959 2.63539
R10890 VDPWR.n2969 VDPWR.n2967 2.63539
R10891 VDPWR.n815 VDPWR.n813 2.63539
R10892 VDPWR.n2633 VDPWR.n2631 2.63539
R10893 VDPWR.n2636 VDPWR.n2634 2.63539
R10894 VDPWR.n828 VDPWR.n826 2.63539
R10895 VDPWR.n832 VDPWR.n830 2.63539
R10896 VDPWR.n2326 VDPWR.n2325 2.62345
R10897 VDPWR.n2041 VDPWR.n2040 2.61352
R10898 VDPWR.n2378 VDPWR.n2377 2.56175
R10899 VDPWR.n576 VDPWR.n575 2.54018
R10900 VDPWR.n555 VDPWR.n554 2.54018
R10901 VDPWR.n296 VDPWR.n295 2.54018
R10902 VDPWR.n275 VDPWR.n274 2.54018
R10903 VDPWR.n792 VDPWR.n789 2.54018
R10904 VDPWR.n39 VDPWR.n38 2.54018
R10905 VDPWR.n18 VDPWR.n17 2.54018
R10906 VDPWR.n3023 VDPWR.n793 2.3878
R10907 VDPWR.n818 VDPWR.n817 2.37764
R10908 VDPWR.n1483 VDPWR.n1482 2.37495
R10909 VDPWR.n1513 VDPWR.n1512 2.37495
R10910 VDPWR.n1510 VDPWR.n1509 2.37495
R10911 VDPWR.n1522 VDPWR.n1521 2.37495
R10912 VDPWR.n1517 VDPWR.n1516 2.37495
R10913 VDPWR.n1722 VDPWR.n1721 2.37495
R10914 VDPWR.n1439 VDPWR.n1438 2.37495
R10915 VDPWR.n1288 VDPWR.n1287 2.37495
R10916 VDPWR.n1285 VDPWR.n1284 2.37495
R10917 VDPWR.n1297 VDPWR.n1296 2.37495
R10918 VDPWR.n1292 VDPWR.n1291 2.37495
R10919 VDPWR.n1428 VDPWR.n1427 2.37495
R10920 VDPWR.n1423 VDPWR.n1422 2.37495
R10921 VDPWR.n1911 VDPWR.n1910 2.37495
R10922 VDPWR.n1905 VDPWR.n1904 2.37495
R10923 VDPWR.n1918 VDPWR.n1917 2.37495
R10924 VDPWR.n1914 VDPWR.n1913 2.37495
R10925 VDPWR.n2056 VDPWR.n2055 2.37495
R10926 VDPWR.n2053 VDPWR.n2052 2.37495
R10927 VDPWR.n2215 VDPWR.n2214 2.37495
R10928 VDPWR.n2212 VDPWR.n2211 2.37495
R10929 VDPWR.n2444 VDPWR.n2443 2.37495
R10930 VDPWR.n1175 VDPWR.n1174 2.37495
R10931 VDPWR.n966 VDPWR.n965 2.37495
R10932 VDPWR.n963 VDPWR.n962 2.37495
R10933 VDPWR.n2467 VDPWR.n2466 2.37495
R10934 VDPWR.n2464 VDPWR.n2463 2.37495
R10935 VDPWR.n2599 VDPWR.n2598 2.37495
R10936 VDPWR.n2596 VDPWR.n2595 2.37495
R10937 VDPWR.n926 VDPWR.n925 2.37495
R10938 VDPWR.n2922 VDPWR.n2921 2.37495
R10939 VDPWR.n2968 VDPWR.n2967 2.37495
R10940 VDPWR.n2960 VDPWR.n2959 2.37495
R10941 VDPWR.n814 VDPWR.n813 2.37495
R10942 VDPWR.n2635 VDPWR.n2634 2.37495
R10943 VDPWR.n2632 VDPWR.n2631 2.37495
R10944 VDPWR.n831 VDPWR.n830 2.37495
R10945 VDPWR.n827 VDPWR.n826 2.37495
R10946 VDPWR.n601 VDPWR.n597 2.33701
R10947 VDPWR.n589 VDPWR.n588 2.33701
R10948 VDPWR.n575 VDPWR.n574 2.33701
R10949 VDPWR.n555 VDPWR.n549 2.33701
R10950 VDPWR.n321 VDPWR.n317 2.33701
R10951 VDPWR.n309 VDPWR.n308 2.33701
R10952 VDPWR.n295 VDPWR.n294 2.33701
R10953 VDPWR.n275 VDPWR.n269 2.33701
R10954 VDPWR.n1246 VDPWR.n1245 2.33701
R10955 VDPWR.n1119 VDPWR.n1118 2.33701
R10956 VDPWR.n2909 VDPWR.n2902 2.33701
R10957 VDPWR.n2797 VDPWR.n2654 2.33701
R10958 VDPWR.n64 VDPWR.n60 2.33701
R10959 VDPWR.n52 VDPWR.n51 2.33701
R10960 VDPWR.n38 VDPWR.n37 2.33701
R10961 VDPWR.n18 VDPWR.n12 2.33701
R10962 VDPWR.n1592 VDPWR.n1485 2.32777
R10963 VDPWR.n1965 VDPWR.n1964 2.32777
R10964 VDPWR.n1383 VDPWR.n1382 2.28432
R10965 VDPWR.n2576 VDPWR.n960 2.28407
R10966 VDPWR.n2576 VDPWR.n961 2.28407
R10967 VDPWR.n2209 VDPWR.n2207 2.28374
R10968 VDPWR.n1992 VDPWR.n1991 2.27742
R10969 VDPWR.n2035 VDPWR.n2034 2.25932
R10970 VDPWR.n2101 VDPWR.n2018 2.25932
R10971 VDPWR.n2603 VDPWR.n2594 2.25293
R10972 VDPWR.n3030 VDPWR.n3029 2.23542
R10973 VDPWR.n2524 VDPWR.n2523 2.22199
R10974 VDPWR.n3056 VDPWR.n3055 2.16151
R10975 VDPWR.n401 VDPWR.n400 2.13883
R10976 VDPWR.n482 VDPWR.n481 2.13544
R10977 VDPWR.n583 VDPWR.n576 2.13383
R10978 VDPWR.n554 VDPWR.n553 2.13383
R10979 VDPWR.n303 VDPWR.n296 2.13383
R10980 VDPWR.n274 VDPWR.n273 2.13383
R10981 VDPWR.n3025 VDPWR.n792 2.13383
R10982 VDPWR.n46 VDPWR.n39 2.13383
R10983 VDPWR.n17 VDPWR.n16 2.13383
R10984 VDPWR.n2408 VDPWR.n2407 2.0932
R10985 VDPWR.n973 VDPWR.n972 2.07374
R10986 VDPWR.n984 VDPWR.n983 2.07374
R10987 VDPWR.n597 VDPWR.n595 2.03225
R10988 VDPWR.n588 VDPWR.n587 2.03225
R10989 VDPWR.n574 VDPWR.n573 2.03225
R10990 VDPWR.n549 VDPWR.n547 2.03225
R10991 VDPWR.n317 VDPWR.n315 2.03225
R10992 VDPWR.n308 VDPWR.n307 2.03225
R10993 VDPWR.n294 VDPWR.n293 2.03225
R10994 VDPWR.n269 VDPWR.n267 2.03225
R10995 VDPWR.n1118 VDPWR.n1117 2.03225
R10996 VDPWR.n2654 VDPWR.n2653 2.03225
R10997 VDPWR.n60 VDPWR.n58 2.03225
R10998 VDPWR.n51 VDPWR.n50 2.03225
R10999 VDPWR.n37 VDPWR.n36 2.03225
R11000 VDPWR.n12 VDPWR.n10 2.03225
R11001 VDPWR.n1416 VDPWR.n1414 2.01703
R11002 VDPWR.n1421 VDPWR.n1419 2.01703
R11003 VDPWR.n2590 VDPWR.n2588 2.01703
R11004 VDPWR.n2593 VDPWR.n2591 2.01703
R11005 VDPWR.n3032 VDPWR.n3031 1.98145
R11006 VDPWR.n794 VDPWR.n793 1.98145
R11007 VDPWR.n481 VDPWR.n466 1.95379
R11008 VDPWR.n2302 VDPWR.n2301 1.88902
R11009 VDPWR.n2377 VDPWR.n1200 1.88902
R11010 VDPWR.n1420 VDPWR.n1419 1.88416
R11011 VDPWR.n1415 VDPWR.n1414 1.88416
R11012 VDPWR.n2592 VDPWR.n2591 1.88416
R11013 VDPWR.n2589 VDPWR.n2588 1.88416
R11014 VDPWR.n1952 VDPWR.n1951 1.88325
R11015 VDPWR.n1561 VDPWR.n1560 1.88295
R11016 VDPWR.n1865 VDPWR.n1311 1.88295
R11017 VDPWR.n660 VDPWR.n656 1.88285
R11018 VDPWR.n477 VDPWR.n476 1.88285
R11019 VDPWR.n417 VDPWR.n413 1.88285
R11020 VDPWR.n3067 VDPWR.n3066 1.88285
R11021 VDPWR.n1085 VDPWR.n1034 1.88285
R11022 VDPWR.n1535 VDPWR.n1534 1.85065
R11023 VDPWR.n1537 VDPWR.n1501 1.85065
R11024 VDPWR.n1667 VDPWR.n1666 1.85065
R11025 VDPWR.n1305 VDPWR.n1304 1.85065
R11026 VDPWR.n1887 VDPWR.n1306 1.85065
R11027 VDPWR.n1969 VDPWR.n1968 1.85065
R11028 VDPWR.n1924 VDPWR.n1901 1.85065
R11029 VDPWR.n1926 VDPWR.n1272 1.85065
R11030 VDPWR.n2233 VDPWR.n2232 1.85065
R11031 VDPWR.n2698 VDPWR.n2696 1.85065
R11032 VDPWR.n2534 VDPWR.n1017 1.82907
R11033 VDPWR.n2901 VDPWR.n2900 1.82907
R11034 VDPWR.n1665 VDPWR.n1664 1.81289
R11035 VDPWR.n2231 VDPWR.n2230 1.81289
R11036 VDPWR.n653 VDPWR.n652 1.753
R11037 VDPWR.n373 VDPWR.n372 1.753
R11038 VDPWR.n116 VDPWR.n115 1.753
R11039 VDPWR.n2112 VDPWR.n2015 1.73737
R11040 VDPWR.n2353 VDPWR.n2350 1.73737
R11041 VDPWR.n2431 VDPWR.n2430 1.73737
R11042 VDPWR.n2344 VDPWR.n2343 1.69306
R11043 VDPWR.n2423 VDPWR.n1178 1.69306
R11044 VDPWR.n3011 VDPWR.n868 1.69188
R11045 VDPWR.n3011 VDPWR.n3010 1.69188
R11046 VDPWR.n2504 VDPWR.n867 1.69188
R11047 VDPWR.n2506 VDPWR.n867 1.69188
R11048 VDPWR.n2088 VDPWR.n1191 1.69188
R11049 VDPWR.n2090 VDPWR.n1191 1.69188
R11050 VDPWR.n1769 VDPWR.n1768 1.69188
R11051 VDPWR.n1770 VDPWR.n1769 1.69188
R11052 VDPWR.n1689 VDPWR.n1392 1.69188
R11053 VDPWR.n1678 VDPWR.n1392 1.69188
R11054 VDPWR.n2401 VDPWR.n1192 1.69188
R11055 VDPWR.n2916 VDPWR.n2915 1.69188
R11056 VDPWR.n2915 VDPWR.n2914 1.69188
R11057 VDPWR.n1129 VDPWR.n887 1.69188
R11058 VDPWR.n1112 VDPWR.n887 1.69188
R11059 VDPWR.n2360 VDPWR.n2359 1.69188
R11060 VDPWR.n2359 VDPWR.n2358 1.69188
R11061 VDPWR.n2120 VDPWR.n1210 1.69188
R11062 VDPWR.n2123 VDPWR.n1210 1.69188
R11063 VDPWR.n1794 VDPWR.n1793 1.69188
R11064 VDPWR.n1795 VDPWR.n1794 1.69188
R11065 VDPWR.n1653 VDPWR.n1363 1.69188
R11066 VDPWR.n1639 VDPWR.n1363 1.69188
R11067 VDPWR.n2880 VDPWR.n2879 1.69188
R11068 VDPWR.n2879 VDPWR.n2878 1.69188
R11069 VDPWR.n2320 VDPWR.n2319 1.69188
R11070 VDPWR.n2319 VDPWR.n2318 1.69188
R11071 VDPWR.n2149 VDPWR.n1230 1.69188
R11072 VDPWR.n2152 VDPWR.n1230 1.69188
R11073 VDPWR.n1823 VDPWR.n1822 1.69188
R11074 VDPWR.n1824 VDPWR.n1823 1.69188
R11075 VDPWR.n1615 VDPWR.n1339 1.69188
R11076 VDPWR.n1606 VDPWR.n1339 1.69188
R11077 VDPWR.n1076 VDPWR.n913 1.69188
R11078 VDPWR.n2582 VDPWR.n955 1.69188
R11079 VDPWR.n2582 VDPWR.n2581 1.69188
R11080 VDPWR.n2240 VDPWR.n954 1.69188
R11081 VDPWR.n2226 VDPWR.n954 1.69188
R11082 VDPWR.n1934 VDPWR.n1933 1.69188
R11083 VDPWR.n1933 VDPWR.n1932 1.69188
R11084 VDPWR.n1894 VDPWR.n1277 1.69188
R11085 VDPWR.n1894 VDPWR.n1893 1.69188
R11086 VDPWR.n1543 VDPWR.n1276 1.69188
R11087 VDPWR.n1530 VDPWR.n1276 1.69188
R11088 VDPWR.n2803 VDPWR.n2583 1.69188
R11089 VDPWR.n2977 VDPWR.n774 1.69188
R11090 VDPWR.n2974 VDPWR.n774 1.69188
R11091 VDPWR.n2480 VDPWR.n2455 1.69188
R11092 VDPWR.n2470 VDPWR.n2455 1.69188
R11093 VDPWR.n2454 VDPWR.n1168 1.69188
R11094 VDPWR.n2454 VDPWR.n2453 1.69188
R11095 VDPWR.n2069 VDPWR.n1167 1.69188
R11096 VDPWR.n2059 VDPWR.n1167 1.69188
R11097 VDPWR.n1736 VDPWR.n1733 1.69188
R11098 VDPWR.n1745 VDPWR.n1733 1.69188
R11099 VDPWR.n1732 VDPWR.n1432 1.69188
R11100 VDPWR.n1732 VDPWR.n1731 1.69188
R11101 VDPWR.n2842 VDPWR.n2841 1.69188
R11102 VDPWR.n2841 VDPWR.n2840 1.69188
R11103 VDPWR.n2538 VDPWR.n933 1.69188
R11104 VDPWR.n2540 VDPWR.n933 1.69188
R11105 VDPWR.n2275 VDPWR.n2274 1.69188
R11106 VDPWR.n2274 VDPWR.n2273 1.69188
R11107 VDPWR.n2188 VDPWR.n1258 1.69188
R11108 VDPWR.n2188 VDPWR.n2187 1.69188
R11109 VDPWR.n1851 VDPWR.n1257 1.69188
R11110 VDPWR.n1854 VDPWR.n1257 1.69188
R11111 VDPWR.n1582 VDPWR.n1581 1.69188
R11112 VDPWR.n1581 VDPWR.n1580 1.69188
R11113 VDPWR.t185 VDPWR 1.67895
R11114 VDPWR.t747 VDPWR 1.67895
R11115 VDPWR.n2905 VDPWR.n2904 1.67669
R11116 VDPWR.n1667 VDPWR.n1665 1.66186
R11117 VDPWR.n2233 VDPWR.n2231 1.66186
R11118 VDPWR.n2733 VDPWR.n2695 1.64857
R11119 VDPWR.n1536 VDPWR.n1535 1.6241
R11120 VDPWR.n1547 VDPWR.n1501 1.6241
R11121 VDPWR.n1666 VDPWR.n1456 1.6241
R11122 VDPWR.n1888 VDPWR.n1305 1.6241
R11123 VDPWR.n1877 VDPWR.n1306 1.6241
R11124 VDPWR.n1927 VDPWR.n1924 1.6241
R11125 VDPWR.n1938 VDPWR.n1272 1.6241
R11126 VDPWR.n2232 VDPWR.n2199 1.6241
R11127 VDPWR.n2728 VDPWR.n2698 1.6241
R11128 VDPWR.n1562 VDPWR.n1561 1.62167
R11129 VDPWR.n1862 VDPWR.n1311 1.62167
R11130 VDPWR.n1953 VDPWR.n1952 1.62136
R11131 VDPWR.n3110 VDPWR.n117 1.59405
R11132 VDPWR.n753 VDPWR.n752 1.57294
R11133 VDPWR.n746 VDPWR.t174 1.53603
R11134 VDPWR.n743 VDPWR.t174 1.53603
R11135 VDPWR.n530 VDPWR.n529 1.51493
R11136 VDPWR.n2015 VDPWR.n2013 1.51082
R11137 VDPWR.n2350 VDPWR.n2349 1.51082
R11138 VDPWR.n2430 VDPWR.n2429 1.51082
R11139 VDPWR.n757 VDPWR 1.48239
R11140 VDPWR.n572 VDPWR.n570 1.46504
R11141 VDPWR.n292 VDPWR.n290 1.46504
R11142 VDPWR.n35 VDPWR.n33 1.46504
R11143 VDPWR.n531 VDPWR.n253 1.42384
R11144 VDPWR.n645 VDPWR.n545 1.4005
R11145 VDPWR.n365 VDPWR.n265 1.4005
R11146 VDPWR.n1108 VDPWR.n1107 1.4005
R11147 VDPWR.n2563 VDPWR.n988 1.4005
R11148 VDPWR.n108 VDPWR.n8 1.4005
R11149 VDPWR.n1970 VDPWR.n1969 1.39755
R11150 VDPWR.n2330 VDPWR.n2329 1.36443
R11151 VDPWR.n2413 VDPWR.n2412 1.36443
R11152 VDPWR.n757 VDPWR.n756 1.34339
R11153 VDPWR.n1116 VDPWR.n1028 1.3232
R11154 VDPWR.n401 VDPWR.n388 1.28133
R11155 VDPWR.n2041 VDPWR.n2039 1.2502
R11156 VDPWR.n256 VDPWR.n253 1.22948
R11157 VDPWR.n3071 VDPWR.n3070 1.16528
R11158 VDPWR.n754 VDPWR.n118 1.15151
R11159 VDPWR.n702 VDPWR.n701 1.143
R11160 VDPWR.n686 VDPWR.n685 1.143
R11161 VDPWR.n513 VDPWR.n512 1.143
R11162 VDPWR.n497 VDPWR.n496 1.143
R11163 VDPWR.n459 VDPWR.n458 1.143
R11164 VDPWR.n443 VDPWR.n442 1.143
R11165 VDPWR.n3103 VDPWR.n3102 1.143
R11166 VDPWR.n3087 VDPWR.n3086 1.143
R11167 VDPWR.n718 VDPWR.n717 1.13925
R11168 VDPWR.n529 VDPWR.n528 1.13925
R11169 VDPWR.n465 VDPWR.n464 1.13925
R11170 VDPWR.n3109 VDPWR.n3108 1.13925
R11171 VDPWR.n3051 VDPWR.n3050 1.13717
R11172 VDPWR.n670 VDPWR.n669 1.13675
R11173 VDPWR.n481 VDPWR.n480 1.13675
R11174 VDPWR.n427 VDPWR.n426 1.13675
R11175 VDPWR.n714 VDPWR.n713 1.12991
R11176 VDPWR.n690 VDPWR.n688 1.12991
R11177 VDPWR.n682 VDPWR.n674 1.12991
R11178 VDPWR.n525 VDPWR.n524 1.12991
R11179 VDPWR.n501 VDPWR.n499 1.12991
R11180 VDPWR.n493 VDPWR.n485 1.12991
R11181 VDPWR.n461 VDPWR.n412 1.12991
R11182 VDPWR.n447 VDPWR.n445 1.12991
R11183 VDPWR.n439 VDPWR.n431 1.12991
R11184 VDPWR.n3105 VDPWR.n768 1.12991
R11185 VDPWR.n3091 VDPWR.n3089 1.12991
R11186 VDPWR.n3083 VDPWR.n3075 1.12991
R11187 VDPWR.n2714 VDPWR.n2713 1.11173
R11188 VDPWR.n2652 VDPWR.n2622 1.08324
R11189 VDPWR.n720 VDPWR.n719 1.06914
R11190 VDPWR.n594 VDPWR 1.06099
R11191 VDPWR.n314 VDPWR 1.06099
R11192 VDPWR.n57 VDPWR 1.06099
R11193 VDPWR.n1526 VDPWR.n1525 1.05773
R11194 VDPWR.n1301 VDPWR.n1300 1.05773
R11195 VDPWR.n1922 VDPWR.n1903 1.05773
R11196 VDPWR.n2694 VDPWR.n2693 1.05773
R11197 VDPWR.n2340 VDPWR.n1220 1.04968
R11198 VDPWR.n2422 VDPWR.n2421 1.04968
R11199 VDPWR.n972 VDPWR.n960 0.992049
R11200 VDPWR.n984 VDPWR.n961 0.992049
R11201 VDPWR.n2165 VDPWR.n1967 0.899674
R11202 VDPWR VDPWR.n118 0.891339
R11203 VDPWR.n755 VDPWR.n754 0.884173
R11204 VDPWR.n2291 VDPWR.n1245 0.863992
R11205 VDPWR.n375 VDPWR.n374 0.853
R11206 VDPWR.n3042 VDPWR.n778 0.853
R11207 VDPWR.n2741 VDPWR.n914 0.853
R11208 VDPWR.n2769 VDPWR.n934 0.853
R11209 VDPWR.n2802 VDPWR.n2801 0.853
R11210 VDPWR.n3014 VDPWR.n3013 0.853
R11211 VDPWR.n687 VDPWR.n686 0.849559
R11212 VDPWR.n444 VDPWR.n443 0.849559
R11213 VDPWR.n498 VDPWR.n497 0.849559
R11214 VDPWR.n530 VDPWR.n376 0.843267
R11215 VDPWR.n2777 VDPWR.n2776 0.813198
R11216 VDPWR.n2753 VDPWR.n2752 0.813198
R11217 VDPWR.n531 VDPWR.n530 0.810458
R11218 VDPWR VDPWR.n3053 0.778686
R11219 VDPWR.n738 VDPWR.n737 0.7755
R11220 VDPWR.n671 VDPWR.n670 0.770881
R11221 VDPWR.n428 VDPWR.n427 0.770881
R11222 VDPWR.n402 VDPWR.n401 0.767167
R11223 VDPWR.n374 VDPWR.n373 0.763912
R11224 VDPWR.n632 VDPWR.n561 0.753441
R11225 VDPWR.n352 VDPWR.n281 0.753441
R11226 VDPWR.n1758 VDPWR.n1757 0.753441
R11227 VDPWR.n95 VDPWR.n24 0.753441
R11228 VDPWR.n1776 VDPWR.n1387 0.740996
R11229 VDPWR.n460 VDPWR.n459 0.73614
R11230 VDPWR.n703 VDPWR.n702 0.717512
R11231 VDPWR.n514 VDPWR.n513 0.717512
R11232 VDPWR.n1156 VDPWR.n1155 0.706789
R11233 VDPWR.n757 VDPWR.n118 0.70421
R11234 VDPWR.n255 VDPWR 0.659186
R11235 VDPWR.n3055 VDPWR.n3054 0.65336
R11236 VDPWR.n862 VDPWR.n810 0.65125
R11237 VDPWR.n1659 VDPWR.n1458 0.635211
R11238 VDPWR.n1693 VDPWR.n1447 0.635211
R11239 VDPWR.n1408 VDPWR.n1396 0.635211
R11240 VDPWR.n2300 VDPWR.n2299 0.635211
R11241 VDPWR.n2368 VDPWR.n1204 0.635211
R11242 VDPWR.n2375 VDPWR.n2374 0.635211
R11243 VDPWR.n1136 VDPWR.n1133 0.635211
R11244 VDPWR.n1155 VDPWR.n1151 0.635211
R11245 VDPWR.n2500 VDPWR.n2499 0.635211
R11246 VDPWR.n1160 VDPWR.n1158 0.635211
R11247 VDPWR.n2333 VDPWR.n1223 0.630008
R11248 VDPWR.n2407 VDPWR.n1187 0.630008
R11249 VDPWR.n2409 VDPWR.n1184 0.630008
R11250 VDPWR.n655 VDPWR.n536 0.624567
R11251 VDPWR.n542 VDPWR.n540 0.6005
R11252 VDPWR.n262 VDPWR.n260 0.6005
R11253 VDPWR.n5 VDPWR.n3 0.6005
R11254 VDPWR.n2336 VDPWR.n2335 0.52509
R11255 VDPWR.n466 VDPWR.n465 0.518882
R11256 VDPWR.n654 VDPWR.n653 0.511794
R11257 VDPWR.n3116 VDPWR.n116 0.511794
R11258 VDPWR.n142 VDPWR.n141 0.465384
R11259 VDPWR.n653 VDPWR 0.460219
R11260 VDPWR.n373 VDPWR 0.460219
R11261 VDPWR.n116 VDPWR 0.460219
R11262 VDPWR.n3031 VDPWR.n3030 0.457643
R11263 VDPWR.n375 VDPWR.n256 0.45408
R11264 VDPWR.n718 VDPWR.n703 0.405788
R11265 VDPWR.n648 VDPWR.n540 0.4005
R11266 VDPWR.n368 VDPWR.n260 0.4005
R11267 VDPWR.n111 VDPWR.n3 0.4005
R11268 VDPWR.n686 VDPWR.n671 0.379066
R11269 VDPWR.n443 VDPWR.n428 0.379066
R11270 VDPWR.n497 VDPWR.n482 0.379066
R11271 VDPWR.n720 VDPWR.n253 0.375001
R11272 VDPWR.n376 VDPWR 0.36983
R11273 VDPWR.n1594 VDPWR.n1593 0.369731
R11274 VDPWR.n1623 VDPWR.n1471 0.369731
R11275 VDPWR.n1624 VDPWR.n1470 0.369731
R11276 VDPWR.n1646 VDPWR.n1645 0.369731
R11277 VDPWR.n1555 VDPWR.n1554 0.369731
R11278 VDPWR.n1560 VDPWR.n1497 0.369731
R11279 VDPWR.n1563 VDPWR.n1562 0.369731
R11280 VDPWR.n1586 VDPWR.n1486 0.369731
R11281 VDPWR.n1694 VDPWR.n1446 0.369731
R11282 VDPWR.n1710 VDPWR.n1437 0.369731
R11283 VDPWR.n1871 VDPWR.n1309 0.369731
R11284 VDPWR.n1866 VDPWR.n1865 0.369731
R11285 VDPWR.n1862 VDPWR.n1861 0.369731
R11286 VDPWR.n1847 VDPWR.n1329 0.369731
R11287 VDPWR.n1834 VDPWR.n1333 0.369731
R11288 VDPWR.n1816 VDPWR.n1815 0.369731
R11289 VDPWR.n1810 VDPWR.n1355 0.369731
R11290 VDPWR.n1377 VDPWR.n1376 0.369731
R11291 VDPWR.n2132 VDPWR.n1993 0.369731
R11292 VDPWR.n2012 VDPWR.n2011 0.369731
R11293 VDPWR.n1990 VDPWR.n1988 0.369731
R11294 VDPWR.n2133 VDPWR.n1992 0.369731
R11295 VDPWR.n2156 VDPWR.n1971 0.369731
R11296 VDPWR.n2143 VDPWR.n2142 0.369731
R11297 VDPWR.n1954 VDPWR.n1953 0.369731
R11298 VDPWR.n2175 VDPWR.n2174 0.369731
R11299 VDPWR.n1946 VDPWR.n1945 0.369731
R11300 VDPWR.n1951 VDPWR.n1268 0.369731
R11301 VDPWR.n2251 VDPWR.n2250 0.369731
R11302 VDPWR.n2255 VDPWR.n2195 0.369731
R11303 VDPWR.n2257 VDPWR.n2256 0.369731
R11304 VDPWR.n2282 VDPWR.n2281 0.369731
R11305 VDPWR.n529 VDPWR.n514 0.360095
R11306 VDPWR.n702 VDPWR.n687 0.348599
R11307 VDPWR.n459 VDPWR.n444 0.348599
R11308 VDPWR.n513 VDPWR.n498 0.348599
R11309 VDPWR.n3054 VDPWR.n117 0.320594
R11310 VDPWR.n2370 VDPWR.n2369 0.317855
R11311 VDPWR.n2369 VDPWR.n1203 0.317855
R11312 VDPWR.n750 VDPWR.n738 0.310024
R11313 VDPWR.n3048 VDPWR 0.306
R11314 VDPWR.n604 VDPWR.n595 0.305262
R11315 VDPWR.n623 VDPWR.n622 0.305262
R11316 VDPWR.n573 VDPWR.n572 0.305262
R11317 VDPWR.n582 VDPWR.n581 0.305262
R11318 VDPWR.n558 VDPWR.n547 0.305262
R11319 VDPWR.n324 VDPWR.n315 0.305262
R11320 VDPWR.n343 VDPWR.n342 0.305262
R11321 VDPWR.n293 VDPWR.n292 0.305262
R11322 VDPWR.n302 VDPWR.n301 0.305262
R11323 VDPWR.n278 VDPWR.n267 0.305262
R11324 VDPWR.n749 VDPWR.n739 0.305262
R11325 VDPWR.n2051 VDPWR.n2043 0.305262
R11326 VDPWR.n2294 VDPWR.n1244 0.305262
R11327 VDPWR.n1117 VDPWR.n1116 0.305262
R11328 VDPWR.n1121 VDPWR.n1021 0.305262
R11329 VDPWR.n2565 VDPWR.n986 0.305262
R11330 VDPWR.n2900 VDPWR.n2899 0.305262
R11331 VDPWR.n2904 VDPWR.n2903 0.305262
R11332 VDPWR.n2988 VDPWR.n2947 0.305262
R11333 VDPWR.n2958 VDPWR.n2957 0.305262
R11334 VDPWR.n2659 VDPWR.n2658 0.305262
R11335 VDPWR.n2781 VDPWR.n2660 0.305262
R11336 VDPWR.n2775 VDPWR.n2774 0.305262
R11337 VDPWR.n2653 VDPWR.n2652 0.305262
R11338 VDPWR.n2795 VDPWR.n2794 0.305262
R11339 VDPWR.n2759 VDPWR.n2758 0.305262
R11340 VDPWR.n2757 VDPWR.n2676 0.305262
R11341 VDPWR.n2748 VDPWR.n2679 0.305262
R11342 VDPWR.n3035 VDPWR.n788 0.305262
R11343 VDPWR.n3020 VDPWR.n794 0.305262
R11344 VDPWR.n862 VDPWR.n861 0.305262
R11345 VDPWR.n825 VDPWR.n824 0.305262
R11346 VDPWR.n67 VDPWR.n58 0.305262
R11347 VDPWR.n86 VDPWR.n85 0.305262
R11348 VDPWR.n36 VDPWR.n35 0.305262
R11349 VDPWR.n45 VDPWR.n44 0.305262
R11350 VDPWR.n21 VDPWR.n10 0.305262
R11351 VDPWR.n2801 VDPWR.n2618 0.297373
R11352 VDPWR.n383 VDPWR.t362 0.27666
R11353 VDPWR.t362 VDPWR.n382 0.27666
R11354 VDPWR.n395 VDPWR.t547 0.27666
R11355 VDPWR.t547 VDPWR.n394 0.27666
R11356 VDPWR.n755 VDPWR.n720 0.262659
R11357 VDPWR.n737 VDPWR.n728 0.2565
R11358 VDPWR.n2560 VDPWR.n2557 0.25148
R11359 VDPWR.n1047 VDPWR.n1045 0.246654
R11360 VDPWR.n2603 VDPWR 0.237784
R11361 VDPWR.n1735 VDPWR.n1418 0.231913
R11362 VDPWR.n1526 VDPWR.n1508 0.227049
R11363 VDPWR.n1549 VDPWR.n1499 0.227049
R11364 VDPWR.n1663 VDPWR.n1662 0.227049
R11365 VDPWR.n1673 VDPWR.n1454 0.227049
R11366 VDPWR.n1301 VDPWR.n1283 0.227049
R11367 VDPWR.n1872 VDPWR.n1308 0.227049
R11368 VDPWR.n2115 VDPWR.n2013 0.227049
R11369 VDPWR.n2110 VDPWR.n2109 0.227049
R11370 VDPWR.n2157 VDPWR.n1970 0.227049
R11371 VDPWR.n1903 VDPWR.n1902 0.227049
R11372 VDPWR.n1940 VDPWR.n1270 0.227049
R11373 VDPWR.n2223 VDPWR.n2205 0.227049
R11374 VDPWR.n2249 VDPWR.n2197 0.227049
R11375 VDPWR.n2349 VDPWR.n2348 0.227049
R11376 VDPWR.n2364 VDPWR.n1206 0.227049
R11377 VDPWR.n2429 VDPWR.n2428 0.227049
R11378 VDPWR.n2432 VDPWR.n1173 0.227049
R11379 VDPWR.n2490 VDPWR.n1162 0.227049
R11380 VDPWR.n2462 VDPWR.n2461 0.227049
R11381 VDPWR.n2693 VDPWR.n2692 0.227049
R11382 VDPWR.n2727 VDPWR.n2726 0.227049
R11383 VDPWR VDPWR.n1785 0.217591
R11384 VDPWR.n1781 VDPWR.n1780 0.21207
R11385 VDPWR.n1137 VDPWR.n1136 0.21207
R11386 VDPWR.n2498 VDPWR.n2497 0.21207
R11387 VDPWR VDPWR.n2613 0.209323
R11388 VDPWR.n3104 VDPWR.n3103 0.209134
R11389 VDPWR.n3088 VDPWR.n3087 0.206276
R11390 VDPWR.n3048 VDPWR.n3047 0.206051
R11391 VDPWR.n2902 VDPWR.n2901 0.203675
R11392 VDPWR VDPWR.n2603 0.200023
R11393 VDPWR.n3053 VDPWR.n769 0.197315
R11394 VDPWR.n3043 VDPWR.n769 0.196829
R11395 VDPWR.n3047 VDPWR.n3046 0.196829
R11396 VDPWR.n2618 VDPWR.n776 0.195044
R11397 VDPWR.n2613 VDPWR.n775 0.195044
R11398 VDPWR.n2555 VDPWR.n992 0.194439
R11399 VDPWR.n3114 VDPWR 0.189894
R11400 VDPWR.n2085 VDPWR.n2030 0.180304
R11401 VDPWR.n2896 VDPWR.n896 0.180304
R11402 VDPWR.n1591 VDPWR 0.17983
R11403 VDPWR VDPWR.n2171 0.17983
R11404 VDPWR VDPWR.n2079 0.17983
R11405 VDPWR.n979 VDPWR 0.17983
R11406 VDPWR.n1520 VDPWR 0.179485
R11407 VDPWR.n1295 VDPWR 0.179485
R11408 VDPWR.n1418 VDPWR 0.179485
R11409 VDPWR VDPWR.n1909 0.179485
R11410 VDPWR.n2079 VDPWR 0.179485
R11411 VDPWR.n2920 VDPWR 0.179485
R11412 VDPWR.n738 VDPWR.n727 0.176553
R11413 VDPWR VDPWR.n1519 0.172576
R11414 VDPWR VDPWR.n1294 0.172576
R11415 VDPWR.n1916 VDPWR 0.172576
R11416 VDPWR VDPWR.n2218 0.172576
R11417 VDPWR VDPWR.n969 0.172576
R11418 VDPWR VDPWR.n2602 0.172576
R11419 VDPWR VDPWR.n2638 0.172576
R11420 VDPWR.n535 VDPWR 0.163379
R11421 VDPWR.n1769 VDPWR.n1392 0.1603
R11422 VDPWR.n1769 VDPWR.n1191 0.1603
R11423 VDPWR.n2401 VDPWR.n1191 0.1603
R11424 VDPWR.n2401 VDPWR.n867 0.1603
R11425 VDPWR.n3011 VDPWR.n867 0.1603
R11426 VDPWR.n3013 VDPWR.n3011 0.1603
R11427 VDPWR.n1794 VDPWR.n1363 0.1603
R11428 VDPWR.n1794 VDPWR.n1210 0.1603
R11429 VDPWR.n2359 VDPWR.n1210 0.1603
R11430 VDPWR.n2359 VDPWR.n887 0.1603
R11431 VDPWR.n2915 VDPWR.n887 0.1603
R11432 VDPWR.n2915 VDPWR.n778 0.1603
R11433 VDPWR.n1823 VDPWR.n1339 0.1603
R11434 VDPWR.n1823 VDPWR.n1230 0.1603
R11435 VDPWR.n2319 VDPWR.n1230 0.1603
R11436 VDPWR.n2319 VDPWR.n913 0.1603
R11437 VDPWR.n2879 VDPWR.n913 0.1603
R11438 VDPWR.n2879 VDPWR.n914 0.1603
R11439 VDPWR.n1894 VDPWR.n1276 0.1603
R11440 VDPWR.n1933 VDPWR.n1894 0.1603
R11441 VDPWR.n1933 VDPWR.n954 0.1603
R11442 VDPWR.n2582 VDPWR.n954 0.1603
R11443 VDPWR.n2803 VDPWR.n2582 0.1603
R11444 VDPWR.n2803 VDPWR.n2802 0.1603
R11445 VDPWR.n1581 VDPWR.n1257 0.1603
R11446 VDPWR.n2188 VDPWR.n1257 0.1603
R11447 VDPWR.n2274 VDPWR.n2188 0.1603
R11448 VDPWR.n2274 VDPWR.n933 0.1603
R11449 VDPWR.n2841 VDPWR.n933 0.1603
R11450 VDPWR.n2841 VDPWR.n934 0.1603
R11451 VDPWR.n1733 VDPWR.n1732 0.158327
R11452 VDPWR.n1733 VDPWR.n1167 0.158327
R11453 VDPWR.n2454 VDPWR.n1167 0.158327
R11454 VDPWR.n2455 VDPWR.n2454 0.158327
R11455 VDPWR.n2455 VDPWR.n774 0.158327
R11456 VDPWR.n3050 VDPWR.n774 0.158327
R11457 VDPWR.n1332 VDPWR 0.158169
R11458 VDPWR VDPWR.n1813 0.158169
R11459 VDPWR.n2702 VDPWR 0.158169
R11460 VDPWR.n848 VDPWR 0.158169
R11461 VDPWR.n203 VDPWR.n202 0.155911
R11462 VDPWR.n2292 VDPWR.n2291 0.152881
R11463 VDPWR.n3072 VDPWR.n3071 0.152187
R11464 VDPWR.n756 VDPWR.n755 0.150053
R11465 VDPWR.n979 VDPWR.n957 0.143027
R11466 VDPWR.n1520 VDPWR 0.14207
R11467 VDPWR.n1295 VDPWR 0.14207
R11468 VDPWR.n1909 VDPWR 0.14207
R11469 VDPWR.n2920 VDPWR 0.14207
R11470 VDPWR.n1591 VDPWR 0.141725
R11471 VDPWR.n1785 VDPWR 0.141725
R11472 VDPWR.n2171 VDPWR 0.141725
R11473 VDPWR VDPWR.n1843 0.120408
R11474 VDPWR.n2219 VDPWR 0.120408
R11475 VDPWR VDPWR.n2718 0.120408
R11476 VDPWR.n848 VDPWR 0.120408
R11477 VDPWR.n586 VDPWR.n565 0.120292
R11478 VDPWR.n625 VDPWR.n566 0.120292
R11479 VDPWR.n618 VDPWR.n617 0.120292
R11480 VDPWR.n617 VDPWR.n591 0.120292
R11481 VDPWR.n613 VDPWR.n612 0.120292
R11482 VDPWR.n612 VDPWR.n611 0.120292
R11483 VDPWR.n608 VDPWR.n607 0.120292
R11484 VDPWR.n607 VDPWR.n606 0.120292
R11485 VDPWR.n603 VDPWR.n602 0.120292
R11486 VDPWR.n602 VDPWR.n596 0.120292
R11487 VDPWR.n598 VDPWR.n596 0.120292
R11488 VDPWR.n571 VDPWR.n567 0.120292
R11489 VDPWR.n584 VDPWR.n568 0.120292
R11490 VDPWR.n635 VDPWR.n562 0.120292
R11491 VDPWR.n636 VDPWR.n635 0.120292
R11492 VDPWR.n651 VDPWR.n537 0.120292
R11493 VDPWR.n647 VDPWR.n646 0.120292
R11494 VDPWR.n646 VDPWR.n541 0.120292
R11495 VDPWR.n557 VDPWR.n556 0.120292
R11496 VDPWR.n556 VDPWR.n548 0.120292
R11497 VDPWR.n551 VDPWR.n548 0.120292
R11498 VDPWR.n306 VDPWR.n285 0.120292
R11499 VDPWR.n345 VDPWR.n286 0.120292
R11500 VDPWR.n338 VDPWR.n337 0.120292
R11501 VDPWR.n337 VDPWR.n311 0.120292
R11502 VDPWR.n333 VDPWR.n332 0.120292
R11503 VDPWR.n332 VDPWR.n331 0.120292
R11504 VDPWR.n328 VDPWR.n327 0.120292
R11505 VDPWR.n327 VDPWR.n326 0.120292
R11506 VDPWR.n323 VDPWR.n322 0.120292
R11507 VDPWR.n322 VDPWR.n316 0.120292
R11508 VDPWR.n318 VDPWR.n316 0.120292
R11509 VDPWR.n291 VDPWR.n287 0.120292
R11510 VDPWR.n304 VDPWR.n288 0.120292
R11511 VDPWR.n355 VDPWR.n282 0.120292
R11512 VDPWR.n356 VDPWR.n355 0.120292
R11513 VDPWR.n371 VDPWR.n257 0.120292
R11514 VDPWR.n367 VDPWR.n366 0.120292
R11515 VDPWR.n366 VDPWR.n261 0.120292
R11516 VDPWR.n277 VDPWR.n276 0.120292
R11517 VDPWR.n276 VDPWR.n268 0.120292
R11518 VDPWR.n271 VDPWR.n268 0.120292
R11519 VDPWR.n1533 VDPWR.n1527 0.120292
R11520 VDPWR.n1546 VDPWR.n1500 0.120292
R11521 VDPWR.n1551 VDPWR.n1500 0.120292
R11522 VDPWR.n1552 VDPWR.n1551 0.120292
R11523 VDPWR.n1553 VDPWR.n1498 0.120292
R11524 VDPWR.n1558 VDPWR.n1498 0.120292
R11525 VDPWR.n1559 VDPWR.n1558 0.120292
R11526 VDPWR.n1565 VDPWR.n1496 0.120292
R11527 VDPWR.n1566 VDPWR.n1565 0.120292
R11528 VDPWR.n1567 VDPWR.n1566 0.120292
R11529 VDPWR.n1596 VDPWR.n1481 0.120292
R11530 VDPWR.n1597 VDPWR.n1596 0.120292
R11531 VDPWR.n1598 VDPWR.n1597 0.120292
R11532 VDPWR.n1598 VDPWR.n1479 0.120292
R11533 VDPWR.n1604 VDPWR.n1479 0.120292
R11534 VDPWR.n1622 VDPWR.n1472 0.120292
R11535 VDPWR VDPWR.n1622 0.120292
R11536 VDPWR.n1626 VDPWR.n1625 0.120292
R11537 VDPWR.n1626 VDPWR.n1469 0.120292
R11538 VDPWR.n1630 VDPWR.n1469 0.120292
R11539 VDPWR.n1631 VDPWR.n1630 0.120292
R11540 VDPWR.n1631 VDPWR.n1467 0.120292
R11541 VDPWR.n1635 VDPWR.n1467 0.120292
R11542 VDPWR.n1636 VDPWR.n1635 0.120292
R11543 VDPWR.n1642 VDPWR.n1636 0.120292
R11544 VDPWR.n1661 VDPWR.n1457 0.120292
R11545 VDPWR.n1668 VDPWR.n1457 0.120292
R11546 VDPWR.n1669 VDPWR.n1668 0.120292
R11547 VDPWR.n1670 VDPWR.n1669 0.120292
R11548 VDPWR.n1670 VDPWR.n1455 0.120292
R11549 VDPWR.n1675 VDPWR.n1455 0.120292
R11550 VDPWR.n1676 VDPWR.n1675 0.120292
R11551 VDPWR.n1696 VDPWR.n1695 0.120292
R11552 VDPWR.n1696 VDPWR.n1445 0.120292
R11553 VDPWR.n1700 VDPWR.n1445 0.120292
R11554 VDPWR.n1701 VDPWR.n1700 0.120292
R11555 VDPWR.n1701 VDPWR.n1443 0.120292
R11556 VDPWR.n1705 VDPWR.n1443 0.120292
R11557 VDPWR.n1706 VDPWR.n1705 0.120292
R11558 VDPWR.n1707 VDPWR.n1706 0.120292
R11559 VDPWR.n1707 VDPWR.n1441 0.120292
R11560 VDPWR.n1712 VDPWR.n1441 0.120292
R11561 VDPWR.n1303 VDPWR.n1302 0.120292
R11562 VDPWR.n1878 VDPWR.n1307 0.120292
R11563 VDPWR.n1874 VDPWR.n1307 0.120292
R11564 VDPWR.n1874 VDPWR.n1873 0.120292
R11565 VDPWR.n1870 VDPWR.n1869 0.120292
R11566 VDPWR.n1869 VDPWR.n1310 0.120292
R11567 VDPWR.n1864 VDPWR.n1310 0.120292
R11568 VDPWR.n1863 VDPWR.n1312 0.120292
R11569 VDPWR.n1858 VDPWR.n1312 0.120292
R11570 VDPWR.n1858 VDPWR.n1857 0.120292
R11571 VDPWR.n1833 VDPWR.n1832 0.120292
R11572 VDPWR.n1832 VDPWR.n1334 0.120292
R11573 VDPWR.n1827 VDPWR.n1334 0.120292
R11574 VDPWR.n1819 VDPWR.n1343 0.120292
R11575 VDPWR.n1814 VDPWR.n1343 0.120292
R11576 VDPWR.n1809 VDPWR.n1808 0.120292
R11577 VDPWR.n1808 VDPWR.n1356 0.120292
R11578 VDPWR.n1803 VDPWR.n1356 0.120292
R11579 VDPWR.n1803 VDPWR.n1802 0.120292
R11580 VDPWR.n1802 VDPWR.n1358 0.120292
R11581 VDPWR.n1798 VDPWR.n1358 0.120292
R11582 VDPWR.n1779 VDPWR.n1778 0.120292
R11583 VDPWR.n1778 VDPWR.n1777 0.120292
R11584 VDPWR.n1777 VDPWR.n1386 0.120292
R11585 VDPWR.n1773 VDPWR.n1386 0.120292
R11586 VDPWR.n1765 VDPWR.n1395 0.120292
R11587 VDPWR.n1761 VDPWR.n1395 0.120292
R11588 VDPWR.n1761 VDPWR.n1760 0.120292
R11589 VDPWR.n1760 VDPWR.n1410 0.120292
R11590 VDPWR.n1754 VDPWR.n1410 0.120292
R11591 VDPWR.n1754 VDPWR.n1753 0.120292
R11592 VDPWR.n1908 VDPWR.n1907 0.120292
R11593 VDPWR.n1937 VDPWR.n1271 0.120292
R11594 VDPWR.n1942 VDPWR.n1271 0.120292
R11595 VDPWR.n1943 VDPWR.n1942 0.120292
R11596 VDPWR.n1944 VDPWR.n1269 0.120292
R11597 VDPWR.n1949 VDPWR.n1269 0.120292
R11598 VDPWR.n1950 VDPWR.n1949 0.120292
R11599 VDPWR.n1956 VDPWR.n1267 0.120292
R11600 VDPWR.n1957 VDPWR.n1956 0.120292
R11601 VDPWR.n1958 VDPWR.n1957 0.120292
R11602 VDPWR.n2170 VDPWR.n1966 0.120292
R11603 VDPWR.n2160 VDPWR.n1966 0.120292
R11604 VDPWR.n2160 VDPWR.n2159 0.120292
R11605 VDPWR.n2159 VDPWR.n2158 0.120292
R11606 VDPWR.n2146 VDPWR.n1978 0.120292
R11607 VDPWR.n2141 VDPWR.n1978 0.120292
R11608 VDPWR.n2140 VDPWR.n2139 0.120292
R11609 VDPWR.n2139 VDPWR.n1989 0.120292
R11610 VDPWR.n2135 VDPWR.n1989 0.120292
R11611 VDPWR.n2135 VDPWR.n2134 0.120292
R11612 VDPWR.n2131 VDPWR.n2130 0.120292
R11613 VDPWR.n2130 VDPWR.n1994 0.120292
R11614 VDPWR.n2126 VDPWR.n1994 0.120292
R11615 VDPWR.n2114 VDPWR.n2113 0.120292
R11616 VDPWR.n2113 VDPWR.n2014 0.120292
R11617 VDPWR.n2108 VDPWR.n2014 0.120292
R11618 VDPWR.n2106 VDPWR.n2017 0.120292
R11619 VDPWR.n2100 VDPWR.n2099 0.120292
R11620 VDPWR.n2099 VDPWR.n2019 0.120292
R11621 VDPWR.n2077 VDPWR.n2038 0.120292
R11622 VDPWR.n2072 VDPWR.n2038 0.120292
R11623 VDPWR.n2229 VDPWR.n2224 0.120292
R11624 VDPWR.n2243 VDPWR.n2198 0.120292
R11625 VDPWR.n2247 VDPWR.n2198 0.120292
R11626 VDPWR.n2248 VDPWR.n2247 0.120292
R11627 VDPWR.n2253 VDPWR.n2196 0.120292
R11628 VDPWR.n2254 VDPWR.n2253 0.120292
R11629 VDPWR.n2259 VDPWR.n2258 0.120292
R11630 VDPWR.n2259 VDPWR.n2193 0.120292
R11631 VDPWR.n2263 VDPWR.n2193 0.120292
R11632 VDPWR.n2264 VDPWR.n2263 0.120292
R11633 VDPWR.n2297 VDPWR.n2296 0.120292
R11634 VDPWR.n2298 VDPWR.n1242 0.120292
R11635 VDPWR.n2304 VDPWR.n1242 0.120292
R11636 VDPWR.n2305 VDPWR.n2304 0.120292
R11637 VDPWR.n2324 VDPWR.n2323 0.120292
R11638 VDPWR.n2324 VDPWR.n1224 0.120292
R11639 VDPWR.n2331 VDPWR.n1224 0.120292
R11640 VDPWR.n2332 VDPWR.n2331 0.120292
R11641 VDPWR.n2338 VDPWR.n1221 0.120292
R11642 VDPWR.n2339 VDPWR.n2338 0.120292
R11643 VDPWR.n2339 VDPWR.n1218 0.120292
R11644 VDPWR.n2345 VDPWR.n1218 0.120292
R11645 VDPWR.n2372 VDPWR.n1201 0.120292
R11646 VDPWR.n2380 VDPWR.n1201 0.120292
R11647 VDPWR.n2381 VDPWR.n2380 0.120292
R11648 VDPWR.n2382 VDPWR.n2381 0.120292
R11649 VDPWR.n2382 VDPWR.n1198 0.120292
R11650 VDPWR.n2387 VDPWR.n1198 0.120292
R11651 VDPWR.n2388 VDPWR.n2387 0.120292
R11652 VDPWR.n2411 VDPWR.n2410 0.120292
R11653 VDPWR.n2411 VDPWR.n1182 0.120292
R11654 VDPWR.n2418 VDPWR.n1182 0.120292
R11655 VDPWR.n2419 VDPWR.n2418 0.120292
R11656 VDPWR.n2419 VDPWR.n1179 0.120292
R11657 VDPWR.n2425 VDPWR.n1179 0.120292
R11658 VDPWR.n2426 VDPWR.n2425 0.120292
R11659 VDPWR.n2427 VDPWR.n1177 0.120292
R11660 VDPWR.n2434 VDPWR.n1177 0.120292
R11661 VDPWR.n2567 VDPWR.n2566 0.120292
R11662 VDPWR.n2562 VDPWR.n987 0.120292
R11663 VDPWR.n2562 VDPWR.n2561 0.120292
R11664 VDPWR.n2561 VDPWR.n989 0.120292
R11665 VDPWR.n996 VDPWR.n989 0.120292
R11666 VDPWR.n2553 VDPWR.n996 0.120292
R11667 VDPWR.n2552 VDPWR.n2551 0.120292
R11668 VDPWR.n2551 VDPWR.n997 0.120292
R11669 VDPWR.n1050 VDPWR.n1049 0.120292
R11670 VDPWR.n1057 VDPWR.n1056 0.120292
R11671 VDPWR.n1064 VDPWR.n1063 0.120292
R11672 VDPWR.n1089 VDPWR.n1088 0.120292
R11673 VDPWR.n1095 VDPWR.n1033 0.120292
R11674 VDPWR.n1096 VDPWR.n1095 0.120292
R11675 VDPWR.n1097 VDPWR.n1096 0.120292
R11676 VDPWR.n1097 VDPWR.n1030 0.120292
R11677 VDPWR.n1102 VDPWR.n1030 0.120292
R11678 VDPWR.n2527 VDPWR.n2526 0.120292
R11679 VDPWR.n2526 VDPWR.n1134 0.120292
R11680 VDPWR.n2521 VDPWR.n1134 0.120292
R11681 VDPWR.n2521 VDPWR.n2520 0.120292
R11682 VDPWR.n2520 VDPWR.n1139 0.120292
R11683 VDPWR.n2516 VDPWR.n1139 0.120292
R11684 VDPWR.n2516 VDPWR.n2515 0.120292
R11685 VDPWR.n2515 VDPWR.n1142 0.120292
R11686 VDPWR.n2501 VDPWR.n1150 0.120292
R11687 VDPWR.n2495 VDPWR.n1150 0.120292
R11688 VDPWR.n2494 VDPWR.n2493 0.120292
R11689 VDPWR.n2493 VDPWR.n1159 0.120292
R11690 VDPWR.n2489 VDPWR.n2488 0.120292
R11691 VDPWR.n2488 VDPWR.n1163 0.120292
R11692 VDPWR.n2484 VDPWR.n1163 0.120292
R11693 VDPWR.n2484 VDPWR.n2483 0.120292
R11694 VDPWR.n2812 VDPWR.n946 0.120292
R11695 VDPWR.n2813 VDPWR.n2812 0.120292
R11696 VDPWR.n2814 VDPWR.n2813 0.120292
R11697 VDPWR.n2814 VDPWR.n942 0.120292
R11698 VDPWR.n2819 VDPWR.n942 0.120292
R11699 VDPWR.n2820 VDPWR.n2819 0.120292
R11700 VDPWR.n2821 VDPWR.n2820 0.120292
R11701 VDPWR.n2821 VDPWR.n940 0.120292
R11702 VDPWR.n2825 VDPWR.n940 0.120292
R11703 VDPWR.n2826 VDPWR.n2825 0.120292
R11704 VDPWR.n2827 VDPWR.n2826 0.120292
R11705 VDPWR.n2855 VDPWR.n924 0.120292
R11706 VDPWR.n2856 VDPWR.n2855 0.120292
R11707 VDPWR.n2857 VDPWR.n2856 0.120292
R11708 VDPWR.n2857 VDPWR.n921 0.120292
R11709 VDPWR.n2863 VDPWR.n921 0.120292
R11710 VDPWR.n2864 VDPWR.n2863 0.120292
R11711 VDPWR.n2865 VDPWR.n2864 0.120292
R11712 VDPWR.n2865 VDPWR.n918 0.120292
R11713 VDPWR.n905 VDPWR.n902 0.120292
R11714 VDPWR.n2888 VDPWR.n902 0.120292
R11715 VDPWR.n2890 VDPWR.n899 0.120292
R11716 VDPWR.n899 VDPWR.n896 0.120292
R11717 VDPWR.n2928 VDPWR.n881 0.120292
R11718 VDPWR.n2929 VDPWR.n2928 0.120292
R11719 VDPWR.n2935 VDPWR.n878 0.120292
R11720 VDPWR.n2936 VDPWR.n2935 0.120292
R11721 VDPWR.n2937 VDPWR.n2936 0.120292
R11722 VDPWR.n2997 VDPWR.n2996 0.120292
R11723 VDPWR.n2996 VDPWR.n2944 0.120292
R11724 VDPWR.n2992 VDPWR.n2944 0.120292
R11725 VDPWR.n2992 VDPWR.n2991 0.120292
R11726 VDPWR.n2991 VDPWR.n2990 0.120292
R11727 VDPWR.n2987 VDPWR.n2986 0.120292
R11728 VDPWR.n2986 VDPWR.n2948 0.120292
R11729 VDPWR.n2644 VDPWR.n2627 0.120292
R11730 VDPWR.n2798 VDPWR.n2621 0.120292
R11731 VDPWR.n2791 VDPWR.n2657 0.120292
R11732 VDPWR.n2784 VDPWR.n2783 0.120292
R11733 VDPWR.n2779 VDPWR.n2661 0.120292
R11734 VDPWR.n2755 VDPWR.n2677 0.120292
R11735 VDPWR.n2750 VDPWR.n2677 0.120292
R11736 VDPWR.n2750 VDPWR.n2749 0.120292
R11737 VDPWR.n2731 VDPWR.n2730 0.120292
R11738 VDPWR.n2730 VDPWR.n2729 0.120292
R11739 VDPWR.n2729 VDPWR.n2697 0.120292
R11740 VDPWR.n2723 VDPWR.n2722 0.120292
R11741 VDPWR.n3028 VDPWR.n3027 0.120292
R11742 VDPWR.n3027 VDPWR.n3026 0.120292
R11743 VDPWR.n3026 VDPWR.n790 0.120292
R11744 VDPWR.n3022 VDPWR.n3021 0.120292
R11745 VDPWR.n858 VDPWR.n857 0.120292
R11746 VDPWR.n857 VDPWR.n812 0.120292
R11747 VDPWR.n49 VDPWR.n28 0.120292
R11748 VDPWR.n88 VDPWR.n29 0.120292
R11749 VDPWR.n81 VDPWR.n80 0.120292
R11750 VDPWR.n80 VDPWR.n54 0.120292
R11751 VDPWR.n76 VDPWR.n75 0.120292
R11752 VDPWR.n75 VDPWR.n74 0.120292
R11753 VDPWR.n71 VDPWR.n70 0.120292
R11754 VDPWR.n70 VDPWR.n69 0.120292
R11755 VDPWR.n66 VDPWR.n65 0.120292
R11756 VDPWR.n65 VDPWR.n59 0.120292
R11757 VDPWR.n61 VDPWR.n59 0.120292
R11758 VDPWR.n34 VDPWR.n30 0.120292
R11759 VDPWR.n47 VDPWR.n31 0.120292
R11760 VDPWR.n98 VDPWR.n25 0.120292
R11761 VDPWR.n99 VDPWR.n98 0.120292
R11762 VDPWR.n114 VDPWR.n0 0.120292
R11763 VDPWR.n110 VDPWR.n109 0.120292
R11764 VDPWR.n109 VDPWR.n4 0.120292
R11765 VDPWR.n20 VDPWR.n19 0.120292
R11766 VDPWR.n19 VDPWR.n11 0.120292
R11767 VDPWR.n14 VDPWR.n11 0.120292
R11768 VDPWR.n626 VDPWR.n565 0.11899
R11769 VDPWR.n346 VDPWR.n285 0.11899
R11770 VDPWR.n89 VDPWR.n28 0.11899
R11771 VDPWR.n3052 VDPWR.n770 0.116902
R11772 VDPWR.n3054 VDPWR 0.115443
R11773 VDPWR.n2169 VDPWR.n2168 0.113774
R11774 VDPWR.n2168 VDPWR.n2163 0.113774
R11775 VDPWR.n756 VDPWR.n117 0.113371
R11776 VDPWR.n460 VDPWR.n402 0.1125
R11777 VDPWR.n1714 VDPWR.n1712 0.112479
R11778 VDPWR.n2436 VDPWR.n2434 0.112479
R11779 VDPWR.n2483 VDPWR.n2482 0.112479
R11780 VDPWR.n2980 VDPWR.n2979 0.112479
R11781 VDPWR.n843 VDPWR.n842 0.112479
R11782 VDPWR.n1605 VDPWR.n1604 0.107271
R11783 VDPWR.n1827 VDPWR.n1826 0.107271
R11784 VDPWR.n2155 VDPWR.n2154 0.107271
R11785 VDPWR.n2305 VDPWR.n1232 0.107271
R11786 VDPWR.n1064 VDPWR.n1041 0.107271
R11787 VDPWR.n918 VDPWR.n916 0.107271
R11788 VDPWR.n3044 VDPWR.n776 0.10625
R11789 VDPWR.n3045 VDPWR.n775 0.10625
R11790 VDPWR.n2335 VDPWR.n2334 0.105418
R11791 VDPWR.n2417 VDPWR.n2416 0.105418
R11792 VDPWR.n1519 VDPWR 0.105238
R11793 VDPWR.n1294 VDPWR 0.105238
R11794 VDPWR.n1916 VDPWR 0.105238
R11795 VDPWR.n2218 VDPWR 0.105238
R11796 VDPWR.n969 VDPWR 0.105238
R11797 VDPWR.n2602 VDPWR 0.105238
R11798 VDPWR.n2638 VDPWR 0.105238
R11799 VDPWR.n376 VDPWR.n254 0.103147
R11800 VDPWR.n2075 VDPWR.n2074 0.102087
R11801 VDPWR.n1123 VDPWR.n1122 0.102087
R11802 VDPWR.n2985 VDPWR.n2984 0.102087
R11803 VDPWR.n571 VDPWR 0.0981562
R11804 VDPWR.n291 VDPWR 0.0981562
R11805 VDPWR VDPWR.n1496 0.0981562
R11806 VDPWR.n1590 VDPWR 0.0981562
R11807 VDPWR.n1625 VDPWR 0.0981562
R11808 VDPWR.n1656 VDPWR 0.0981562
R11809 VDPWR VDPWR.n1863 0.0981562
R11810 VDPWR.n1845 VDPWR 0.0981562
R11811 VDPWR.n1809 VDPWR 0.0981562
R11812 VDPWR VDPWR.n1790 0.0981562
R11813 VDPWR.n1779 VDPWR 0.0981562
R11814 VDPWR VDPWR.n1267 0.0981562
R11815 VDPWR VDPWR.n2172 0.0981562
R11816 VDPWR VDPWR.n2170 0.0981562
R11817 VDPWR VDPWR.n2140 0.0981562
R11818 VDPWR.n2131 VDPWR 0.0981562
R11819 VDPWR VDPWR.n2117 0.0981562
R11820 VDPWR VDPWR.n2106 0.0981562
R11821 VDPWR VDPWR.n2077 0.0981562
R11822 VDPWR.n2258 VDPWR 0.0981562
R11823 VDPWR.n2284 VDPWR 0.0981562
R11824 VDPWR.n2290 VDPWR 0.0981562
R11825 VDPWR.n2296 VDPWR 0.0981562
R11826 VDPWR VDPWR.n1221 0.0981562
R11827 VDPWR.n2372 VDPWR 0.0981562
R11828 VDPWR.n2567 VDPWR 0.0981562
R11829 VDPWR.n1056 VDPWR 0.0981562
R11830 VDPWR VDPWR.n1033 0.0981562
R11831 VDPWR VDPWR.n905 0.0981562
R11832 VDPWR.n2642 VDPWR 0.0981562
R11833 VDPWR VDPWR.n2791 0.0981562
R11834 VDPWR VDPWR.n2779 0.0981562
R11835 VDPWR VDPWR.n2755 0.0981562
R11836 VDPWR.n2682 VDPWR 0.0981562
R11837 VDPWR VDPWR.n2723 0.0981562
R11838 VDPWR.n3028 VDPWR 0.0981562
R11839 VDPWR VDPWR.n3017 0.0981562
R11840 VDPWR VDPWR.n843 0.0981562
R11841 VDPWR.n34 VDPWR 0.0981562
R11842 VDPWR.n3043 VDPWR.n3042 0.0977722
R11843 VDPWR.n2741 VDPWR.n776 0.0977722
R11844 VDPWR.n2769 VDPWR.n2618 0.0977722
R11845 VDPWR.n3014 VDPWR.n769 0.0977722
R11846 VDPWR.n1063 VDPWR 0.0968542
R11847 VDPWR VDPWR.n2980 0.0968542
R11848 VDPWR.n627 VDPWR 0.0955521
R11849 VDPWR.n347 VDPWR 0.0955521
R11850 VDPWR.n90 VDPWR 0.0955521
R11851 VDPWR.n2839 VDPWR.n2838 0.0950946
R11852 VDPWR.n2843 VDPWR.n931 0.0950946
R11853 VDPWR.n2877 VDPWR.n2876 0.0950946
R11854 VDPWR.n2881 VDPWR.n911 0.0950946
R11855 VDPWR.n2742 VDPWR.n2686 0.0950946
R11856 VDPWR.n2736 VDPWR.n2688 0.0950946
R11857 VDPWR.n1640 VDPWR.n1638 0.0950946
R11858 VDPWR.n1654 VDPWR.n1461 0.0950946
R11859 VDPWR.n1608 VDPWR.n1607 0.0950946
R11860 VDPWR.n1616 VDPWR.n1475 0.0950946
R11861 VDPWR.n1579 VDPWR.n1578 0.0950946
R11862 VDPWR.n1583 VDPWR.n1488 0.0950946
R11863 VDPWR.n1531 VDPWR.n1529 0.0950946
R11864 VDPWR.n1544 VDPWR.n1503 0.0950946
R11865 VDPWR.n1717 VDPWR.n1715 0.0950946
R11866 VDPWR.n1728 VDPWR.n1433 0.0950946
R11867 VDPWR.n1679 VDPWR.n1677 0.0950946
R11868 VDPWR.n1690 VDPWR.n1449 0.0950946
R11869 VDPWR.n1796 VDPWR.n1361 0.0950946
R11870 VDPWR.n1792 VDPWR.n1365 0.0950946
R11871 VDPWR.n1825 VDPWR.n1337 0.0950946
R11872 VDPWR.n1821 VDPWR.n1341 0.0950946
R11873 VDPWR.n1855 VDPWR.n1315 0.0950946
R11874 VDPWR.n1850 VDPWR.n1318 0.0950946
R11875 VDPWR.n1892 VDPWR.n1891 0.0950946
R11876 VDPWR.n1884 VDPWR.n1883 0.0950946
R11877 VDPWR.n1739 VDPWR.n1737 0.0950946
R11878 VDPWR.n1746 VDPWR.n1431 0.0950946
R11879 VDPWR.n1771 VDPWR.n1390 0.0950946
R11880 VDPWR.n1767 VDPWR.n1394 0.0950946
R11881 VDPWR.n2124 VDPWR.n1997 0.0950946
R11882 VDPWR.n2119 VDPWR.n2000 0.0950946
R11883 VDPWR.n2153 VDPWR.n1973 0.0950946
R11884 VDPWR.n2148 VDPWR.n1976 0.0950946
R11885 VDPWR.n2186 VDPWR.n2185 0.0950946
R11886 VDPWR.n2179 VDPWR.n1264 0.0950946
R11887 VDPWR.n1931 VDPWR.n1930 0.0950946
R11888 VDPWR.n1935 VDPWR.n1274 0.0950946
R11889 VDPWR.n2070 VDPWR.n2045 0.0950946
R11890 VDPWR.n2060 VDPWR.n2058 0.0950946
R11891 VDPWR.n2093 VDPWR.n2022 0.0950946
R11892 VDPWR.n2087 VDPWR.n2025 0.0950946
R11893 VDPWR.n2509 VDPWR.n1146 0.0950946
R11894 VDPWR.n2503 VDPWR.n1149 0.0950946
R11895 VDPWR.n3009 VDPWR.n3008 0.0950946
R11896 VDPWR.n3002 VDPWR.n874 0.0950946
R11897 VDPWR.n2399 VDPWR.n2398 0.0950946
R11898 VDPWR.n2404 VDPWR.n2403 0.0950946
R11899 VDPWR.n2317 VDPWR.n2316 0.0950946
R11900 VDPWR.n2321 VDPWR.n1228 0.0950946
R11901 VDPWR.n2272 VDPWR.n2271 0.0950946
R11902 VDPWR.n2277 VDPWR.n2276 0.0950946
R11903 VDPWR.n2227 VDPWR.n2225 0.0950946
R11904 VDPWR.n2241 VDPWR.n2201 0.0950946
R11905 VDPWR.n2439 VDPWR.n2437 0.0950946
R11906 VDPWR.n2450 VDPWR.n1169 0.0950946
R11907 VDPWR.n2357 VDPWR.n2356 0.0950946
R11908 VDPWR.n2361 VDPWR.n1208 0.0950946
R11909 VDPWR.n1113 VDPWR.n1111 0.0950946
R11910 VDPWR.n1130 VDPWR.n1023 0.0950946
R11911 VDPWR.n2913 VDPWR.n2912 0.0950946
R11912 VDPWR.n2917 VDPWR.n885 0.0950946
R11913 VDPWR.n2707 VDPWR.n781 0.0950946
R11914 VDPWR.n3040 VDPWR.n780 0.0950946
R11915 VDPWR.n1072 VDPWR.n1040 0.0950946
R11916 VDPWR.n1080 VDPWR.n1079 0.0950946
R11917 VDPWR.n2543 VDPWR.n1004 0.0950946
R11918 VDPWR.n2537 VDPWR.n1007 0.0950946
R11919 VDPWR.n2481 VDPWR.n1166 0.0950946
R11920 VDPWR.n2471 VDPWR.n2469 0.0950946
R11921 VDPWR.n2580 VDPWR.n2579 0.0950946
R11922 VDPWR.n2573 VDPWR.n2572 0.0950946
R11923 VDPWR.n2610 VDPWR.n2609 0.0950946
R11924 VDPWR.n2806 VDPWR.n2805 0.0950946
R11925 VDPWR.n2978 VDPWR.n2952 0.0950946
R11926 VDPWR.n2973 VDPWR.n2955 0.0950946
R11927 VDPWR.n2771 VDPWR.n2665 0.0950946
R11928 VDPWR.n2767 VDPWR.n2667 0.0950946
R11929 VDPWR.n2623 VDPWR.n2617 0.0950946
R11930 VDPWR.n2800 VDPWR.n2619 0.0950946
R11931 VDPWR.n841 VDPWR.n840 0.0950946
R11932 VDPWR.n833 VDPWR.n771 0.0950946
R11933 VDPWR.n3015 VDPWR.n798 0.0950946
R11934 VDPWR.n865 VDPWR.n800 0.0950946
R11935 VDPWR VDPWR.n2219 0.0930646
R11936 VDPWR.n585 VDPWR.n567 0.0916458
R11937 VDPWR.n305 VDPWR.n287 0.0916458
R11938 VDPWR.n48 VDPWR.n30 0.0916458
R11939 VDPWR.n3044 VDPWR.n3043 0.0913766
R11940 VDPWR.n3046 VDPWR.n3045 0.0913766
R11941 VDPWR.n914 VDPWR 0.08745
R11942 VDPWR.n3109 VDPWR.n758 0.08675
R11943 VDPWR.n3087 VDPWR.n3072 0.0848934
R11944 VDPWR.n3103 VDPWR.n3088 0.0844041
R11945 VDPWR.n1532 VDPWR.n1528 0.0838333
R11946 VDPWR.n1545 VDPWR.n1502 0.0838333
R11947 VDPWR.n1577 VDPWR.n1576 0.0838333
R11948 VDPWR.n1611 VDPWR.n1474 0.0838333
R11949 VDPWR.n1641 VDPWR.n1637 0.0838333
R11950 VDPWR.n1685 VDPWR.n1452 0.0838333
R11951 VDPWR.n1727 VDPWR.n1726 0.0838333
R11952 VDPWR.n1890 VDPWR.n1279 0.0838333
R11953 VDPWR.n1885 VDPWR.n1879 0.0838333
R11954 VDPWR.n1324 VDPWR.n1322 0.0838333
R11955 VDPWR.n1350 VDPWR.n1346 0.0838333
R11956 VDPWR.n1797 VDPWR.n1360 0.0838333
R11957 VDPWR.n1401 VDPWR.n1397 0.0838333
R11958 VDPWR.n1747 VDPWR.n1430 0.0838333
R11959 VDPWR.n1929 VDPWR.n1896 0.0838333
R11960 VDPWR.n1936 VDPWR.n1273 0.0838333
R11961 VDPWR.n2184 VDPWR.n2183 0.0838333
R11962 VDPWR.n1983 VDPWR.n1981 0.0838333
R11963 VDPWR.n2125 VDPWR.n1996 0.0838333
R11964 VDPWR.n2061 VDPWR.n2050 0.0838333
R11965 VDPWR.n2228 VDPWR.n2204 0.0838333
R11966 VDPWR.n2242 VDPWR.n2200 0.0838333
R11967 VDPWR.n2270 VDPWR.n2269 0.0838333
R11968 VDPWR.n1238 VDPWR.n1235 0.0838333
R11969 VDPWR.n2355 VDPWR.n1212 0.0838333
R11970 VDPWR.n2397 VDPWR.n2396 0.0838333
R11971 VDPWR.n2449 VDPWR.n2448 0.0838333
R11972 VDPWR.n2578 VDPWR.n957 0.0838333
R11973 VDPWR.n2544 VDPWR.n1003 0.0838333
R11974 VDPWR.n1081 VDPWR.n1037 0.0838333
R11975 VDPWR.n1114 VDPWR.n1110 0.0838333
R11976 VDPWR.n2510 VDPWR.n1145 0.0838333
R11977 VDPWR.n2472 VDPWR.n2460 0.0838333
R11978 VDPWR.n2608 VDPWR.n2585 0.0838333
R11979 VDPWR.n2807 VDPWR.n951 0.0838333
R11980 VDPWR.n2873 VDPWR.n910 0.0838333
R11981 VDPWR.n2911 VDPWR.n889 0.0838333
R11982 VDPWR.n3007 VDPWR.n3006 0.0838333
R11983 VDPWR.n2972 VDPWR.n2956 0.0838333
R11984 VDPWR.n2626 VDPWR.n2624 0.0838333
R11985 VDPWR.n2799 VDPWR.n2620 0.0838333
R11986 VDPWR.n2738 VDPWR.n2737 0.0838333
R11987 VDPWR.n835 VDPWR.n834 0.0838333
R11988 VDPWR.n3050 VDPWR.n3049 0.0828951
R11989 VDPWR.n3012 VDPWR 0.08275
R11990 VDPWR.n777 VDPWR 0.08275
R11991 VDPWR.n2614 VDPWR 0.08275
R11992 VDPWR.n2612 VDPWR 0.08275
R11993 VDPWR VDPWR.n2030 0.082648
R11994 VDPWR VDPWR.n2896 0.082648
R11995 VDPWR.n1843 VDPWR 0.082648
R11996 VDPWR VDPWR.n1332 0.082648
R11997 VDPWR.n1813 VDPWR 0.082648
R11998 VDPWR.n2718 VDPWR 0.082648
R11999 VDPWR VDPWR.n2702 0.082648
R12000 VDPWR.n3012 VDPWR 0.0822391
R12001 VDPWR.n777 VDPWR 0.0822391
R12002 VDPWR.n2614 VDPWR 0.0812362
R12003 VDPWR.n1585 VDPWR.n1584 0.0812292
R12004 VDPWR.n1618 VDPWR.n1617 0.0812292
R12005 VDPWR.n1465 VDPWR.n1460 0.0812292
R12006 VDPWR.n1684 VDPWR.n1448 0.0812292
R12007 VDPWR.n1719 VDPWR.n1436 0.0812292
R12008 VDPWR.n1849 VDPWR.n1848 0.0812292
R12009 VDPWR.n1820 VDPWR.n1342 0.0812292
R12010 VDPWR.n1373 VDPWR.n1366 0.0812292
R12011 VDPWR.n1406 VDPWR.n1405 0.0812292
R12012 VDPWR.n1741 VDPWR.n1426 0.0812292
R12013 VDPWR.n2173 VDPWR.n1265 0.0812292
R12014 VDPWR.n2147 VDPWR.n1977 0.0812292
R12015 VDPWR.n2008 VDPWR.n2001 0.0812292
R12016 VDPWR.n2028 VDPWR.n2027 0.0812292
R12017 VDPWR.n2065 VDPWR.n2064 0.0812292
R12018 VDPWR.n2283 VDPWR.n1252 0.0812292
R12019 VDPWR.n2322 VDPWR.n1227 0.0812292
R12020 VDPWR.n2363 VDPWR.n1207 0.0812292
R12021 VDPWR.n2405 VDPWR.n1188 0.0812292
R12022 VDPWR.n2441 VDPWR.n1172 0.0812292
R12023 VDPWR.n2536 VDPWR.n2535 0.0812292
R12024 VDPWR.n1082 VDPWR.n1035 0.0812292
R12025 VDPWR.n1027 VDPWR.n1022 0.0812292
R12026 VDPWR.n1153 VDPWR.n1152 0.0812292
R12027 VDPWR.n2476 VDPWR.n2475 0.0812292
R12028 VDPWR.n2845 VDPWR.n2844 0.0812292
R12029 VDPWR.n2906 VDPWR.n884 0.0812292
R12030 VDPWR.n3001 VDPWR.n873 0.0812292
R12031 VDPWR.n2966 VDPWR.n2965 0.0812292
R12032 VDPWR.n2762 VDPWR.n2670 0.0812292
R12033 VDPWR.n2735 VDPWR.n2691 0.0812292
R12034 VDPWR.n3039 VDPWR.n3038 0.0812292
R12035 VDPWR.n829 VDPWR.n823 0.0812292
R12036 VDPWR.n535 VDPWR 0.0800455
R12037 VDPWR VDPWR.n2612 0.0797771
R12038 VDPWR.n1573 VDPWR.n1494 0.0760208
R12039 VDPWR.n1649 VDPWR.n1464 0.0760208
R12040 VDPWR.n1326 VDPWR.n1325 0.0760208
R12041 VDPWR.n1372 VDPWR.n1368 0.0760208
R12042 VDPWR.n1766 VDPWR.n1765 0.0760208
R12043 VDPWR.n2178 VDPWR.n1263 0.0760208
R12044 VDPWR.n2007 VDPWR.n2005 0.0760208
R12045 VDPWR.n2086 VDPWR.n2085 0.0760208
R12046 VDPWR.n2278 VDPWR.n1254 0.0760208
R12047 VDPWR.n2354 VDPWR.n1216 0.0760208
R12048 VDPWR.n2410 VDPWR.n1185 0.0760208
R12049 VDPWR.n1013 VDPWR.n1012 0.0760208
R12050 VDPWR.n1125 VDPWR.n1026 0.0760208
R12051 VDPWR.n2502 VDPWR.n2501 0.0760208
R12052 VDPWR.n2833 VDPWR.n2832 0.0760208
R12053 VDPWR.n2910 VDPWR.n893 0.0760208
R12054 VDPWR.n2997 VDPWR.n875 0.0760208
R12055 VDPWR.n859 VDPWR.n802 0.0760208
R12056 VDPWR.n752 VDPWR 0.0710357
R12057 VDPWR.n1539 VDPWR.n1506 0.0708125
R12058 VDPWR.n1609 VDPWR.n1478 0.0708125
R12059 VDPWR.n1889 VDPWR.n1281 0.0708125
R12060 VDPWR.n1345 VDPWR.n1336 0.0708125
R12061 VDPWR.n1773 VDPWR.n1772 0.0708125
R12062 VDPWR.n1928 VDPWR.n1900 0.0708125
R12063 VDPWR.n1980 VDPWR.n1972 0.0708125
R12064 VDPWR.n2021 VDPWR.n2019 0.0708125
R12065 VDPWR.n2236 VDPWR.n2234 0.0708125
R12066 VDPWR.n2315 VDPWR.n1234 0.0708125
R12067 VDPWR.n2388 VDPWR.n1194 0.0708125
R12068 VDPWR.n2577 VDPWR.n959 0.0708125
R12069 VDPWR.n1071 VDPWR.n1069 0.0708125
R12070 VDPWR.n1144 VDPWR.n1142 0.0708125
R12071 VDPWR.n2607 VDPWR.n950 0.0708125
R12072 VDPWR.n2875 VDPWR.n2870 0.0708125
R12073 VDPWR.n2937 VDPWR.n870 0.0708125
R12074 VDPWR.n3017 VDPWR.n3016 0.0708125
R12075 VDPWR.n2835 VDPWR.n937 0.0680676
R12076 VDPWR.n2835 VDPWR.n2834 0.0680676
R12077 VDPWR.n2872 VDPWR.n917 0.0680676
R12078 VDPWR.n2872 VDPWR.n2871 0.0680676
R12079 VDPWR.n2740 VDPWR.n2739 0.0680676
R12080 VDPWR.n2739 VDPWR.n2687 0.0680676
R12081 VDPWR.n1650 VDPWR.n1463 0.0680676
R12082 VDPWR.n1651 VDPWR.n1650 0.0680676
R12083 VDPWR.n1612 VDPWR.n1477 0.0680676
R12084 VDPWR.n1613 VDPWR.n1612 0.0680676
R12085 VDPWR.n1575 VDPWR.n1492 0.0680676
R12086 VDPWR.n1575 VDPWR.n1574 0.0680676
R12087 VDPWR.n1540 VDPWR.n1505 0.0680676
R12088 VDPWR.n1541 VDPWR.n1540 0.0680676
R12089 VDPWR.n1716 VDPWR.n1435 0.0680676
R12090 VDPWR.n1729 VDPWR.n1435 0.0680676
R12091 VDPWR.n1686 VDPWR.n1451 0.0680676
R12092 VDPWR.n1687 VDPWR.n1686 0.0680676
R12093 VDPWR.n1371 VDPWR.n1369 0.0680676
R12094 VDPWR.n1371 VDPWR.n1370 0.0680676
R12095 VDPWR.n1349 VDPWR.n1347 0.0680676
R12096 VDPWR.n1349 VDPWR.n1348 0.0680676
R12097 VDPWR.n1323 VDPWR.n1316 0.0680676
R12098 VDPWR.n1323 VDPWR.n1317 0.0680676
R12099 VDPWR.n1880 VDPWR.n1280 0.0680676
R12100 VDPWR.n1882 VDPWR.n1880 0.0680676
R12101 VDPWR.n1742 VDPWR.n1740 0.0680676
R12102 VDPWR.n1743 VDPWR.n1742 0.0680676
R12103 VDPWR.n1400 VDPWR.n1398 0.0680676
R12104 VDPWR.n1400 VDPWR.n1399 0.0680676
R12105 VDPWR.n2006 VDPWR.n1998 0.0680676
R12106 VDPWR.n2006 VDPWR.n1999 0.0680676
R12107 VDPWR.n1982 VDPWR.n1974 0.0680676
R12108 VDPWR.n1982 VDPWR.n1975 0.0680676
R12109 VDPWR.n2182 VDPWR.n1261 0.0680676
R12110 VDPWR.n2182 VDPWR.n2181 0.0680676
R12111 VDPWR.n1899 VDPWR.n1897 0.0680676
R12112 VDPWR.n1899 VDPWR.n1898 0.0680676
R12113 VDPWR.n2067 VDPWR.n2066 0.0680676
R12114 VDPWR.n2066 VDPWR.n2047 0.0680676
R12115 VDPWR.n2092 VDPWR.n2023 0.0680676
R12116 VDPWR.n2024 VDPWR.n2023 0.0680676
R12117 VDPWR.n2508 VDPWR.n1147 0.0680676
R12118 VDPWR.n1148 VDPWR.n1147 0.0680676
R12119 VDPWR.n3005 VDPWR.n871 0.0680676
R12120 VDPWR.n3005 VDPWR.n3004 0.0680676
R12121 VDPWR.n2395 VDPWR.n1195 0.0680676
R12122 VDPWR.n2395 VDPWR.n1189 0.0680676
R12123 VDPWR.n1237 VDPWR.n1233 0.0680676
R12124 VDPWR.n1237 VDPWR.n1236 0.0680676
R12125 VDPWR.n2268 VDPWR.n2191 0.0680676
R12126 VDPWR.n2268 VDPWR.n1255 0.0680676
R12127 VDPWR.n2237 VDPWR.n2203 0.0680676
R12128 VDPWR.n2238 VDPWR.n2237 0.0680676
R12129 VDPWR.n2438 VDPWR.n1171 0.0680676
R12130 VDPWR.n2451 VDPWR.n1171 0.0680676
R12131 VDPWR.n1215 VDPWR.n1213 0.0680676
R12132 VDPWR.n1215 VDPWR.n1214 0.0680676
R12133 VDPWR.n1126 VDPWR.n1025 0.0680676
R12134 VDPWR.n1127 VDPWR.n1126 0.0680676
R12135 VDPWR.n892 VDPWR.n890 0.0680676
R12136 VDPWR.n892 VDPWR.n891 0.0680676
R12137 VDPWR.n782 VDPWR.n779 0.0680676
R12138 VDPWR.n3041 VDPWR.n782 0.0680676
R12139 VDPWR.n1074 VDPWR.n1073 0.0680676
R12140 VDPWR.n1073 VDPWR.n1038 0.0680676
R12141 VDPWR.n2542 VDPWR.n1005 0.0680676
R12142 VDPWR.n1006 VDPWR.n1005 0.0680676
R12143 VDPWR.n2478 VDPWR.n2477 0.0680676
R12144 VDPWR.n2477 VDPWR.n2457 0.0680676
R12145 VDPWR.n980 VDPWR.n958 0.0680676
R12146 VDPWR.n982 VDPWR.n980 0.0680676
R12147 VDPWR.n2587 VDPWR.n2586 0.0680676
R12148 VDPWR.n2586 VDPWR.n952 0.0680676
R12149 VDPWR.n2964 VDPWR.n2953 0.0680676
R12150 VDPWR.n2964 VDPWR.n2954 0.0680676
R12151 VDPWR.n2770 VDPWR.n2666 0.0680676
R12152 VDPWR.n2768 VDPWR.n2666 0.0680676
R12153 VDPWR.n2649 VDPWR.n2616 0.0680676
R12154 VDPWR.n2649 VDPWR.n2615 0.0680676
R12155 VDPWR.n822 VDPWR.n772 0.0680676
R12156 VDPWR.n822 VDPWR.n773 0.0680676
R12157 VDPWR.n801 VDPWR.n799 0.0680676
R12158 VDPWR.n866 VDPWR.n801 0.0680676
R12159 VDPWR.n1567 VDPWR.n1491 0.0656042
R12160 VDPWR.n1857 VDPWR.n1856 0.0656042
R12161 VDPWR.n1958 VDPWR.n1260 0.0656042
R12162 VDPWR.n2264 VDPWR.n2190 0.0656042
R12163 VDPWR.n1002 VDPWR.n997 0.0656042
R12164 VDPWR.n2827 VDPWR.n936 0.0656042
R12165 VDPWR.n2664 VDPWR.n2661 0.0656042
R12166 VDPWR.n717 VDPWR 0.06425
R12167 VDPWR.n701 VDPWR 0.06425
R12168 VDPWR.n685 VDPWR 0.06425
R12169 VDPWR.n669 VDPWR 0.06425
R12170 VDPWR.n528 VDPWR 0.06425
R12171 VDPWR.n512 VDPWR 0.06425
R12172 VDPWR.n496 VDPWR 0.06425
R12173 VDPWR.n480 VDPWR 0.06425
R12174 VDPWR.n464 VDPWR 0.06425
R12175 VDPWR.n388 VDPWR 0.06425
R12176 VDPWR.n400 VDPWR 0.06425
R12177 VDPWR.n458 VDPWR 0.06425
R12178 VDPWR.n442 VDPWR 0.06425
R12179 VDPWR.n426 VDPWR 0.06425
R12180 VDPWR.n3108 VDPWR 0.06425
R12181 VDPWR.n3102 VDPWR 0.06425
R12182 VDPWR.n3086 VDPWR 0.06425
R12183 VDPWR.n3070 VDPWR 0.06425
R12184 VDPWR.n753 VDPWR 0.0615066
R12185 VDPWR.n619 VDPWR 0.0603958
R12186 VDPWR VDPWR.n618 0.0603958
R12187 VDPWR.n613 VDPWR 0.0603958
R12188 VDPWR.n608 VDPWR 0.0603958
R12189 VDPWR.n603 VDPWR 0.0603958
R12190 VDPWR.n579 VDPWR 0.0603958
R12191 VDPWR VDPWR.n578 0.0603958
R12192 VDPWR VDPWR.n562 0.0603958
R12193 VDPWR.n638 VDPWR 0.0603958
R12194 VDPWR VDPWR.n637 0.0603958
R12195 VDPWR.n647 VDPWR 0.0603958
R12196 VDPWR.n557 VDPWR 0.0603958
R12197 VDPWR.n339 VDPWR 0.0603958
R12198 VDPWR VDPWR.n338 0.0603958
R12199 VDPWR.n333 VDPWR 0.0603958
R12200 VDPWR.n328 VDPWR 0.0603958
R12201 VDPWR.n323 VDPWR 0.0603958
R12202 VDPWR.n299 VDPWR 0.0603958
R12203 VDPWR VDPWR.n298 0.0603958
R12204 VDPWR VDPWR.n282 0.0603958
R12205 VDPWR.n358 VDPWR 0.0603958
R12206 VDPWR VDPWR.n357 0.0603958
R12207 VDPWR.n367 VDPWR 0.0603958
R12208 VDPWR.n277 VDPWR 0.0603958
R12209 VDPWR.n1527 VDPWR 0.0603958
R12210 VDPWR.n1553 VDPWR 0.0603958
R12211 VDPWR VDPWR.n1481 0.0603958
R12212 VDPWR.n1657 VDPWR 0.0603958
R12213 VDPWR.n1660 VDPWR 0.0603958
R12214 VDPWR.n1661 VDPWR 0.0603958
R12215 VDPWR.n1695 VDPWR 0.0603958
R12216 VDPWR.n1302 VDPWR 0.0603958
R12217 VDPWR.n1870 VDPWR 0.0603958
R12218 VDPWR VDPWR.n1844 0.0603958
R12219 VDPWR.n1833 VDPWR 0.0603958
R12220 VDPWR.n1786 VDPWR 0.0603958
R12221 VDPWR VDPWR.n1784 0.0603958
R12222 VDPWR VDPWR.n1752 0.0603958
R12223 VDPWR VDPWR.n1908 0.0603958
R12224 VDPWR.n1944 VDPWR 0.0603958
R12225 VDPWR.n2155 VDPWR 0.0603958
R12226 VDPWR.n2114 VDPWR 0.0603958
R12227 VDPWR VDPWR.n2107 0.0603958
R12228 VDPWR.n2100 VDPWR 0.0603958
R12229 VDPWR.n2080 VDPWR 0.0603958
R12230 VDPWR VDPWR.n2078 0.0603958
R12231 VDPWR.n2072 VDPWR 0.0603958
R12232 VDPWR.n2220 VDPWR 0.0603958
R12233 VDPWR.n2224 VDPWR 0.0603958
R12234 VDPWR VDPWR.n2196 0.0603958
R12235 VDPWR.n2285 VDPWR 0.0603958
R12236 VDPWR.n2289 VDPWR 0.0603958
R12237 VDPWR.n2298 VDPWR 0.0603958
R12238 VDPWR VDPWR.n2345 0.0603958
R12239 VDPWR.n2346 VDPWR 0.0603958
R12240 VDPWR.n2347 VDPWR 0.0603958
R12241 VDPWR.n2366 VDPWR 0.0603958
R12242 VDPWR.n2367 VDPWR 0.0603958
R12243 VDPWR.n2371 VDPWR 0.0603958
R12244 VDPWR VDPWR.n2426 0.0603958
R12245 VDPWR.n2427 VDPWR 0.0603958
R12246 VDPWR.n970 VDPWR 0.0603958
R12247 VDPWR.n978 VDPWR 0.0603958
R12248 VDPWR.n987 VDPWR 0.0603958
R12249 VDPWR VDPWR.n2552 0.0603958
R12250 VDPWR.n1018 VDPWR 0.0603958
R12251 VDPWR.n1049 VDPWR 0.0603958
R12252 VDPWR.n1051 VDPWR 0.0603958
R12253 VDPWR VDPWR.n1057 0.0603958
R12254 VDPWR.n1058 VDPWR 0.0603958
R12255 VDPWR.n1062 VDPWR 0.0603958
R12256 VDPWR VDPWR.n1089 0.0603958
R12257 VDPWR.n1090 VDPWR 0.0603958
R12258 VDPWR VDPWR.n1102 0.0603958
R12259 VDPWR.n1103 VDPWR 0.0603958
R12260 VDPWR.n1103 VDPWR 0.0603958
R12261 VDPWR.n1109 VDPWR 0.0603958
R12262 VDPWR.n1115 VDPWR 0.0603958
R12263 VDPWR.n1132 VDPWR 0.0603958
R12264 VDPWR.n2528 VDPWR 0.0603958
R12265 VDPWR VDPWR.n2527 0.0603958
R12266 VDPWR VDPWR.n2494 0.0603958
R12267 VDPWR.n2489 VDPWR 0.0603958
R12268 VDPWR.n2604 VDPWR 0.0603958
R12269 VDPWR.n2846 VDPWR 0.0603958
R12270 VDPWR VDPWR.n924 0.0603958
R12271 VDPWR.n2889 VDPWR 0.0603958
R12272 VDPWR VDPWR.n2889 0.0603958
R12273 VDPWR.n2890 VDPWR 0.0603958
R12274 VDPWR.n2897 VDPWR 0.0603958
R12275 VDPWR.n2898 VDPWR 0.0603958
R12276 VDPWR.n2919 VDPWR 0.0603958
R12277 VDPWR VDPWR.n881 0.0603958
R12278 VDPWR.n2929 VDPWR 0.0603958
R12279 VDPWR VDPWR.n878 0.0603958
R12280 VDPWR.n2987 VDPWR 0.0603958
R12281 VDPWR.n2981 VDPWR 0.0603958
R12282 VDPWR.n2639 VDPWR 0.0603958
R12283 VDPWR.n2643 VDPWR 0.0603958
R12284 VDPWR.n2644 VDPWR 0.0603958
R12285 VDPWR VDPWR.n2621 0.0603958
R12286 VDPWR.n2793 VDPWR 0.0603958
R12287 VDPWR VDPWR.n2792 0.0603958
R12288 VDPWR VDPWR.n2657 0.0603958
R12289 VDPWR.n2785 VDPWR 0.0603958
R12290 VDPWR VDPWR.n2784 0.0603958
R12291 VDPWR.n2783 VDPWR 0.0603958
R12292 VDPWR.n2780 VDPWR 0.0603958
R12293 VDPWR.n2762 VDPWR 0.0603958
R12294 VDPWR VDPWR.n2761 0.0603958
R12295 VDPWR VDPWR.n2760 0.0603958
R12296 VDPWR.n2756 VDPWR 0.0603958
R12297 VDPWR.n2681 VDPWR 0.0603958
R12298 VDPWR VDPWR.n2682 0.0603958
R12299 VDPWR.n2744 VDPWR 0.0603958
R12300 VDPWR.n2744 VDPWR 0.0603958
R12301 VDPWR.n2724 VDPWR 0.0603958
R12302 VDPWR.n2722 VDPWR 0.0603958
R12303 VDPWR.n2719 VDPWR 0.0603958
R12304 VDPWR.n786 VDPWR 0.0603958
R12305 VDPWR.n3034 VDPWR 0.0603958
R12306 VDPWR VDPWR.n3033 0.0603958
R12307 VDPWR VDPWR.n790 0.0603958
R12308 VDPWR.n3022 VDPWR 0.0603958
R12309 VDPWR.n3018 VDPWR 0.0603958
R12310 VDPWR VDPWR.n858 0.0603958
R12311 VDPWR.n852 VDPWR 0.0603958
R12312 VDPWR VDPWR.n851 0.0603958
R12313 VDPWR VDPWR.n847 0.0603958
R12314 VDPWR.n844 VDPWR 0.0603958
R12315 VDPWR.n82 VDPWR 0.0603958
R12316 VDPWR VDPWR.n81 0.0603958
R12317 VDPWR.n76 VDPWR 0.0603958
R12318 VDPWR.n71 VDPWR 0.0603958
R12319 VDPWR.n66 VDPWR 0.0603958
R12320 VDPWR.n42 VDPWR 0.0603958
R12321 VDPWR VDPWR.n41 0.0603958
R12322 VDPWR VDPWR.n25 0.0603958
R12323 VDPWR.n101 VDPWR 0.0603958
R12324 VDPWR VDPWR.n100 0.0603958
R12325 VDPWR.n110 VDPWR 0.0603958
R12326 VDPWR.n20 VDPWR 0.0603958
R12327 VDPWR.n3052 VDPWR.n3051 0.0600933
R12328 VDPWR.n560 VDPWR 0.0590938
R12329 VDPWR.n280 VDPWR 0.0590938
R12330 VDPWR.n23 VDPWR 0.0590938
R12331 VDPWR.n3104 VDPWR.n758 0.0589638
R12332 VDPWR.n2026 VDPWR 0.0577917
R12333 VDPWR.n2571 VDPWR 0.0577917
R12334 VDPWR.n806 VDPWR 0.0577917
R12335 VDPWR.n935 VDPWR.n932 0.0574697
R12336 VDPWR.n915 VDPWR.n912 0.0574697
R12337 VDPWR.n1652 VDPWR.n1462 0.0574697
R12338 VDPWR.n1614 VDPWR.n1476 0.0574697
R12339 VDPWR.n1490 VDPWR.n1489 0.0574697
R12340 VDPWR.n1542 VDPWR.n1504 0.0574697
R12341 VDPWR.n1730 VDPWR.n1434 0.0574697
R12342 VDPWR.n1688 VDPWR.n1450 0.0574697
R12343 VDPWR.n1364 VDPWR.n1362 0.0574697
R12344 VDPWR.n1340 VDPWR.n1338 0.0574697
R12345 VDPWR.n1853 VDPWR.n1852 0.0574697
R12346 VDPWR.n1881 VDPWR.n1278 0.0574697
R12347 VDPWR.n1744 VDPWR.n1734 0.0574697
R12348 VDPWR.n1393 VDPWR.n1391 0.0574697
R12349 VDPWR.n2122 VDPWR.n2121 0.0574697
R12350 VDPWR.n2151 VDPWR.n2150 0.0574697
R12351 VDPWR.n2180 VDPWR.n1259 0.0574697
R12352 VDPWR.n1895 VDPWR.n1275 0.0574697
R12353 VDPWR.n2068 VDPWR.n2046 0.0574697
R12354 VDPWR.n2091 VDPWR.n2089 0.0574697
R12355 VDPWR.n2507 VDPWR.n2505 0.0574697
R12356 VDPWR.n3003 VDPWR.n869 0.0574697
R12357 VDPWR.n2400 VDPWR.n1193 0.0574697
R12358 VDPWR.n2402 VDPWR.n1190 0.0574697
R12359 VDPWR.n1231 VDPWR.n1229 0.0574697
R12360 VDPWR.n2189 VDPWR.n1256 0.0574697
R12361 VDPWR.n2239 VDPWR.n2202 0.0574697
R12362 VDPWR.n2452 VDPWR.n1170 0.0574697
R12363 VDPWR.n1211 VDPWR.n1209 0.0574697
R12364 VDPWR.n1128 VDPWR.n1024 0.0574697
R12365 VDPWR.n888 VDPWR.n886 0.0574697
R12366 VDPWR.n1075 VDPWR.n1039 0.0574697
R12367 VDPWR.n1078 VDPWR.n1077 0.0574697
R12368 VDPWR.n2541 VDPWR.n2539 0.0574697
R12369 VDPWR.n2479 VDPWR.n2456 0.0574697
R12370 VDPWR.n981 VDPWR.n956 0.0574697
R12371 VDPWR.n2611 VDPWR.n2584 0.0574697
R12372 VDPWR.n2804 VDPWR.n953 0.0574697
R12373 VDPWR.n2976 VDPWR.n2975 0.0574697
R12374 VDPWR.n1493 VDPWR.n1491 0.0551875
R12375 VDPWR.n1856 VDPWR.n1314 0.0551875
R12376 VDPWR.n1262 VDPWR.n1260 0.0551875
R12377 VDPWR.n2267 VDPWR.n2190 0.0551875
R12378 VDPWR.n2545 VDPWR.n1002 0.0551875
R12379 VDPWR.n2831 VDPWR.n936 0.0551875
R12380 VDPWR.n2773 VDPWR.n2664 0.0551875
R12381 VDPWR.n751 VDPWR.n750 0.0540714
R12382 VDPWR.n465 VDPWR.n402 0.054
R12383 VDPWR.n1718 VDPWR 0.0538854
R12384 VDPWR.n2766 VDPWR 0.0538854
R12385 VDPWR VDPWR.n2709 0.0538854
R12386 VDPWR.n3114 VDPWR 0.0535303
R12387 VDPWR.n3053 VDPWR.n3052 0.0529556
R12388 VDPWR.n652 VDPWR 0.0525833
R12389 VDPWR.n372 VDPWR 0.0525833
R12390 VDPWR VDPWR.n2071 0.0525833
R12391 VDPWR VDPWR.n2836 0.0525833
R12392 VDPWR.n2668 VDPWR 0.0525833
R12393 VDPWR.n2708 VDPWR 0.0525833
R12394 VDPWR.n115 VDPWR 0.0525833
R12395 VDPWR VDPWR.n753 0.0500269
R12396 VDPWR.n1539 VDPWR.n1538 0.0499792
R12397 VDPWR.n1610 VDPWR.n1609 0.0499792
R12398 VDPWR.n1681 VDPWR.n1680 0.0499792
R12399 VDPWR.n1886 VDPWR.n1281 0.0499792
R12400 VDPWR.n1351 VDPWR.n1345 0.0499792
R12401 VDPWR.n1772 VDPWR.n1389 0.0499792
R12402 VDPWR.n1925 VDPWR.n1900 0.0499792
R12403 VDPWR.n1984 VDPWR.n1980 0.0499792
R12404 VDPWR VDPWR.n2021 0.0499792
R12405 VDPWR.n2236 VDPWR.n2235 0.0499792
R12406 VDPWR.n2315 VDPWR.n2314 0.0499792
R12407 VDPWR.n2394 VDPWR.n1194 0.0499792
R12408 VDPWR.n2575 VDPWR.n959 0.0499792
R12409 VDPWR.n1071 VDPWR.n1070 0.0499792
R12410 VDPWR.n2511 VDPWR.n1144 0.0499792
R12411 VDPWR.n2808 VDPWR.n950 0.0499792
R12412 VDPWR.n2875 VDPWR.n2874 0.0499792
R12413 VDPWR.n872 VDPWR.n870 0.0499792
R12414 VDPWR.n2651 VDPWR.n2650 0.0499792
R12415 VDPWR.n2690 VDPWR.n2689 0.0499792
R12416 VDPWR.n3016 VDPWR.n797 0.0499792
R12417 VDPWR VDPWR.n2743 0.047375
R12418 VDPWR.n652 VDPWR.n651 0.0460729
R12419 VDPWR.n372 VDPWR.n371 0.0460729
R12420 VDPWR.n115 VDPWR.n114 0.0460729
R12421 VDPWR.n1494 VDPWR.n1487 0.0447708
R12422 VDPWR.n1649 VDPWR.n1648 0.0447708
R12423 VDPWR.n1720 VDPWR.n1718 0.0447708
R12424 VDPWR.n1325 VDPWR.n1319 0.0447708
R12425 VDPWR.n1374 VDPWR.n1372 0.0447708
R12426 VDPWR.n1738 VDPWR.n1425 0.0447708
R12427 VDPWR.n2178 VDPWR.n2177 0.0447708
R12428 VDPWR.n2009 VDPWR.n2007 0.0447708
R12429 VDPWR.n2086 VDPWR.n2029 0.0447708
R12430 VDPWR.n2049 VDPWR.n2048 0.0447708
R12431 VDPWR.n2279 VDPWR.n2278 0.0447708
R12432 VDPWR.n2351 VDPWR.n1216 0.0447708
R12433 VDPWR.n2442 VDPWR.n2440 0.0447708
R12434 VDPWR.n1012 VDPWR.n1008 0.0447708
R12435 VDPWR.n1125 VDPWR.n1124 0.0447708
R12436 VDPWR.n2459 VDPWR.n2458 0.0447708
R12437 VDPWR.n2832 VDPWR.n930 0.0447708
R12438 VDPWR.n2907 VDPWR.n893 0.0447708
R12439 VDPWR.n3000 VDPWR.n875 0.0447708
R12440 VDPWR.n2963 VDPWR.n2962 0.0447708
R12441 VDPWR.n2766 VDPWR.n2765 0.0447708
R12442 VDPWR.n2709 VDPWR.n783 0.0447708
R12443 VDPWR.n863 VDPWR.n802 0.0447708
R12444 VDPWR.n839 VDPWR.n838 0.0447708
R12445 VDPWR.n2838 VDPWR.n937 0.0410405
R12446 VDPWR.n2834 VDPWR.n931 0.0410405
R12447 VDPWR.n2876 VDPWR.n917 0.0410405
R12448 VDPWR.n2871 VDPWR.n911 0.0410405
R12449 VDPWR.n2740 VDPWR.n2686 0.0410405
R12450 VDPWR.n2736 VDPWR.n2687 0.0410405
R12451 VDPWR.n1638 VDPWR.n1463 0.0410405
R12452 VDPWR.n1651 VDPWR.n1461 0.0410405
R12453 VDPWR.n1608 VDPWR.n1477 0.0410405
R12454 VDPWR.n1613 VDPWR.n1475 0.0410405
R12455 VDPWR.n1578 VDPWR.n1492 0.0410405
R12456 VDPWR.n1574 VDPWR.n1488 0.0410405
R12457 VDPWR.n1529 VDPWR.n1505 0.0410405
R12458 VDPWR.n1541 VDPWR.n1503 0.0410405
R12459 VDPWR.n1717 VDPWR.n1716 0.0410405
R12460 VDPWR.n1729 VDPWR.n1728 0.0410405
R12461 VDPWR.n1677 VDPWR.n1451 0.0410405
R12462 VDPWR.n1687 VDPWR.n1449 0.0410405
R12463 VDPWR.n1369 VDPWR.n1361 0.0410405
R12464 VDPWR.n1370 VDPWR.n1365 0.0410405
R12465 VDPWR.n1347 VDPWR.n1337 0.0410405
R12466 VDPWR.n1348 VDPWR.n1341 0.0410405
R12467 VDPWR.n1316 VDPWR.n1315 0.0410405
R12468 VDPWR.n1318 VDPWR.n1317 0.0410405
R12469 VDPWR.n1891 VDPWR.n1280 0.0410405
R12470 VDPWR.n1884 VDPWR.n1882 0.0410405
R12471 VDPWR.n1740 VDPWR.n1739 0.0410405
R12472 VDPWR.n1743 VDPWR.n1431 0.0410405
R12473 VDPWR.n1398 VDPWR.n1390 0.0410405
R12474 VDPWR.n1399 VDPWR.n1394 0.0410405
R12475 VDPWR.n1998 VDPWR.n1997 0.0410405
R12476 VDPWR.n2000 VDPWR.n1999 0.0410405
R12477 VDPWR.n1974 VDPWR.n1973 0.0410405
R12478 VDPWR.n1976 VDPWR.n1975 0.0410405
R12479 VDPWR.n2185 VDPWR.n1261 0.0410405
R12480 VDPWR.n2181 VDPWR.n2179 0.0410405
R12481 VDPWR.n1930 VDPWR.n1897 0.0410405
R12482 VDPWR.n1898 VDPWR.n1274 0.0410405
R12483 VDPWR.n2067 VDPWR.n2045 0.0410405
R12484 VDPWR.n2058 VDPWR.n2047 0.0410405
R12485 VDPWR.n2093 VDPWR.n2092 0.0410405
R12486 VDPWR.n2025 VDPWR.n2024 0.0410405
R12487 VDPWR.n2509 VDPWR.n2508 0.0410405
R12488 VDPWR.n1149 VDPWR.n1148 0.0410405
R12489 VDPWR.n3008 VDPWR.n871 0.0410405
R12490 VDPWR.n3004 VDPWR.n3002 0.0410405
R12491 VDPWR.n2398 VDPWR.n1195 0.0410405
R12492 VDPWR.n2404 VDPWR.n1189 0.0410405
R12493 VDPWR.n2316 VDPWR.n1233 0.0410405
R12494 VDPWR.n1236 VDPWR.n1228 0.0410405
R12495 VDPWR.n2271 VDPWR.n2191 0.0410405
R12496 VDPWR.n2277 VDPWR.n1255 0.0410405
R12497 VDPWR.n2225 VDPWR.n2203 0.0410405
R12498 VDPWR.n2238 VDPWR.n2201 0.0410405
R12499 VDPWR.n2439 VDPWR.n2438 0.0410405
R12500 VDPWR.n2451 VDPWR.n2450 0.0410405
R12501 VDPWR.n2356 VDPWR.n1213 0.0410405
R12502 VDPWR.n1214 VDPWR.n1208 0.0410405
R12503 VDPWR.n1111 VDPWR.n1025 0.0410405
R12504 VDPWR.n1127 VDPWR.n1023 0.0410405
R12505 VDPWR.n2912 VDPWR.n890 0.0410405
R12506 VDPWR.n891 VDPWR.n885 0.0410405
R12507 VDPWR.n2707 VDPWR.n779 0.0410405
R12508 VDPWR.n3041 VDPWR.n3040 0.0410405
R12509 VDPWR.n1074 VDPWR.n1072 0.0410405
R12510 VDPWR.n1080 VDPWR.n1038 0.0410405
R12511 VDPWR.n2543 VDPWR.n2542 0.0410405
R12512 VDPWR.n1007 VDPWR.n1006 0.0410405
R12513 VDPWR.n2478 VDPWR.n1166 0.0410405
R12514 VDPWR.n2469 VDPWR.n2457 0.0410405
R12515 VDPWR.n2579 VDPWR.n958 0.0410405
R12516 VDPWR.n2573 VDPWR.n982 0.0410405
R12517 VDPWR.n2609 VDPWR.n2587 0.0410405
R12518 VDPWR.n2806 VDPWR.n952 0.0410405
R12519 VDPWR.n2953 VDPWR.n2952 0.0410405
R12520 VDPWR.n2955 VDPWR.n2954 0.0410405
R12521 VDPWR.n2771 VDPWR.n2770 0.0410405
R12522 VDPWR.n2768 VDPWR.n2767 0.0410405
R12523 VDPWR.n2623 VDPWR.n2616 0.0410405
R12524 VDPWR.n2619 VDPWR.n2615 0.0410405
R12525 VDPWR.n840 VDPWR.n772 0.0410405
R12526 VDPWR.n833 VDPWR.n773 0.0410405
R12527 VDPWR.n799 VDPWR.n798 0.0410405
R12528 VDPWR.n866 VDPWR.n865 0.0410405
R12529 VDPWR.n255 VDPWR.n254 0.0403788
R12530 VDPWR VDPWR.n375 0.0403708
R12531 VDPWR.n1584 VDPWR.n1487 0.0395625
R12532 VDPWR.n1617 VDPWR.n1472 0.0395625
R12533 VDPWR.n1648 VDPWR.n1465 0.0395625
R12534 VDPWR.n1692 VDPWR.n1448 0.0395625
R12535 VDPWR.n1720 VDPWR.n1719 0.0395625
R12536 VDPWR.n1849 VDPWR.n1319 0.0395625
R12537 VDPWR.n1820 VDPWR.n1819 0.0395625
R12538 VDPWR.n1374 VDPWR.n1373 0.0395625
R12539 VDPWR.n1407 VDPWR.n1406 0.0395625
R12540 VDPWR.n1741 VDPWR.n1425 0.0395625
R12541 VDPWR.n2177 VDPWR.n1265 0.0395625
R12542 VDPWR.n2147 VDPWR.n2146 0.0395625
R12543 VDPWR.n2009 VDPWR.n2008 0.0395625
R12544 VDPWR.n2029 VDPWR.n2028 0.0395625
R12545 VDPWR.n2065 VDPWR.n2049 0.0395625
R12546 VDPWR.n2279 VDPWR.n1252 0.0395625
R12547 VDPWR.n2323 VDPWR.n2322 0.0395625
R12548 VDPWR.n2351 VDPWR.n1207 0.0395625
R12549 VDPWR.n2406 VDPWR.n2405 0.0395625
R12550 VDPWR.n2442 VDPWR.n2441 0.0395625
R12551 VDPWR.n2536 VDPWR.n1008 0.0395625
R12552 VDPWR.n1088 VDPWR.n1035 0.0395625
R12553 VDPWR.n1124 VDPWR.n1027 0.0395625
R12554 VDPWR.n1154 VDPWR.n1153 0.0395625
R12555 VDPWR.n2476 VDPWR.n2459 0.0395625
R12556 VDPWR.n2844 VDPWR.n930 0.0395625
R12557 VDPWR.n2882 VDPWR.n906 0.0395625
R12558 VDPWR.n2907 VDPWR.n2906 0.0395625
R12559 VDPWR.n3001 VDPWR.n3000 0.0395625
R12560 VDPWR.n2965 VDPWR.n2963 0.0395625
R12561 VDPWR.n2765 VDPWR.n2670 0.0395625
R12562 VDPWR.n2731 VDPWR.n2691 0.0395625
R12563 VDPWR.n3039 VDPWR.n783 0.0395625
R12564 VDPWR.n864 VDPWR.n863 0.0395625
R12565 VDPWR.n838 VDPWR.n823 0.0395625
R12566 VDPWR.n579 VDPWR 0.0382604
R12567 VDPWR.n299 VDPWR 0.0382604
R12568 VDPWR.n42 VDPWR 0.0382604
R12569 VDPWR.n2734 VDPWR.n2733 0.0382581
R12570 VDPWR.n754 VDPWR 0.0376452
R12571 VDPWR VDPWR.n594 0.0369583
R12572 VDPWR VDPWR.n314 0.0369583
R12573 VDPWR VDPWR.n57 0.0369583
R12574 VDPWR.n1538 VDPWR.n1502 0.0343542
R12575 VDPWR.n1611 VDPWR.n1610 0.0343542
R12576 VDPWR.n1726 VDPWR.n1725 0.0343542
R12577 VDPWR.n1886 VDPWR.n1885 0.0343542
R12578 VDPWR.n1351 VDPWR.n1350 0.0343542
R12579 VDPWR.n1397 VDPWR.n1389 0.0343542
R12580 VDPWR.n1748 VDPWR.n1747 0.0343542
R12581 VDPWR.n1925 VDPWR.n1273 0.0343542
R12582 VDPWR.n1984 VDPWR.n1983 0.0343542
R12583 VDPWR.n2062 VDPWR.n2061 0.0343542
R12584 VDPWR.n2235 VDPWR.n2200 0.0343542
R12585 VDPWR.n2314 VDPWR.n1238 0.0343542
R12586 VDPWR.n2397 VDPWR.n2394 0.0343542
R12587 VDPWR.n2448 VDPWR.n2447 0.0343542
R12588 VDPWR.n1070 VDPWR.n1037 0.0343542
R12589 VDPWR.n2511 VDPWR.n2510 0.0343542
R12590 VDPWR.n2473 VDPWR.n2472 0.0343542
R12591 VDPWR.n2808 VDPWR.n2807 0.0343542
R12592 VDPWR.n2874 VDPWR.n2873 0.0343542
R12593 VDPWR.n3007 VDPWR.n872 0.0343542
R12594 VDPWR.n2972 VDPWR.n2971 0.0343542
R12595 VDPWR.n2651 VDPWR.n2620 0.0343542
R12596 VDPWR.n2738 VDPWR.n2690 0.0343542
R12597 VDPWR.n805 VDPWR.n797 0.0343542
R12598 VDPWR.n836 VDPWR.n835 0.0343542
R12599 VDPWR VDPWR.n1660 0.0330521
R12600 VDPWR VDPWR.n978 0.0330521
R12601 VDPWR VDPWR.n1050 0.0330521
R12602 VDPWR.n2528 VDPWR 0.0330521
R12603 VDPWR VDPWR.n2642 0.0330521
R12604 VDPWR.n3034 VDPWR 0.0330521
R12605 VDPWR.n619 VDPWR 0.03175
R12606 VDPWR.n638 VDPWR 0.03175
R12607 VDPWR.n339 VDPWR 0.03175
R12608 VDPWR.n358 VDPWR 0.03175
R12609 VDPWR.n142 VDPWR.n138 0.03175
R12610 VDPWR.n173 VDPWR.n172 0.03175
R12611 VDPWR.n172 VDPWR.n151 0.03175
R12612 VDPWR.n168 VDPWR.n167 0.03175
R12613 VDPWR.n167 VDPWR.n166 0.03175
R12614 VDPWR.n163 VDPWR.n162 0.03175
R12615 VDPWR.n162 VDPWR.n161 0.03175
R12616 VDPWR.n158 VDPWR.n157 0.03175
R12617 VDPWR.n157 VDPWR.n156 0.03175
R12618 VDPWR.n201 VDPWR.n128 0.03175
R12619 VDPWR.n197 VDPWR.n196 0.03175
R12620 VDPWR.n196 VDPWR.n195 0.03175
R12621 VDPWR.n192 VDPWR.n191 0.03175
R12622 VDPWR.n191 VDPWR.n190 0.03175
R12623 VDPWR.n187 VDPWR.n186 0.03175
R12624 VDPWR.n186 VDPWR.n185 0.03175
R12625 VDPWR.n182 VDPWR.n181 0.03175
R12626 VDPWR.n181 VDPWR.n180 0.03175
R12627 VDPWR VDPWR.n1590 0.03175
R12628 VDPWR VDPWR.n1656 0.03175
R12629 VDPWR.n1657 VDPWR 0.03175
R12630 VDPWR.n1845 VDPWR 0.03175
R12631 VDPWR.n1844 VDPWR 0.03175
R12632 VDPWR.n1790 VDPWR 0.03175
R12633 VDPWR.n1752 VDPWR 0.03175
R12634 VDPWR.n2172 VDPWR 0.03175
R12635 VDPWR.n2117 VDPWR 0.03175
R12636 VDPWR.n2080 VDPWR 0.03175
R12637 VDPWR VDPWR.n2284 0.03175
R12638 VDPWR.n2285 VDPWR 0.03175
R12639 VDPWR VDPWR.n2346 0.03175
R12640 VDPWR VDPWR.n2366 0.03175
R12641 VDPWR.n970 VDPWR 0.03175
R12642 VDPWR VDPWR.n1018 0.03175
R12643 VDPWR VDPWR.n1109 0.03175
R12644 VDPWR VDPWR.n1132 0.03175
R12645 VDPWR.n2837 VDPWR 0.03175
R12646 VDPWR.n2846 VDPWR 0.03175
R12647 VDPWR.n2785 VDPWR 0.03175
R12648 VDPWR.n2772 VDPWR 0.03175
R12649 VDPWR.n2761 VDPWR 0.03175
R12650 VDPWR.n2760 VDPWR 0.03175
R12651 VDPWR VDPWR.n2685 0.03175
R12652 VDPWR.n2719 VDPWR 0.03175
R12653 VDPWR VDPWR.n2706 0.03175
R12654 VDPWR VDPWR.n786 0.03175
R12655 VDPWR.n807 VDPWR 0.03175
R12656 VDPWR.n847 VDPWR 0.03175
R12657 VDPWR.n82 VDPWR 0.03175
R12658 VDPWR.n101 VDPWR 0.03175
R12659 VDPWR.n1434 VDPWR.n1432 0.0292489
R12660 VDPWR.n1731 VDPWR.n1730 0.0292489
R12661 VDPWR.n1736 VDPWR.n1734 0.0292489
R12662 VDPWR.n1745 VDPWR.n1744 0.0292489
R12663 VDPWR.n2069 VDPWR.n2068 0.0292489
R12664 VDPWR.n2059 VDPWR.n2046 0.0292489
R12665 VDPWR.n3010 VDPWR.n869 0.0292489
R12666 VDPWR.n3003 VDPWR.n868 0.0292489
R12667 VDPWR.n2507 VDPWR.n2506 0.0292489
R12668 VDPWR.n2505 VDPWR.n2504 0.0292489
R12669 VDPWR.n2091 VDPWR.n2090 0.0292489
R12670 VDPWR.n2089 VDPWR.n2088 0.0292489
R12671 VDPWR.n1770 VDPWR.n1391 0.0292489
R12672 VDPWR.n1768 VDPWR.n1393 0.0292489
R12673 VDPWR.n1678 VDPWR.n1450 0.0292489
R12674 VDPWR.n1689 VDPWR.n1688 0.0292489
R12675 VDPWR.n1192 VDPWR.n1190 0.0292489
R12676 VDPWR.n1193 VDPWR.n1192 0.0292489
R12677 VDPWR.n1170 VDPWR.n1168 0.0292489
R12678 VDPWR.n2453 VDPWR.n2452 0.0292489
R12679 VDPWR.n2914 VDPWR.n888 0.0292489
R12680 VDPWR.n2916 VDPWR.n886 0.0292489
R12681 VDPWR.n1112 VDPWR.n1024 0.0292489
R12682 VDPWR.n1129 VDPWR.n1128 0.0292489
R12683 VDPWR.n2358 VDPWR.n1211 0.0292489
R12684 VDPWR.n2360 VDPWR.n1209 0.0292489
R12685 VDPWR.n2123 VDPWR.n2122 0.0292489
R12686 VDPWR.n2121 VDPWR.n2120 0.0292489
R12687 VDPWR.n1795 VDPWR.n1362 0.0292489
R12688 VDPWR.n1793 VDPWR.n1364 0.0292489
R12689 VDPWR.n1639 VDPWR.n1462 0.0292489
R12690 VDPWR.n1653 VDPWR.n1652 0.0292489
R12691 VDPWR.n2878 VDPWR.n915 0.0292489
R12692 VDPWR.n2880 VDPWR.n912 0.0292489
R12693 VDPWR.n2318 VDPWR.n1231 0.0292489
R12694 VDPWR.n2320 VDPWR.n1229 0.0292489
R12695 VDPWR.n2152 VDPWR.n2151 0.0292489
R12696 VDPWR.n2150 VDPWR.n2149 0.0292489
R12697 VDPWR.n1824 VDPWR.n1338 0.0292489
R12698 VDPWR.n1822 VDPWR.n1340 0.0292489
R12699 VDPWR.n1606 VDPWR.n1476 0.0292489
R12700 VDPWR.n1615 VDPWR.n1614 0.0292489
R12701 VDPWR.n1077 VDPWR.n1076 0.0292489
R12702 VDPWR.n1076 VDPWR.n1075 0.0292489
R12703 VDPWR.n2480 VDPWR.n2479 0.0292489
R12704 VDPWR.n2470 VDPWR.n2456 0.0292489
R12705 VDPWR.n2581 VDPWR.n956 0.0292489
R12706 VDPWR.n981 VDPWR.n955 0.0292489
R12707 VDPWR.n2226 VDPWR.n2202 0.0292489
R12708 VDPWR.n2240 VDPWR.n2239 0.0292489
R12709 VDPWR.n1932 VDPWR.n1895 0.0292489
R12710 VDPWR.n1934 VDPWR.n1275 0.0292489
R12711 VDPWR.n1893 VDPWR.n1278 0.0292489
R12712 VDPWR.n1881 VDPWR.n1277 0.0292489
R12713 VDPWR.n1530 VDPWR.n1504 0.0292489
R12714 VDPWR.n1543 VDPWR.n1542 0.0292489
R12715 VDPWR.n2583 VDPWR.n953 0.0292489
R12716 VDPWR.n2584 VDPWR.n2583 0.0292489
R12717 VDPWR.n2977 VDPWR.n2976 0.0292489
R12718 VDPWR.n2975 VDPWR.n2974 0.0292489
R12719 VDPWR.n2840 VDPWR.n935 0.0292489
R12720 VDPWR.n2842 VDPWR.n932 0.0292489
R12721 VDPWR.n2541 VDPWR.n2540 0.0292489
R12722 VDPWR.n2539 VDPWR.n2538 0.0292489
R12723 VDPWR.n2273 VDPWR.n2189 0.0292489
R12724 VDPWR.n2275 VDPWR.n1256 0.0292489
R12725 VDPWR.n2187 VDPWR.n1259 0.0292489
R12726 VDPWR.n2180 VDPWR.n1258 0.0292489
R12727 VDPWR.n1854 VDPWR.n1853 0.0292489
R12728 VDPWR.n1852 VDPWR.n1851 0.0292489
R12729 VDPWR.n1580 VDPWR.n1490 0.0292489
R12730 VDPWR.n1582 VDPWR.n1489 0.0292489
R12731 VDPWR.n585 VDPWR.n584 0.0291458
R12732 VDPWR.n305 VDPWR.n304 0.0291458
R12733 VDPWR.n1577 VDPWR.n1493 0.0291458
R12734 VDPWR.n1642 VDPWR.n1641 0.0291458
R12735 VDPWR.n1322 VDPWR.n1314 0.0291458
R12736 VDPWR.n1798 VDPWR.n1797 0.0291458
R12737 VDPWR.n2184 VDPWR.n1262 0.0291458
R12738 VDPWR.n2126 VDPWR.n2125 0.0291458
R12739 VDPWR.n2270 VDPWR.n2267 0.0291458
R12740 VDPWR.n2347 VDPWR.n1212 0.0291458
R12741 VDPWR.n2545 VDPWR.n2544 0.0291458
R12742 VDPWR.n1115 VDPWR.n1114 0.0291458
R12743 VDPWR.n2898 VDPWR.n889 0.0291458
R12744 VDPWR.n48 VDPWR.n47 0.0291458
R12745 VDPWR.n752 VDPWR.n751 0.0281786
R12746 VDPWR.n2094 VDPWR 0.0265417
R12747 VDPWR.n2574 VDPWR 0.0265417
R12748 VDPWR VDPWR.n805 0.0265417
R12749 VDPWR.n202 VDPWR.n127 0.0249565
R12750 VDPWR.n726 VDPWR.n724 0.0247347
R12751 VDPWR.n1533 VDPWR.n1532 0.0239375
R12752 VDPWR.n1303 VDPWR.n1279 0.0239375
R12753 VDPWR.n1907 VDPWR.n1896 0.0239375
R12754 VDPWR.n2229 VDPWR.n2228 0.0239375
R12755 VDPWR VDPWR.n1062 0.0239375
R12756 VDPWR.n2604 VDPWR.n2585 0.0239375
R12757 VDPWR.n2981 VDPWR 0.0239375
R12758 VDPWR.n2627 VDPWR.n2626 0.0239375
R12759 VDPWR.n654 VDPWR 0.0236148
R12760 VDPWR VDPWR.n3116 0.0236148
R12761 VDPWR.n727 VDPWR.n722 0.0234592
R12762 VDPWR VDPWR.n566 0.0226354
R12763 VDPWR VDPWR.n591 0.0226354
R12764 VDPWR.n611 VDPWR 0.0226354
R12765 VDPWR.n606 VDPWR 0.0226354
R12766 VDPWR.n598 VDPWR 0.0226354
R12767 VDPWR VDPWR.n568 0.0226354
R12768 VDPWR.n578 VDPWR 0.0226354
R12769 VDPWR.n628 VDPWR 0.0226354
R12770 VDPWR VDPWR.n636 0.0226354
R12771 VDPWR.n637 VDPWR 0.0226354
R12772 VDPWR VDPWR.n537 0.0226354
R12773 VDPWR VDPWR.n541 0.0226354
R12774 VDPWR VDPWR.n546 0.0226354
R12775 VDPWR.n551 VDPWR 0.0226354
R12776 VDPWR VDPWR.n286 0.0226354
R12777 VDPWR VDPWR.n311 0.0226354
R12778 VDPWR.n331 VDPWR 0.0226354
R12779 VDPWR.n326 VDPWR 0.0226354
R12780 VDPWR.n318 VDPWR 0.0226354
R12781 VDPWR VDPWR.n288 0.0226354
R12782 VDPWR.n298 VDPWR 0.0226354
R12783 VDPWR.n348 VDPWR 0.0226354
R12784 VDPWR VDPWR.n356 0.0226354
R12785 VDPWR.n357 VDPWR 0.0226354
R12786 VDPWR VDPWR.n257 0.0226354
R12787 VDPWR VDPWR.n261 0.0226354
R12788 VDPWR VDPWR.n266 0.0226354
R12789 VDPWR.n271 VDPWR 0.0226354
R12790 VDPWR VDPWR.n1552 0.0226354
R12791 VDPWR.n1559 VDPWR 0.0226354
R12792 VDPWR.n1585 VDPWR 0.0226354
R12793 VDPWR VDPWR.n1676 0.0226354
R12794 VDPWR.n1681 VDPWR 0.0226354
R12795 VDPWR.n1692 VDPWR 0.0226354
R12796 VDPWR VDPWR.n1691 0.0226354
R12797 VDPWR.n1713 VDPWR 0.0226354
R12798 VDPWR.n1725 VDPWR 0.0226354
R12799 VDPWR.n1873 VDPWR 0.0226354
R12800 VDPWR.n1864 VDPWR 0.0226354
R12801 VDPWR.n1848 VDPWR 0.0226354
R12802 VDPWR.n1814 VDPWR 0.0226354
R12803 VDPWR.n1786 VDPWR 0.0226354
R12804 VDPWR.n1784 VDPWR 0.0226354
R12805 VDPWR.n1407 VDPWR 0.0226354
R12806 VDPWR.n1766 VDPWR 0.0226354
R12807 VDPWR.n1753 VDPWR 0.0226354
R12808 VDPWR VDPWR.n1417 0.0226354
R12809 VDPWR.n1748 VDPWR 0.0226354
R12810 VDPWR VDPWR.n1943 0.0226354
R12811 VDPWR.n1950 VDPWR 0.0226354
R12812 VDPWR.n2173 VDPWR 0.0226354
R12813 VDPWR.n2158 VDPWR 0.0226354
R12814 VDPWR.n2141 VDPWR 0.0226354
R12815 VDPWR.n2134 VDPWR 0.0226354
R12816 VDPWR.n2108 VDPWR 0.0226354
R12817 VDPWR.n2107 VDPWR 0.0226354
R12818 VDPWR.n2078 VDPWR 0.0226354
R12819 VDPWR VDPWR.n2044 0.0226354
R12820 VDPWR.n2062 VDPWR 0.0226354
R12821 VDPWR.n2220 VDPWR 0.0226354
R12822 VDPWR.n2248 VDPWR 0.0226354
R12823 VDPWR.n2254 VDPWR 0.0226354
R12824 VDPWR VDPWR.n2283 0.0226354
R12825 VDPWR VDPWR.n2289 0.0226354
R12826 VDPWR.n2290 VDPWR 0.0226354
R12827 VDPWR VDPWR.n2297 0.0226354
R12828 VDPWR.n2332 VDPWR 0.0226354
R12829 VDPWR.n2367 VDPWR 0.0226354
R12830 VDPWR VDPWR.n2371 0.0226354
R12831 VDPWR.n2406 VDPWR 0.0226354
R12832 VDPWR VDPWR.n1185 0.0226354
R12833 VDPWR.n2435 VDPWR 0.0226354
R12834 VDPWR.n2447 VDPWR 0.0226354
R12835 VDPWR.n2575 VDPWR 0.0226354
R12836 VDPWR.n2570 VDPWR 0.0226354
R12837 VDPWR.n2566 VDPWR 0.0226354
R12838 VDPWR.n2553 VDPWR 0.0226354
R12839 VDPWR.n2535 VDPWR 0.0226354
R12840 VDPWR.n1051 VDPWR 0.0226354
R12841 VDPWR.n1058 VDPWR 0.0226354
R12842 VDPWR.n1090 VDPWR 0.0226354
R12843 VDPWR.n1154 VDPWR 0.0226354
R12844 VDPWR.n2502 VDPWR 0.0226354
R12845 VDPWR.n2495 VDPWR 0.0226354
R12846 VDPWR VDPWR.n1165 0.0226354
R12847 VDPWR.n2473 VDPWR 0.0226354
R12848 VDPWR VDPWR.n2831 0.0226354
R12849 VDPWR VDPWR.n2845 0.0226354
R12850 VDPWR.n2883 VDPWR 0.0226354
R12851 VDPWR.n906 VDPWR 0.0226354
R12852 VDPWR VDPWR.n2888 0.0226354
R12853 VDPWR VDPWR.n2919 0.0226354
R12854 VDPWR.n2990 VDPWR 0.0226354
R12855 VDPWR VDPWR.n2948 0.0226354
R12856 VDPWR VDPWR.n2951 0.0226354
R12857 VDPWR.n2971 VDPWR 0.0226354
R12858 VDPWR.n2639 VDPWR 0.0226354
R12859 VDPWR VDPWR.n2643 0.0226354
R12860 VDPWR VDPWR.n2648 0.0226354
R12861 VDPWR.n2793 VDPWR 0.0226354
R12862 VDPWR.n2792 VDPWR 0.0226354
R12863 VDPWR.n2780 VDPWR 0.0226354
R12864 VDPWR.n2773 VDPWR 0.0226354
R12865 VDPWR VDPWR.n2669 0.0226354
R12866 VDPWR.n2756 VDPWR 0.0226354
R12867 VDPWR.n2749 VDPWR 0.0226354
R12868 VDPWR VDPWR.n2681 0.0226354
R12869 VDPWR VDPWR.n2697 0.0226354
R12870 VDPWR.n2724 VDPWR 0.0226354
R12871 VDPWR.n2710 VDPWR 0.0226354
R12872 VDPWR.n3033 VDPWR 0.0226354
R12873 VDPWR.n3021 VDPWR 0.0226354
R12874 VDPWR.n3018 VDPWR 0.0226354
R12875 VDPWR.n859 VDPWR 0.0226354
R12876 VDPWR VDPWR.n812 0.0226354
R12877 VDPWR.n852 VDPWR 0.0226354
R12878 VDPWR.n851 VDPWR 0.0226354
R12879 VDPWR.n844 VDPWR 0.0226354
R12880 VDPWR VDPWR.n821 0.0226354
R12881 VDPWR.n836 VDPWR 0.0226354
R12882 VDPWR VDPWR.n29 0.0226354
R12883 VDPWR VDPWR.n54 0.0226354
R12884 VDPWR.n74 VDPWR 0.0226354
R12885 VDPWR.n69 VDPWR 0.0226354
R12886 VDPWR.n61 VDPWR 0.0226354
R12887 VDPWR VDPWR.n31 0.0226354
R12888 VDPWR.n41 VDPWR 0.0226354
R12889 VDPWR.n91 VDPWR 0.0226354
R12890 VDPWR VDPWR.n99 0.0226354
R12891 VDPWR.n100 VDPWR 0.0226354
R12892 VDPWR VDPWR.n0 0.0226354
R12893 VDPWR VDPWR.n4 0.0226354
R12894 VDPWR VDPWR.n9 0.0226354
R12895 VDPWR.n14 VDPWR 0.0226354
R12896 VDPWR.n248 VDPWR.n121 0.0226154
R12897 VDPWR.n243 VDPWR.n242 0.0226154
R12898 VDPWR.n238 VDPWR.n237 0.0226154
R12899 VDPWR.n233 VDPWR.n232 0.0226154
R12900 VDPWR.n228 VDPWR.n227 0.0226154
R12901 VDPWR.n223 VDPWR.n222 0.0226154
R12902 VDPWR.n218 VDPWR.n217 0.0226154
R12903 VDPWR.n213 VDPWR.n212 0.0226154
R12904 VDPWR.n208 VDPWR.n207 0.0226154
R12905 VDPWR.n3045 VDPWR.n3044 0.0218125
R12906 VDPWR VDPWR.n2017 0.0213333
R12907 VDPWR VDPWR.n1159 0.0213333
R12908 VDPWR VDPWR.n2882 0.0213333
R12909 VDPWR VDPWR.n2897 0.0213333
R12910 VDPWR.n864 VDPWR 0.0213333
R12911 VDPWR VDPWR.n1655 0.0200312
R12912 VDPWR.n1791 VDPWR 0.0200312
R12913 VDPWR.n2118 VDPWR 0.0200312
R12914 VDPWR.n2362 VDPWR 0.0200312
R12915 VDPWR VDPWR.n1131 0.0200312
R12916 VDPWR VDPWR.n2918 0.0200312
R12917 VDPWR VDPWR.n784 0.0200312
R12918 VDPWR VDPWR.n248 0.0185288
R12919 VDPWR.n243 VDPWR 0.0185288
R12920 VDPWR.n238 VDPWR 0.0185288
R12921 VDPWR.n233 VDPWR 0.0185288
R12922 VDPWR.n223 VDPWR 0.0185288
R12923 VDPWR.n218 VDPWR 0.0185288
R12924 VDPWR.n213 VDPWR 0.0185288
R12925 VDPWR.n208 VDPWR 0.0185288
R12926 VDPWR VDPWR.n137 0.016125
R12927 VDPWR.n149 VDPWR 0.016125
R12928 VDPWR.n150 VDPWR 0.016125
R12929 VDPWR.n174 VDPWR 0.016125
R12930 VDPWR VDPWR.n173 0.016125
R12931 VDPWR.n168 VDPWR 0.016125
R12932 VDPWR.n163 VDPWR 0.016125
R12933 VDPWR.n158 VDPWR 0.016125
R12934 VDPWR VDPWR.n127 0.016125
R12935 VDPWR.n197 VDPWR 0.016125
R12936 VDPWR.n192 VDPWR 0.016125
R12937 VDPWR.n187 VDPWR 0.016125
R12938 VDPWR.n182 VDPWR 0.016125
R12939 VDPWR.n177 VDPWR 0.016125
R12940 VDPWR.n1691 VDPWR 0.016125
R12941 VDPWR.n1738 VDPWR 0.016125
R12942 VDPWR.n2048 VDPWR 0.016125
R12943 VDPWR.n2440 VDPWR 0.016125
R12944 VDPWR.n2458 VDPWR 0.016125
R12945 VDPWR.n2962 VDPWR 0.016125
R12946 VDPWR.n839 VDPWR 0.016125
R12947 VDPWR.n203 VDPWR 0.0137212
R12948 VDPWR.n1528 VDPWR.n1506 0.0135208
R12949 VDPWR.n1605 VDPWR.n1478 0.0135208
R12950 VDPWR.n1890 VDPWR.n1889 0.0135208
R12951 VDPWR.n1826 VDPWR.n1336 0.0135208
R12952 VDPWR.n1929 VDPWR.n1928 0.0135208
R12953 VDPWR.n2154 VDPWR.n1972 0.0135208
R12954 VDPWR.n2234 VDPWR.n2204 0.0135208
R12955 VDPWR.n1234 VDPWR.n1232 0.0135208
R12956 VDPWR.n2578 VDPWR.n2577 0.0135208
R12957 VDPWR.n1069 VDPWR.n1041 0.0135208
R12958 VDPWR.n2608 VDPWR.n2607 0.0135208
R12959 VDPWR.n2870 VDPWR.n916 0.0135208
R12960 VDPWR.n2648 VDPWR.n2624 0.0135208
R12961 VDPWR.n2743 VDPWR.n2685 0.0135208
R12962 VDPWR.n3055 VDPWR 0.0122968
R12963 VDPWR VDPWR.n1452 0.0122188
R12964 VDPWR VDPWR.n2094 0.0122188
R12965 VDPWR VDPWR.n2574 0.0122188
R12966 VDPWR VDPWR.n249 0.0115577
R12967 VDPWR VDPWR.n121 0.0115577
R12968 VDPWR.n122 VDPWR 0.0115577
R12969 VDPWR.n242 VDPWR 0.0115577
R12970 VDPWR VDPWR.n241 0.0115577
R12971 VDPWR.n237 VDPWR 0.0115577
R12972 VDPWR VDPWR.n236 0.0115577
R12973 VDPWR.n232 VDPWR 0.0115577
R12974 VDPWR VDPWR.n231 0.0115577
R12975 VDPWR.n227 VDPWR 0.0115577
R12976 VDPWR VDPWR.n226 0.0115577
R12977 VDPWR.n222 VDPWR 0.0115577
R12978 VDPWR VDPWR.n221 0.0115577
R12979 VDPWR.n217 VDPWR 0.0115577
R12980 VDPWR VDPWR.n216 0.0115577
R12981 VDPWR.n212 VDPWR 0.0115577
R12982 VDPWR VDPWR.n211 0.0115577
R12983 VDPWR.n207 VDPWR 0.0115577
R12984 VDPWR.n252 VDPWR 0.0115577
R12985 VDPWR.n1680 VDPWR 0.0109167
R12986 VDPWR.n2650 VDPWR 0.0109167
R12987 VDPWR.n2689 VDPWR 0.0109167
R12988 VDPWR.n3047 VDPWR 0.00972152
R12989 VDPWR.n3046 VDPWR 0.00972152
R12990 VDPWR VDPWR.n775 0.00972152
R12991 VDPWR.n2613 VDPWR 0.00972152
R12992 VDPWR.n374 VDPWR.n254 0.00887356
R12993 VDPWR.n137 VDPWR 0.00865217
R12994 VDPWR VDPWR.n149 0.00865217
R12995 VDPWR VDPWR.n150 0.00865217
R12996 VDPWR.n174 VDPWR 0.00865217
R12997 VDPWR.n177 VDPWR 0.00865217
R12998 VDPWR.n1576 VDPWR.n1573 0.0083125
R12999 VDPWR.n1637 VDPWR.n1464 0.0083125
R13000 VDPWR.n1714 VDPWR.n1713 0.0083125
R13001 VDPWR.n1326 VDPWR.n1324 0.0083125
R13002 VDPWR.n1368 VDPWR.n1360 0.0083125
R13003 VDPWR.n1735 VDPWR.n1417 0.0083125
R13004 VDPWR.n2183 VDPWR.n1263 0.0083125
R13005 VDPWR.n2005 VDPWR.n1996 0.0083125
R13006 VDPWR.n2071 VDPWR.n2044 0.0083125
R13007 VDPWR.n2269 VDPWR.n1254 0.0083125
R13008 VDPWR.n2355 VDPWR.n2354 0.0083125
R13009 VDPWR.n2436 VDPWR.n2435 0.0083125
R13010 VDPWR.n1013 VDPWR.n1003 0.0083125
R13011 VDPWR.n1110 VDPWR.n1026 0.0083125
R13012 VDPWR.n2482 VDPWR.n1165 0.0083125
R13013 VDPWR.n2836 VDPWR.n2833 0.0083125
R13014 VDPWR.n2911 VDPWR.n2910 0.0083125
R13015 VDPWR.n2979 VDPWR.n2951 0.0083125
R13016 VDPWR.n2669 VDPWR.n2668 0.0083125
R13017 VDPWR.n2710 VDPWR.n2708 0.0083125
R13018 VDPWR.n842 VDPWR.n821 0.0083125
R13019 VDPWR.n202 VDPWR.n201 0.00729348
R13020 VDPWR.n2837 VDPWR 0.00701042
R13021 VDPWR VDPWR.n2772 0.00701042
R13022 VDPWR.n2706 VDPWR 0.00701042
R13023 VDPWR.n3049 VDPWR.n3048 0.006375
R13024 VDPWR VDPWR.n151 0.00627446
R13025 VDPWR.n166 VDPWR 0.00627446
R13026 VDPWR.n161 VDPWR 0.00627446
R13027 VDPWR.n156 VDPWR 0.00627446
R13028 VDPWR VDPWR.n128 0.00627446
R13029 VDPWR.n195 VDPWR 0.00627446
R13030 VDPWR.n190 VDPWR 0.00627446
R13031 VDPWR.n185 VDPWR 0.00627446
R13032 VDPWR.n180 VDPWR 0.00627446
R13033 VDPWR VDPWR.n252 0.00626923
R13034 VDPWR.n138 VDPWR 0.00593478
R13035 VDPWR.n228 VDPWR.n203 0.00530769
R13036 VDPWR.n3013 VDPWR.n3012 0.0052
R13037 VDPWR.n778 VDPWR.n777 0.0052
R13038 VDPWR.n2802 VDPWR.n2614 0.0052
R13039 VDPWR.n2612 VDPWR.n934 0.0052
R13040 VDPWR.n249 VDPWR 0.00458654
R13041 VDPWR VDPWR.n122 0.00458654
R13042 VDPWR.n241 VDPWR 0.00458654
R13043 VDPWR.n236 VDPWR 0.00458654
R13044 VDPWR.n231 VDPWR 0.00458654
R13045 VDPWR.n226 VDPWR 0.00458654
R13046 VDPWR.n221 VDPWR 0.00458654
R13047 VDPWR.n216 VDPWR 0.00458654
R13048 VDPWR.n211 VDPWR 0.00458654
R13049 VDPWR.n3049 VDPWR 0.00398148
R13050 VDPWR.n628 VDPWR.n627 0.00310417
R13051 VDPWR.n348 VDPWR.n347 0.00310417
R13052 VDPWR.n1546 VDPWR.n1545 0.00310417
R13053 VDPWR.n1618 VDPWR.n1474 0.00310417
R13054 VDPWR.n1655 VDPWR.n1460 0.00310417
R13055 VDPWR.n1685 VDPWR.n1684 0.00310417
R13056 VDPWR.n1727 VDPWR.n1436 0.00310417
R13057 VDPWR.n1879 VDPWR.n1878 0.00310417
R13058 VDPWR.n1346 VDPWR.n1342 0.00310417
R13059 VDPWR.n1791 VDPWR.n1366 0.00310417
R13060 VDPWR.n1405 VDPWR.n1401 0.00310417
R13061 VDPWR.n1430 VDPWR.n1426 0.00310417
R13062 VDPWR.n1937 VDPWR.n1936 0.00310417
R13063 VDPWR.n1981 VDPWR.n1977 0.00310417
R13064 VDPWR.n2118 VDPWR.n2001 0.00310417
R13065 VDPWR.n2027 VDPWR.n2026 0.00310417
R13066 VDPWR.n2064 VDPWR.n2050 0.00310417
R13067 VDPWR.n2243 VDPWR.n2242 0.00310417
R13068 VDPWR.n1235 VDPWR.n1227 0.00310417
R13069 VDPWR.n2363 VDPWR.n2362 0.00310417
R13070 VDPWR.n2396 VDPWR.n1188 0.00310417
R13071 VDPWR.n2449 VDPWR.n1172 0.00310417
R13072 VDPWR.n2571 VDPWR.n2570 0.00310417
R13073 VDPWR.n1082 VDPWR.n1081 0.00310417
R13074 VDPWR.n1131 VDPWR.n1022 0.00310417
R13075 VDPWR.n1152 VDPWR.n1145 0.00310417
R13076 VDPWR.n2475 VDPWR.n2460 0.00310417
R13077 VDPWR.n951 VDPWR.n946 0.00310417
R13078 VDPWR.n2883 VDPWR.n910 0.00310417
R13079 VDPWR.n2918 VDPWR.n884 0.00310417
R13080 VDPWR.n3006 VDPWR.n873 0.00310417
R13081 VDPWR.n2966 VDPWR.n2956 0.00310417
R13082 VDPWR.n2799 VDPWR.n2798 0.00310417
R13083 VDPWR.n2737 VDPWR.n2735 0.00310417
R13084 VDPWR.n3038 VDPWR.n784 0.00310417
R13085 VDPWR.n807 VDPWR.n806 0.00310417
R13086 VDPWR.n834 VDPWR.n829 0.00310417
R13087 VDPWR.n91 VDPWR.n90 0.00310417
R13088 VDPWR.n626 VDPWR.n625 0.00180208
R13089 VDPWR.n594 VDPWR 0.00180208
R13090 VDPWR.n560 VDPWR.n546 0.00180208
R13091 VDPWR.n346 VDPWR.n345 0.00180208
R13092 VDPWR.n314 VDPWR 0.00180208
R13093 VDPWR.n280 VDPWR.n266 0.00180208
R13094 VDPWR.n89 VDPWR.n88 0.00180208
R13095 VDPWR.n57 VDPWR 0.00180208
R13096 VDPWR.n23 VDPWR.n9 0.00180208
R13097 VDPWR.n727 VDPWR.n726 0.00177551
R13098 VDPWR.n256 VDPWR.n255 0.00105731
R13099 muxtest_0.x2.x2.GP1.n2 muxtest_0.x2.x2.GP1.t4 450.938
R13100 muxtest_0.x2.x2.GP1.n2 muxtest_0.x2.x2.GP1.t5 445.666
R13101 muxtest_0.x2.x2.GP1.n4 muxtest_0.x2.x2.GP1.n3 195.832
R13102 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n0 96.8352
R13103 muxtest_0.x2.x2.GP1.n3 muxtest_0.x2.x2.GP1.t1 26.5955
R13104 muxtest_0.x2.x2.GP1.n3 muxtest_0.x2.x2.GP1.t0 26.5955
R13105 muxtest_0.x2.x2.GP1.n0 muxtest_0.x2.x2.GP1.t3 24.9236
R13106 muxtest_0.x2.x2.GP1.n0 muxtest_0.x2.x2.GP1.t2 24.9236
R13107 muxtest_0.x2.x2.GP1.n5 muxtest_0.x2.x2.GP1.n4 13.1346
R13108 muxtest_0.x2.x2.GP1.n4 muxtest_0.x2.x2.GP1 12.2007
R13109 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n1 11.2645
R13110 muxtest_0.x2.x2.GP1.n1 muxtest_0.x2.x2.GP1 6.1445
R13111 muxtest_0.x2.x2.GP1.n1 muxtest_0.x2.x2.GP1 4.65505
R13112 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n2 3.07707
R13113 muxtest_0.x2.x2.GP1.n5 muxtest_0.x2.x2.GP1 2.0485
R13114 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP1.n5 1.55202
R13115 ua[3].n10 ua[3].t9 26.3998
R13116 ua[3].n6 ua[3].t0 23.6581
R13117 ua[3].n1 ua[3].t5 23.6581
R13118 ua[3].n10 ua[3].t8 23.5483
R13119 ua[3].n8 ua[3].t10 23.3739
R13120 ua[3].n3 ua[3].t4 23.3739
R13121 ua[3].n11 ua[3].t7 12.9758
R13122 ua[3].n11 ua[3].t6 10.8618
R13123 ua[3].n6 ua[3].t3 10.7528
R13124 ua[3].n1 ua[3].t11 10.7528
R13125 ua[3].n5 ua[3].t2 10.6417
R13126 ua[3].n0 ua[3].t1 10.6417
R13127 ua[3].n15 ua[3] 4.48702
R13128 ua[3].n12 ua[3].n10 3.06895
R13129 ua[3].n12 ua[3].n11 2.14822
R13130 ua[3].n14 ua[3] 1.938
R13131 ua[3].n7 ua[3].n6 1.30064
R13132 ua[3].n2 ua[3].n1 1.30064
R13133 ua[3].n13 ua[3].n12 1.12636
R13134 ua[3] ua[3].n9 0.983856
R13135 ua[3] ua[3].n4 0.966624
R13136 ua[3].n8 ua[3].n7 0.726502
R13137 ua[3].n3 ua[3].n2 0.726502
R13138 ua[3].n17 ua[3].n16 0.683625
R13139 ua[3].n7 ua[3].n5 0.512491
R13140 ua[3].n2 ua[3].n0 0.512491
R13141 ua[3].n15 ua[3] 0.398
R13142 ua[3] ua[3].n15 0.398
R13143 ua[3].n16 ua[3] 0.37425
R13144 ua[3].n9 ua[3].n5 0.359663
R13145 ua[3].n4 ua[3].n0 0.359663
R13146 ua[3].n16 ua[3] 0.2705
R13147 ua[3].n9 ua[3].n8 0.216071
R13148 ua[3].n4 ua[3].n3 0.216071
R13149 ua[3].n14 ua[3].n13 0.148615
R13150 ua[3] ua[3].n14 0.146333
R13151 ua[3].n17 ua[3] 0.124875
R13152 ua[3].n13 ua[3] 0.0655
R13153 ua[3] ua[3].n17 0.063
R13154 ua[2].n6 ua[2].t14 23.6581
R13155 ua[2].n15 ua[2].t5 23.6581
R13156 ua[2].n22 ua[2].t2 23.6581
R13157 ua[2].n1 ua[2].t1 23.6581
R13158 ua[2].n5 ua[2].t15 23.3739
R13159 ua[2].n14 ua[2].t4 23.3739
R13160 ua[2].n21 ua[2].t3 23.3739
R13161 ua[2].n0 ua[2].t0 23.3739
R13162 ua[2].n28 ua[2] 21.5313
R13163 ua[2].n6 ua[2].t13 10.7528
R13164 ua[2].n15 ua[2].t11 10.7528
R13165 ua[2].n22 ua[2].t8 10.7528
R13166 ua[2].n1 ua[2].t6 10.7528
R13167 ua[2].n8 ua[2].t12 10.6417
R13168 ua[2].n17 ua[2].t10 10.6417
R13169 ua[2].n24 ua[2].t9 10.6417
R13170 ua[2].n3 ua[2].t7 10.6417
R13171 ua[2].n7 ua[2].n6 1.30064
R13172 ua[2].n16 ua[2].n15 1.30064
R13173 ua[2].n23 ua[2].n22 1.30064
R13174 ua[2].n2 ua[2].n1 1.30064
R13175 ua[2] ua[2].n4 0.983856
R13176 ua[2].n10 ua[2].n9 0.956356
R13177 ua[2].n26 ua[2].n25 0.946356
R13178 ua[2].n19 ua[2].n18 0.927606
R13179 ua[2].n7 ua[2].n5 0.726502
R13180 ua[2].n16 ua[2].n14 0.726502
R13181 ua[2].n23 ua[2].n21 0.726502
R13182 ua[2].n2 ua[2].n0 0.726502
R13183 ua[2].n11 ua[2] 0.681056
R13184 ua[2].n20 ua[2].n13 0.54925
R13185 ua[2].n27 ua[2].n20 0.54425
R13186 ua[2].n28 ua[2].n27 0.53675
R13187 ua[2].n8 ua[2].n7 0.512491
R13188 ua[2].n17 ua[2].n16 0.512491
R13189 ua[2].n24 ua[2].n23 0.512491
R13190 ua[2].n3 ua[2].n2 0.512491
R13191 ua[2].n9 ua[2].n8 0.359663
R13192 ua[2].n18 ua[2].n17 0.359663
R13193 ua[2].n25 ua[2].n24 0.359663
R13194 ua[2].n4 ua[2].n3 0.359663
R13195 ua[2].n9 ua[2].n5 0.216071
R13196 ua[2].n18 ua[2].n14 0.216071
R13197 ua[2].n25 ua[2].n21 0.216071
R13198 ua[2].n4 ua[2].n0 0.216071
R13199 ua[2].n20 ua[2] 0.18675
R13200 ua[2].n13 ua[2] 0.18425
R13201 ua[2].n27 ua[2] 0.16425
R13202 ua[2] ua[2].n28 0.163
R13203 ua[2].n12 ua[2] 0.135115
R13204 ua[2].n19 ua[2] 0.05675
R13205 ua[2] ua[2].n19 0.0561931
R13206 ua[2].n12 ua[2].n11 0.0530774
R13207 ua[2].n26 ua[2] 0.038
R13208 ua[2] ua[2].n26 0.0376287
R13209 ua[2].n10 ua[2] 0.028
R13210 ua[2] ua[2].n10 0.0266905
R13211 ua[2].n11 ua[2] 0.01175
R13212 ua[2].n13 ua[2].n12 0.006125
R13213 ringtest_0.x4.clknet_0_clk.n33 ringtest_0.x4.clknet_0_clk.n31 333.392
R13214 ringtest_0.x4.clknet_0_clk.n38 ringtest_0.x4.clknet_0_clk.n26 301.392
R13215 ringtest_0.x4.clknet_0_clk.n37 ringtest_0.x4.clknet_0_clk.n27 301.392
R13216 ringtest_0.x4.clknet_0_clk.n36 ringtest_0.x4.clknet_0_clk.n28 301.392
R13217 ringtest_0.x4.clknet_0_clk.n35 ringtest_0.x4.clknet_0_clk.n29 301.392
R13218 ringtest_0.x4.clknet_0_clk.n34 ringtest_0.x4.clknet_0_clk.n30 301.392
R13219 ringtest_0.x4.clknet_0_clk.n33 ringtest_0.x4.clknet_0_clk.n32 301.392
R13220 ringtest_0.x4.clknet_0_clk.n39 ringtest_0.x4.clknet_0_clk.n25 297.863
R13221 ringtest_0.x4.clknet_0_clk.n2 ringtest_0.x4.clknet_0_clk.n0 248.638
R13222 ringtest_0.x4.clknet_0_clk.n2 ringtest_0.x4.clknet_0_clk.n1 203.463
R13223 ringtest_0.x4.clknet_0_clk.n4 ringtest_0.x4.clknet_0_clk.n3 203.463
R13224 ringtest_0.x4.clknet_0_clk.n8 ringtest_0.x4.clknet_0_clk.n7 203.463
R13225 ringtest_0.x4.clknet_0_clk.n24 ringtest_0.x4.clknet_0_clk.n23 203.463
R13226 ringtest_0.x4.clknet_0_clk.n6 ringtest_0.x4.clknet_0_clk.n5 202.456
R13227 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n41 199.607
R13228 ringtest_0.x4.clknet_0_clk.n21 ringtest_0.x4.clknet_0_clk.n9 188.201
R13229 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.t46 184.768
R13230 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.t43 184.768
R13231 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.t42 184.768
R13232 ringtest_0.x4.clknet_0_clk.n15 ringtest_0.x4.clknet_0_clk.t45 184.768
R13233 ringtest_0.x4.clknet_0_clk.n10 ringtest_0.x4.clknet_0_clk.t41 184.768
R13234 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.t37 184.768
R13235 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.t40 184.768
R13236 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.t39 184.768
R13237 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n18 173.609
R13238 ringtest_0.x4.clknet_0_clk.n14 ringtest_0.x4.clknet_0_clk.n13 171.375
R13239 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.t38 146.208
R13240 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.t35 146.208
R13241 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.t34 146.208
R13242 ringtest_0.x4.clknet_0_clk.n15 ringtest_0.x4.clknet_0_clk.t36 146.208
R13243 ringtest_0.x4.clknet_0_clk.n10 ringtest_0.x4.clknet_0_clk.t33 146.208
R13244 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.t44 146.208
R13245 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.t32 146.208
R13246 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.t47 146.208
R13247 ringtest_0.x4.clknet_0_clk.n4 ringtest_0.x4.clknet_0_clk.n2 45.177
R13248 ringtest_0.x4.clknet_0_clk.n22 ringtest_0.x4.clknet_0_clk.n8 45.177
R13249 ringtest_0.x4.clknet_0_clk.n24 ringtest_0.x4.clknet_0_clk.n22 45.177
R13250 ringtest_0.x4.clknet_0_clk.n6 ringtest_0.x4.clknet_0_clk.n4 44.0476
R13251 ringtest_0.x4.clknet_0_clk.n8 ringtest_0.x4.clknet_0_clk.n6 44.0476
R13252 ringtest_0.x4.clknet_0_clk.n18 ringtest_0.x4.clknet_0_clk.n17 40.6397
R13253 ringtest_0.x4.clknet_0_clk.n17 ringtest_0.x4.clknet_0_clk.n16 40.6397
R13254 ringtest_0.x4.clknet_0_clk.n16 ringtest_0.x4.clknet_0_clk.n15 40.6397
R13255 ringtest_0.x4.clknet_0_clk.n11 ringtest_0.x4.clknet_0_clk.n10 40.6397
R13256 ringtest_0.x4.clknet_0_clk.n12 ringtest_0.x4.clknet_0_clk.n11 40.6397
R13257 ringtest_0.x4.clknet_0_clk.n13 ringtest_0.x4.clknet_0_clk.n12 40.6397
R13258 ringtest_0.x4.clknet_0_clk.n0 ringtest_0.x4.clknet_0_clk.t18 40.0005
R13259 ringtest_0.x4.clknet_0_clk.n0 ringtest_0.x4.clknet_0_clk.t31 40.0005
R13260 ringtest_0.x4.clknet_0_clk.n1 ringtest_0.x4.clknet_0_clk.t20 40.0005
R13261 ringtest_0.x4.clknet_0_clk.n1 ringtest_0.x4.clknet_0_clk.t22 40.0005
R13262 ringtest_0.x4.clknet_0_clk.n3 ringtest_0.x4.clknet_0_clk.t24 40.0005
R13263 ringtest_0.x4.clknet_0_clk.n3 ringtest_0.x4.clknet_0_clk.t26 40.0005
R13264 ringtest_0.x4.clknet_0_clk.n5 ringtest_0.x4.clknet_0_clk.t21 40.0005
R13265 ringtest_0.x4.clknet_0_clk.n5 ringtest_0.x4.clknet_0_clk.t23 40.0005
R13266 ringtest_0.x4.clknet_0_clk.n7 ringtest_0.x4.clknet_0_clk.t25 40.0005
R13267 ringtest_0.x4.clknet_0_clk.n7 ringtest_0.x4.clknet_0_clk.t27 40.0005
R13268 ringtest_0.x4.clknet_0_clk.n9 ringtest_0.x4.clknet_0_clk.t16 40.0005
R13269 ringtest_0.x4.clknet_0_clk.n9 ringtest_0.x4.clknet_0_clk.t29 40.0005
R13270 ringtest_0.x4.clknet_0_clk.n23 ringtest_0.x4.clknet_0_clk.t30 40.0005
R13271 ringtest_0.x4.clknet_0_clk.n23 ringtest_0.x4.clknet_0_clk.t28 40.0005
R13272 ringtest_0.x4.clknet_0_clk.n41 ringtest_0.x4.clknet_0_clk.t17 40.0005
R13273 ringtest_0.x4.clknet_0_clk.n41 ringtest_0.x4.clknet_0_clk.t19 40.0005
R13274 ringtest_0.x4.clknet_0_clk.n38 ringtest_0.x4.clknet_0_clk.n37 32.0005
R13275 ringtest_0.x4.clknet_0_clk.n37 ringtest_0.x4.clknet_0_clk.n36 32.0005
R13276 ringtest_0.x4.clknet_0_clk.n35 ringtest_0.x4.clknet_0_clk.n34 32.0005
R13277 ringtest_0.x4.clknet_0_clk.n34 ringtest_0.x4.clknet_0_clk.n33 32.0005
R13278 ringtest_0.x4.clknet_0_clk.n36 ringtest_0.x4.clknet_0_clk.n35 31.2005
R13279 ringtest_0.x4.clknet_0_clk.n31 ringtest_0.x4.clknet_0_clk.t11 27.5805
R13280 ringtest_0.x4.clknet_0_clk.n31 ringtest_0.x4.clknet_0_clk.t8 27.5805
R13281 ringtest_0.x4.clknet_0_clk.n26 ringtest_0.x4.clknet_0_clk.t7 27.5805
R13282 ringtest_0.x4.clknet_0_clk.n26 ringtest_0.x4.clknet_0_clk.t5 27.5805
R13283 ringtest_0.x4.clknet_0_clk.n25 ringtest_0.x4.clknet_0_clk.t10 27.5805
R13284 ringtest_0.x4.clknet_0_clk.n25 ringtest_0.x4.clknet_0_clk.t12 27.5805
R13285 ringtest_0.x4.clknet_0_clk.n27 ringtest_0.x4.clknet_0_clk.t9 27.5805
R13286 ringtest_0.x4.clknet_0_clk.n27 ringtest_0.x4.clknet_0_clk.t6 27.5805
R13287 ringtest_0.x4.clknet_0_clk.n28 ringtest_0.x4.clknet_0_clk.t2 27.5805
R13288 ringtest_0.x4.clknet_0_clk.n28 ringtest_0.x4.clknet_0_clk.t4 27.5805
R13289 ringtest_0.x4.clknet_0_clk.n29 ringtest_0.x4.clknet_0_clk.t14 27.5805
R13290 ringtest_0.x4.clknet_0_clk.n29 ringtest_0.x4.clknet_0_clk.t0 27.5805
R13291 ringtest_0.x4.clknet_0_clk.n30 ringtest_0.x4.clknet_0_clk.t1 27.5805
R13292 ringtest_0.x4.clknet_0_clk.n30 ringtest_0.x4.clknet_0_clk.t3 27.5805
R13293 ringtest_0.x4.clknet_0_clk.n32 ringtest_0.x4.clknet_0_clk.t13 27.5805
R13294 ringtest_0.x4.clknet_0_clk.n32 ringtest_0.x4.clknet_0_clk.t15 27.5805
R13295 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n14 25.9814
R13296 ringtest_0.x4.clknet_0_clk.n22 ringtest_0.x4.clknet_0_clk.n21 15.262
R13297 ringtest_0.x4.clknet_0_clk.n20 ringtest_0.x4.clknet_0_clk.n19 14.7771
R13298 ringtest_0.x4.clknet_0_clk.n40 ringtest_0.x4.clknet_0_clk.n24 13.177
R13299 ringtest_0.x4.clknet_0_clk.n39 ringtest_0.x4.clknet_0_clk.n38 10.4484
R13300 ringtest_0.x4.clknet_0_clk.n19 ringtest_0.x4.clknet_0_clk 10.3624
R13301 ringtest_0.x4.clknet_0_clk.n21 ringtest_0.x4.clknet_0_clk.n20 9.3005
R13302 ringtest_0.x4.clknet_0_clk.n19 ringtest_0.x4.clknet_0_clk 3.45447
R13303 ringtest_0.x4.clknet_0_clk.n40 ringtest_0.x4.clknet_0_clk 3.13183
R13304 ringtest_0.x4.clknet_0_clk.n14 ringtest_0.x4.clknet_0_clk 2.23542
R13305 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n39 1.75844
R13306 ringtest_0.x4.clknet_0_clk.n20 ringtest_0.x4.clknet_0_clk 1.5927
R13307 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_0_clk.n40 0.604792
R13308 ringtest_0.x4.net6.n3 ringtest_0.x4.net6.t13 323.342
R13309 ringtest_0.x4.net6.n0 ringtest_0.x4.net6.t4 323.342
R13310 ringtest_0.x4.net6.n1 ringtest_0.x4.net6.t2 260.322
R13311 ringtest_0.x4.net6.n8 ringtest_0.x4.net6.t5 241.536
R13312 ringtest_0.x4.net6.n17 ringtest_0.x4.net6.t0 222.679
R13313 ringtest_0.x4.net6.n12 ringtest_0.x4.net6.t14 212.081
R13314 ringtest_0.x4.net6.n13 ringtest_0.x4.net6.t7 212.081
R13315 ringtest_0.x4.net6.n3 ringtest_0.x4.net6.t6 194.809
R13316 ringtest_0.x4.net6.n0 ringtest_0.x4.net6.t8 194.809
R13317 ringtest_0.x4.net6.n5 ringtest_0.x4.net6.t10 183.505
R13318 ringtest_0.x4.net6.n1 ringtest_0.x4.net6.t12 175.169
R13319 ringtest_0.x4.net6.n8 ringtest_0.x4.net6.t11 169.237
R13320 ringtest_0.x4.net6 ringtest_0.x4.net6.n3 158.133
R13321 ringtest_0.x4.net6 ringtest_0.x4.net6.n0 158.133
R13322 ringtest_0.x4.net6 ringtest_0.x4.net6.n8 157.555
R13323 ringtest_0.x4.net6.n15 ringtest_0.x4.net6.n14 155.52
R13324 ringtest_0.x4.net6.n6 ringtest_0.x4.net6.n5 153.863
R13325 ringtest_0.x4.net6.n2 ringtest_0.x4.net6.n1 152
R13326 ringtest_0.x4.net6.n12 ringtest_0.x4.net6.t9 139.78
R13327 ringtest_0.x4.net6.n13 ringtest_0.x4.net6.t15 139.78
R13328 ringtest_0.x4.net6.n18 ringtest_0.x4.net6.t1 129.078
R13329 ringtest_0.x4.net6.n5 ringtest_0.x4.net6.t3 114.532
R13330 ringtest_0.x4.net6.n18 ringtest_0.x4.net6.n17 96.7191
R13331 ringtest_0.x4.net6.n11 ringtest_0.x4.net6 55.2785
R13332 ringtest_0.x4.net6.n14 ringtest_0.x4.net6.n13 37.246
R13333 ringtest_0.x4.net6.n14 ringtest_0.x4.net6.n12 24.1005
R13334 ringtest_0.x4.net6.n10 ringtest_0.x4.net6.n9 21.4124
R13335 ringtest_0.x4.net6.n16 ringtest_0.x4.net6.n15 21.1949
R13336 ringtest_0.x4.net6.n4 ringtest_0.x4.net6.n2 20.043
R13337 ringtest_0.x4.net6.n7 ringtest_0.x4.net6.n6 15.2615
R13338 ringtest_0.x4.net6.n17 ringtest_0.x4.net6.n16 12.4213
R13339 ringtest_0.x4.net6.n9 ringtest_0.x4.net6 12.3175
R13340 ringtest_0.x4.net6.n16 ringtest_0.x4.net6.n11 8.09819
R13341 ringtest_0.x4.net6.n11 ringtest_0.x4.net6.n10 7.53948
R13342 ringtest_0.x4.net6.n4 ringtest_0.x4.net6 7.39885
R13343 ringtest_0.x4.net6 ringtest_0.x4.net6.n18 5.84085
R13344 ringtest_0.x4.net6.n15 ringtest_0.x4.net6 5.4405
R13345 ringtest_0.x4.net6.n9 ringtest_0.x4.net6 4.10616
R13346 ringtest_0.x4.net6.n7 ringtest_0.x4.net6.n4 2.60421
R13347 ringtest_0.x4.net6.n10 ringtest_0.x4.net6.n7 2.43577
R13348 ringtest_0.x4.net6.n6 ringtest_0.x4.net6 1.97868
R13349 ringtest_0.x4.net6.n2 ringtest_0.x4.net6 1.55726
R13350 ringtest_0.x4.clknet_1_1__leaf_clk.n29 ringtest_0.x4.clknet_1_1__leaf_clk.n27 333.392
R13351 ringtest_0.x4.clknet_1_1__leaf_clk.n29 ringtest_0.x4.clknet_1_1__leaf_clk.n28 301.392
R13352 ringtest_0.x4.clknet_1_1__leaf_clk.n31 ringtest_0.x4.clknet_1_1__leaf_clk.n30 301.392
R13353 ringtest_0.x4.clknet_1_1__leaf_clk.n33 ringtest_0.x4.clknet_1_1__leaf_clk.n32 301.392
R13354 ringtest_0.x4.clknet_1_1__leaf_clk.n35 ringtest_0.x4.clknet_1_1__leaf_clk.n34 301.392
R13355 ringtest_0.x4.clknet_1_1__leaf_clk.n37 ringtest_0.x4.clknet_1_1__leaf_clk.n36 301.392
R13356 ringtest_0.x4.clknet_1_1__leaf_clk.n39 ringtest_0.x4.clknet_1_1__leaf_clk.n38 301.392
R13357 ringtest_0.x4.clknet_1_1__leaf_clk.n40 ringtest_0.x4.clknet_1_1__leaf_clk.n26 297.863
R13358 ringtest_0.x4.clknet_1_1__leaf_clk.n18 ringtest_0.x4.clknet_1_1__leaf_clk.t36 294.557
R13359 ringtest_0.x4.clknet_1_1__leaf_clk.n15 ringtest_0.x4.clknet_1_1__leaf_clk.t33 294.557
R13360 ringtest_0.x4.clknet_1_1__leaf_clk.n13 ringtest_0.x4.clknet_1_1__leaf_clk.t34 294.557
R13361 ringtest_0.x4.clknet_1_1__leaf_clk.n11 ringtest_0.x4.clknet_1_1__leaf_clk.t41 294.557
R13362 ringtest_0.x4.clknet_1_1__leaf_clk.n10 ringtest_0.x4.clknet_1_1__leaf_clk.t32 294.557
R13363 ringtest_0.x4.clknet_1_1__leaf_clk.n2 ringtest_0.x4.clknet_1_1__leaf_clk.n0 248.638
R13364 ringtest_0.x4.clknet_1_1__leaf_clk.n18 ringtest_0.x4.clknet_1_1__leaf_clk.t39 211.01
R13365 ringtest_0.x4.clknet_1_1__leaf_clk.n15 ringtest_0.x4.clknet_1_1__leaf_clk.t40 211.01
R13366 ringtest_0.x4.clknet_1_1__leaf_clk.n13 ringtest_0.x4.clknet_1_1__leaf_clk.t38 211.01
R13367 ringtest_0.x4.clknet_1_1__leaf_clk.n11 ringtest_0.x4.clknet_1_1__leaf_clk.t35 211.01
R13368 ringtest_0.x4.clknet_1_1__leaf_clk.n10 ringtest_0.x4.clknet_1_1__leaf_clk.t37 211.01
R13369 ringtest_0.x4.clknet_1_1__leaf_clk.n2 ringtest_0.x4.clknet_1_1__leaf_clk.n1 203.463
R13370 ringtest_0.x4.clknet_1_1__leaf_clk.n4 ringtest_0.x4.clknet_1_1__leaf_clk.n3 203.463
R13371 ringtest_0.x4.clknet_1_1__leaf_clk.n8 ringtest_0.x4.clknet_1_1__leaf_clk.n7 203.463
R13372 ringtest_0.x4.clknet_1_1__leaf_clk.n25 ringtest_0.x4.clknet_1_1__leaf_clk.n24 203.463
R13373 ringtest_0.x4.clknet_1_1__leaf_clk.n6 ringtest_0.x4.clknet_1_1__leaf_clk.n5 202.456
R13374 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n42 199.607
R13375 ringtest_0.x4.clknet_1_1__leaf_clk.n22 ringtest_0.x4.clknet_1_1__leaf_clk.n9 188.201
R13376 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n13 156.207
R13377 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n10 156.207
R13378 ringtest_0.x4.clknet_1_1__leaf_clk.n19 ringtest_0.x4.clknet_1_1__leaf_clk.n18 153.097
R13379 ringtest_0.x4.clknet_1_1__leaf_clk.n16 ringtest_0.x4.clknet_1_1__leaf_clk.n15 152.296
R13380 ringtest_0.x4.clknet_1_1__leaf_clk.n12 ringtest_0.x4.clknet_1_1__leaf_clk.n11 152.296
R13381 ringtest_0.x4.clknet_1_1__leaf_clk.n4 ringtest_0.x4.clknet_1_1__leaf_clk.n2 45.177
R13382 ringtest_0.x4.clknet_1_1__leaf_clk.n23 ringtest_0.x4.clknet_1_1__leaf_clk.n8 45.177
R13383 ringtest_0.x4.clknet_1_1__leaf_clk.n25 ringtest_0.x4.clknet_1_1__leaf_clk.n23 45.177
R13384 ringtest_0.x4.clknet_1_1__leaf_clk.n6 ringtest_0.x4.clknet_1_1__leaf_clk.n4 44.0476
R13385 ringtest_0.x4.clknet_1_1__leaf_clk.n8 ringtest_0.x4.clknet_1_1__leaf_clk.n6 44.0476
R13386 ringtest_0.x4.clknet_1_1__leaf_clk.n0 ringtest_0.x4.clknet_1_1__leaf_clk.t29 40.0005
R13387 ringtest_0.x4.clknet_1_1__leaf_clk.n0 ringtest_0.x4.clknet_1_1__leaf_clk.t30 40.0005
R13388 ringtest_0.x4.clknet_1_1__leaf_clk.n1 ringtest_0.x4.clknet_1_1__leaf_clk.t31 40.0005
R13389 ringtest_0.x4.clknet_1_1__leaf_clk.n1 ringtest_0.x4.clknet_1_1__leaf_clk.t28 40.0005
R13390 ringtest_0.x4.clknet_1_1__leaf_clk.n3 ringtest_0.x4.clknet_1_1__leaf_clk.t27 40.0005
R13391 ringtest_0.x4.clknet_1_1__leaf_clk.n3 ringtest_0.x4.clknet_1_1__leaf_clk.t26 40.0005
R13392 ringtest_0.x4.clknet_1_1__leaf_clk.n5 ringtest_0.x4.clknet_1_1__leaf_clk.t22 40.0005
R13393 ringtest_0.x4.clknet_1_1__leaf_clk.n5 ringtest_0.x4.clknet_1_1__leaf_clk.t24 40.0005
R13394 ringtest_0.x4.clknet_1_1__leaf_clk.n7 ringtest_0.x4.clknet_1_1__leaf_clk.t18 40.0005
R13395 ringtest_0.x4.clknet_1_1__leaf_clk.n7 ringtest_0.x4.clknet_1_1__leaf_clk.t20 40.0005
R13396 ringtest_0.x4.clknet_1_1__leaf_clk.n9 ringtest_0.x4.clknet_1_1__leaf_clk.t21 40.0005
R13397 ringtest_0.x4.clknet_1_1__leaf_clk.n9 ringtest_0.x4.clknet_1_1__leaf_clk.t23 40.0005
R13398 ringtest_0.x4.clknet_1_1__leaf_clk.n24 ringtest_0.x4.clknet_1_1__leaf_clk.t17 40.0005
R13399 ringtest_0.x4.clknet_1_1__leaf_clk.n24 ringtest_0.x4.clknet_1_1__leaf_clk.t25 40.0005
R13400 ringtest_0.x4.clknet_1_1__leaf_clk.n42 ringtest_0.x4.clknet_1_1__leaf_clk.t19 40.0005
R13401 ringtest_0.x4.clknet_1_1__leaf_clk.n42 ringtest_0.x4.clknet_1_1__leaf_clk.t16 40.0005
R13402 ringtest_0.x4.clknet_1_1__leaf_clk.n21 ringtest_0.x4.clknet_1_1__leaf_clk 34.5053
R13403 ringtest_0.x4.clknet_1_1__leaf_clk.n14 ringtest_0.x4.clknet_1_1__leaf_clk 33.8485
R13404 ringtest_0.x4.clknet_1_1__leaf_clk.n31 ringtest_0.x4.clknet_1_1__leaf_clk.n29 32.0005
R13405 ringtest_0.x4.clknet_1_1__leaf_clk.n33 ringtest_0.x4.clknet_1_1__leaf_clk.n31 32.0005
R13406 ringtest_0.x4.clknet_1_1__leaf_clk.n37 ringtest_0.x4.clknet_1_1__leaf_clk.n35 32.0005
R13407 ringtest_0.x4.clknet_1_1__leaf_clk.n39 ringtest_0.x4.clknet_1_1__leaf_clk.n37 32.0005
R13408 ringtest_0.x4.clknet_1_1__leaf_clk.n35 ringtest_0.x4.clknet_1_1__leaf_clk.n33 31.2005
R13409 ringtest_0.x4.clknet_1_1__leaf_clk.n27 ringtest_0.x4.clknet_1_1__leaf_clk.t3 27.5805
R13410 ringtest_0.x4.clknet_1_1__leaf_clk.n27 ringtest_0.x4.clknet_1_1__leaf_clk.t4 27.5805
R13411 ringtest_0.x4.clknet_1_1__leaf_clk.n28 ringtest_0.x4.clknet_1_1__leaf_clk.t5 27.5805
R13412 ringtest_0.x4.clknet_1_1__leaf_clk.n28 ringtest_0.x4.clknet_1_1__leaf_clk.t2 27.5805
R13413 ringtest_0.x4.clknet_1_1__leaf_clk.n30 ringtest_0.x4.clknet_1_1__leaf_clk.t1 27.5805
R13414 ringtest_0.x4.clknet_1_1__leaf_clk.n30 ringtest_0.x4.clknet_1_1__leaf_clk.t0 27.5805
R13415 ringtest_0.x4.clknet_1_1__leaf_clk.n32 ringtest_0.x4.clknet_1_1__leaf_clk.t12 27.5805
R13416 ringtest_0.x4.clknet_1_1__leaf_clk.n32 ringtest_0.x4.clknet_1_1__leaf_clk.t14 27.5805
R13417 ringtest_0.x4.clknet_1_1__leaf_clk.n34 ringtest_0.x4.clknet_1_1__leaf_clk.t8 27.5805
R13418 ringtest_0.x4.clknet_1_1__leaf_clk.n34 ringtest_0.x4.clknet_1_1__leaf_clk.t10 27.5805
R13419 ringtest_0.x4.clknet_1_1__leaf_clk.n36 ringtest_0.x4.clknet_1_1__leaf_clk.t11 27.5805
R13420 ringtest_0.x4.clknet_1_1__leaf_clk.n36 ringtest_0.x4.clknet_1_1__leaf_clk.t13 27.5805
R13421 ringtest_0.x4.clknet_1_1__leaf_clk.n26 ringtest_0.x4.clknet_1_1__leaf_clk.t9 27.5805
R13422 ringtest_0.x4.clknet_1_1__leaf_clk.n26 ringtest_0.x4.clknet_1_1__leaf_clk.t6 27.5805
R13423 ringtest_0.x4.clknet_1_1__leaf_clk.n38 ringtest_0.x4.clknet_1_1__leaf_clk.t7 27.5805
R13424 ringtest_0.x4.clknet_1_1__leaf_clk.n38 ringtest_0.x4.clknet_1_1__leaf_clk.t15 27.5805
R13425 ringtest_0.x4.clknet_1_1__leaf_clk.n23 ringtest_0.x4.clknet_1_1__leaf_clk.n22 15.262
R13426 ringtest_0.x4.clknet_1_1__leaf_clk.n20 ringtest_0.x4.clknet_1_1__leaf_clk.n19 13.8005
R13427 ringtest_0.x4.clknet_1_1__leaf_clk.n41 ringtest_0.x4.clknet_1_1__leaf_clk.n25 13.177
R13428 ringtest_0.x4.clknet_1_1__leaf_clk.n14 ringtest_0.x4.clknet_1_1__leaf_clk.n12 11.6482
R13429 ringtest_0.x4.clknet_1_1__leaf_clk.n22 ringtest_0.x4.clknet_1_1__leaf_clk.n21 10.8268
R13430 ringtest_0.x4.clknet_1_1__leaf_clk.n40 ringtest_0.x4.clknet_1_1__leaf_clk.n39 10.4484
R13431 ringtest_0.x4.clknet_1_1__leaf_clk.n17 ringtest_0.x4.clknet_1_1__leaf_clk.n16 9.3005
R13432 ringtest_0.x4.clknet_1_1__leaf_clk.n20 ringtest_0.x4.clknet_1_1__leaf_clk.n17 8.37704
R13433 ringtest_0.x4.clknet_1_1__leaf_clk.n21 ringtest_0.x4.clknet_1_1__leaf_clk 5.19349
R13434 ringtest_0.x4.clknet_1_1__leaf_clk.n17 ringtest_0.x4.clknet_1_1__leaf_clk.n14 3.99105
R13435 ringtest_0.x4.clknet_1_1__leaf_clk.n41 ringtest_0.x4.clknet_1_1__leaf_clk 3.13183
R13436 ringtest_0.x4.clknet_1_1__leaf_clk.n19 ringtest_0.x4.clknet_1_1__leaf_clk 3.10907
R13437 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n40 1.75844
R13438 ringtest_0.x4.clknet_1_1__leaf_clk.n16 ringtest_0.x4.clknet_1_1__leaf_clk 1.67435
R13439 ringtest_0.x4.clknet_1_1__leaf_clk.n12 ringtest_0.x4.clknet_1_1__leaf_clk 1.67435
R13440 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n20 0.693495
R13441 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.clknet_1_1__leaf_clk.n41 0.604792
R13442 ui_in[1].n10 ui_in[1].t8 327.99
R13443 ui_in[1].n3 ui_in[1].t1 293.969
R13444 ui_in[1].n6 ui_in[1].t7 256.07
R13445 ui_in[1].n0 ui_in[1].t0 212.081
R13446 ui_in[1].n1 ui_in[1].t2 212.081
R13447 ui_in[1].n10 ui_in[1].t9 199.457
R13448 ui_in[1].n2 ui_in[1].n1 182.929
R13449 ui_in[1] ui_in[1].n3 154.065
R13450 ui_in[1].n11 ui_in[1].n10 152
R13451 ui_in[1].n7 ui_in[1].n6 152
R13452 ui_in[1].n6 ui_in[1].t3 150.03
R13453 ui_in[1].n0 ui_in[1].t5 139.78
R13454 ui_in[1].n1 ui_in[1].t6 139.78
R13455 ui_in[1].n3 ui_in[1].t4 138.338
R13456 ui_in[1].n1 ui_in[1].n0 61.346
R13457 ui_in[1].n16 ui_in[1] 30.7401
R13458 ui_in[1].n5 ui_in[1] 17.455
R13459 ui_in[1].n14 ui_in[1].n13 14.6836
R13460 ui_in[1].n13 ui_in[1].n12 14.6704
R13461 ui_in[1].n4 ui_in[1] 13.8328
R13462 ui_in[1].n14 ui_in[1].n2 10.6811
R13463 ui_in[1].n7 ui_in[1].n5 10.4374
R13464 ui_in[1].n9 ui_in[1].n8 8.15776
R13465 ui_in[1].n12 ui_in[1] 6.61383
R13466 ui_in[1].n2 ui_in[1] 6.1445
R13467 ui_in[1].n4 ui_in[1] 5.16179
R13468 ui_in[1].n11 ui_in[1] 4.90717
R13469 ui_in[1].n9 ui_in[1].n4 4.65206
R13470 ui_in[1].n15 ui_in[1] 4.54217
R13471 ui_in[1].n8 ui_in[1] 3.93896
R13472 ui_in[1].n12 ui_in[1].n11 2.98717
R13473 ui_in[1].n5 ui_in[1] 2.16665
R13474 ui_in[1].n8 ui_in[1].n7 1.57588
R13475 ui_in[1].n13 ui_in[1].n9 0.79438
R13476 ui_in[1].n15 ui_in[1] 0.606561
R13477 ui_in[1] ui_in[1].n14 0.248606
R13478 ui_in[1] ui_in[1].n15 0.222091
R13479 ui_in[1] ui_in[1].n16 0.122375
R13480 ui_in[1].n16 ui_in[1] 0.121168
R13481 muxtest_0.x1.x3.GP1.n3 muxtest_0.x1.x3.GP1.t4 450.938
R13482 muxtest_0.x1.x3.GP1.n2 muxtest_0.x1.x3.GP1.t6 450.938
R13483 muxtest_0.x1.x3.GP1.n3 muxtest_0.x1.x3.GP1.t5 445.666
R13484 muxtest_0.x1.x3.GP1.n2 muxtest_0.x1.x3.GP1.t7 445.666
R13485 muxtest_0.x1.x3.GP1.n6 muxtest_0.x1.x3.GP1.n5 195.832
R13486 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n0 96.8352
R13487 muxtest_0.x1.x3.GP1.n5 muxtest_0.x1.x3.GP1.t0 26.5955
R13488 muxtest_0.x1.x3.GP1.n5 muxtest_0.x1.x3.GP1.t1 26.5955
R13489 muxtest_0.x1.x3.GP1.n0 muxtest_0.x1.x3.GP1.t3 24.9236
R13490 muxtest_0.x1.x3.GP1.n0 muxtest_0.x1.x3.GP1.t2 24.9236
R13491 muxtest_0.x1.x3.GP1.n4 muxtest_0.x1.x3.GP1 13.257
R13492 muxtest_0.x1.x3.GP1.n7 muxtest_0.x1.x3.GP1.n6 13.1346
R13493 muxtest_0.x1.x3.GP1.n6 muxtest_0.x1.x3.GP1 11.8965
R13494 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n1 11.2645
R13495 muxtest_0.x1.x3.GP1.n1 muxtest_0.x1.x3.GP1 6.1445
R13496 muxtest_0.x1.x3.GP1.n4 muxtest_0.x1.x3.GP1 5.31412
R13497 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n4 5.26828
R13498 muxtest_0.x1.x3.GP1.n1 muxtest_0.x1.x3.GP1 4.65505
R13499 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n2 3.07895
R13500 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n3 2.90754
R13501 muxtest_0.x1.x3.GP1.n7 muxtest_0.x1.x3.GP1 2.0485
R13502 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP1.n7 1.55202
R13503 muxtest_0.x1.x3.GP4.n3 muxtest_0.x1.x3.GP4.t5 450.938
R13504 muxtest_0.x1.x3.GP4.n2 muxtest_0.x1.x3.GP4.t7 450.938
R13505 muxtest_0.x1.x3.GP4.n3 muxtest_0.x1.x3.GP4.t4 445.666
R13506 muxtest_0.x1.x3.GP4.n2 muxtest_0.x1.x3.GP4.t6 445.666
R13507 muxtest_0.x1.x3.GP4.n7 muxtest_0.x1.x3.GP4.n6 208.965
R13508 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n0 96.8352
R13509 muxtest_0.x1.x3.GP4.n6 muxtest_0.x1.x3.GP4.t0 26.5955
R13510 muxtest_0.x1.x3.GP4.n6 muxtest_0.x1.x3.GP4.t1 26.5955
R13511 muxtest_0.x1.x3.GP4.n0 muxtest_0.x1.x3.GP4.t3 24.9236
R13512 muxtest_0.x1.x3.GP4.n0 muxtest_0.x1.x3.GP4.t2 24.9236
R13513 muxtest_0.x1.x3.GP4.n4 muxtest_0.x1.x3.x4.GP 10.9863
R13514 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n5 10.2405
R13515 muxtest_0.x1.x1.gpo3 muxtest_0.x1.x3.GP4.n4 9.34192
R13516 muxtest_0.x1.x3.GP4.n5 muxtest_0.x1.x1.gpo3 7.73829
R13517 muxtest_0.x1.x3.GP4.n1 muxtest_0.x1.x1.x14.Y 6.1445
R13518 muxtest_0.x1.x3.GP4.n4 muxtest_0.x1.x2.x4.GP 5.84951
R13519 muxtest_0.x1.x3.GP4.n1 muxtest_0.x1.x1.x14.Y 4.65505
R13520 muxtest_0.x1.x2.x4.GP muxtest_0.x1.x3.GP4.n3 2.95993
R13521 muxtest_0.x1.x3.x4.GP muxtest_0.x1.x3.GP4.n2 2.95993
R13522 muxtest_0.x1.x3.GP4.n7 muxtest_0.x1.x1.x14.Y 2.0485
R13523 muxtest_0.x1.x1.x14.Y muxtest_0.x1.x3.GP4.n7 1.55202
R13524 muxtest_0.x1.x3.GP4.n5 muxtest_0.x1.x3.GP4.n1 1.0245
R13525 ringtest_0.x4._11_ ringtest_0.x4._11_.n0 623.909
R13526 ringtest_0.x4._11_.n24 ringtest_0.x4._11_.t6 334.723
R13527 ringtest_0.x4._11_.n5 ringtest_0.x4._11_.t5 334.723
R13528 ringtest_0.x4._11_.n18 ringtest_0.x4._11_.t19 261.887
R13529 ringtest_0.x4._11_.n14 ringtest_0.x4._11_.t14 256.07
R13530 ringtest_0.x4._11_.n8 ringtest_0.x4._11_.t10 241.536
R13531 ringtest_0.x4._11_.n3 ringtest_0.x4._11_.t13 241.536
R13532 ringtest_0.x4._11_.n1 ringtest_0.x4._11_.t12 231.835
R13533 ringtest_0.x4._11_.n21 ringtest_0.x4._11_.t8 230.363
R13534 ringtest_0.x4._11_ ringtest_0.x4._11_.n30 216.464
R13535 ringtest_0.x4._11_.n24 ringtest_0.x4._11_.t20 206.19
R13536 ringtest_0.x4._11_.n5 ringtest_0.x4._11_.t17 206.19
R13537 ringtest_0.x4._11_.n11 ringtest_0.x4._11_.t11 183.505
R13538 ringtest_0.x4._11_.n8 ringtest_0.x4._11_.t21 169.237
R13539 ringtest_0.x4._11_.n3 ringtest_0.x4._11_.t7 169.237
R13540 ringtest_0.x4._11_.n21 ringtest_0.x4._11_.t16 158.064
R13541 ringtest_0.x4._11_ ringtest_0.x4._11_.n3 157.555
R13542 ringtest_0.x4._11_ ringtest_0.x4._11_.n8 157.166
R13543 ringtest_0.x4._11_.n1 ringtest_0.x4._11_.t9 157.07
R13544 ringtest_0.x4._11_.n18 ringtest_0.x4._11_.t15 155.847
R13545 ringtest_0.x4._11_.n22 ringtest_0.x4._11_.n21 154.048
R13546 ringtest_0.x4._11_.n12 ringtest_0.x4._11_.n11 153.863
R13547 ringtest_0.x4._11_.n19 ringtest_0.x4._11_.n18 153.13
R13548 ringtest_0.x4._11_.n25 ringtest_0.x4._11_.n24 152
R13549 ringtest_0.x4._11_.n15 ringtest_0.x4._11_.n14 152
R13550 ringtest_0.x4._11_.n6 ringtest_0.x4._11_.n5 152
R13551 ringtest_0.x4._11_.n2 ringtest_0.x4._11_.n1 152
R13552 ringtest_0.x4._11_.n14 ringtest_0.x4._11_.t4 150.03
R13553 ringtest_0.x4._11_.n11 ringtest_0.x4._11_.t18 114.532
R13554 ringtest_0.x4._11_.n27 ringtest_0.x4._11_.n26 41.0809
R13555 ringtest_0.x4._11_.n30 ringtest_0.x4._11_.t2 38.5719
R13556 ringtest_0.x4._11_.n30 ringtest_0.x4._11_.t3 38.5719
R13557 ringtest_0.x4._11_.n0 ringtest_0.x4._11_.t1 26.5955
R13558 ringtest_0.x4._11_.n0 ringtest_0.x4._11_.t0 26.5955
R13559 ringtest_0.x4._11_.n17 ringtest_0.x4._11_.n16 25.2401
R13560 ringtest_0.x4._11_.n20 ringtest_0.x4._11_.n19 22.3199
R13561 ringtest_0.x4._11_.n10 ringtest_0.x4._11_.n9 21.8442
R13562 ringtest_0.x4._11_.n10 ringtest_0.x4._11_.n7 20.8523
R13563 ringtest_0.x4._11_.n28 ringtest_0.x4._11_.n27 13.7699
R13564 ringtest_0.x4._11_.n28 ringtest_0.x4._11_.n2 12.7179
R13565 ringtest_0.x4._11_.n4 ringtest_0.x4._11_ 12.3175
R13566 ringtest_0.x4._11_.n9 ringtest_0.x4._11_ 11.4531
R13567 ringtest_0.x4._11_.n7 ringtest_0.x4._11_.n4 11.4418
R13568 ringtest_0.x4._11_.n23 ringtest_0.x4._11_.n20 10.8618
R13569 ringtest_0.x4._11_.n7 ringtest_0.x4._11_.n6 10.3976
R13570 ringtest_0.x4._11_.n25 ringtest_0.x4._11_ 9.6005
R13571 ringtest_0.x4._11_.n29 ringtest_0.x4._11_ 9.6005
R13572 ringtest_0.x4._11_ ringtest_0.x4._11_.n22 9.39918
R13573 ringtest_0.x4._11_.n13 ringtest_0.x4._11_.n12 9.3005
R13574 ringtest_0.x4._11_.n29 ringtest_0.x4._11_.n28 9.3005
R13575 ringtest_0.x4._11_.n23 ringtest_0.x4._11_ 8.80957
R13576 ringtest_0.x4._11_.n6 ringtest_0.x4._11_ 8.22907
R13577 ringtest_0.x4._11_.n15 ringtest_0.x4._11_ 7.6805
R13578 ringtest_0.x4._11_.n16 ringtest_0.x4._11_.n15 4.6085
R13579 ringtest_0.x4._11_.n16 ringtest_0.x4._11_ 4.58918
R13580 ringtest_0.x4._11_.n22 ringtest_0.x4._11_ 4.3525
R13581 ringtest_0.x4._11_.n4 ringtest_0.x4._11_ 4.10616
R13582 ringtest_0.x4._11_.n9 ringtest_0.x4._11_ 3.81804
R13583 ringtest_0.x4._11_.n26 ringtest_0.x4._11_ 3.62717
R13584 ringtest_0.x4._11_.n19 ringtest_0.x4._11_ 3.2005
R13585 ringtest_0.x4._11_ ringtest_0.x4._11_.n29 3.2005
R13586 ringtest_0.x4._11_.n17 ringtest_0.x4._11_.n13 2.49494
R13587 ringtest_0.x4._11_.n2 ringtest_0.x4._11_ 2.3045
R13588 ringtest_0.x4._11_.n12 ringtest_0.x4._11_ 1.97868
R13589 ringtest_0.x4._11_.n13 ringtest_0.x4._11_.n10 1.71582
R13590 ringtest_0.x4._11_.n27 ringtest_0.x4._11_.n23 1.38649
R13591 ringtest_0.x4._11_.n26 ringtest_0.x4._11_.n25 1.2805
R13592 ringtest_0.x4._11_.n20 ringtest_0.x4._11_.n17 1.24753
R13593 ui_in[0].n5 ui_in[0].t7 327.99
R13594 ui_in[0].n9 ui_in[0].t4 293.969
R13595 ui_in[0].n3 ui_in[0].t5 261.887
R13596 ui_in[0].n0 ui_in[0].t8 212.081
R13597 ui_in[0].n1 ui_in[0].t6 212.081
R13598 ui_in[0].n5 ui_in[0].t1 199.457
R13599 ui_in[0].n2 ui_in[0].n1 183.185
R13600 ui_in[0].n3 ui_in[0].t9 155.847
R13601 ui_in[0] ui_in[0].n9 154.065
R13602 ui_in[0].n4 ui_in[0].n3 153.506
R13603 ui_in[0].n6 ui_in[0].n5 152
R13604 ui_in[0].n0 ui_in[0].t3 139.78
R13605 ui_in[0].n1 ui_in[0].t0 139.78
R13606 ui_in[0].n9 ui_in[0].t2 138.338
R13607 ui_in[0].n1 ui_in[0].n0 61.346
R13608 ui_in[0].n13 ui_in[0] 38.2119
R13609 ui_in[0].n10 ui_in[0] 13.4199
R13610 ui_in[0].n11 ui_in[0].n8 11.7395
R13611 ui_in[0].n12 ui_in[0].n11 11.5949
R13612 ui_in[0].n8 ui_in[0].n4 10.4004
R13613 ui_in[0].n12 ui_in[0].n2 9.68118
R13614 ui_in[0].n6 ui_in[0] 9.6005
R13615 ui_in[0].n2 ui_in[0] 5.8885
R13616 ui_in[0].n10 ui_in[0] 5.57469
R13617 ui_in[0].n13 ui_in[0] 4.74482
R13618 ui_in[0].n8 ui_in[0].n7 4.6505
R13619 ui_in[0].n11 ui_in[0].n10 4.6505
R13620 ui_in[0].n7 ui_in[0].n6 2.98717
R13621 ui_in[0].n4 ui_in[0] 2.82403
R13622 ui_in[0].n7 ui_in[0] 1.9205
R13623 ui_in[0] ui_in[0].n12 0.559212
R13624 ui_in[0] ui_in[0].n13 0.02675
R13625 muxtest_0.R3R4.n5 muxtest_0.R3R4.t1 26.3998
R13626 muxtest_0.R3R4.n0 muxtest_0.R3R4.t9 26.3998
R13627 muxtest_0.R3R4.n5 muxtest_0.R3R4.t0 23.5483
R13628 muxtest_0.R3R4.n0 muxtest_0.R3R4.t8 23.5483
R13629 muxtest_0.R3R4.n6 muxtest_0.R3R4.t7 12.9758
R13630 muxtest_0.R3R4.n1 muxtest_0.R3R4.t4 12.9758
R13631 muxtest_0.R3R4.n6 muxtest_0.R3R4.t6 10.8618
R13632 muxtest_0.R3R4.n1 muxtest_0.R3R4.t5 10.8618
R13633 muxtest_0.R3R4.n4 muxtest_0.R3R4.t3 10.5285
R13634 muxtest_0.R3R4.n11 muxtest_0.R3R4.n10 7.08509
R13635 muxtest_0.R3R4.n7 muxtest_0.R3R4.n5 3.06895
R13636 muxtest_0.R3R4.n2 muxtest_0.R3R4.n0 3.06895
R13637 muxtest_0.R3R4.n7 muxtest_0.R3R4.n6 2.14822
R13638 muxtest_0.R3R4.n2 muxtest_0.R3R4.n1 2.14822
R13639 muxtest_0.R3R4.n8 muxtest_0.R3R4.n7 1.12636
R13640 muxtest_0.R3R4.n3 muxtest_0.R3R4.n2 1.12636
R13641 muxtest_0.R3R4.n4 muxtest_0.R3R4.t2 1.06523
R13642 muxtest_0.R3R4.n12 muxtest_0.R3R4 0.893
R13643 muxtest_0.R3R4.n9 muxtest_0.R3R4 0.670143
R13644 muxtest_0.R3R4.n12 muxtest_0.R3R4.n11 0.40675
R13645 muxtest_0.R3R4.n10 muxtest_0.R3R4.n9 0.223714
R13646 muxtest_0.R3R4.n11 muxtest_0.R3R4.n4 0.183423
R13647 muxtest_0.R3R4 muxtest_0.R3R4.n3 0.148615
R13648 muxtest_0.R3R4.n9 muxtest_0.R3R4.n8 0.132418
R13649 muxtest_0.R3R4.n12 muxtest_0.R3R4 0.08425
R13650 muxtest_0.R3R4.n8 muxtest_0.R3R4 0.0655
R13651 muxtest_0.R3R4.n3 muxtest_0.R3R4 0.0655
R13652 muxtest_0.R3R4 muxtest_0.R3R4.n12 0.04425
R13653 muxtest_0.R3R4.n10 muxtest_0.R3R4 0.00907843
R13654 ui_in[4].n26 ui_in[4].t3 327.99
R13655 ui_in[4].n10 ui_in[4].t0 327.99
R13656 ui_in[4].n19 ui_in[4].t1 293.969
R13657 ui_in[4].n3 ui_in[4].t19 293.969
R13658 ui_in[4].n22 ui_in[4].t14 256.07
R13659 ui_in[4].n6 ui_in[4].t12 256.07
R13660 ui_in[4].n16 ui_in[4].t9 212.081
R13661 ui_in[4].n17 ui_in[4].t15 212.081
R13662 ui_in[4].n0 ui_in[4].t6 212.081
R13663 ui_in[4].n1 ui_in[4].t4 212.081
R13664 ui_in[4].n26 ui_in[4].t8 199.457
R13665 ui_in[4].n10 ui_in[4].t5 199.457
R13666 ui_in[4].n18 ui_in[4].n17 182.929
R13667 ui_in[4].n2 ui_in[4].n1 182.929
R13668 ui_in[4] ui_in[4].n19 154.065
R13669 ui_in[4] ui_in[4].n3 154.065
R13670 ui_in[4].n27 ui_in[4].n26 152
R13671 ui_in[4].n23 ui_in[4].n22 152
R13672 ui_in[4].n11 ui_in[4].n10 152
R13673 ui_in[4].n7 ui_in[4].n6 152
R13674 ui_in[4].n22 ui_in[4].t11 150.03
R13675 ui_in[4].n6 ui_in[4].t7 150.03
R13676 ui_in[4].n16 ui_in[4].t18 139.78
R13677 ui_in[4].n17 ui_in[4].t2 139.78
R13678 ui_in[4].n0 ui_in[4].t16 139.78
R13679 ui_in[4].n1 ui_in[4].t10 139.78
R13680 ui_in[4].n19 ui_in[4].t17 138.338
R13681 ui_in[4].n3 ui_in[4].t13 138.338
R13682 ui_in[4].n17 ui_in[4].n16 61.346
R13683 ui_in[4].n1 ui_in[4].n0 61.346
R13684 ui_in[4].n31 ui_in[4] 31.335
R13685 ui_in[4].n21 ui_in[4] 17.455
R13686 ui_in[4].n5 ui_in[4] 17.455
R13687 ui_in[4].n30 ui_in[4].n29 14.6836
R13688 ui_in[4].n14 ui_in[4].n13 14.6836
R13689 ui_in[4].n29 ui_in[4].n28 14.6704
R13690 ui_in[4].n13 ui_in[4].n12 14.6704
R13691 ui_in[4].n20 ui_in[4] 13.8328
R13692 ui_in[4].n4 ui_in[4] 13.8328
R13693 ui_in[4].n31 ui_in[4] 12.499
R13694 ui_in[4].n30 ui_in[4].n18 10.6811
R13695 ui_in[4].n14 ui_in[4].n2 10.6811
R13696 ui_in[4].n23 ui_in[4].n21 10.4374
R13697 ui_in[4].n7 ui_in[4].n5 10.4374
R13698 ui_in[4].n25 ui_in[4].n24 8.15776
R13699 ui_in[4].n9 ui_in[4].n8 8.15776
R13700 ui_in[4].n28 ui_in[4] 6.61383
R13701 ui_in[4].n12 ui_in[4] 6.61383
R13702 ui_in[4].n18 ui_in[4] 6.1445
R13703 ui_in[4].n2 ui_in[4] 6.1445
R13704 ui_in[4].n20 ui_in[4] 5.16179
R13705 ui_in[4].n4 ui_in[4] 5.16179
R13706 ui_in[4].n27 ui_in[4] 4.90717
R13707 ui_in[4].n11 ui_in[4] 4.90717
R13708 ui_in[4].n25 ui_in[4].n20 4.65206
R13709 ui_in[4].n9 ui_in[4].n4 4.65206
R13710 ui_in[4].n24 ui_in[4] 3.93896
R13711 ui_in[4].n8 ui_in[4] 3.93896
R13712 ui_in[4].n28 ui_in[4].n27 2.98717
R13713 ui_in[4].n12 ui_in[4].n11 2.98717
R13714 ui_in[4].n21 ui_in[4] 2.16665
R13715 ui_in[4].n5 ui_in[4] 2.16665
R13716 ui_in[4].n24 ui_in[4].n23 1.57588
R13717 ui_in[4].n8 ui_in[4].n7 1.57588
R13718 ui_in[4].n29 ui_in[4].n25 0.79438
R13719 ui_in[4].n13 ui_in[4].n9 0.79438
R13720 ui_in[4] ui_in[4].n15 0.287559
R13721 ui_in[4] ui_in[4].n31 0.28675
R13722 ui_in[4] ui_in[4].n30 0.248606
R13723 ui_in[4] ui_in[4].n14 0.248606
R13724 ui_in[4].n15 ui_in[4] 0.11603
R13725 ui_in[4].n15 ui_in[4] 0.0460882
R13726 muxtest_0.R1R2.n0 muxtest_0.R1R2.t3 26.3998
R13727 muxtest_0.R1R2.n0 muxtest_0.R1R2.t2 23.5483
R13728 muxtest_0.R1R2.n1 muxtest_0.R1R2.t5 12.9758
R13729 muxtest_0.R1R2.n1 muxtest_0.R1R2.t4 10.8618
R13730 muxtest_0.R1R2.n4 muxtest_0.R1R2.t1 10.5285
R13731 muxtest_0.R1R2.n2 muxtest_0.R1R2.n0 3.06895
R13732 muxtest_0.R1R2.n2 muxtest_0.R1R2.n1 2.14822
R13733 muxtest_0.R1R2.n3 muxtest_0.R1R2.n2 1.12636
R13734 muxtest_0.R1R2.n4 muxtest_0.R1R2.t0 1.06052
R13735 muxtest_0.R1R2.n5 muxtest_0.R1R2 0.96675
R13736 muxtest_0.R1R2.n5 muxtest_0.R1R2.n4 0.494965
R13737 muxtest_0.R1R2 muxtest_0.R1R2.n3 0.132418
R13738 muxtest_0.R1R2.n5 muxtest_0.R1R2 0.06925
R13739 muxtest_0.R1R2.n3 muxtest_0.R1R2 0.0655
R13740 muxtest_0.R1R2 muxtest_0.R1R2.n5 0.04425
R13741 a_19289_13081.n0 a_19289_13081.t12 1681.78
R13742 a_19289_13081.n2 a_19289_13081.t7 1681.21
R13743 a_19289_13081.n1 a_19289_13081.t13 1681.21
R13744 a_19289_13081.n0 a_19289_13081.t2 1681.21
R13745 a_19289_13081.n13 a_19289_13081.t14 1681.21
R13746 a_19289_13081.n11 a_19289_13081.t10 1681.21
R13747 a_19289_13081.n9 a_19289_13081.t17 1681.21
R13748 a_19289_13081.n7 a_19289_13081.t9 1681.21
R13749 a_19289_13081.n3 a_19289_13081.t4 703.317
R13750 a_19289_13081.n7 a_19289_13081.t6 702.768
R13751 a_19289_13081.n5 a_19289_13081.t11 702.747
R13752 a_19289_13081.n4 a_19289_13081.t5 702.747
R13753 a_19289_13081.n3 a_19289_13081.t15 702.747
R13754 a_19289_13081.n12 a_19289_13081.t3 702.747
R13755 a_19289_13081.n10 a_19289_13081.t8 702.747
R13756 a_19289_13081.n8 a_19289_13081.t16 702.747
R13757 a_19289_13081.n6 a_19289_13081.t0 30.088
R13758 a_19289_13081.t1 a_19289_13081.n15 26.0464
R13759 a_19289_13081.n15 a_19289_13081.n2 20.0759
R13760 a_19289_13081.n6 a_19289_13081.n5 0.875353
R13761 a_19289_13081.n1 a_19289_13081.n0 0.576859
R13762 a_19289_13081.n2 a_19289_13081.n1 0.576859
R13763 a_19289_13081.n4 a_19289_13081.n3 0.570292
R13764 a_19289_13081.n5 a_19289_13081.n4 0.570292
R13765 a_19289_13081.n15 a_19289_13081.n14 0.267403
R13766 a_19289_13081.n14 a_19289_13081.n6 0.10833
R13767 a_19289_13081.n14 a_19289_13081.n13 0.0744583
R13768 a_19289_13081.n8 a_19289_13081.n7 0.0205
R13769 a_19289_13081.n9 a_19289_13081.n8 0.0205
R13770 a_19289_13081.n10 a_19289_13081.n9 0.0205
R13771 a_19289_13081.n11 a_19289_13081.n10 0.0205
R13772 a_19289_13081.n12 a_19289_13081.n11 0.0205
R13773 a_19289_13081.n13 a_19289_13081.n12 0.0205
R13774 ringtest_0.drv_out.n7 ringtest_0.drv_out.t21 184.768
R13775 ringtest_0.drv_out.n6 ringtest_0.drv_out.t20 184.768
R13776 ringtest_0.drv_out.n5 ringtest_0.drv_out.t23 184.768
R13777 ringtest_0.drv_out.n4 ringtest_0.drv_out.t22 184.768
R13778 ringtest_0.drv_out.n8 ringtest_0.drv_out.n7 171.375
R13779 ringtest_0.drv_out.n7 ringtest_0.drv_out.t25 146.208
R13780 ringtest_0.drv_out.n6 ringtest_0.drv_out.t24 146.208
R13781 ringtest_0.drv_out.n5 ringtest_0.drv_out.t27 146.208
R13782 ringtest_0.drv_out.n4 ringtest_0.drv_out.t26 146.208
R13783 ringtest_0.drv_out.n7 ringtest_0.drv_out.n6 40.6397
R13784 ringtest_0.drv_out.n6 ringtest_0.drv_out.n5 40.6397
R13785 ringtest_0.drv_out.n5 ringtest_0.drv_out.n4 40.6397
R13786 ringtest_0.drv_out.n0 ringtest_0.drv_out.t0 26.3998
R13787 ringtest_0.drv_out.n21 ringtest_0.drv_out.n20 26.0838
R13788 ringtest_0.drv_out.n21 ringtest_0.drv_out.n17 26.0838
R13789 ringtest_0.drv_out.n21 ringtest_0.drv_out.n19 26.0838
R13790 ringtest_0.drv_out.n21 ringtest_0.drv_out.n18 26.0838
R13791 ringtest_0.drv_out.n16 ringtest_0.drv_out.n12 24.902
R13792 ringtest_0.drv_out.n16 ringtest_0.drv_out.n14 24.902
R13793 ringtest_0.drv_out.n16 ringtest_0.drv_out.n13 24.902
R13794 ringtest_0.drv_out.n16 ringtest_0.drv_out.n15 24.902
R13795 ringtest_0.drv_out.n0 ringtest_0.drv_out.t17 23.5483
R13796 ringtest_0.drv_out.n1 ringtest_0.drv_out.t18 12.9758
R13797 ringtest_0.drv_out ringtest_0.drv_out.n8 12.3171
R13798 ringtest_0.drv_out.n1 ringtest_0.drv_out.t19 10.8618
R13799 ringtest_0.drv_out.n20 ringtest_0.drv_out.t16 6.6005
R13800 ringtest_0.drv_out.n20 ringtest_0.drv_out.t11 6.6005
R13801 ringtest_0.drv_out.n17 ringtest_0.drv_out.t12 6.6005
R13802 ringtest_0.drv_out.n17 ringtest_0.drv_out.t14 6.6005
R13803 ringtest_0.drv_out.n19 ringtest_0.drv_out.t9 6.6005
R13804 ringtest_0.drv_out.n19 ringtest_0.drv_out.t10 6.6005
R13805 ringtest_0.drv_out.n18 ringtest_0.drv_out.t13 6.6005
R13806 ringtest_0.drv_out.n18 ringtest_0.drv_out.t15 6.6005
R13807 ringtest_0.drv_out.n11 ringtest_0.drv_out 5.69273
R13808 ringtest_0.drv_out.n12 ringtest_0.drv_out.t7 3.61217
R13809 ringtest_0.drv_out.n12 ringtest_0.drv_out.t2 3.61217
R13810 ringtest_0.drv_out.n14 ringtest_0.drv_out.t3 3.61217
R13811 ringtest_0.drv_out.n14 ringtest_0.drv_out.t5 3.61217
R13812 ringtest_0.drv_out.n13 ringtest_0.drv_out.t4 3.61217
R13813 ringtest_0.drv_out.n13 ringtest_0.drv_out.t6 3.61217
R13814 ringtest_0.drv_out.n15 ringtest_0.drv_out.t8 3.61217
R13815 ringtest_0.drv_out.n15 ringtest_0.drv_out.t1 3.61217
R13816 ringtest_0.drv_out.n2 ringtest_0.drv_out.n0 3.06895
R13817 ringtest_0.drv_out.n11 ringtest_0.drv_out 2.87193
R13818 ringtest_0.drv_out.n8 ringtest_0.drv_out 2.23542
R13819 ringtest_0.drv_out.n2 ringtest_0.drv_out.n1 2.14822
R13820 ringtest_0.drv_out.n10 ringtest_0.drv_out 1.7806
R13821 ringtest_0.drv_out ringtest_0.drv_out.n10 1.54574
R13822 ringtest_0.drv_out.n9 ringtest_0.drv_out 1.25273
R13823 ringtest_0.drv_out.n3 ringtest_0.drv_out.n2 1.12636
R13824 ringtest_0.drv_out ringtest_0.drv_out.n22 0.461707
R13825 ringtest_0.drv_out.n9 ringtest_0.drv_out 0.316378
R13826 ringtest_0.drv_out ringtest_0.drv_out.n11 0.188041
R13827 ringtest_0.drv_out ringtest_0.drv_out.n3 0.138152
R13828 ringtest_0.drv_out.n22 ringtest_0.drv_out.n16 0.0921193
R13829 ringtest_0.drv_out.n22 ringtest_0.drv_out.n21 0.069392
R13830 ringtest_0.drv_out.n3 ringtest_0.drv_out 0.0655
R13831 ringtest_0.drv_out.n10 ringtest_0.drv_out.n9 0.0596216
R13832 ringtest_0.x4.net3.t3 ringtest_0.x4.net3.t4 395.01
R13833 ringtest_0.x4.net3 ringtest_0.x4.net3.t3 320.745
R13834 ringtest_0.x4.net3.n3 ringtest_0.x4.net3.t6 260.322
R13835 ringtest_0.x4.net3.n0 ringtest_0.x4.net3.t7 229.369
R13836 ringtest_0.x4.net3.n7 ringtest_0.x4.net3.t0 222.68
R13837 ringtest_0.x4.net3.n3 ringtest_0.x4.net3.t5 175.169
R13838 ringtest_0.x4.net3.n0 ringtest_0.x4.net3.t2 157.07
R13839 ringtest_0.x4.net3.n4 ringtest_0.x4.net3.n3 152
R13840 ringtest_0.x4.net3.n1 ringtest_0.x4.net3.n0 152
R13841 ringtest_0.x4.net3.n8 ringtest_0.x4.net3.t1 132.322
R13842 ringtest_0.x4.net3.n8 ringtest_0.x4.net3.n7 95.0273
R13843 ringtest_0.x4.net3.n5 ringtest_0.x4.net3 25.2581
R13844 ringtest_0.x4.net3.n5 ringtest_0.x4.net3 20.1696
R13845 ringtest_0.x4.net3.n7 ringtest_0.x4.net3.n6 12.7813
R13846 ringtest_0.x4.net3.n1 ringtest_0.x4.net3 12.0005
R13847 ringtest_0.x4.net3 ringtest_0.x4.net3.n4 11.2497
R13848 ringtest_0.x4.net3.n6 ringtest_0.x4.net3.n2 9.79203
R13849 ringtest_0.x4.net3.n6 ringtest_0.x4.net3.n5 5.9277
R13850 ringtest_0.x4.net3.n2 ringtest_0.x4.net3 4.53383
R13851 ringtest_0.x4.net3 ringtest_0.x4.net3.n8 2.70465
R13852 ringtest_0.x4.net3.n2 ringtest_0.x4.net3.n1 1.6005
R13853 ringtest_0.x4.net3.n4 ringtest_0.x4.net3 1.55726
R13854 ui_in[2].n2 ui_in[2].t0 450.938
R13855 ui_in[2].n2 ui_in[2].t6 445.666
R13856 ui_in[2].n0 ui_in[2].t7 377.486
R13857 ui_in[2].n0 ui_in[2].t1 374.202
R13858 ui_in[2].n5 ui_in[2].t2 212.081
R13859 ui_in[2].n6 ui_in[2].t3 212.081
R13860 ui_in[2].n7 ui_in[2].n6 183.441
R13861 ui_in[2].n5 ui_in[2].t4 139.78
R13862 ui_in[2].n6 ui_in[2].t5 139.78
R13863 ui_in[2].n6 ui_in[2].n5 61.346
R13864 ui_in[2].n4 ui_in[2].n1 12.4088
R13865 ui_in[2] ui_in[2].n7 11.4331
R13866 ui_in[2].n4 ui_in[2].n3 9.10647
R13867 ui_in[2].n8 ui_in[2].n4 8.98648
R13868 ui_in[2].n7 ui_in[2] 5.6325
R13869 ui_in[2].n8 ui_in[2] 5.02323
R13870 ui_in[2].n3 ui_in[2].n2 3.1748
R13871 ui_in[2] ui_in[2].n0 2.04102
R13872 ui_in[2] ui_in[2].n8 0.888758
R13873 ui_in[2].n1 ui_in[2] 0.412375
R13874 ui_in[2].n3 ui_in[2] 0.063625
R13875 ui_in[2].n1 ui_in[2] 0.061125
R13876 ringtest_0.x3.x2.GP4.n2 ringtest_0.x3.x2.GP4.t5 450.938
R13877 ringtest_0.x3.x2.GP4.n2 ringtest_0.x3.x2.GP4.t4 445.666
R13878 ringtest_0.x3.x2.GP4.n5 ringtest_0.x3.x2.GP4.n4 208.965
R13879 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n0 96.8352
R13880 ringtest_0.x3.x2.GP4.n4 ringtest_0.x3.x2.GP4.t1 26.5955
R13881 ringtest_0.x3.x2.GP4.n4 ringtest_0.x3.x2.GP4.t0 26.5955
R13882 ringtest_0.x3.x2.GP4.n0 ringtest_0.x3.x2.GP4.t3 24.9236
R13883 ringtest_0.x3.x2.GP4.n0 ringtest_0.x3.x2.GP4.t2 24.9236
R13884 ringtest_0.x3.x1.gpo3 ringtest_0.x3.x2.x4.GP 16.5032
R13885 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n3 10.2405
R13886 ringtest_0.x3.x2.GP4.n3 ringtest_0.x3.x1.gpo3 7.76481
R13887 ringtest_0.x3.x2.GP4.n1 ringtest_0.x3.x1.x14.Y 6.1445
R13888 ringtest_0.x3.x2.GP4.n1 ringtest_0.x3.x1.x14.Y 4.65505
R13889 ringtest_0.x3.x2.x4.GP ringtest_0.x3.x2.GP4.n2 2.95993
R13890 ringtest_0.x3.x2.GP4.n5 ringtest_0.x3.x1.x14.Y 2.0485
R13891 ringtest_0.x3.x1.x14.Y ringtest_0.x3.x2.GP4.n5 1.55202
R13892 ringtest_0.x3.x2.GP4.n3 ringtest_0.x3.x2.GP4.n1 1.0245
R13893 ringtest_0.counter7.n0 ringtest_0.counter7.t2 368.521
R13894 ringtest_0.counter7.n1 ringtest_0.counter7.t3 216.155
R13895 ringtest_0.counter7.n1 ringtest_0.counter7 78.8791
R13896 ringtest_0.counter7.n4 ringtest_0.counter7.t4 26.3998
R13897 ringtest_0.counter7.n4 ringtest_0.counter7.t5 23.5483
R13898 ringtest_0.counter7.n3 ringtest_0.counter7.n2 18.2765
R13899 ringtest_0.counter7.n5 ringtest_0.counter7.t1 12.9758
R13900 ringtest_0.counter7.n5 ringtest_0.counter7.t0 10.8618
R13901 ringtest_0.counter7 ringtest_0.counter7.n0 10.5563
R13902 ringtest_0.counter7.n0 ringtest_0.counter7 5.48477
R13903 ringtest_0.counter7.n2 ringtest_0.counter7 4.18512
R13904 ringtest_0.counter7.n6 ringtest_0.counter7.n4 3.06895
R13905 ringtest_0.counter7.n6 ringtest_0.counter7.n5 2.14822
R13906 ringtest_0.counter7 ringtest_0.counter7.n6 1.27287
R13907 ringtest_0.counter7.n3 ringtest_0.counter7 1.27059
R13908 ringtest_0.counter7.n2 ringtest_0.counter7.n1 0.985115
R13909 ringtest_0.counter7 ringtest_0.counter7.n3 0.647091
R13910 ua[1].n6 ua[1].t11 23.6581
R13911 ua[1].n12 ua[1].t6 23.6581
R13912 ua[1].n19 ua[1].t7 23.6581
R13913 ua[1].n1 ua[1].t5 23.6581
R13914 ua[1].n5 ua[1].t3 23.3739
R13915 ua[1].n11 ua[1].t0 23.3739
R13916 ua[1].n18 ua[1].t8 23.3739
R13917 ua[1].n0 ua[1].t4 23.3739
R13918 ua[1].n25 ua[1] 15.3856
R13919 ua[1].n6 ua[1].t12 10.7528
R13920 ua[1].n12 ua[1].t10 10.7528
R13921 ua[1].n19 ua[1].t14 10.7528
R13922 ua[1].n1 ua[1].t1 10.7528
R13923 ua[1].n8 ua[1].t13 10.6417
R13924 ua[1].n14 ua[1].t9 10.6417
R13925 ua[1].n21 ua[1].t15 10.6417
R13926 ua[1].n3 ua[1].t2 10.6417
R13927 ua[1].n7 ua[1].n6 1.30064
R13928 ua[1].n13 ua[1].n12 1.30064
R13929 ua[1].n20 ua[1].n19 1.30064
R13930 ua[1].n2 ua[1].n1 1.30064
R13931 ua[1] ua[1].n4 0.983856
R13932 ua[1].n23 ua[1].n22 0.946356
R13933 ua[1].n16 ua[1].n15 0.927606
R13934 ua[1].n10 ua[1].n9 0.925106
R13935 ua[1].n17 ua[1] 0.748625
R13936 ua[1].n7 ua[1].n5 0.726502
R13937 ua[1].n13 ua[1].n11 0.726502
R13938 ua[1].n20 ua[1].n18 0.726502
R13939 ua[1].n2 ua[1].n0 0.726502
R13940 ua[1].n24 ua[1].n17 0.54425
R13941 ua[1].n25 ua[1] 0.532375
R13942 ua[1].n8 ua[1].n7 0.512491
R13943 ua[1].n14 ua[1].n13 0.512491
R13944 ua[1].n21 ua[1].n20 0.512491
R13945 ua[1].n3 ua[1].n2 0.512491
R13946 ua[1].n9 ua[1].n8 0.359663
R13947 ua[1].n15 ua[1].n14 0.359663
R13948 ua[1].n22 ua[1].n21 0.359663
R13949 ua[1].n4 ua[1].n3 0.359663
R13950 ua[1].n9 ua[1].n5 0.216071
R13951 ua[1].n15 ua[1].n11 0.216071
R13952 ua[1].n22 ua[1].n18 0.216071
R13953 ua[1].n4 ua[1].n0 0.216071
R13954 ua[1].n17 ua[1] 0.20175
R13955 ua[1].n24 ua[1] 0.17925
R13956 ua[1] ua[1].n25 0.178
R13957 ua[1].n24 ua[1] 0.063
R13958 ua[1].n10 ua[1] 0.05925
R13959 ua[1].n16 ua[1] 0.05675
R13960 ua[1] ua[1].n16 0.0561931
R13961 ua[1] ua[1].n10 0.0561872
R13962 ua[1].n23 ua[1] 0.038
R13963 ua[1] ua[1].n23 0.0376287
R13964 ua[1] ua[1].n24 0.004875
R13965 ringtest_0.x4.clknet_1_0__leaf_clk.n25 ringtest_0.x4.clknet_1_0__leaf_clk.n23 333.392
R13966 ringtest_0.x4.clknet_1_0__leaf_clk.n25 ringtest_0.x4.clknet_1_0__leaf_clk.n24 301.392
R13967 ringtest_0.x4.clknet_1_0__leaf_clk.n27 ringtest_0.x4.clknet_1_0__leaf_clk.n26 301.392
R13968 ringtest_0.x4.clknet_1_0__leaf_clk.n29 ringtest_0.x4.clknet_1_0__leaf_clk.n28 301.392
R13969 ringtest_0.x4.clknet_1_0__leaf_clk.n22 ringtest_0.x4.clknet_1_0__leaf_clk.n4 301.392
R13970 ringtest_0.x4.clknet_1_0__leaf_clk.n31 ringtest_0.x4.clknet_1_0__leaf_clk.n30 301.392
R13971 ringtest_0.x4.clknet_1_0__leaf_clk.n21 ringtest_0.x4.clknet_1_0__leaf_clk.n5 297.863
R13972 ringtest_0.x4.clknet_1_0__leaf_clk.n2 ringtest_0.x4.clknet_1_0__leaf_clk.t32 294.557
R13973 ringtest_0.x4.clknet_1_0__leaf_clk.n0 ringtest_0.x4.clknet_1_0__leaf_clk.t38 294.557
R13974 ringtest_0.x4.clknet_1_0__leaf_clk.n41 ringtest_0.x4.clknet_1_0__leaf_clk.t35 294.557
R13975 ringtest_0.x4.clknet_1_0__leaf_clk.n38 ringtest_0.x4.clknet_1_0__leaf_clk.t33 294.557
R13976 ringtest_0.x4.clknet_1_0__leaf_clk.n36 ringtest_0.x4.clknet_1_0__leaf_clk.t36 294.557
R13977 ringtest_0.x4.clknet_1_0__leaf_clk.n34 ringtest_0.x4.clknet_1_0__leaf_clk.n33 287.303
R13978 ringtest_0.x4.clknet_1_0__leaf_clk.n8 ringtest_0.x4.clknet_1_0__leaf_clk.n6 248.638
R13979 ringtest_0.x4.clknet_1_0__leaf_clk.n2 ringtest_0.x4.clknet_1_0__leaf_clk.t37 211.01
R13980 ringtest_0.x4.clknet_1_0__leaf_clk.n0 ringtest_0.x4.clknet_1_0__leaf_clk.t41 211.01
R13981 ringtest_0.x4.clknet_1_0__leaf_clk.n41 ringtest_0.x4.clknet_1_0__leaf_clk.t34 211.01
R13982 ringtest_0.x4.clknet_1_0__leaf_clk.n38 ringtest_0.x4.clknet_1_0__leaf_clk.t40 211.01
R13983 ringtest_0.x4.clknet_1_0__leaf_clk.n36 ringtest_0.x4.clknet_1_0__leaf_clk.t39 211.01
R13984 ringtest_0.x4.clknet_1_0__leaf_clk.n8 ringtest_0.x4.clknet_1_0__leaf_clk.n7 203.463
R13985 ringtest_0.x4.clknet_1_0__leaf_clk.n10 ringtest_0.x4.clknet_1_0__leaf_clk.n9 203.463
R13986 ringtest_0.x4.clknet_1_0__leaf_clk.n14 ringtest_0.x4.clknet_1_0__leaf_clk.n13 203.463
R13987 ringtest_0.x4.clknet_1_0__leaf_clk.n16 ringtest_0.x4.clknet_1_0__leaf_clk.n15 203.463
R13988 ringtest_0.x4.clknet_1_0__leaf_clk.n18 ringtest_0.x4.clknet_1_0__leaf_clk.n17 203.463
R13989 ringtest_0.x4.clknet_1_0__leaf_clk.n12 ringtest_0.x4.clknet_1_0__leaf_clk.n11 202.456
R13990 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n19 199.607
R13991 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n2 156.207
R13992 ringtest_0.x4.clknet_1_0__leaf_clk.n37 ringtest_0.x4.clknet_1_0__leaf_clk.n36 153.097
R13993 ringtest_0.x4.clknet_1_0__leaf_clk.n39 ringtest_0.x4.clknet_1_0__leaf_clk.n38 152.296
R13994 ringtest_0.x4.clknet_1_0__leaf_clk.n1 ringtest_0.x4.clknet_1_0__leaf_clk.n0 152
R13995 ringtest_0.x4.clknet_1_0__leaf_clk.n42 ringtest_0.x4.clknet_1_0__leaf_clk.n41 152
R13996 ringtest_0.x4.clknet_1_0__leaf_clk.n10 ringtest_0.x4.clknet_1_0__leaf_clk.n8 45.177
R13997 ringtest_0.x4.clknet_1_0__leaf_clk.n16 ringtest_0.x4.clknet_1_0__leaf_clk.n14 45.177
R13998 ringtest_0.x4.clknet_1_0__leaf_clk.n18 ringtest_0.x4.clknet_1_0__leaf_clk.n16 45.177
R13999 ringtest_0.x4.clknet_1_0__leaf_clk.n12 ringtest_0.x4.clknet_1_0__leaf_clk.n10 44.0476
R14000 ringtest_0.x4.clknet_1_0__leaf_clk.n14 ringtest_0.x4.clknet_1_0__leaf_clk.n12 44.0476
R14001 ringtest_0.x4.clknet_1_0__leaf_clk.n6 ringtest_0.x4.clknet_1_0__leaf_clk.t24 40.0005
R14002 ringtest_0.x4.clknet_1_0__leaf_clk.n6 ringtest_0.x4.clknet_1_0__leaf_clk.t27 40.0005
R14003 ringtest_0.x4.clknet_1_0__leaf_clk.n7 ringtest_0.x4.clknet_1_0__leaf_clk.t29 40.0005
R14004 ringtest_0.x4.clknet_1_0__leaf_clk.n7 ringtest_0.x4.clknet_1_0__leaf_clk.t31 40.0005
R14005 ringtest_0.x4.clknet_1_0__leaf_clk.n9 ringtest_0.x4.clknet_1_0__leaf_clk.t26 40.0005
R14006 ringtest_0.x4.clknet_1_0__leaf_clk.n9 ringtest_0.x4.clknet_1_0__leaf_clk.t28 40.0005
R14007 ringtest_0.x4.clknet_1_0__leaf_clk.n11 ringtest_0.x4.clknet_1_0__leaf_clk.t30 40.0005
R14008 ringtest_0.x4.clknet_1_0__leaf_clk.n11 ringtest_0.x4.clknet_1_0__leaf_clk.t25 40.0005
R14009 ringtest_0.x4.clknet_1_0__leaf_clk.n13 ringtest_0.x4.clknet_1_0__leaf_clk.t17 40.0005
R14010 ringtest_0.x4.clknet_1_0__leaf_clk.n13 ringtest_0.x4.clknet_1_0__leaf_clk.t20 40.0005
R14011 ringtest_0.x4.clknet_1_0__leaf_clk.n15 ringtest_0.x4.clknet_1_0__leaf_clk.t22 40.0005
R14012 ringtest_0.x4.clknet_1_0__leaf_clk.n15 ringtest_0.x4.clknet_1_0__leaf_clk.t23 40.0005
R14013 ringtest_0.x4.clknet_1_0__leaf_clk.n17 ringtest_0.x4.clknet_1_0__leaf_clk.t19 40.0005
R14014 ringtest_0.x4.clknet_1_0__leaf_clk.n17 ringtest_0.x4.clknet_1_0__leaf_clk.t21 40.0005
R14015 ringtest_0.x4.clknet_1_0__leaf_clk.n19 ringtest_0.x4.clknet_1_0__leaf_clk.t16 40.0005
R14016 ringtest_0.x4.clknet_1_0__leaf_clk.n19 ringtest_0.x4.clknet_1_0__leaf_clk.t18 40.0005
R14017 ringtest_0.x4.clknet_1_0__leaf_clk.n27 ringtest_0.x4.clknet_1_0__leaf_clk.n25 32.0005
R14018 ringtest_0.x4.clknet_1_0__leaf_clk.n29 ringtest_0.x4.clknet_1_0__leaf_clk.n27 32.0005
R14019 ringtest_0.x4.clknet_1_0__leaf_clk.n32 ringtest_0.x4.clknet_1_0__leaf_clk.n22 32.0005
R14020 ringtest_0.x4.clknet_1_0__leaf_clk.n32 ringtest_0.x4.clknet_1_0__leaf_clk.n31 32.0005
R14021 ringtest_0.x4.clknet_1_0__leaf_clk.n31 ringtest_0.x4.clknet_1_0__leaf_clk.n29 31.2005
R14022 ringtest_0.x4.clknet_1_0__leaf_clk.n35 ringtest_0.x4.clknet_1_0__leaf_clk.n34 28.6283
R14023 ringtest_0.x4.clknet_1_0__leaf_clk.n3 ringtest_0.x4.clknet_1_0__leaf_clk 28.0697
R14024 ringtest_0.x4.clknet_1_0__leaf_clk.n23 ringtest_0.x4.clknet_1_0__leaf_clk.t3 27.5805
R14025 ringtest_0.x4.clknet_1_0__leaf_clk.n23 ringtest_0.x4.clknet_1_0__leaf_clk.t6 27.5805
R14026 ringtest_0.x4.clknet_1_0__leaf_clk.n24 ringtest_0.x4.clknet_1_0__leaf_clk.t8 27.5805
R14027 ringtest_0.x4.clknet_1_0__leaf_clk.n24 ringtest_0.x4.clknet_1_0__leaf_clk.t10 27.5805
R14028 ringtest_0.x4.clknet_1_0__leaf_clk.n26 ringtest_0.x4.clknet_1_0__leaf_clk.t5 27.5805
R14029 ringtest_0.x4.clknet_1_0__leaf_clk.n26 ringtest_0.x4.clknet_1_0__leaf_clk.t7 27.5805
R14030 ringtest_0.x4.clknet_1_0__leaf_clk.n28 ringtest_0.x4.clknet_1_0__leaf_clk.t9 27.5805
R14031 ringtest_0.x4.clknet_1_0__leaf_clk.n28 ringtest_0.x4.clknet_1_0__leaf_clk.t4 27.5805
R14032 ringtest_0.x4.clknet_1_0__leaf_clk.n4 ringtest_0.x4.clknet_1_0__leaf_clk.t14 27.5805
R14033 ringtest_0.x4.clknet_1_0__leaf_clk.n4 ringtest_0.x4.clknet_1_0__leaf_clk.t0 27.5805
R14034 ringtest_0.x4.clknet_1_0__leaf_clk.n5 ringtest_0.x4.clknet_1_0__leaf_clk.t11 27.5805
R14035 ringtest_0.x4.clknet_1_0__leaf_clk.n5 ringtest_0.x4.clknet_1_0__leaf_clk.t13 27.5805
R14036 ringtest_0.x4.clknet_1_0__leaf_clk.n33 ringtest_0.x4.clknet_1_0__leaf_clk.t1 27.5805
R14037 ringtest_0.x4.clknet_1_0__leaf_clk.n33 ringtest_0.x4.clknet_1_0__leaf_clk.t2 27.5805
R14038 ringtest_0.x4.clknet_1_0__leaf_clk.n30 ringtest_0.x4.clknet_1_0__leaf_clk.t12 27.5805
R14039 ringtest_0.x4.clknet_1_0__leaf_clk.n30 ringtest_0.x4.clknet_1_0__leaf_clk.t15 27.5805
R14040 ringtest_0.x4.clknet_1_0__leaf_clk.n43 ringtest_0.x4.clknet_1_0__leaf_clk.n42 27.3319
R14041 ringtest_0.x4.clknet_1_0__leaf_clk.n40 ringtest_0.x4.clknet_1_0__leaf_clk.n39 21.4985
R14042 ringtest_0.x4.clknet_1_0__leaf_clk.n3 ringtest_0.x4.clknet_1_0__leaf_clk.n1 21.401
R14043 ringtest_0.x4.clknet_1_0__leaf_clk.n34 ringtest_0.x4.clknet_1_0__leaf_clk.n32 14.0898
R14044 ringtest_0.x4.clknet_1_0__leaf_clk.n20 ringtest_0.x4.clknet_1_0__leaf_clk.n18 13.177
R14045 ringtest_0.x4.clknet_1_0__leaf_clk.n40 ringtest_0.x4.clknet_1_0__leaf_clk.n37 11.0654
R14046 ringtest_0.x4.clknet_1_0__leaf_clk.n22 ringtest_0.x4.clknet_1_0__leaf_clk.n21 10.4484
R14047 ringtest_0.x4.clknet_1_0__leaf_clk.n43 ringtest_0.x4.clknet_1_0__leaf_clk.n40 7.18319
R14048 ringtest_0.x4.clknet_1_0__leaf_clk.n35 ringtest_0.x4.clknet_1_0__leaf_clk.n3 5.63649
R14049 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n20 3.13183
R14050 ringtest_0.x4.clknet_1_0__leaf_clk.n37 ringtest_0.x4.clknet_1_0__leaf_clk 3.10907
R14051 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n43 2.66671
R14052 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_1_0__leaf_clk.n35 2.66671
R14053 ringtest_0.x4.clknet_1_0__leaf_clk.n42 ringtest_0.x4.clknet_1_0__leaf_clk 2.01193
R14054 ringtest_0.x4.clknet_1_0__leaf_clk.n21 ringtest_0.x4.clknet_1_0__leaf_clk 1.75844
R14055 ringtest_0.x4.clknet_1_0__leaf_clk.n39 ringtest_0.x4.clknet_1_0__leaf_clk 1.67435
R14056 ringtest_0.x4.clknet_1_0__leaf_clk.n1 ringtest_0.x4.clknet_1_0__leaf_clk 1.37896
R14057 ringtest_0.x4.clknet_1_0__leaf_clk.n20 ringtest_0.x4.clknet_1_0__leaf_clk 0.604792
R14058 ringtest_0.counter3.n0 ringtest_0.counter3.t0 368.521
R14059 ringtest_0.counter3.n1 ringtest_0.counter3.t1 216.155
R14060 ringtest_0.counter3.n1 ringtest_0.counter3 78.8791
R14061 ringtest_0.counter3.n4 ringtest_0.counter3.t3 26.3998
R14062 ringtest_0.counter3.n4 ringtest_0.counter3.t2 23.5483
R14063 ringtest_0.counter3.n3 ringtest_0.counter3.n2 17.5689
R14064 ringtest_0.counter3.n5 ringtest_0.counter3.t5 12.9693
R14065 ringtest_0.counter3.n5 ringtest_0.counter3.t4 10.8444
R14066 ringtest_0.counter3 ringtest_0.counter3.n0 10.5563
R14067 ringtest_0.counter3.n0 ringtest_0.counter3 5.48477
R14068 ringtest_0.counter3.n2 ringtest_0.counter3 4.18512
R14069 ringtest_0.counter3.n6 ringtest_0.counter3.n4 3.06895
R14070 ringtest_0.counter3.n6 ringtest_0.counter3.n5 2.14822
R14071 ringtest_0.counter3.n3 ringtest_0.counter3 1.28175
R14072 ringtest_0.counter3 ringtest_0.counter3.n6 1.25828
R14073 ringtest_0.counter3.n2 ringtest_0.counter3.n1 0.985115
R14074 ringtest_0.counter3 ringtest_0.counter3.n3 0.688
R14075 muxtest_0.x1.x3.GP2.n3 muxtest_0.x1.x3.GP2.t4 450.938
R14076 muxtest_0.x1.x3.GP2.n2 muxtest_0.x1.x3.GP2.t7 450.938
R14077 muxtest_0.x1.x3.GP2.n3 muxtest_0.x1.x3.GP2.t5 445.666
R14078 muxtest_0.x1.x3.GP2.n2 muxtest_0.x1.x3.GP2.t6 445.666
R14079 muxtest_0.x1.x3.GP2.n6 muxtest_0.x1.x3.GP2.n5 195.958
R14080 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n0 96.8352
R14081 muxtest_0.x1.x3.GP2.n5 muxtest_0.x1.x3.GP2.t0 26.5955
R14082 muxtest_0.x1.x3.GP2.n5 muxtest_0.x1.x3.GP2.t1 26.5955
R14083 muxtest_0.x1.x3.GP2.n0 muxtest_0.x1.x3.GP2.t2 24.9236
R14084 muxtest_0.x1.x3.GP2.n0 muxtest_0.x1.x3.GP2.t3 24.9236
R14085 muxtest_0.x1.x3.GP2.n4 muxtest_0.x1.x3.GP2 14.8953
R14086 muxtest_0.x1.x3.GP2.n7 muxtest_0.x1.x3.GP2.n6 13.0077
R14087 muxtest_0.x1.x3.GP2.n6 muxtest_0.x1.x3.GP2 11.8741
R14088 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n1 11.2645
R14089 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n4 8.64182
R14090 muxtest_0.x1.x3.GP2.n1 muxtest_0.x1.x3.GP2 6.1445
R14091 muxtest_0.x1.x3.GP2.n4 muxtest_0.x1.x3.GP2 5.75481
R14092 muxtest_0.x1.x3.GP2.n1 muxtest_0.x1.x3.GP2 4.65505
R14093 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n2 3.12276
R14094 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n3 2.94361
R14095 muxtest_0.x1.x3.GP2.n7 muxtest_0.x1.x3.GP2 2.0485
R14096 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP2.n7 1.55202
R14097 muxtest_0.R5R6.n0 muxtest_0.R5R6.t1 26.3998
R14098 muxtest_0.R5R6.n0 muxtest_0.R5R6.t2 23.5483
R14099 muxtest_0.R5R6.n1 muxtest_0.R5R6.t4 12.9758
R14100 muxtest_0.R5R6.n1 muxtest_0.R5R6.t5 10.8618
R14101 muxtest_0.R5R6.n4 muxtest_0.R5R6.t3 10.55
R14102 muxtest_0.R5R6.n2 muxtest_0.R5R6.n0 3.06895
R14103 muxtest_0.R5R6.n2 muxtest_0.R5R6.n1 2.14822
R14104 muxtest_0.R5R6.n3 muxtest_0.R5R6.n2 1.12636
R14105 muxtest_0.R5R6.n4 muxtest_0.R5R6.t0 1.11543
R14106 muxtest_0.R5R6 muxtest_0.R5R6.n4 0.694875
R14107 muxtest_0.R5R6 muxtest_0.R5R6.n3 0.132418
R14108 muxtest_0.R5R6.n3 muxtest_0.R5R6 0.0655
R14109 ringtest_0.x4._16_.n12 ringtest_0.x4._16_.t0 339.418
R14110 ringtest_0.x4._16_ ringtest_0.x4._16_.t1 269.426
R14111 ringtest_0.x4._16_.n1 ringtest_0.x4._16_.t7 264.029
R14112 ringtest_0.x4._16_ ringtest_0.x4._16_.n5 241.976
R14113 ringtest_0.x4._16_.n3 ringtest_0.x4._16_.t3 241.536
R14114 ringtest_0.x4._16_.n5 ringtest_0.x4._16_.t8 241.536
R14115 ringtest_0.x4._16_.n1 ringtest_0.x4._16_.t2 206.19
R14116 ringtest_0.x4._16_.n4 ringtest_0.x4._16_.n3 171.332
R14117 ringtest_0.x4._16_.n3 ringtest_0.x4._16_.t9 169.237
R14118 ringtest_0.x4._16_.n5 ringtest_0.x4._16_.t4 169.237
R14119 ringtest_0.x4._16_.n2 ringtest_0.x4._16_.n1 160.96
R14120 ringtest_0.x4._16_.n9 ringtest_0.x4._16_.n8 153.165
R14121 ringtest_0.x4._16_.n8 ringtest_0.x4._16_.t6 144.548
R14122 ringtest_0.x4._16_.n8 ringtest_0.x4._16_.t5 128.482
R14123 ringtest_0.x4._16_.n7 ringtest_0.x4._16_.n2 21.45
R14124 ringtest_0.x4._16_.n7 ringtest_0.x4._16_.n6 16.7975
R14125 ringtest_0.x4._16_.n10 ringtest_0.x4._16_ 15.8161
R14126 ringtest_0.x4._16_.n11 ringtest_0.x4._16_.n10 14.0946
R14127 ringtest_0.x4._16_ ringtest_0.x4._16_.n0 11.2645
R14128 ringtest_0.x4._16_ ringtest_0.x4._16_.n9 9.55788
R14129 ringtest_0.x4._16_.n6 ringtest_0.x4._16_ 6.4005
R14130 ringtest_0.x4._16_.n0 ringtest_0.x4._16_ 6.1445
R14131 ringtest_0.x4._16_.n2 ringtest_0.x4._16_ 5.4405
R14132 ringtest_0.x4._16_.n0 ringtest_0.x4._16_ 4.63498
R14133 ringtest_0.x4._16_.n4 ringtest_0.x4._16_ 4.44132
R14134 ringtest_0.x4._16_.n11 ringtest_0.x4._16_ 4.3525
R14135 ringtest_0.x4._16_.n13 ringtest_0.x4._16_.n12 4.0914
R14136 ringtest_0.x4._16_ ringtest_0.x4._16_.n13 3.61789
R14137 ringtest_0.x4._16_.n9 ringtest_0.x4._16_ 3.29747
R14138 ringtest_0.x4._16_.n13 ringtest_0.x4._16_.n11 2.3045
R14139 ringtest_0.x4._16_.n12 ringtest_0.x4._16_ 1.74382
R14140 ringtest_0.x4._16_.n6 ringtest_0.x4._16_.n4 1.50638
R14141 ringtest_0.x4._16_.n10 ringtest_0.x4._16_.n7 1.38649
R14142 muxtest_0.x2.x2.GP2.n2 muxtest_0.x2.x2.GP2.t4 450.938
R14143 muxtest_0.x2.x2.GP2.n2 muxtest_0.x2.x2.GP2.t5 445.666
R14144 muxtest_0.x2.x2.GP2.n4 muxtest_0.x2.x2.GP2.n3 195.958
R14145 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n0 96.8352
R14146 muxtest_0.x2.x2.GP2.n3 muxtest_0.x2.x2.GP2.t1 26.5955
R14147 muxtest_0.x2.x2.GP2.n3 muxtest_0.x2.x2.GP2.t0 26.5955
R14148 muxtest_0.x2.x2.GP2.n0 muxtest_0.x2.x2.GP2.t2 24.9236
R14149 muxtest_0.x2.x2.GP2.n0 muxtest_0.x2.x2.GP2.t3 24.9236
R14150 muxtest_0.x2.x2.GP2.n5 muxtest_0.x2.x2.GP2.n4 13.0077
R14151 muxtest_0.x2.x2.GP2.n4 muxtest_0.x2.x2.GP2 11.995
R14152 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n1 11.2645
R14153 muxtest_0.x2.x2.GP2.n1 muxtest_0.x2.x2.GP2 6.1445
R14154 muxtest_0.x2.x2.GP2.n1 muxtest_0.x2.x2.GP2 4.65505
R14155 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n2 3.12839
R14156 muxtest_0.x2.x2.GP2.n5 muxtest_0.x2.x2.GP2 2.0485
R14157 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP2.n5 1.55202
R14158 muxtest_0.R6R7.n0 muxtest_0.R6R7.t3 26.3998
R14159 muxtest_0.R6R7.n0 muxtest_0.R6R7.t2 23.5483
R14160 muxtest_0.R6R7.n4 muxtest_0.R6R7.t4 17.4454
R14161 muxtest_0.R6R7.n1 muxtest_0.R6R7.t1 12.9758
R14162 muxtest_0.R6R7.n1 muxtest_0.R6R7.t0 10.8618
R14163 muxtest_0.R6R7.n4 muxtest_0.R6R7.t5 10.5739
R14164 muxtest_0.R6R7.n2 muxtest_0.R6R7.n0 3.06895
R14165 muxtest_0.R6R7.n2 muxtest_0.R6R7.n1 2.14822
R14166 muxtest_0.R6R7.n3 muxtest_0.R6R7.n2 1.12636
R14167 muxtest_0.R6R7.n5 muxtest_0.R6R7 1.11925
R14168 muxtest_0.R6R7.n5 muxtest_0.R6R7.n4 0.370193
R14169 muxtest_0.R6R7 muxtest_0.R6R7.n3 0.138152
R14170 muxtest_0.R6R7.n5 muxtest_0.R6R7 0.073
R14171 muxtest_0.R6R7.n3 muxtest_0.R6R7 0.0655
R14172 muxtest_0.R6R7 muxtest_0.R6R7.n5 0.04925
R14173 ua[0].n6 ua[0].t6 26.3998
R14174 ua[0].n0 ua[0].t0 26.3998
R14175 ua[0].n6 ua[0].t5 23.5483
R14176 ua[0].n0 ua[0].t1 23.5483
R14177 ua[0].n7 ua[0].t3 12.9758
R14178 ua[0].n1 ua[0].t7 12.9758
R14179 ua[0].n5 ua[0] 12.8371
R14180 ua[0].n7 ua[0].t4 10.8618
R14181 ua[0].n1 ua[0].t8 10.8618
R14182 ua[0].n4 ua[0].t2 10.5739
R14183 ua[0].n8 ua[0].n6 3.06895
R14184 ua[0].n2 ua[0].n0 3.06895
R14185 ua[0].n8 ua[0].n7 2.14822
R14186 ua[0].n2 ua[0].n1 2.14822
R14187 ua[0].n4 ua[0] 1.39577
R14188 ua[0].n9 ua[0].n8 1.12636
R14189 ua[0].n3 ua[0].n2 1.12636
R14190 ua[0].n5 ua[0].n4 0.545106
R14191 ua[0] ua[0].n9 0.138152
R14192 ua[0] ua[0].n3 0.134513
R14193 ua[0].n9 ua[0] 0.0655
R14194 ua[0].n3 ua[0] 0.0655
R14195 ua[0] ua[0].n5 0.0579534
R14196 ua[0].n5 ua[0] 0.0532872
R14197 muxtest_0.R7R8.n5 muxtest_0.R7R8.t0 26.3998
R14198 muxtest_0.R7R8.n0 muxtest_0.R7R8.t8 26.3998
R14199 muxtest_0.R7R8.n5 muxtest_0.R7R8.t1 23.5483
R14200 muxtest_0.R7R8.n0 muxtest_0.R7R8.t7 23.5483
R14201 muxtest_0.R7R8.n6 muxtest_0.R7R8.t4 12.9758
R14202 muxtest_0.R7R8.n1 muxtest_0.R7R8.t6 12.9758
R14203 muxtest_0.R7R8.n6 muxtest_0.R7R8.t3 10.8618
R14204 muxtest_0.R7R8.n1 muxtest_0.R7R8.t5 10.8618
R14205 muxtest_0.R7R8.n4 muxtest_0.R7R8.t9 10.5709
R14206 muxtest_0.R7R8.n9 muxtest_0.R7R8 8.65896
R14207 muxtest_0.R7R8.n7 muxtest_0.R7R8.n5 3.06895
R14208 muxtest_0.R7R8.n2 muxtest_0.R7R8.n0 3.06895
R14209 muxtest_0.R7R8.n7 muxtest_0.R7R8.n6 2.14822
R14210 muxtest_0.R7R8.n2 muxtest_0.R7R8.n1 2.14822
R14211 muxtest_0.R7R8.n8 muxtest_0.R7R8.n7 1.12636
R14212 muxtest_0.R7R8.n3 muxtest_0.R7R8.n2 1.12636
R14213 muxtest_0.R7R8.n4 muxtest_0.R7R8.t2 1.01856
R14214 muxtest_0.R7R8 muxtest_0.R7R8.n9 0.32175
R14215 muxtest_0.R7R8.n9 muxtest_0.R7R8.n4 0.230945
R14216 muxtest_0.R7R8 muxtest_0.R7R8.n3 0.148615
R14217 muxtest_0.R7R8 muxtest_0.R7R8.n8 0.134513
R14218 muxtest_0.R7R8.n8 muxtest_0.R7R8 0.0655
R14219 muxtest_0.R7R8.n3 muxtest_0.R7R8 0.0655
R14220 ui_in[3].n18 ui_in[3].t0 327.99
R14221 ui_in[3].n5 ui_in[3].t19 327.99
R14222 ui_in[3].n22 ui_in[3].t4 293.969
R14223 ui_in[3].n9 ui_in[3].t17 293.969
R14224 ui_in[3].n16 ui_in[3].t11 261.887
R14225 ui_in[3].n3 ui_in[3].t10 261.887
R14226 ui_in[3].n13 ui_in[3].t5 212.081
R14227 ui_in[3].n14 ui_in[3].t8 212.081
R14228 ui_in[3].n0 ui_in[3].t18 212.081
R14229 ui_in[3].n1 ui_in[3].t3 212.081
R14230 ui_in[3].n18 ui_in[3].t14 199.457
R14231 ui_in[3].n5 ui_in[3].t9 199.457
R14232 ui_in[3].n15 ui_in[3].n14 183.185
R14233 ui_in[3].n2 ui_in[3].n1 183.185
R14234 ui_in[3].n16 ui_in[3].t7 155.847
R14235 ui_in[3].n3 ui_in[3].t6 155.847
R14236 ui_in[3] ui_in[3].n22 154.065
R14237 ui_in[3] ui_in[3].n9 154.065
R14238 ui_in[3].n17 ui_in[3].n16 153.506
R14239 ui_in[3].n4 ui_in[3].n3 153.506
R14240 ui_in[3].n19 ui_in[3].n18 152
R14241 ui_in[3].n6 ui_in[3].n5 152
R14242 ui_in[3].n13 ui_in[3].t13 139.78
R14243 ui_in[3].n14 ui_in[3].t16 139.78
R14244 ui_in[3].n0 ui_in[3].t2 139.78
R14245 ui_in[3].n1 ui_in[3].t12 139.78
R14246 ui_in[3].n22 ui_in[3].t1 138.338
R14247 ui_in[3].n9 ui_in[3].t15 138.338
R14248 ui_in[3].n14 ui_in[3].n13 61.346
R14249 ui_in[3].n1 ui_in[3].n0 61.346
R14250 ui_in[3].n26 ui_in[3] 36.5723
R14251 ui_in[3].n23 ui_in[3] 13.4199
R14252 ui_in[3].n10 ui_in[3] 13.4199
R14253 ui_in[3].n26 ui_in[3] 12.2088
R14254 ui_in[3].n24 ui_in[3].n21 11.7395
R14255 ui_in[3].n11 ui_in[3].n8 11.7395
R14256 ui_in[3].n25 ui_in[3].n24 11.5949
R14257 ui_in[3].n12 ui_in[3].n11 11.5949
R14258 ui_in[3].n21 ui_in[3].n17 10.4004
R14259 ui_in[3].n8 ui_in[3].n4 10.4004
R14260 ui_in[3].n25 ui_in[3].n15 9.68118
R14261 ui_in[3].n12 ui_in[3].n2 9.68118
R14262 ui_in[3].n19 ui_in[3] 9.6005
R14263 ui_in[3].n6 ui_in[3] 9.6005
R14264 ui_in[3].n15 ui_in[3] 5.8885
R14265 ui_in[3].n2 ui_in[3] 5.8885
R14266 ui_in[3].n23 ui_in[3] 5.57469
R14267 ui_in[3].n10 ui_in[3] 5.57469
R14268 ui_in[3].n21 ui_in[3].n20 4.6505
R14269 ui_in[3].n24 ui_in[3].n23 4.6505
R14270 ui_in[3].n8 ui_in[3].n7 4.6505
R14271 ui_in[3].n11 ui_in[3].n10 4.6505
R14272 ui_in[3].n20 ui_in[3].n19 2.98717
R14273 ui_in[3].n7 ui_in[3].n6 2.98717
R14274 ui_in[3].n17 ui_in[3] 2.82403
R14275 ui_in[3].n4 ui_in[3] 2.82403
R14276 ui_in[3].n20 ui_in[3] 1.9205
R14277 ui_in[3].n7 ui_in[3] 1.9205
R14278 ui_in[3] ui_in[3].n25 0.559212
R14279 ui_in[3] ui_in[3].n12 0.559212
R14280 ui_in[3] ui_in[3].n26 0.47425
R14281 ringtest_0.x3.x2.GP1.n2 ringtest_0.x3.x2.GP1.t5 450.938
R14282 ringtest_0.x3.x2.GP1.n2 ringtest_0.x3.x2.GP1.t4 445.666
R14283 ringtest_0.x3.x2.GP1.n4 ringtest_0.x3.x2.GP1.n3 195.832
R14284 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n0 96.8352
R14285 ringtest_0.x3.x2.GP1.n3 ringtest_0.x3.x2.GP1.t1 26.5955
R14286 ringtest_0.x3.x2.GP1.n3 ringtest_0.x3.x2.GP1.t0 26.5955
R14287 ringtest_0.x3.x2.GP1.n0 ringtest_0.x3.x2.GP1.t3 24.9236
R14288 ringtest_0.x3.x2.GP1.n0 ringtest_0.x3.x2.GP1.t2 24.9236
R14289 ringtest_0.x3.x2.GP1.n5 ringtest_0.x3.x2.GP1.n4 13.1346
R14290 ringtest_0.x3.x2.GP1.n4 ringtest_0.x3.x2.GP1 12.2007
R14291 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n1 11.2645
R14292 ringtest_0.x3.x2.GP1.n1 ringtest_0.x3.x2.GP1 6.1445
R14293 ringtest_0.x3.x2.GP1.n1 ringtest_0.x3.x2.GP1 4.65505
R14294 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n2 3.07707
R14295 ringtest_0.x3.x2.GP1.n5 ringtest_0.x3.x2.GP1 2.0485
R14296 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP1.n5 1.55202
R14297 ringtest_0.ring_out.n0 ringtest_0.ring_out.t13 844.321
R14298 ringtest_0.ring_out.n0 ringtest_0.ring_out.t12 354.322
R14299 ringtest_0.ring_out.n3 ringtest_0.ring_out.n1 243.68
R14300 ringtest_0.ring_out.n8 ringtest_0.ring_out.t10 212.081
R14301 ringtest_0.ring_out.n7 ringtest_0.ring_out.t11 212.081
R14302 ringtest_0.ring_out.n5 ringtest_0.ring_out.n4 206.249
R14303 ringtest_0.ring_out.n3 ringtest_0.ring_out.n2 205.28
R14304 ringtest_0.ring_out.n9 ringtest_0.ring_out.n8 184.806
R14305 ringtest_0.ring_out.n8 ringtest_0.ring_out.t14 139.78
R14306 ringtest_0.ring_out.n7 ringtest_0.ring_out.t15 139.78
R14307 ringtest_0.ring_out.n8 ringtest_0.ring_out.n7 61.346
R14308 ringtest_0.ring_out.n1 ringtest_0.ring_out.t1 26.5955
R14309 ringtest_0.ring_out.n1 ringtest_0.ring_out.t0 26.5955
R14310 ringtest_0.ring_out.n2 ringtest_0.ring_out.t6 26.5955
R14311 ringtest_0.ring_out.n2 ringtest_0.ring_out.t7 26.5955
R14312 ringtest_0.ring_out.n11 ringtest_0.ring_out.t4 26.3998
R14313 ringtest_0.ring_out ringtest_0.ring_out.n3 24.9955
R14314 ringtest_0.ring_out.n4 ringtest_0.ring_out.t8 24.9236
R14315 ringtest_0.ring_out.n4 ringtest_0.ring_out.t9 24.9236
R14316 ringtest_0.ring_out.n11 ringtest_0.ring_out.t5 23.5483
R14317 ringtest_0.ring_out.n10 ringtest_0.ring_out.n9 21.363
R14318 ringtest_0.ring_out ringtest_0.ring_out.n5 14.8576
R14319 ringtest_0.ring_out.n12 ringtest_0.ring_out.t3 12.9758
R14320 ringtest_0.ring_out.n6 ringtest_0.ring_out 10.9719
R14321 ringtest_0.ring_out.n12 ringtest_0.ring_out.t2 10.8618
R14322 ringtest_0.ring_out.n10 ringtest_0.ring_out.n6 9.53262
R14323 ringtest_0.ring_out.n6 ringtest_0.ring_out 4.57193
R14324 ringtest_0.ring_out.n13 ringtest_0.ring_out.n11 3.06895
R14325 ringtest_0.ring_out.n9 ringtest_0.ring_out 2.32777
R14326 ringtest_0.ring_out.n13 ringtest_0.ring_out.n12 2.14822
R14327 ringtest_0.ring_out ringtest_0.ring_out.n13 1.12636
R14328 ringtest_0.ring_out.n5 ringtest_0.ring_out 0.686214
R14329 ringtest_0.ring_out ringtest_0.ring_out.n10 0.631142
R14330 ringtest_0.ring_out ringtest_0.ring_out.n0 0.354518
R14331 ringtest_0.x3.x2.GP2.n2 ringtest_0.x3.x2.GP2.t4 450.938
R14332 ringtest_0.x3.x2.GP2.n2 ringtest_0.x3.x2.GP2.t5 445.666
R14333 ringtest_0.x3.x2.GP2.n4 ringtest_0.x3.x2.GP2.n3 195.958
R14334 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n0 96.8352
R14335 ringtest_0.x3.x2.GP2.n3 ringtest_0.x3.x2.GP2.t1 26.5955
R14336 ringtest_0.x3.x2.GP2.n3 ringtest_0.x3.x2.GP2.t0 26.5955
R14337 ringtest_0.x3.x2.GP2.n0 ringtest_0.x3.x2.GP2.t3 24.9236
R14338 ringtest_0.x3.x2.GP2.n0 ringtest_0.x3.x2.GP2.t2 24.9236
R14339 ringtest_0.x3.x2.GP2.n5 ringtest_0.x3.x2.GP2.n4 13.0077
R14340 ringtest_0.x3.x2.GP2.n4 ringtest_0.x3.x2.GP2 11.995
R14341 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n1 11.2645
R14342 ringtest_0.x3.x2.GP2.n1 ringtest_0.x3.x2.GP2 6.1445
R14343 ringtest_0.x3.x2.GP2.n1 ringtest_0.x3.x2.GP2 4.65505
R14344 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n2 3.12839
R14345 ringtest_0.x3.x2.GP2.n5 ringtest_0.x3.x2.GP2 2.0485
R14346 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP2.n5 1.55202
R14347 muxtest_0.x2.x2.GP4.n2 muxtest_0.x2.x2.GP4.t4 450.938
R14348 muxtest_0.x2.x2.GP4.n2 muxtest_0.x2.x2.GP4.t5 445.666
R14349 muxtest_0.x2.x2.GP4.n5 muxtest_0.x2.x2.GP4.n4 208.965
R14350 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n0 96.8352
R14351 muxtest_0.x2.x2.GP4.n4 muxtest_0.x2.x2.GP4.t1 26.5955
R14352 muxtest_0.x2.x2.GP4.n4 muxtest_0.x2.x2.GP4.t0 26.5955
R14353 muxtest_0.x2.x2.GP4.n0 muxtest_0.x2.x2.GP4.t3 24.9236
R14354 muxtest_0.x2.x2.GP4.n0 muxtest_0.x2.x2.GP4.t2 24.9236
R14355 muxtest_0.x2.x1.gpo3 muxtest_0.x2.x2.x4.GP 16.5032
R14356 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n3 10.2405
R14357 muxtest_0.x2.x2.GP4.n3 muxtest_0.x2.x1.gpo3 7.76481
R14358 muxtest_0.x2.x2.GP4.n1 muxtest_0.x2.x1.x14.Y 6.1445
R14359 muxtest_0.x2.x2.GP4.n1 muxtest_0.x2.x1.x14.Y 4.65505
R14360 muxtest_0.x2.x2.x4.GP muxtest_0.x2.x2.GP4.n2 2.95993
R14361 muxtest_0.x2.x2.GP4.n5 muxtest_0.x2.x1.x14.Y 2.0485
R14362 muxtest_0.x2.x1.x14.Y muxtest_0.x2.x2.GP4.n5 1.55202
R14363 muxtest_0.x2.x2.GP4.n3 muxtest_0.x2.x2.GP4.n1 1.0245
R14364 muxtest_0.R4R5.n0 muxtest_0.R4R5.t1 26.3998
R14365 muxtest_0.R4R5.n0 muxtest_0.R4R5.t2 23.5483
R14366 muxtest_0.R4R5.n1 muxtest_0.R4R5.t5 12.9758
R14367 muxtest_0.R4R5.n1 muxtest_0.R4R5.t4 10.8618
R14368 muxtest_0.R4R5.n4 muxtest_0.R4R5.t0 10.8231
R14369 muxtest_0.R4R5.n4 muxtest_0.R4R5.t3 10.5739
R14370 muxtest_0.R4R5.n2 muxtest_0.R4R5.n0 3.06895
R14371 muxtest_0.R4R5.n2 muxtest_0.R4R5.n1 2.14822
R14372 muxtest_0.R4R5.n3 muxtest_0.R4R5.n2 1.12636
R14373 muxtest_0.R4R5 muxtest_0.R4R5.n4 0.790021
R14374 muxtest_0.R4R5 muxtest_0.R4R5.n3 0.134513
R14375 muxtest_0.R4R5.n3 muxtest_0.R4R5 0.0655
R14376 muxtest_0.R2R3.n0 muxtest_0.R2R3.t4 26.3998
R14377 muxtest_0.R2R3.n0 muxtest_0.R2R3.t5 23.5483
R14378 muxtest_0.R2R3.n1 muxtest_0.R2R3.t2 12.9758
R14379 muxtest_0.R2R3.n1 muxtest_0.R2R3.t1 10.8618
R14380 muxtest_0.R2R3.n4 muxtest_0.R2R3.t0 10.8167
R14381 muxtest_0.R2R3.n4 muxtest_0.R2R3.t3 10.5739
R14382 muxtest_0.R2R3.n2 muxtest_0.R2R3.n0 3.06895
R14383 muxtest_0.R2R3.n2 muxtest_0.R2R3.n1 2.14822
R14384 muxtest_0.R2R3.n3 muxtest_0.R2R3.n2 1.12636
R14385 muxtest_0.R2R3 muxtest_0.R2R3.n4 0.71627
R14386 muxtest_0.R2R3 muxtest_0.R2R3.n3 0.138152
R14387 muxtest_0.R2R3.n3 muxtest_0.R2R3 0.0655
R14388 ui_in[6].n0 ui_in[6].t0 212.081
R14389 ui_in[6].n1 ui_in[6].t1 212.081
R14390 ui_in[6] ui_in[6].n2 152.512
R14391 ui_in[6].n0 ui_in[6].t2 139.78
R14392 ui_in[6].n1 ui_in[6].t3 139.78
R14393 ui_in[6].n2 ui_in[6].n0 30.6732
R14394 ui_in[6].n2 ui_in[6].n1 30.6732
R14395 ui_in[6].n3 ui_in[6] 16.4378
R14396 ui_in[6] ui_in[6].n3 0.7505
R14397 ui_in[6].n3 ui_in[6] 0.0808571
R14398 ui_in[5].n0 ui_in[5].t0 260.322
R14399 ui_in[5].n0 ui_in[5].t1 175.169
R14400 ui_in[5].n1 ui_in[5].n0 153.13
R14401 ui_in[5].n3 ui_in[5] 22.4521
R14402 ui_in[5] ui_in[5].n1 9.86591
R14403 ui_in[5].n3 ui_in[5].n2 4.07076
R14404 ui_in[5].n1 ui_in[5] 3.2005
R14405 ui_in[5].n2 ui_in[5] 0.960321
R14406 ui_in[5].n2 ui_in[5] 0.392836
R14407 ui_in[5] ui_in[5].n3 0.0499792
C0 ringtest_0.x4.net1 ringtest_0.x4._01_ 1.96e-19
C1 a_25925_6788# ringtest_0.x4._24_ 4.18e-19
C2 ringtest_0.x4._23_ a_26569_6422# 0.213625f
C3 ringtest_0.x4._09_ a_27273_4220# 0.17213f
C4 ringtest_0.x4.net2 ringtest_0.x4.clknet_1_0__leaf_clk 0.026712f
C5 ringtest_0.x4._00_ a_21675_9686# 0.07841f
C6 a_21425_9686# a_21561_9116# 7.31e-19
C7 a_26749_6422# a_26201_4790# 3.35e-21
C8 a_26201_4790# ringtest_0.x4.net11 3.07e-19
C9 ringtest_0.x4._09_ a_26766_4790# 3.07e-19
C10 ringtest_0.x4._02_ a_21840_5308# 4.65e-19
C11 a_21233_5340# a_21672_5334# 0.273138f
C12 ringtest_0.x4._22_ a_26367_5340# 4.96e-21
C13 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x3.nselect2 5.69e-21
C14 ringtest_0.x4._08_ a_27149_5334# 2.34e-19
C15 ringtest_0.x4.counter[9] VDPWR 0.438942f
C16 ringtest_0.x4._18_ a_24329_6640# 6.58e-19
C17 a_21785_8054# VDPWR 0.264209f
C18 ringtest_0.x4.net8 a_23770_5308# 2.76e-19
C19 a_23879_6940# a_24336_6544# 0.016444f
C20 ringtest_0.x4._20_ a_25593_5156# 1.2e-20
C21 ringtest_0.x4.clknet_1_0__leaf_clk a_22181_5334# 3.7e-19
C22 ringtest_0.x4._11_ a_21672_5334# 0.003174f
C23 ringtest_0.x4._07_ ringtest_0.x4.counter[5] 1.62e-19
C24 a_27491_4566# VDPWR 0.003335f
C25 ringtest_0.counter3 m3_17046_7066# 8.01e-20
C26 ringtest_0.x4.clknet_0_clk a_22817_6146# 3.43e-19
C27 a_25055_3867# ringtest_0.x4.counter[5] 0.1107f
C28 muxtest_0.R7R8 ui_in[4] 0.104361f
C29 ringtest_0.drv_out m3_17036_9140# 0.132758f
C30 ringtest_0.x4.clknet_1_1__leaf_clk a_26640_5334# 0.001015f
C31 ringtest_0.x4.net6 a_22765_5308# 0.080758f
C32 ringtest_0.x4.clknet_0_clk a_26095_6788# 9.17e-20
C33 a_12019_24012# VDPWR 9.09e-19
C34 ringtest_0.x4._11_ ringtest_0.x4._24_ 4.57e-19
C35 a_27273_4220# a_27659_4246# 0.006406f
C36 a_23949_6654# a_23837_5878# 2.76e-20
C37 ringtest_0.x4.clknet_1_0__leaf_clk a_22399_8976# 0.018091f
C38 ringtest_0.x4._23_ a_27489_3702# 9.55e-20
C39 ringtest_0.x4._14_ ringtest_0.x4.net5 0.258421f
C40 a_24329_6640# a_24763_6143# 0.00484f
C41 a_27149_5334# VDPWR 0.005027f
C42 ringtest_0.x4._16_ a_25336_4902# 8.82e-22
C43 a_21399_5340# a_21948_5156# 0.002f
C44 ringtest_0.x4.net9 a_25168_5156# 0.003585f
C45 ringtest_0.x4.net11 a_27303_4246# 0.01512f
C46 a_26808_4902# a_26895_3867# 2.21e-20
C47 a_21672_5334# a_21675_4790# 0.004962f
C48 ringtest_0.x4.net1 a_21785_8054# 0.232539f
C49 ringtest_0.x4.net6 ringtest_0.x4._13_ 2.81e-21
C50 a_25925_6788# a_26007_6788# 0.005781f
C51 ringtest_0.x4.net2 ringtest_0.x4.net4 8.49e-21
C52 a_25225_5334# a_26367_5340# 8.68e-20
C53 a_22097_5334# a_22223_5712# 0.006169f
C54 a_22097_5334# VDPWR 0.22678f
C55 ringtest_0.x4.clknet_1_1__leaf_clk a_25149_4220# 1.84e-19
C56 muxtest_0.x1.x1.nSEL1 a_19842_32287# 1.59e-19
C57 ringtest_0.x4.net4 a_23381_4818# 4.87e-19
C58 ringtest_0.x4._16_ VDPWR 2.15022f
C59 a_26201_4790# ringtest_0.x4._09_ 0.098799f
C60 ringtest_0.x4.net7 a_25168_5156# 0.005696f
C61 a_24329_6640# ringtest_0.x4.clknet_1_1__leaf_clk 0.228247f
C62 ringtest_0.x4._03_ a_22390_4566# 9.33e-19
C63 a_22695_8304# VDPWR 0.006514f
C64 ringtest_0.x3.x2.GN4 ua[1] 0.446629f
C65 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.025028f
C66 muxtest_0.x1.x3.GN2 ui_in[2] 0.001516f
C67 a_24763_6143# a_24545_5878# 0.004465f
C68 ringtest_0.x4._06_ ringtest_0.x4._07_ 5.11e-20
C69 a_11845_23906# a_12297_23648# 0.002207f
C70 a_16755_12091# ringtest_0.x3.x2.GN4 0.003699f
C71 ringtest_0.x3.x2.GN1 a_15749_12123# 0.001144f
C72 ringtest_0.x4._04_ a_21840_5308# 8.38e-20
C73 a_24004_6128# a_23837_5878# 0.046138f
C74 a_17231_12017# ringtest_0.x3.x2.GN2 7.58e-21
C75 a_21785_5878# a_21672_5334# 0.002054f
C76 ringtest_0.x4._14_ a_21007_3867# 0.001394f
C77 ringtest_0.x4._23_ a_26640_5334# 0.012578f
C78 ringtest_0.x4.clknet_1_0__leaf_clk a_21840_5308# 0.01796f
C79 a_26367_5340# a_26640_5156# 1.54e-19
C80 ringtest_0.x4._18_ a_23151_5334# 2.06e-20
C81 a_26808_5308# a_26808_4902# 0.012451f
C82 a_26640_5334# a_26367_4790# 1.54e-19
C83 ringtest_0.x4._16_ a_23467_4584# 8.82e-20
C84 ringtest_0.x4._11_ a_22224_6244# 0.054008f
C85 a_21852_9416# ui_in[5] 4.56e-21
C86 muxtest_0.x1.x4.A muxtest_0.R4R5 0.003925f
C87 ringtest_0.x4.net3 a_21395_6940# 0.011213f
C88 a_24536_6699# a_24527_5340# 8.21e-21
C89 a_24329_6640# a_24800_5334# 8.34e-21
C90 a_24465_6800# a_24361_5340# 5.48e-20
C91 ringtest_0.x4._11_ a_26007_6788# 2.28e-19
C92 ringtest_0.x4.clknet_1_1__leaf_clk a_24545_5878# 3.57e-20
C93 VDPWR ui_in[4] 9.576571f
C94 ringtest_0.x4.net11 ringtest_0.x4.counter[8] 0.024563f
C95 ringtest_0.x4.clknet_0_clk a_24536_6699# 0.004436f
C96 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VDPWR 0.636224f
C97 ringtest_0.x4.net6 ringtest_0.x4.net8 0.806426f
C98 a_21852_9416# ringtest_0.x4._12_ 0.003541f
C99 ringtest_0.x4.clknet_1_1__leaf_clk a_25364_5878# 1.80017f
C100 a_21425_9686# a_21785_8054# 2.44e-21
C101 ringtest_0.x4._09_ a_27303_4246# 0.07143f
C102 muxtest_0.x2.nselect2 ui_in[3] 1.88e-19
C103 ringtest_0.x4.net8 a_24895_4790# 0.003497f
C104 a_17231_12017# ui_in[3] 0.220366f
C105 ringtest_0.x4._23_ a_25149_4220# 2.79e-19
C106 a_23809_4790# ringtest_0.x4.counter[4] 2.6e-19
C107 ringtest_0.x4._23_ a_26735_5156# 8.32e-19
C108 a_26808_4902# a_26555_4790# 3.39e-19
C109 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP1 8.08e-19
C110 muxtest_0.R7R8 ui_in[0] 2.25e-21
C111 ringtest_0.x4._06_ a_26201_5340# 4.19e-21
C112 ringtest_0.x4.net10 a_26817_4566# 8.38e-19
C113 ringtest_0.x4.net6 a_24729_4790# 0.083542f
C114 ringtest_0.x4._18_ ringtest_0.x4._19_ 0.036736f
C115 a_12473_23980# muxtest_0.x2.x2.GN2 0.017071f
C116 a_22649_6244# VDPWR 0.169028f
C117 ringtest_0.x4.clknet_1_1__leaf_clk a_24317_4942# 0.050301f
C118 a_24729_4790# a_24895_4790# 0.966391f
C119 ringtest_0.x4._21_ ringtest_0.x4._16_ 0.249175f
C120 ringtest_0.x4._16_ ringtest_0.x4.counter[2] 3.86e-19
C121 a_26201_6788# VDPWR 0.002272f
C122 ringtest_0.x4.net4 a_21840_5308# 5.24e-19
C123 ringtest_0.x4.clknet_1_1__leaf_clk a_23151_5334# 8.24e-20
C124 ringtest_0.x4._03_ a_22074_4790# 0.001074f
C125 a_21509_4790# ringtest_0.x4.net5 8.46e-19
C126 ringtest_0.x4._15_ a_26367_5340# 0.058771f
C127 ringtest_0.x3.x1.nSEL0 a_16203_12091# 0.001174f
C128 ringtest_0.x4._22_ a_26375_4612# 2.76e-20
C129 ringtest_0.x3.x2.GP1 VDPWR 1.86466f
C130 ringtest_0.x4._04_ a_22392_5990# 0.04931f
C131 a_21785_5878# a_22224_6244# 0.269567f
C132 a_23467_4818# VDPWR 0.00273f
C133 ringtest_0.x4._18_ a_22265_5308# 3.26e-20
C134 ringtest_0.x4._11_ a_25977_4220# 0.19543f
C135 a_22765_5308# ringtest_0.x4.net5 0.001034f
C136 ringtest_0.x4._23_ a_25364_5878# 0.042503f
C137 ringtest_0.x4.clknet_1_0__leaf_clk a_22392_5990# 5.16e-19
C138 muxtest_0.x1.x3.GN1 ua[3] 4.34e-20
C139 a_21852_9416# a_22245_8054# 6.42e-21
C140 ringtest_0.x4._11_ a_25719_4790# 2.44e-19
C141 ringtest_0.x3.x2.GN4 m3_17046_7066# 0.084813f
C142 a_25364_5878# a_26367_4790# 2.14e-19
C143 a_23837_5878# ringtest_0.x4._20_ 6.22e-20
C144 ringtest_0.x4._22_ ringtest_0.x4._20_ 2.69e-20
C145 a_19114_31955# ui_in[1] 0.03417f
C146 a_23879_6940# ringtest_0.x4._16_ 4.51e-19
C147 a_24361_5340# a_26555_5334# 2.33e-21
C148 ringtest_0.counter7 ringtest_0.x4.net9 0.006102f
C149 ringtest_0.x4._11_ a_24336_6544# 3.7e-19
C150 muxtest_0.x1.x5.GN muxtest_0.x1.x5.A 4.01025f
C151 muxtest_0.x1.x3.GN2 a_19794_32347# 3.11e-20
C152 a_19242_32347# muxtest_0.x1.x3.GN3 5.17e-20
C153 a_21587_5334# VDPWR 0.075425f
C154 ringtest_0.ring_out ringtest_0.x3.x2.GP2 0.080385f
C155 ringtest_0.x4._15_ a_22765_4478# 1.84e-19
C156 ringtest_0.x4.net6 a_26749_6422# 7.38e-20
C157 a_19842_32287# muxtest_0.x1.x3.GN1 1.69e-20
C158 a_25761_5058# a_25977_4220# 0.001105f
C159 muxtest_0.x1.x5.GN a_19114_31955# 3.56e-19
C160 muxtest_0.x1.x4.A ui_in[2] 4.96786f
C161 ringtest_0.x4._05_ ringtest_0.x4.net6 0.03493f
C162 a_23949_6654# ringtest_0.x4._15_ 1.78e-19
C163 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ui_in[4] 4.96e-21
C164 a_25761_5058# a_25719_4790# 7.84e-20
C165 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._19_ 0.060342f
C166 ringtest_0.x4._18_ ringtest_0.x4.net7 0.004371f
C167 ringtest_0.counter7 ringtest_0.x4.net7 6.88e-20
C168 a_22541_5058# a_22765_4478# 0.001036f
C169 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 3.14e-21
C170 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.001676f
C171 ringtest_0.x4._24_ ringtest_0.x4.net10 0.13484f
C172 a_19666_31955# ui_in[2] 0.009143f
C173 VDPWR ui_in[0] 1.24711f
C174 ringtest_0.x4._17_ ringtest_0.x4._18_ 0.181987f
C175 a_22139_5878# a_21233_5340# 3.23e-19
C176 muxtest_0.R3R4 muxtest_0.x2.x2.GN2 0.015374f
C177 ringtest_0.x4.net9 a_24763_6143# 0.122363f
C178 a_12849_23648# ui_in[4] 0.261734f
C179 ringtest_0.x4.net3 VDPWR 2.09599f
C180 a_27273_4220# VDPWR 0.229336f
C181 a_24070_5852# ringtest_0.x4._06_ 0.004838f
C182 a_21845_9116# VDPWR 0.716493f
C183 ringtest_0.x4.net8 a_23932_6128# 0.001644f
C184 a_22649_6244# ringtest_0.x4._21_ 8.88e-21
C185 ringtest_0.x4._11_ a_22139_5878# 0.020189f
C186 a_27659_4246# ringtest_0.x4.counter[8] 1.28e-20
C187 ringtest_0.x4._19_ a_24800_5334# 6.46e-21
C188 a_24465_6800# VDPWR 0.187397f
C189 ringtest_0.x4._01_ ringtest_0.x4._11_ 0.20957f
C190 ringtest_0.x4._12_ ringtest_0.x4._10_ 0.002721f
C191 ringtest_0.x4.net4 a_22392_5990# 0.034264f
C192 ringtest_0.x4.net7 a_24763_6143# 1.85e-20
C193 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net9 0.461828f
C194 a_21561_8830# a_21852_8720# 0.192341f
C195 ringtest_0.x4._15_ a_24004_6128# 5.11e-20
C196 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VDPWR 0.636188f
C197 a_25149_4220# a_25441_4612# 0.001675f
C198 ringtest_0.x4._23_ a_26913_4566# 2.44e-19
C199 ringtest_0.x4._17_ a_24763_6143# 2.72e-19
C200 a_25364_5878# a_25593_5156# 0.001605f
C201 muxtest_0.x1.x1.nSEL0 ui_in[1] 0.137587f
C202 a_26749_6422# a_27169_6641# 0.017591f
C203 ringtest_0.counter7 ringtest_0.x4.counter[0] 0.003899f
C204 a_22052_9116# a_21981_9142# 0.239923f
C205 ringtest_0.x4.net2 a_21561_8830# 0.00144f
C206 ringtest_0.drv_out ua[1] 4.52048f
C207 a_21465_9294# ringtest_0.x4.clknet_1_0__leaf_clk 0.007095f
C208 ringtest_0.x4._18_ a_22817_6146# 0.001543f
C209 ringtest_0.x4._08_ a_26201_4790# 1.13e-19
C210 ringtest_0.x4.net8 ringtest_0.x4.net5 0.002187f
C211 ringtest_0.x4.net1 ringtest_0.x4.net3 0.313425f
C212 ringtest_0.x4._11_ a_21863_4790# 4.78e-19
C213 ringtest_0.ring_out a_16707_12151# 2.99e-20
C214 ringtest_0.x4.net1 a_21845_9116# 0.003904f
C215 a_22111_10993# a_22052_9116# 2.02e-20
C216 ringtest_0.ring_out ringtest_0.x3.x2.GN2 0.23158f
C217 a_23770_5308# a_24361_5340# 0.044245f
C218 ringtest_0.x4._19_ ringtest_0.x4._23_ 2.58e-20
C219 ringtest_0.x4.net10 a_27815_3867# 0.219068f
C220 ringtest_0.x4.net8 a_24895_5334# 4.84e-19
C221 ringtest_0.x4.net6 ringtest_0.x4._09_ 1.5e-20
C222 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net7 0.397702f
C223 ringtest_0.x4._15_ a_23963_4790# 2.18e-19
C224 ringtest_0.x4._11_ a_23899_5334# 0.07562f
C225 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x5.GN 0.043714f
C226 ringtest_0.x4._16_ a_24968_5308# 0.001117f
C227 muxtest_0.x2.x2.GP3 ua[2] 0.357853f
C228 ringtest_0.x4.net9 a_24800_5334# 6.38e-21
C229 ringtest_0.x4._08_ a_26555_5334# 0.134213f
C230 a_25168_5156# a_25294_4790# 0.005525f
C231 a_22733_6244# VDPWR 0.004177f
C232 ringtest_0.x4.clknet_0_clk a_22765_5308# 4.87e-21
C233 ringtest_0.x4._15_ a_23381_4818# 0.22097f
C234 ringtest_0.x4._17_ ringtest_0.x4.clknet_1_1__leaf_clk 0.044595f
C235 ringtest_0.x4._23_ a_26735_5334# 8.32e-19
C236 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN2 0.154394f
C237 ringtest_0.x3.x2.GN3 ringtest_0.counter7 0.005062f
C238 muxtest_0.R7R8 muxtest_0.x2.x2.GN4 3.97956f
C239 a_22541_5058# a_23381_4818# 7.43e-20
C240 ringtest_0.x4._14_ a_22486_4246# 0.003598f
C241 a_21675_4790# a_21863_4790# 0.097994f
C242 ringtest_0.x4.net7 a_24800_5334# 0.034093f
C243 a_21785_8054# ringtest_0.x4._11_ 0.005192f
C244 a_21785_5878# a_22139_5878# 0.062224f
C245 a_26201_4790# VDPWR 0.658381f
C246 ringtest_0.x4._10_ a_22245_8054# 0.423817f
C247 uio_in[5] uio_in[4] 0.031023f
C248 ringtest_0.ring_out ui_in[3] 3.69e-19
C249 muxtest_0.x1.x3.GP3 ua[3] 0.023203f
C250 ringtest_0.x4.net3 ringtest_0.x4.counter[2] 7.38e-19
C251 ringtest_0.x4._17_ a_24800_5334# 9.6e-21
C252 ringtest_0.x4._23_ ringtest_0.x4.net9 0.065132f
C253 a_11845_23906# VDPWR 0.211573f
C254 a_22457_5156# VDPWR 0.004413f
C255 ua[3] ua[5] 0.008019f
C256 ringtest_0.x4.net9 a_26367_4790# 0.047741f
C257 a_27233_5308# ringtest_0.x4.net10 0.084593f
C258 a_23899_5654# a_23899_5334# 6.96e-20
C259 a_27065_5334# a_27191_5712# 0.006169f
C260 ringtest_0.x4.clknet_1_0__leaf_clk a_21981_8976# 0.024273f
C261 a_24465_6800# ringtest_0.x4._21_ 1.21e-19
C262 a_26555_5334# VDPWR 0.077172f
C263 ringtest_0.x4.net2 a_21049_8598# 0.07281f
C264 ringtest_0.x4._15_ a_26375_4612# 0.002119f
C265 a_19842_32287# muxtest_0.x1.x3.GP3 4.69e-19
C266 a_19666_31955# a_19794_32347# 0.004764f
C267 muxtest_0.x2.x1.nSEL1 ui_in[2] 8.19e-21
C268 ringtest_0.x4._00_ a_21561_9116# 0.001635f
C269 a_21425_9686# a_21845_9116# 0.001828f
C270 ringtest_0.x4._24_ a_26808_4902# 0.014122f
C271 ringtest_0.x4.net7 ringtest_0.x4._23_ 0.074369f
C272 ringtest_0.x4.net7 a_26367_4790# 0.001362f
C273 ringtest_0.x4._02_ a_22265_5308# 1.8e-19
C274 ringtest_0.x4.net5 a_22390_4566# 0.075434f
C275 a_21233_5340# a_22097_5334# 0.032244f
C276 ringtest_0.counter7 a_26627_4246# 1.91e-19
C277 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ui_in[4] 4.96e-21
C278 ringtest_0.x4._17_ ringtest_0.x4._23_ 0.082072f
C279 ringtest_0.x4._04_ a_23151_5334# 2.55e-19
C280 ringtest_0.x4._15_ ringtest_0.x4._20_ 0.093509f
C281 ringtest_0.x4._16_ a_21233_5340# 0.001516f
C282 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP2 2.65608f
C283 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.025028f
C284 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 7.08e-21
C285 ringtest_0.x4.net10 a_25977_4220# 0.158335f
C286 ringtest_0.x4._18_ a_24536_6699# 5.4e-20
C287 ringtest_0.x4.net8 a_24527_5340# 0.031957f
C288 muxtest_0.R1R2 ua[3] 0.017912f
C289 a_23879_6940# a_24465_6800# 0.013455f
C290 ringtest_0.x4._11_ a_22097_5334# 0.017838f
C291 a_27303_4246# VDPWR 0.283149f
C292 ringtest_0.x3.x1.nSEL1 a_16707_12151# 4.08e-19
C293 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN2 0.209956f
C294 ringtest_0.x4._11_ ringtest_0.x4._16_ 0.223435f
C295 a_15575_12017# ringtest_0.x3.x2.GN1 0.12869f
C296 a_22373_5156# a_22499_4790# 0.006169f
C297 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net8 8.45e-19
C298 ringtest_0.x4._11_ a_22695_8304# 0.002858f
C299 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A a_15575_12017# 6.58e-22
C300 ringtest_0.x4.clknet_1_1__leaf_clk a_27065_5334# 1.84e-19
C301 a_21007_3867# ringtest_0.x4.counter[1] 0.057818f
C302 ringtest_0.x4.net6 a_24361_5340# 0.0618f
C303 muxtest_0.x2.x2.GN4 VDPWR 1.23441f
C304 ringtest_0.x4._22_ a_25149_4220# 0.106132f
C305 a_24527_5340# a_24729_4790# 0.003672f
C306 a_24361_5340# a_24895_4790# 0.003047f
C307 muxtest_0.x1.x3.GN2 muxtest_0.R2R3 3.99837f
C308 ringtest_0.x4.net3 a_21375_3867# 0.233128f
C309 ringtest_0.x4.clknet_1_0__leaf_clk a_22228_8598# 0.002447f
C310 ringtest_0.x4._03_ VDPWR 0.386375f
C311 a_24329_6640# ringtest_0.x4._22_ 1.01e-19
C312 a_24536_6699# a_24763_6143# 3.7e-19
C313 muxtest_0.x1.x3.GN2 ui_in[1] 0.108644f
C314 a_21672_5334# a_21948_5156# 4.47e-19
C315 ringtest_0.x4.net9 a_25593_5156# 0.031858f
C316 a_22265_5308# a_22116_4902# 0.001344f
C317 a_22097_5334# a_21675_4790# 0.003824f
C318 ringtest_0.x4.counter[5] ua[1] 3.21e-19
C319 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VDPWR 0.638508f
C320 ringtest_0.x4.clknet_0_clk a_24729_4790# 1.17e-21
C321 ringtest_0.x4._00_ ringtest_0.x4._01_ 0.014628f
C322 a_25925_6788# a_26201_6788# 0.00119f
C323 m2_11882_23495# ui_in[4] 0.183786f
C324 ringtest_0.x4._16_ a_21675_4790# 2.51e-21
C325 ringtest_0.x3.x1.nSEL1 m2_15612_11606# 0.00815f
C326 a_22765_5308# a_22983_5654# 0.007234f
C327 a_26201_5340# a_26808_5308# 0.141453f
C328 ringtest_0.x3.x1.nSEL1 ui_in[3] 0.168464f
C329 ringtest_0.x4._15_ a_26569_6422# 0.001697f
C330 a_23770_5308# VDPWR 0.169696f
C331 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN2 7.45e-19
C332 ringtest_0.x4._16_ a_23899_5654# 0.001343f
C333 a_24045_6654# a_24264_6788# 0.006169f
C334 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN1 0.034842f
C335 ringtest_0.x4.net7 a_25593_5156# 0.040127f
C336 a_12473_23980# muxtest_0.x2.x2.GP1 2.33e-21
C337 a_24536_6699# ringtest_0.x4.clknet_1_1__leaf_clk 4.65e-20
C338 ringtest_0.x4._03_ a_23467_4584# 5.07e-20
C339 ringtest_0.x4.counter[8] VDPWR 0.211772f
C340 a_21939_8054# VDPWR 1.78e-19
C341 ringtest_0.x4.net4 a_23151_5334# 6.79e-19
C342 ringtest_0.x4._22_ a_24545_5878# 9.75e-19
C343 ringtest_0.x3.x2.GN3 a_16707_12151# 0.001073f
C344 ringtest_0.x3.x2.GN2 a_17405_12123# 8.14e-21
C345 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN4 0.001072f
C346 a_12297_23648# a_12473_23980# 0.185422f
C347 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GN3 0.067463f
C348 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP3 0.005595f
C349 ringtest_0.x4._04_ a_22265_5308# 0.008333f
C350 a_21785_5878# a_22097_5334# 0.001393f
C351 a_24699_6200# ringtest_0.x4._07_ 0.096566f
C352 ringtest_0.x4._14_ a_22295_3867# 4.42e-19
C353 a_25364_5878# ringtest_0.x4._22_ 8.12e-19
C354 a_22074_4790# ringtest_0.x4.net5 3e-19
C355 a_25225_5334# a_25149_4220# 3.32e-21
C356 muxtest_0.x2.nselect2 ua[3] 0.005153f
C357 a_21785_5878# ringtest_0.x4._16_ 6.86e-20
C358 ringtest_0.x4.clknet_1_0__leaf_clk a_22265_5308# 0.002373f
C359 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A a_16203_12091# 2.34e-20
C360 a_26367_5340# a_27065_5156# 1.3e-19
C361 a_25055_3867# ringtest_0.x4.counter[6] 4.98e-19
C362 a_27065_5334# a_26367_4790# 1.3e-19
C363 a_26640_5334# a_26640_5156# 0.013839f
C364 ringtest_0.x4._11_ a_22649_6244# 0.043928f
C365 a_22052_9116# ui_in[5] 1.46e-21
C366 ringtest_0.x4._17_ a_23993_5654# 3.09e-20
C367 a_21951_5878# a_24070_5852# 8.39e-21
C368 ringtest_0.x4.net9 a_25441_4612# 6.97e-19
C369 ringtest_0.x4._05_ a_24527_5340# 2.65e-21
C370 ui_in[6] uio_in[0] 0.001316f
C371 ringtest_0.x4.clknet_0_clk a_26749_6422# 1.5e-20
C372 ringtest_0.x4._11_ a_26201_6788# 0.005861f
C373 muxtest_0.x1.x3.GP1 muxtest_0.R4R5 0.123828f
C374 muxtest_0.x2.x2.GP3 m3_13302_19985# 0.002824f
C375 ringtest_0.x4._13_ a_21591_6128# 0.01129f
C376 ringtest_0.ring_out a_17377_14114# 0.105448f
C377 muxtest_0.x1.x3.GN3 muxtest_0.R7R8 0.129382f
C378 ringtest_0.x4.net1 a_21939_8054# 0.002601f
C379 ringtest_0.x4.clknet_0_clk ringtest_0.x4._05_ 0.067252f
C380 a_22052_9116# ringtest_0.x4._12_ 5.69e-20
C381 ringtest_0.x4._07_ a_23809_4790# 1.81e-20
C382 a_17405_12123# ui_in[3] 1.4e-19
C383 ringtest_0.x3.x2.GN3 ui_in[3] 0.254198f
C384 ringtest_0.drv_out a_25421_6641# 0.012863f
C385 ringtest_0.x4.net7 a_25441_4612# 0.006602f
C386 ringtest_0.x4._23_ a_26627_4246# 0.04546f
C387 ringtest_0.x4.net6 ringtest_0.x4._08_ 5.42e-20
C388 ringtest_0.x4.net8 a_25168_5156# 0.001808f
C389 ringtest_0.x4._11_ a_23467_4818# 0.003027f
C390 ringtest_0.x4._17_ ringtest_0.x4._04_ 6.62e-21
C391 a_26367_4790# a_26627_4246# 0.008374f
C392 muxtest_0.x2.x2.GP2 muxtest_0.x2.x2.GP3 0.031766f
C393 a_21233_5340# a_21587_5334# 0.062224f
C394 ringtest_0.x4.net10 ringtest_0.x4.counter[9] 0.092658f
C395 a_21951_5878# a_22373_5156# 0.001133f
C396 a_26367_4790# a_27149_5156# 6.32e-19
C397 a_22224_6244# a_21948_5156# 9.19e-21
C398 a_26640_5156# a_26735_5156# 0.007724f
C399 a_22392_5990# a_22541_5058# 8.5e-21
C400 a_23899_5334# ringtest_0.x4.counter[4] 4.47e-20
C401 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._17_ 3.38e-20
C402 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ui_in[4] 4.1e-20
C403 ringtest_0.x4.net10 a_27491_4566# 0.002502f
C404 ringtest_0.x4.clknet_1_1__leaf_clk a_25294_4790# 4.82e-19
C405 ringtest_0.x4.net6 a_25336_4902# 6.78e-21
C406 a_12849_23648# muxtest_0.x2.x2.GN4 6.84e-19
C407 ringtest_0.x4._11_ a_21587_5334# 2.52e-19
C408 a_25364_5878# a_25225_5334# 5.73e-19
C409 ringtest_0.x4._21_ a_23770_5308# 0.005326f
C410 muxtest_0.R3R4 muxtest_0.x2.x2.GP1 0.011522f
C411 a_13025_23980# muxtest_0.x2.x2.GN2 5.62e-20
C412 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 1.11e-20
C413 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.001676f
C414 a_24895_4790# a_25336_4902# 0.110715f
C415 a_24729_4790# a_25168_5156# 0.273138f
C416 a_19114_31955# ui_in[0] 0.246193f
C417 a_24712_6422# VDPWR 0.004407f
C418 ringtest_0.counter3 ringtest_0.x4._16_ 1.05e-19
C419 ringtest_0.x4.net4 a_22265_5308# 0.110738f
C420 ringtest_0.x4.counter[5] ringtest_0.x4.counter[6] 0.070133f
C421 ringtest_0.x3.x1.nSEL0 a_16755_12091# 1.21e-20
C422 ringtest_0.x4.net3 a_21233_5340# 0.023332f
C423 ringtest_0.x4._15_ a_26640_5334# 0.001174f
C424 ringtest_0.x4._22_ a_26913_4566# 3.67e-19
C425 ringtest_0.x4.net6 VDPWR 3.03875f
C426 muxtest_0.x1.x4.A muxtest_0.R2R3 4.52053f
C427 a_21785_5878# a_22649_6244# 0.030894f
C428 ringtest_0.x4._04_ a_22817_6146# 0.003723f
C429 ringtest_0.x4.net10 a_27149_5334# 3.67e-19
C430 a_24895_4790# VDPWR 0.315465f
C431 ringtest_0.x4.net3 ringtest_0.x4._11_ 0.005186f
C432 ringtest_0.x4._18_ a_22765_5308# 0.002375f
C433 muxtest_0.x1.x3.GP2 muxtest_0.R7R8 0.131352f
C434 ringtest_0.x4._19_ ringtest_0.x4._22_ 7e-20
C435 a_23879_6940# a_23770_5308# 4.81e-21
C436 ringtest_0.x4._11_ a_27273_4220# 2.01e-20
C437 ringtest_0.x4.clknet_1_0__leaf_clk a_22817_6146# 1.77e-20
C438 muxtest_0.x1.x3.GN3 muxtest_0.R5R6 4.12612f
C439 a_21845_9116# ringtest_0.x4._11_ 8.58e-21
C440 ringtest_0.x4._11_ a_26766_4790# 4.03e-21
C441 a_25364_5878# a_26640_5156# 6.58e-20
C442 a_27169_6641# ringtest_0.x4._08_ 0.109717f
C443 a_19666_31955# ui_in[1] 0.261734f
C444 ringtest_0.x4._11_ a_24465_6800# 5.19e-20
C445 a_24361_5340# a_24895_5334# 0.001632f
C446 a_21465_9294# a_21561_8830# 6.79e-19
C447 a_24045_6654# a_24070_5852# 0.006438f
C448 a_23949_6654# a_24004_6128# 3.4e-19
C449 a_21561_9116# a_21465_8830# 6.79e-19
C450 muxtest_0.x1.x5.GN muxtest_0.x1.x4.A 4.14763f
C451 a_21055_5334# VDPWR 0.0067f
C452 muxtest_0.x1.x3.GN3 VDPWR 0.766397f
C453 ringtest_0.x4._15_ a_25149_4220# 1.2e-20
C454 ringtest_0.x4._19_ a_23619_6788# 8.17e-20
C455 ringtest_0.x4.net6 ringtest_0.x4._25_ 2.22e-20
C456 ringtest_0.x4._17_ ringtest_0.x4.net4 9.08e-20
C457 ringtest_0.x4.net2 a_21507_9686# 0.00492f
C458 muxtest_0.x1.x5.GN a_19666_31955# 3.51e-19
C459 a_21509_4790# a_22295_3867# 8.97e-21
C460 a_24329_6640# ringtest_0.x4._15_ 3.85e-20
C461 ringtest_0.x4.net3 a_21675_4790# 0.00115f
C462 ringtest_0.x4._14_ ringtest_0.x4._02_ 0.166596f
C463 muxtest_0.x1.x3.GP1 ui_in[2] 5.64e-19
C464 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GP1 6.21e-20
C465 ringtest_0.x4._16_ a_22775_5878# 4.87e-20
C466 a_16579_11759# ringtest_0.x3.x2.GP3 0.00144f
C467 ringtest_0.x4.net9 ringtest_0.x4._22_ 0.369389f
C468 ui_in[4] ua[2] 0.936267f
C469 a_13501_23906# ui_in[4] 0.125445f
C470 muxtest_0.x2.x1.nSEL0 a_12297_23648# 0.03096f
C471 a_21951_5878# a_21399_5340# 5.5e-20
C472 muxtest_0.x1.x1.nSEL0 ui_in[0] 0.325407f
C473 a_22939_4584# VDPWR 3.83e-21
C474 a_24699_6200# ringtest_0.x4._06_ 0.003245f
C475 ringtest_0.x4._16_ a_23399_3867# 3.59e-21
C476 a_27169_6641# VDPWR 0.285967f
C477 a_21981_9142# VDPWR 0.210607f
C478 ringtest_0.x4._11_ a_22733_6244# 0.002344f
C479 a_22111_10993# VDPWR 0.305606f
C480 ringtest_0.x4.clknet_1_1__leaf_clk a_22765_5308# 1.5e-19
C481 ringtest_0.x4.net4 a_22817_6146# 7.5e-19
C482 ringtest_0.x4.net7 ringtest_0.x4._22_ 0.179589f
C483 muxtest_0.x2.x2.GP3 ua[0] 0.050476f
C484 muxtest_0.x1.x3.GP2 muxtest_0.R5R6 0.312699f
C485 ringtest_0.x4.net3 a_21785_5878# 1.48e-19
C486 a_21465_8830# ringtest_0.x4._01_ 1.56e-19
C487 ringtest_0.x4._15_ a_25364_5878# 0.047247f
C488 ringtest_0.x3.nselect2 VDPWR 1.23654f
C489 ringtest_0.x4.net6 ringtest_0.x4._21_ 0.083542f
C490 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B a_17377_14114# 0.110771f
C491 a_21845_8816# a_22052_8875# 0.260055f
C492 a_21561_8830# a_21981_8976# 0.036838f
C493 ringtest_0.x4._17_ a_23837_5878# 0.060488f
C494 ringtest_0.x4._17_ ringtest_0.x4._22_ 1.76e-19
C495 a_22390_4566# a_22486_4246# 0.002032f
C496 ringtest_0.x4._23_ a_26721_4246# 0.038842f
C497 ringtest_0.x4._11_ a_26201_4790# 0.012822f
C498 ringtest_0.x4.clknet_1_0__leaf_clk a_22201_9142# 0.002297f
C499 ringtest_0.x3.x2.GP1 ringtest_0.counter3 5.62e-21
C500 a_11845_23906# m2_11882_23495# 0.01297f
C501 ringtest_0.x4._14_ a_22116_4902# 1.1e-19
C502 a_27169_6641# ringtest_0.x4._25_ 0.227897f
C503 muxtest_0.x1.x3.GP2 VDPWR 3.26769f
C504 a_26367_4790# a_26721_4246# 1.65e-19
C505 a_21981_9142# a_21803_9508# 9.73e-19
C506 ringtest_0.x4._18_ ringtest_0.x4.net8 0.01511f
C507 a_21852_9416# ringtest_0.x4.clknet_1_0__leaf_clk 0.470509f
C508 a_22052_9116# a_22228_9508# 0.007724f
C509 a_21845_9116# a_22399_9142# 0.062224f
C510 ringtest_0.x4.net2 a_21852_8720# 8.79e-19
C511 ringtest_0.counter7 ringtest_0.x4.net8 6.32e-19
C512 ringtest_0.x4.net7 a_23619_6788# 5.91e-19
C513 ringtest_0.x4._11_ a_22457_5156# 0.002515f
C514 a_24070_5852# a_23809_4790# 7.94e-19
C515 ringtest_0.x4.net1 a_21981_9142# 0.002441f
C516 ringtest_0.drv_out ringtest_0.x3.x2.GN1 3.11e-19
C517 a_24361_5340# a_24527_5340# 0.961627f
C518 ringtest_0.x4._17_ a_23619_6788# 7.93e-19
C519 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP3 2.86851f
C520 a_22111_10993# ringtest_0.x4.net1 0.10983f
C521 ringtest_0.x4.net9 a_25225_5334# 0.002503f
C522 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ui_in[4] 0.008686f
C523 a_23932_6128# VDPWR 0.011201f
C524 a_25761_5058# a_26201_4790# 0.001745f
C525 ringtest_0.x4.clknet_0_clk a_24361_5340# 0.009291f
C526 ringtest_0.x4._15_ a_24317_4942# 2.8e-19
C527 a_23879_6940# ringtest_0.x4.net6 8.49e-19
C528 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.025028f
C529 ua[0] ui_in[6] 0.619336f
C530 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 1.99e-20
C531 a_23949_6654# ringtest_0.x4._20_ 1.63e-20
C532 a_23809_4790# a_23891_4790# 0.005167f
C533 a_22817_6146# a_23837_5878# 3.28e-20
C534 ringtest_0.x4._04_ ringtest_0.x4._14_ 4.63e-22
C535 a_22649_6244# a_22775_5878# 0.006169f
C536 a_21395_6940# ringtest_0.x4.clknet_0_clk 0.317755f
C537 a_15575_12017# ui_in[4] 0.02803f
C538 ringtest_0.x4.net8 a_24763_6143# 0.003744f
C539 ringtest_0.x4._24_ a_26201_5340# 0.031818f
C540 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A a_16755_12091# 9.97e-21
C541 ringtest_0.x3.x1.nSEL1 a_16027_11759# 0.073392f
C542 a_21948_5156# a_21863_4790# 0.037333f
C543 a_21675_4790# a_22457_5156# 3.14e-19
C544 ringtest_0.x4.net7 a_25225_5334# 0.054488f
C545 a_22265_5308# a_22021_4220# 2.52e-20
C546 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._14_ 0.088295f
C547 ringtest_0.x4._12_ a_21395_6940# 4.42e-19
C548 muxtest_0.R7R8 muxtest_0.R3R4 5.65992f
C549 ringtest_0.x4.net3 ringtest_0.counter3 6.21e-20
C550 a_12473_23980# VDPWR 0.193262f
C551 ringtest_0.x4._17_ a_25225_5334# 8.73e-21
C552 ringtest_0.x4.clknet_1_0__leaf_clk a_22319_6244# 4.17e-19
C553 a_21465_8830# a_21785_8054# 3.66e-19
C554 a_21132_8918# ringtest_0.x4._12_ 0.001776f
C555 a_21852_8720# a_22399_8976# 0.099725f
C556 a_22052_8875# a_22201_8964# 0.005525f
C557 muxtest_0.x1.x3.GN4 ua[3] 0.014367f
C558 ringtest_0.x4.net5 VDPWR 0.910107f
C559 ringtest_0.x3.x2.GP3 m3_17032_8096# 0.002824f
C560 ringtest_0.x4.net9 a_26640_5156# 0.023502f
C561 a_12977_24040# ui_in[3] 0.001558f
C562 a_24895_5334# VDPWR 0.004219f
C563 ringtest_0.x4.net2 a_22399_8976# 1.01e-21
C564 muxtest_0.x2.x2.GN2 ui_in[3] 0.11443f
C565 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net8 0.073766f
C566 muxtest_0.x1.x3.GN4 a_20492_32319# 0.001562f
C567 ringtest_0.x4._15_ a_26913_4566# 0.001637f
C568 a_21233_5340# ringtest_0.x4._03_ 0.001727f
C569 ringtest_0.x4._02_ a_21509_4790# 3.71e-19
C570 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP3 0.075682f
C571 muxtest_0.R2R3 ua[0] 2.39e-19
C572 a_24004_6128# ringtest_0.x4._20_ 4.3e-20
C573 ringtest_0.counter7 ringtest_0.x4.counter[1] 0.003115f
C574 a_19842_32287# muxtest_0.x1.x3.GN4 0.003645f
C575 ringtest_0.x4._00_ a_21845_9116# 0.118744f
C576 ringtest_0.x4._24_ a_27233_5058# 0.009415f
C577 ringtest_0.x4._11_ ringtest_0.x4._03_ 0.00174f
C578 ringtest_0.x4.net7 a_26640_5156# 4.39e-19
C579 ringtest_0.x4._19_ ringtest_0.x4._15_ 6.2e-22
C580 ringtest_0.x4._02_ a_22765_5308# 7.66e-20
C581 ringtest_0.x4.net5 a_23467_4584# 0.001706f
C582 ringtest_0.x4.clknet_1_0__leaf_clk a_22043_5156# 5.04e-19
C583 ringtest_0.counter7 ringtest_0.x4.net11 1.31e-19
C584 ringtest_0.x4.clknet_1_1__leaf_clk a_24729_4790# 0.319108f
C585 ringtest_0.x4._18_ ringtest_0.x4._05_ 1.11e-19
C586 ringtest_0.x4.net10 a_27273_4220# 0.104575f
C587 ringtest_0.x4.net8 a_24800_5334# 0.003635f
C588 ringtest_0.x4._20_ a_23963_4790# 0.001506f
C589 muxtest_0.x1.x3.GN2 ui_in[0] 0.114399f
C590 ringtest_0.x4._11_ a_23770_5308# 0.058411f
C591 a_21007_3867# VDPWR 0.251327f
C592 ringtest_0.x3.x2.GN4 ui_in[4] 0.059808f
C593 a_16027_11759# ringtest_0.x3.x2.GN3 6.68e-19
C594 ringtest_0.x4._08_ a_24527_5340# 8.29e-20
C595 ringtest_0.x4._13_ ringtest_0.x4._02_ 0.053355f
C596 a_16203_12091# ringtest_0.x3.x2.GN1 1.46e-19
C597 a_23381_4818# ringtest_0.x4._20_ 3.41e-19
C598 ringtest_0.x4.net4 ringtest_0.x4._14_ 0.209869f
C599 ringtest_0.x4._11_ a_21939_8054# 2.12e-19
C600 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x1.nSEL0 1.14e-19
C601 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.173286f
C602 ringtest_0.x4._15_ a_22265_5308# 1.37e-19
C603 ringtest_0.x4.net6 a_24968_5308# 0.012704f
C604 ringtest_0.x4._03_ a_21675_4790# 0.260627f
C605 muxtest_0.x1.x4.A ui_in[4] 0.045433f
C606 a_21509_4790# a_22116_4902# 0.141453f
C607 ringtest_0.x4._22_ a_26627_4246# 0.140356f
C608 a_24800_5334# a_24729_4790# 2.14e-19
C609 a_24968_5308# a_24895_4790# 0.001607f
C610 a_24361_5340# a_25168_5156# 4.58e-19
C611 a_24527_5340# a_25336_4902# 6.74e-19
C612 ringtest_0.x4._15_ ringtest_0.x4.net9 0.08758f
C613 muxtest_0.R3R4 VDPWR 3.2635f
C614 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._10_ 0.006812f
C615 ringtest_0.x4._16_ a_25083_4790# 1.98e-21
C616 ringtest_0.x4._23_ ringtest_0.x4.net8 0.011201f
C617 ringtest_0.x4._05_ a_24763_6143# 2.43e-19
C618 a_22265_5308# a_22541_5058# 0.007214f
C619 a_22097_5334# a_21948_5156# 0.001152f
C620 ringtest_0.x4.net8 a_26367_4790# 1.04e-19
C621 ringtest_0.x4.clknet_0_clk a_25336_4902# 8.09e-19
C622 ringtest_0.x4._16_ a_21948_5156# 2.79e-19
C623 ringtest_0.x4._21_ ringtest_0.x4.net5 2.83e-22
C624 a_23770_5308# a_23899_5654# 0.010132f
C625 a_26201_5340# a_27233_5308# 0.048748f
C626 a_21840_5308# a_22181_5334# 9.73e-19
C627 a_26367_5340# a_26640_5334# 0.078545f
C628 a_21672_5334# a_21767_5334# 0.007724f
C629 a_24527_5340# VDPWR 0.297793f
C630 ringtest_0.x4.clknet_1_1__leaf_clk a_26749_6422# 3.65e-19
C631 ringtest_0.x4.net6 a_25925_6788# 0.157729f
C632 ringtest_0.x4.net7 ringtest_0.x4._15_ 0.590844f
C633 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net11 1.82e-20
C634 VDPWR ui_in[5] 0.25433f
C635 ringtest_0.x4._04_ a_21509_4790# 2.08e-19
C636 a_21785_5878# ringtest_0.x4._03_ 4.31e-20
C637 ringtest_0.x4._23_ a_24729_4790# 3.56e-21
C638 ringtest_0.x4.net7 a_25263_5156# 5.23e-19
C639 ringtest_0.x4._17_ ringtest_0.x4._15_ 0.083602f
C640 a_13025_23980# muxtest_0.x2.x2.GP1 2.87e-20
C641 ringtest_0.x4._05_ ringtest_0.x4.clknet_1_1__leaf_clk 0.143201f
C642 ringtest_0.x4.clknet_0_clk VDPWR 2.50725f
C643 muxtest_0.x2.x2.GP2 ui_in[4] 4.34e-19
C644 ringtest_0.x4.clknet_1_0__leaf_clk a_21509_4790# 0.293401f
C645 a_24729_4790# a_26367_4790# 8.05e-21
C646 ua[3] ua[4] 0.008019f
C647 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP1 8.08e-19
C648 ringtest_0.counter7 ringtest_0.x4._09_ 5.27e-21
C649 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 5.48e-19
C650 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y 0.001676f
C651 muxtest_0.x2.x1.nSEL1 a_12019_24012# 0.00175f
C652 a_12473_23980# a_12849_23648# 3.02e-19
C653 ringtest_0.x4._12_ VDPWR 0.293048f
C654 ringtest_0.x4._04_ a_22765_5308# 0.171873f
C655 a_27191_5712# ringtest_0.x4._09_ 1.66e-19
C656 ringtest_0.x4.net10 a_26201_4790# 0.001924f
C657 ringtest_0.x4.counter[9] ua[0] 0.004138f
C658 ringtest_0.x4.net7 a_24926_5712# 2.79e-19
C659 ringtest_0.x4.clknet_1_0__leaf_clk a_22765_5308# 1.95e-19
C660 a_27233_5308# a_27233_5058# 0.026048f
C661 ringtest_0.x4._05_ a_24800_5334# 6.05e-21
C662 ringtest_0.x4.net6 a_21233_5340# 1.88e-19
C663 ringtest_0.x4.clknet_1_0__leaf_clk a_21867_8054# 2.61e-19
C664 a_26555_5334# ringtest_0.x4.net10 6.3e-20
C665 ringtest_0.x4._13_ ringtest_0.x4._04_ 1.41e-19
C666 ringtest_0.x4.net1 ui_in[5] 0.067291f
C667 muxtest_0.x2.x1.nSEL0 VDPWR 0.523833f
C668 ringtest_0.x4._22_ a_25294_4790# 6.82e-19
C669 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._13_ 0.02176f
C670 muxtest_0.x1.x3.GN3 muxtest_0.x1.x5.A 0.429924f
C671 ringtest_0.x4._11_ ringtest_0.x4.net6 2.01574f
C672 ringtest_0.x4.counter[6] ua[1] 3.21e-19
C673 ringtest_0.x3.x2.GN1 m3_17036_9140# 6.03e-20
C674 ringtest_0.x4.net8 a_25593_5156# 0.007067f
C675 ringtest_0.x4.net7 a_26173_4612# 6.49e-19
C676 ringtest_0.x4.net1 ringtest_0.x4._12_ 0.312817f
C677 ringtest_0.x4._11_ a_24895_4790# 0.042209f
C678 ringtest_0.x4._23_ a_26749_6422# 0.007723f
C679 ringtest_0.x4._23_ ringtest_0.x4.net11 0.257634f
C680 a_26640_5156# a_26627_4246# 2.47e-19
C681 a_19114_31955# muxtest_0.x1.x3.GN3 6.68e-19
C682 a_21233_5340# a_21055_5334# 5.87e-19
C683 a_26749_6422# a_26367_4790# 3.03e-21
C684 muxtest_0.R4R5 ui_in[2] 6.76e-20
C685 a_18662_32213# VDPWR 0.213938f
C686 a_22224_6244# a_22373_5156# 1.06e-19
C687 a_26808_4902# a_26766_4790# 4.62e-19
C688 a_26367_4790# ringtest_0.x4.net11 2.58e-19
C689 ringtest_0.x4._05_ ringtest_0.x4._23_ 9.36e-20
C690 a_21399_5340# a_21672_5334# 0.078737f
C691 ringtest_0.x4.net4 a_21509_4790# 0.008383f
C692 ringtest_0.x4.net10 a_27303_4246# 0.001384f
C693 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._09_ 0.003413f
C694 ringtest_0.x4.net6 a_25761_5058# 3.96e-21
C695 m2_18699_31802# VDPWR 0.140918f
C696 a_13501_23906# muxtest_0.x2.x2.GN4 0.134079f
C697 muxtest_0.x2.x2.GN4 ua[2] 0.446579f
C698 a_25364_5878# a_26367_5340# 0.008007f
C699 ringtest_0.x4._21_ a_24527_5340# 0.002388f
C700 muxtest_0.x2.x2.GN2 a_12425_24040# 0.002418f
C701 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN2 0.065156f
C702 a_23949_6654# a_24329_6640# 0.048635f
C703 a_22245_8054# VDPWR 0.291372f
C704 a_24729_4790# a_25593_5156# 0.032244f
C705 a_25336_4902# a_25168_5156# 0.239923f
C706 a_24895_4790# a_25761_5058# 0.034054f
C707 a_19666_31955# ui_in[0] 0.086357f
C708 muxtest_0.x2.x1.nSEL1 ui_in[4] 0.275874f
C709 ringtest_0.x4.net4 a_22765_5308# 0.005124f
C710 ringtest_0.x4.clknet_0_clk ringtest_0.x4._21_ 4.86e-19
C711 muxtest_0.x1.x3.GP3 muxtest_0.R1R2 4.25867f
C712 ringtest_0.x3.x1.nSEL0 a_16155_12151# 2.51e-19
C713 ringtest_0.x4._15_ a_27065_5334# 2.78e-19
C714 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN1 0.004375f
C715 ringtest_0.x4._22_ a_26721_4246# 0.063386f
C716 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 5.04e-19
C717 ringtest_0.x4._14_ a_22021_4220# 0.134293f
C718 ringtest_0.x4._04_ ringtest_0.x4.net8 7.52e-21
C719 muxtest_0.x1.x3.GP1 muxtest_0.R2R3 0.127193f
C720 a_25168_5156# VDPWR 0.254209f
C721 a_21007_3867# a_21375_3867# 2.48e-19
C722 ringtest_0.x4.net8 a_25441_4612# 0.001229f
C723 ringtest_0.x4._18_ a_24361_5340# 5.99e-21
C724 ringtest_0.x4._11_ a_22939_4584# 8.14e-19
C725 ringtest_0.x4.net4 ringtest_0.x4._13_ 0.050083f
C726 muxtest_0.x1.x3.GP1 ui_in[1] 8.43e-19
C727 a_23879_6940# a_24527_5340# 4.98e-20
C728 muxtest_0.x1.x3.GP2 muxtest_0.x1.x5.A 0.350698f
C729 a_20318_32213# ui_in[1] 0.125445f
C730 a_24336_6544# ringtest_0.x4._06_ 1.63e-21
C731 ringtest_0.x4.net3 a_21465_8830# 0.115857f
C732 a_24527_5340# a_25309_5334# 3.14e-19
C733 ringtest_0.x4.net1 a_22245_8054# 4.64e-19
C734 a_25225_5334# a_25351_5712# 0.006169f
C735 ringtest_0.x4.clknet_0_clk a_23349_6422# 2.32e-20
C736 a_21425_9686# ringtest_0.x4._12_ 1.27e-21
C737 ringtest_0.x4.net6 a_21785_5878# 0.006287f
C738 a_21852_9416# a_21561_8830# 1.53e-19
C739 a_21561_9116# a_21845_8816# 9.64e-20
C740 a_24329_6640# a_24004_6128# 0.001895f
C741 ringtest_0.x4.clknet_0_clk a_23879_6940# 1.74729f
C742 a_22983_5654# VDPWR 0.001282f
C743 ringtest_0.x4._15_ a_26627_4246# 0.087822f
C744 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP1 0.041018f
C745 ringtest_0.x4._19_ a_24685_6788# 2.79e-19
C746 ringtest_0.x4.net10 ringtest_0.x4.counter[8] 0.009948f
C747 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN3 4.01e-20
C748 ringtest_0.x4.net2 a_21465_9294# 0.092265f
C749 ringtest_0.drv_out ui_in[4] 1.17e-19
C750 ringtest_0.x4._23_ ringtest_0.x4._09_ 0.130147f
C751 muxtest_0.x1.x5.GN a_20318_32213# 1.19e-19
C752 ringtest_0.ring_out a_16579_11759# 5.47e-20
C753 a_26201_4790# a_26808_4902# 0.141453f
C754 a_24536_6699# ringtest_0.x4._15_ 1.61e-21
C755 ringtest_0.x4._09_ a_26367_4790# 0.413296f
C756 ui_in[6] ui_in[7] 0.03107f
C757 ringtest_0.x4.net3 a_21948_5156# 3.32e-20
C758 a_24763_6143# a_24361_5340# 0.004179f
C759 ringtest_0.x4._16_ ringtest_0.x4._07_ 0.003808f
C760 a_13675_24012# ui_in[4] 8.84e-19
C761 ringtest_0.x4._06_ a_24986_5878# 6.53e-20
C762 muxtest_0.x2.x2.GN3 ui_in[4] 0.273874f
C763 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y 0.174714f
C764 a_21591_6128# VDPWR 0.006535f
C765 ringtest_0.x4._23_ a_26766_5712# 9.59e-19
C766 muxtest_0.x2.x1.nSEL0 a_12849_23648# 1.91e-20
C767 a_24004_6128# a_24545_5878# 4.72e-19
C768 a_21951_5878# a_21672_5334# 0.001124f
C769 ringtest_0.x4.clknet_1_0__leaf_clk a_21798_5712# 0.001807f
C770 a_22486_4246# VDPWR 0.011874f
C771 a_22228_9508# VDPWR 0.005789f
C772 ringtest_0.x4.net9 a_25975_3867# 7.77e-19
C773 ringtest_0.x4._11_ a_23932_6128# 0.002546f
C774 ringtest_0.x4.clknet_1_1__leaf_clk a_24361_5340# 0.670964f
C775 ringtest_0.x4._15_ ringtest_0.x4._14_ 1.65e-19
C776 ringtest_0.x4.net4 ringtest_0.x4.net8 0.001699f
C777 a_21852_8720# a_21981_8976# 0.124967f
C778 ringtest_0.x4._24_ a_26895_3867# 0.00116f
C779 a_21845_8816# ringtest_0.x4._01_ 0.092611f
C780 muxtest_0.x2.x2.GP1 ui_in[3] 9.65e-19
C781 ringtest_0.counter3 ringtest_0.x4.net6 1.1e-21
C782 ringtest_0.x4._23_ a_27659_4246# 0.009249f
C783 muxtest_0.x1.x3.GN1 muxtest_0.R6R7 0.254376f
C784 a_25977_4220# a_26269_4612# 0.001675f
C785 ringtest_0.x4.net7 a_25975_3867# 4.41e-19
C786 ringtest_0.x4._14_ a_22541_5058# 1.14e-20
C787 a_26640_5156# a_26721_4246# 7.6e-20
C788 a_12297_23648# ui_in[3] 0.246189f
C789 ringtest_0.x4.net2 a_21981_8976# 8.2e-21
C790 a_21981_9142# a_22399_9142# 3.39e-19
C791 a_22052_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.040993f
C792 ringtest_0.x4.net7 a_24685_6788# 0.002551f
C793 ringtest_0.x4._11_ ringtest_0.x4.net5 0.388184f
C794 ringtest_0.drv_out ringtest_0.x3.x2.GP1 0.125793f
C795 a_24004_6128# a_24317_4942# 2.49e-20
C796 ringtest_0.x4.net1 a_22228_9508# 4.16e-19
C797 a_24527_5340# a_24968_5308# 0.110715f
C798 a_24361_5340# a_24800_5334# 0.260055f
C799 ringtest_0.x4._06_ a_23899_5334# 2.02e-19
C800 a_24070_5852# a_23899_5334# 1.06e-19
C801 ringtest_0.x4.net9 a_26367_5340# 0.001054f
C802 ringtest_0.counter3 a_21055_5334# 1.26e-20
C803 a_25593_5156# ringtest_0.x4._09_ 1.4e-19
C804 ringtest_0.x4._08_ a_27191_5712# 7.43e-19
C805 a_23949_6654# ringtest_0.x4._19_ 0.065395f
C806 ringtest_0.x4.clknet_0_clk a_24968_5308# 3.18e-19
C807 a_21509_4790# a_22021_4220# 2.64e-19
C808 ringtest_0.x4.net4 a_21798_5712# 1.81e-19
C809 a_12977_24040# ua[3] 1.48e-19
C810 ringtest_0.x4._15_ a_25351_5712# 0.00162f
C811 ringtest_0.x4.net6 ringtest_0.x4.net10 1.08e-19
C812 muxtest_0.x2.x2.GN2 ua[3] 0.234749f
C813 ringtest_0.x4.net8 a_23837_5878# 0.057781f
C814 a_16203_12091# ui_in[4] 0.254026f
C815 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN4 0.011047f
C816 ringtest_0.x4._24_ a_26808_5308# 0.015657f
C817 ringtest_0.x4.net8 ringtest_0.x4._22_ 0.137056f
C818 ringtest_0.x3.x1.nSEL1 a_16579_11759# 7.84e-19
C819 a_22116_4902# a_22074_4790# 4.62e-19
C820 a_21675_4790# ringtest_0.x4.net5 8.3e-19
C821 ringtest_0.x4.net7 a_26367_5340# 2.99e-20
C822 ringtest_0.x4._23_ a_24361_5340# 1.94e-21
C823 a_21675_10006# VDPWR 3.05e-19
C824 ringtest_0.x4._04_ a_22350_5878# 2.91e-19
C825 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.173286f
C826 muxtest_0.x1.x5.A muxtest_0.R3R4 4.07e-21
C827 a_21951_5878# a_22224_6244# 0.074434f
C828 ringtest_0.x4._16_ a_22164_4362# 0.146025f
C829 ringtest_0.x4.net4 ringtest_0.x4.counter[1] 3.68e-19
C830 muxtest_0.x1.x3.GN3 a_13501_23906# 1.84e-20
C831 ringtest_0.x4._18_ VDPWR 0.671209f
C832 a_13025_23980# VDPWR 0.261817f
C833 ringtest_0.x4.clknet_1_0__leaf_clk a_22350_5878# 3.26e-19
C834 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[3] 2.42e-19
C835 a_21981_8976# a_22399_8976# 3.39e-19
C836 ringtest_0.x4.net6 a_22775_5878# 5.88e-19
C837 ringtest_0.counter7 VDPWR 2.38177f
C838 a_21845_8816# a_21785_8054# 4.35e-19
C839 ringtest_0.x4.clknet_0_clk a_25925_6788# 1.5e-19
C840 ringtest_0.x4.net6 a_24627_6200# 4.57e-19
C841 ringtest_0.x4.net9 a_27065_5156# 0.020729f
C842 muxtest_0.x2.x2.GN4 m3_13302_19985# 7.07e-19
C843 ringtest_0.x4.net6 ringtest_0.x4.counter[4] 0.003133f
C844 ringtest_0.x4.net4 a_22390_4566# 0.01239f
C845 a_23529_6422# ringtest_0.x4._16_ 1.86e-20
C846 a_27191_5712# VDPWR 7.83e-19
C847 ringtest_0.x4._22_ a_24729_4790# 0.019806f
C848 ringtest_0.x4.net6 a_23399_3867# 3.58e-19
C849 ringtest_0.x4._15_ a_26721_4246# 0.038186f
C850 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._08_ 0.00277f
C851 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN4 0.141966f
C852 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GN3 0.175252f
C853 a_18836_32319# VDPWR 0.001273f
C854 ringtest_0.x4._00_ a_21981_9142# 0.005564f
C855 ringtest_0.x4._24_ a_26555_4790# 3.3e-19
C856 a_21785_5878# ringtest_0.x4.net5 1.51e-20
C857 ringtest_0.x4.net7 a_27065_5156# 1.49e-19
C858 a_22111_10993# ringtest_0.x4._00_ 4.57e-22
C859 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP2 8.45e-19
C860 ringtest_0.x4.net1 a_21675_10006# 0.003019f
C861 a_24763_6143# VDPWR 0.129618f
C862 a_23949_6654# ringtest_0.x4.net7 0.114197f
C863 ringtest_0.x4.clknet_1_1__leaf_clk a_25336_4902# 0.046669f
C864 ringtest_0.x4.net8 a_25225_5334# 0.00311f
C865 ringtest_0.x4._11_ a_24527_5340# 8.46e-20
C866 ringtest_0.x3.x2.GN1 ua[1] 0.430121f
C867 a_22139_5878# a_21399_5340# 2.83e-19
C868 a_22295_3867# VDPWR 0.312095f
C869 ringtest_0.x4._17_ a_23949_6654# 0.0702f
C870 a_16203_12091# ringtest_0.x3.x2.GP1 2.33e-21
C871 ringtest_0.x4._06_ ringtest_0.x4._16_ 0.064563f
C872 muxtest_0.x2.x1.nSEL1 a_11845_23906# 0.193944f
C873 ringtest_0.x4._08_ a_24800_5334# 1.22e-20
C874 a_16579_11759# ringtest_0.x3.x2.GN3 0.104151f
C875 a_24317_4942# ringtest_0.x4._20_ 0.113204f
C876 a_16755_12091# ringtest_0.x3.x2.GN1 3.78e-20
C877 a_24070_5852# ringtest_0.x4._16_ 0.035189f
C878 ringtest_0.x4._11_ ringtest_0.x4.clknet_0_clk 0.042991f
C879 a_21509_4790# a_22541_5058# 0.048748f
C880 ringtest_0.x4.net6 a_25393_5308# 0.002597f
C881 ringtest_0.x4._03_ a_21948_5156# 0.010537f
C882 ringtest_0.x4._15_ a_22765_5308# 8.84e-19
C883 muxtest_0.x1.x3.GP2 a_13501_23906# 6.46e-20
C884 ringtest_0.x4.clknet_1_1__leaf_clk VDPWR 3.30823f
C885 ringtest_0.x3.x2.GP2 VDPWR 1.81711f
C886 ringtest_0.x4._12_ ringtest_0.x4._11_ 0.214271f
C887 a_22399_8976# a_22228_8598# 0.001229f
C888 a_25393_5308# a_24895_4790# 0.002689f
C889 a_25225_5334# a_24729_4790# 0.004606f
C890 ringtest_0.x4._22_ ringtest_0.x4.net11 1.96e-19
C891 muxtest_0.x1.x3.GP3 muxtest_0.R6R7 0.12263f
C892 a_26569_6422# a_25364_5878# 0.010673f
C893 ringtest_0.x4._16_ a_23891_4790# 0.00109f
C894 ringtest_0.x4._05_ ringtest_0.x4._22_ 0.001519f
C895 a_22765_5308# a_22541_5058# 0.002391f
C896 a_22097_5334# a_22373_5156# 5.06e-19
C897 ringtest_0.x4.net7 a_24004_6128# 3.79e-19
C898 ringtest_0.x4._23_ ringtest_0.x4._08_ 0.030554f
C899 ringtest_0.x4._18_ ringtest_0.x4._21_ 0.005609f
C900 ringtest_0.x4._16_ a_22373_5156# 6.21e-20
C901 muxtest_0.x2.x1.nSEL0 m2_11882_23495# 3.43e-19
C902 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP2 3.78674f
C903 a_26367_5340# a_27065_5334# 0.194892f
C904 ringtest_0.x4._17_ a_24004_6128# 0.076419f
C905 ringtest_0.counter7 ringtest_0.x4.counter[2] 0.003115f
C906 a_26808_5308# a_27233_5308# 1.28e-19
C907 ringtest_0.x4._08_ a_26367_4790# 0.001269f
C908 ringtest_0.counter3 ringtest_0.x4.net5 0.082815f
C909 ringtest_0.ring_out ringtest_0.x3.x2.GP3 0.080819f
C910 a_24800_5334# VDPWR 0.25486f
C911 a_24465_6800# a_24264_6788# 4.67e-20
C912 a_24536_6699# a_24685_6788# 0.005525f
C913 a_24336_6544# a_24883_6800# 0.095025f
C914 muxtest_0.R7R8 ui_in[3] 0.025566f
C915 a_21425_9686# a_21675_10006# 0.007234f
C916 ringtest_0.x4.net4 a_22074_4790# 6.57e-19
C917 a_18662_32213# a_19114_31955# 0.002207f
C918 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP1 1.5157f
C919 a_12297_23648# a_12425_24040# 0.004764f
C920 a_23349_6422# ringtest_0.x4._18_ 0.09549f
C921 a_12849_23648# a_13025_23980# 0.185422f
C922 a_12297_23648# muxtest_0.x2.x2.GN1 0.012445f
C923 ringtest_0.x4._21_ a_24763_6143# 1.69e-19
C924 ringtest_0.x4._17_ a_23381_4818# 6.88e-22
C925 ringtest_0.x3.x1.nSEL0 ui_in[4] 0.137394f
C926 ringtest_0.x4._23_ VDPWR 1.67531f
C927 a_27065_5334# a_27065_5156# 0.01464f
C928 muxtest_0.R4R5 muxtest_0.R2R3 7.85e-20
C929 a_21395_6940# ringtest_0.x4._04_ 0.00168f
C930 a_22817_6146# a_24004_6128# 1.25e-19
C931 a_22295_3867# ringtest_0.x4.counter[2] 0.1107f
C932 a_22245_8054# ringtest_0.x4._11_ 0.201886f
C933 a_26367_4790# VDPWR 0.308998f
C934 a_21951_5878# a_22139_5878# 0.095025f
C935 ringtest_0.counter3 a_21007_3867# 2.11e-19
C936 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C937 a_16707_12151# VDPWR 0.001127f
C938 ringtest_0.x4.clknet_1_0__leaf_clk a_21395_6940# 1.67275f
C939 ringtest_0.x3.x2.GN2 VDPWR 0.602894f
C940 ringtest_0.x4._22_ ringtest_0.x4._09_ 0.009594f
C941 muxtest_0.x2.x2.GN4 ua[0] 0.046938f
C942 ringtest_0.x3.x2.GP1 m3_17036_9140# 5.81e-19
C943 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._21_ 0.038033f
C944 ringtest_0.x4._15_ ringtest_0.x4.net8 0.048599f
C945 ringtest_0.x3.x2.GN3 m3_17032_8096# 0.087318f
C946 ringtest_0.x4.net2 ringtest_0.x4.counter[0] 0.010591f
C947 ringtest_0.x4._24_ a_26817_4566# 9.33e-19
C948 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP3 5.60415f
C949 muxtest_0.x1.x3.GN3 muxtest_0.x1.x4.A 0.429865f
C950 ringtest_0.x4.net9 ringtest_0.x4._20_ 1.35e-20
C951 a_23879_6940# a_24763_6143# 1.03e-20
C952 ringtest_0.x4.net3 a_22164_4362# 8.22e-19
C953 ringtest_0.x4.net7 a_26375_4612# 6.33e-20
C954 a_22021_4220# a_22390_4566# 0.046138f
C955 ringtest_0.x4._11_ a_25168_5156# 0.026293f
C956 ringtest_0.x4.net5 ringtest_0.x4.counter[4] 0.001223f
C957 ringtest_0.x4._23_ ringtest_0.x4._25_ 0.0063f
C958 a_27233_5058# a_27273_4220# 0.005283f
C959 a_27065_5156# a_26627_4246# 2.58e-19
C960 a_19666_31955# muxtest_0.x1.x3.GN3 0.104183f
C961 ringtest_0.counter7 a_21375_3867# 2.81e-20
C962 ringtest_0.x4.net5 a_23399_3867# 0.233889f
C963 a_21675_9686# a_21561_9116# 1.96e-19
C964 a_27065_5156# a_27149_5156# 0.008508f
C965 a_22649_6244# a_22373_5156# 2.6e-20
C966 a_19290_32287# VDPWR 0.194389f
C967 a_25421_6641# ringtest_0.x4._24_ 1.86e-20
C968 ringtest_0.x4._02_ VDPWR 0.323624f
C969 a_21399_5340# a_22097_5334# 0.196846f
C970 a_21840_5308# a_22265_5308# 1.28e-19
C971 muxtest_0.x1.x1.nSEL0 a_18662_32213# 0.081627f
C972 muxtest_0.x2.x2.GN4 a_13675_24012# 0.001562f
C973 ringtest_0.x4._15_ a_24729_4790# 4.49e-20
C974 ringtest_0.x4.net8 a_24926_5712# 4.88e-19
C975 m2_15612_11606# VDPWR 0.14037f
C976 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GN4 0.071281f
C977 ringtest_0.x4.net6 a_25083_4790# 0.00565f
C978 ringtest_0.x4.net7 ringtest_0.x4._20_ 0.035834f
C979 ringtest_0.x4._16_ a_21399_5340# 8.97e-20
C980 a_25364_5878# a_26640_5334# 0.01166f
C981 muxtest_0.x1.x3.GP1 ui_in[0] 8.18e-19
C982 VDPWR ui_in[3] 6.03016f
C983 a_24045_6654# a_24336_6544# 0.192261f
C984 a_24729_4790# a_25263_5156# 0.002698f
C985 a_25336_4902# a_25593_5156# 0.036838f
C986 a_23879_6940# ringtest_0.x4.clknet_1_1__leaf_clk 0.002451f
C987 a_24895_4790# a_25083_4790# 0.095025f
C988 muxtest_0.x1.x1.nSEL0 m2_18699_31802# 3.43e-19
C989 a_20318_32213# ui_in[0] 0.220425f
C990 ringtest_0.x4._17_ ringtest_0.x4._20_ 1.89e-19
C991 muxtest_0.R3R4 ua[2] 4.52137f
C992 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GP1 6.21e-20
C993 ringtest_0.x3.nselect2 ringtest_0.x3.x2.GN4 1.53e-20
C994 ui_in[2] ui_in[6] 0.264066f
C995 ringtest_0.x4.clknet_1_1__leaf_clk a_25309_5334# 0.001538f
C996 ringtest_0.x4.net6 a_24715_5334# 0.008614f
C997 muxtest_0.x1.x3.GN4 muxtest_0.R1R2 0.628977f
C998 a_26895_3867# ringtest_0.x4.counter[9] 2.34e-19
C999 ringtest_0.x4._14_ a_22765_4478# 0.112679f
C1000 a_26201_5340# a_26201_4790# 0.037572f
C1001 a_21395_6940# ringtest_0.x4.net4 4.87e-19
C1002 uio_in[4] uio_in[3] 0.031023f
C1003 ringtest_0.x4._11_ a_21591_6128# 0.002118f
C1004 ringtest_0.x4._00_ ui_in[5] 2.67e-19
C1005 a_21375_3867# a_22295_3867# 1.37e-20
C1006 a_25593_5156# VDPWR 0.185094f
C1007 a_23879_6940# a_24800_5334# 5.07e-19
C1008 muxtest_0.x1.x3.GN2 muxtest_0.R3R4 0.271818f
C1009 a_22399_9142# a_22245_8054# 9.03e-20
C1010 a_24329_6640# a_24545_5878# 2.84e-21
C1011 muxtest_0.x1.x3.GP2 muxtest_0.x1.x4.A 0.350401f
C1012 a_22116_4902# VDPWR 0.219142f
C1013 ringtest_0.x4.net3 a_21845_8816# 0.008811f
C1014 a_24465_6800# ringtest_0.x4._06_ 4.29e-19
C1015 a_26201_5340# a_26555_5334# 0.062224f
C1016 a_21587_5334# a_21767_5334# 0.001229f
C1017 a_21852_9416# a_21852_8720# 0.027204f
C1018 a_21845_9116# a_21845_8816# 0.040702f
C1019 a_24336_6544# a_24699_6200# 6.47e-19
C1020 ringtest_0.x4._00_ ringtest_0.x4._12_ 4.17e-19
C1021 a_23993_5654# VDPWR 2.25e-21
C1022 a_19666_31955# muxtest_0.x1.x3.GP2 2.46e-19
C1023 ringtest_0.x4._15_ a_22390_4566# 8.81e-20
C1024 ringtest_0.x4.net2 a_22201_9142# 1.37e-19
C1025 ringtest_0.x4._19_ a_24287_6422# 1.83e-19
C1026 ringtest_0.x4._15_ a_26749_6422# 0.001357f
C1027 ringtest_0.x4._15_ ringtest_0.x4.net11 1.7e-19
C1028 ringtest_0.x4.net7 a_26569_6422# 6.19e-19
C1029 ringtest_0.x4.net2 a_21852_9416# 4.89e-19
C1030 ui_in[1] ui_in[2] 2.795f
C1031 ringtest_0.ring_out a_17231_12017# 0.001281f
C1032 ringtest_0.x4._09_ a_26640_5156# 0.0221f
C1033 a_26201_4790# a_27233_5058# 0.048748f
C1034 ringtest_0.x4._05_ ringtest_0.x4._15_ 9.02e-20
C1035 ringtest_0.x4._17_ a_26569_6422# 0.056144f
C1036 ringtest_0.x4.net3 a_22373_5156# 1.53e-21
C1037 a_22541_5058# a_22390_4566# 0.001062f
C1038 ringtest_0.x4._22_ a_24361_5340# 0.016414f
C1039 a_24763_6143# a_24968_5308# 1.06e-19
C1040 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP3 2.86851f
C1041 muxtest_0.x2.x2.GP1 ua[3] 4.09825f
C1042 ringtest_0.x4._04_ VDPWR 0.272251f
C1043 muxtest_0.x1.x5.GN ui_in[2] 3.98638f
C1044 a_24329_6640# a_24317_4942# 8.37e-20
C1045 a_24699_6200# a_24986_5878# 3.14e-19
C1046 a_22392_5990# a_22265_5308# 0.002135f
C1047 a_21951_5878# a_22097_5334# 3.42e-19
C1048 ringtest_0.x4.clknet_0_clk a_24627_6200# 2.68e-20
C1049 ringtest_0.x4.clknet_1_0__leaf_clk a_22223_5712# 4.11e-19
C1050 a_12297_23648# ua[3] 1.21e-19
C1051 ringtest_0.x4.clknet_1_0__leaf_clk VDPWR 3.68509f
C1052 ringtest_0.x4.net9 a_27489_3702# 0.003439f
C1053 a_21951_5878# ringtest_0.x4._16_ 1.01e-19
C1054 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ui_in[4] 9.08e-20
C1055 a_24045_6654# a_23899_5334# 4.21e-21
C1056 ringtest_0.x4.clknet_1_1__leaf_clk a_24968_5308# 0.01748f
C1057 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.173286f
C1058 ringtest_0.x4.net2 ringtest_0.x4._14_ 0.45134f
C1059 a_21591_6128# a_21785_5878# 5.05e-19
C1060 a_22052_8875# ringtest_0.x4._01_ 0.004715f
C1061 ringtest_0.x4._18_ a_21233_5340# 3.08e-21
C1062 a_26640_5334# a_26735_5334# 0.007724f
C1063 a_26808_5308# a_27149_5334# 9.73e-19
C1064 a_21852_9416# a_22399_8976# 4.5e-20
C1065 ringtest_0.x4._00_ a_22245_8054# 5.19e-20
C1066 a_27233_5058# a_27303_4246# 1.25e-19
C1067 a_12849_23648# ui_in[3] 0.086353f
C1068 a_21803_9508# ringtest_0.x4.clknet_1_0__leaf_clk 7.44e-19
C1069 a_22228_9508# a_22399_9142# 0.001229f
C1070 ringtest_0.drv_out ringtest_0.x4.net6 2.01e-20
C1071 ringtest_0.x4._11_ ringtest_0.x4._18_ 0.035586f
C1072 ringtest_0.x4.net7 a_24287_6422# 6.13e-20
C1073 ringtest_0.x4._11_ ringtest_0.counter7 2.85e-19
C1074 ringtest_0.x4._17_ a_22392_5990# 2.52e-22
C1075 a_24361_5340# a_25225_5334# 0.030894f
C1076 a_21399_5340# a_21587_5334# 0.097818f
C1077 a_24527_5340# a_25393_5308# 0.034054f
C1078 ringtest_0.x4.net1 ringtest_0.x4.clknet_1_0__leaf_clk 0.561165f
C1079 a_24968_5308# a_24800_5334# 0.239923f
C1080 a_18662_32213# muxtest_0.x1.x3.GN2 0.039612f
C1081 ringtest_0.x4._15_ ringtest_0.x4._09_ 0.030214f
C1082 ringtest_0.x4._17_ a_24287_6422# 0.002375f
C1083 ringtest_0.x4.clknet_1_1__leaf_clk a_25925_6788# 0.001522f
C1084 ringtest_0.x4._21_ a_23993_5654# 4.25e-19
C1085 muxtest_0.x1.x3.GN3 ua[0] 0.007815f
C1086 a_24329_6640# ringtest_0.x4._19_ 0.074331f
C1087 ringtest_0.x4.clknet_0_clk a_25393_5308# 0.01296f
C1088 ringtest_0.x4._03_ a_22164_4362# 0.005187f
C1089 ringtest_0.x4.net4 a_22223_5712# 3.33e-19
C1090 a_24317_4942# a_24551_4790# 0.005167f
C1091 ringtest_0.x4._15_ a_26766_5712# 4.15e-19
C1092 ringtest_0.x4.net4 VDPWR 1.1491f
C1093 a_17377_14114# VDPWR 0.006305f
C1094 a_16755_12091# ui_in[4] 0.127717f
C1095 ringtest_0.x4._24_ a_27233_5308# 0.009415f
C1096 ringtest_0.x4._11_ a_24763_6143# 0.004209f
C1097 a_22373_5156# a_22457_5156# 0.008508f
C1098 a_21948_5156# ringtest_0.x4.net5 4.4e-19
C1099 ringtest_0.x4.net3 a_21399_5340# 0.007798f
C1100 a_22765_5308# a_22765_4478# 8.07e-19
C1101 ringtest_0.x4._08_ ringtest_0.x4._22_ 1.19e-20
C1102 ringtest_0.x4.net8 a_25975_3867# 0.2272f
C1103 ringtest_0.x4._18_ a_23899_5654# 9.76e-19
C1104 ringtest_0.x4._11_ a_22295_3867# 3.83e-19
C1105 muxtest_0.x1.x4.A muxtest_0.R3R4 4.53278f
C1106 ringtest_0.x4._16_ a_23381_4584# 0.039613f
C1107 a_12425_24040# VDPWR 4.32e-19
C1108 a_23899_5334# a_23809_4790# 8.68e-19
C1109 a_21951_5878# a_22649_6244# 0.194203f
C1110 a_22392_5990# a_22817_6146# 1.28e-19
C1111 ringtest_0.x4.net9 a_25149_4220# 0.125008f
C1112 muxtest_0.x2.x2.GN1 VDPWR 1.60341f
C1113 a_22052_8875# a_21785_8054# 0.0033f
C1114 ringtest_0.x4.net6 ringtest_0.x4._07_ 0.066033f
C1115 a_21852_8720# ringtest_0.x4._10_ 6.77e-19
C1116 a_23529_6422# a_23770_5308# 6.83e-19
C1117 ringtest_0.x4._01_ a_21803_8598# 2.39e-19
C1118 a_24715_5334# a_24895_5334# 0.001229f
C1119 a_24045_6654# ringtest_0.x4._16_ 1.29e-20
C1120 ringtest_0.x4._07_ a_24895_4790# 0.195848f
C1121 ringtest_0.x4._22_ a_25336_4902# 0.001181f
C1122 ringtest_0.x4._19_ a_25364_5878# 6.04e-19
C1123 a_24329_6640# ringtest_0.x4.net9 6.06e-20
C1124 ringtest_0.x4.net2 ringtest_0.x4._10_ 0.006086f
C1125 ringtest_0.x4.net6 a_25055_3867# 0.013611f
C1126 ringtest_0.x4._11_ ringtest_0.x4.clknet_1_1__leaf_clk 0.367667f
C1127 muxtest_0.R3R4 m3_13302_19985# 0.136776f
C1128 a_24895_4790# a_25055_3867# 1.2e-20
C1129 a_21425_9686# ringtest_0.x4.clknet_1_0__leaf_clk 3.24e-19
C1130 ringtest_0.x4._00_ a_22228_9508# 8.32e-19
C1131 ringtest_0.x4.net7 a_25149_4220# 0.212284f
C1132 a_25925_6788# ringtest_0.x4._23_ 0.026998f
C1133 ringtest_0.x4._18_ a_21785_5878# 7.56e-20
C1134 ringtest_0.x4.net6 a_24264_6788# 1.91e-20
C1135 muxtest_0.x1.x5.GN a_19794_32347# 9.76e-20
C1136 muxtest_0.x1.x1.nSEL1 a_19242_32347# 9.57e-19
C1137 ringtest_0.x4.net7 a_26735_5156# 1.13e-19
C1138 muxtest_0.x1.x3.GP2 ua[0] 1.13e-20
C1139 a_21675_4790# a_22295_3867# 7.04e-21
C1140 a_23837_5878# VDPWR 0.004487f
C1141 a_24329_6640# ringtest_0.x4.net7 0.035144f
C1142 ringtest_0.x4._22_ VDPWR 0.552873f
C1143 ringtest_0.x4._14_ a_21840_5308# 8.48e-21
C1144 ringtest_0.x3.x2.GP1 ua[1] 0.352376f
C1145 ringtest_0.x4.clknet_1_1__leaf_clk a_25761_5058# 0.084941f
C1146 ringtest_0.x4._06_ a_23770_5308# 0.002127f
C1147 muxtest_0.R3R4 muxtest_0.x2.x2.GP2 0.171364f
C1148 ringtest_0.x4.net8 a_26367_5340# 5.19e-19
C1149 ringtest_0.x4._11_ a_24800_5334# 2.99e-20
C1150 a_24135_3867# VDPWR 0.286734f
C1151 ringtest_0.x4._17_ a_24329_6640# 0.42661f
C1152 ringtest_0.x4.net9 a_24545_5878# 0.063508f
C1153 a_24070_5852# a_23770_5308# 8.74e-19
C1154 ringtest_0.x4._19_ a_24317_4942# 4.85e-22
C1155 a_17231_12017# a_17405_12123# 0.006584f
C1156 a_16755_12091# ringtest_0.x3.x2.GP1 2.87e-20
C1157 ringtest_0.x4.net2 a_21509_4790# 5.19e-20
C1158 muxtest_0.x2.x1.nSEL1 a_12473_23980# 0.041068f
C1159 a_15749_12123# ringtest_0.x3.x2.GN2 8.86e-19
C1160 ringtest_0.x3.x2.GN1 a_16155_12151# 1.22e-20
C1161 a_17231_12017# ringtest_0.x3.x2.GN3 1.07e-20
C1162 ringtest_0.x4._08_ a_25225_5334# 7.33e-20
C1163 a_24699_6200# ringtest_0.x4._16_ 0.113309f
C1164 a_23619_6788# VDPWR 0.002065f
C1165 a_25364_5878# ringtest_0.x4.net9 0.111158f
C1166 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ui_in[4] 0.001652f
C1167 ringtest_0.x4.net6 a_26201_5340# 2.14e-19
C1168 ringtest_0.x4._03_ a_22373_5156# 0.001345f
C1169 ringtest_0.x4._15_ a_24361_5340# 0.034785f
C1170 a_21509_4790# a_23381_4818# 7.98e-21
C1171 muxtest_0.x1.x4.A muxtest_0.x2.x1.nSEL0 4.83e-20
C1172 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 5.04e-19
C1173 ringtest_0.x4.net4 ringtest_0.x4.counter[2] 0.006188f
C1174 a_25225_5334# a_25336_4902# 0.001204f
C1175 a_25393_5308# a_25168_5156# 0.003655f
C1176 ringtest_0.x4.net7 a_24545_5878# 2.13e-20
C1177 a_16027_11759# VDPWR 0.161536f
C1178 muxtest_0.x1.x3.GN4 muxtest_0.R6R7 0.156481f
C1179 a_21465_8830# ringtest_0.x4._12_ 0.027335f
C1180 ringtest_0.x4._16_ a_24479_4790# 7.06e-20
C1181 ringtest_0.x4._11_ ringtest_0.x4._23_ 0.090724f
C1182 ringtest_0.x4.net7 a_25364_5878# 0.037674f
C1183 ringtest_0.x4.net2 a_21867_8054# 6.45e-19
C1184 ringtest_0.x4.net6 ringtest_0.x4.counter[5] 0.080069f
C1185 ringtest_0.x4._11_ a_26367_4790# 7.13e-19
C1186 a_19842_32287# muxtest_0.R7R8 7.47e-21
C1187 ringtest_0.x4._16_ a_23809_4790# 0.105405f
C1188 ringtest_0.x4.net2 ringtest_0.x4._13_ 0.197255f
C1189 ringtest_0.x4.net9 a_24317_4942# 3.24e-20
C1190 a_23949_6654# ringtest_0.x4.net8 1.16e-19
C1191 ringtest_0.x4._17_ a_25364_5878# 0.002308f
C1192 a_15749_12123# ui_in[3] 9.55e-19
C1193 a_24527_5340# a_24715_5334# 0.095025f
C1194 ringtest_0.counter3 ringtest_0.counter7 3.44556f
C1195 ui_in[2] ui_in[4] 0.020899f
C1196 muxtest_0.R7R8 m3_13316_18955# 0.131878f
C1197 a_25225_5334# VDPWR 0.181757f
C1198 a_24465_6800# a_24883_6800# 3.39e-19
C1199 ringtest_0.x4._16_ a_22795_5334# 0.059496f
C1200 a_21675_10006# ringtest_0.x4._00_ 0.002065f
C1201 a_19114_31955# a_19290_32287# 0.185422f
C1202 ringtest_0.x4._23_ a_25761_5058# 1.37e-20
C1203 a_21233_5340# ringtest_0.x4._02_ 0.184941f
C1204 a_25761_5058# a_26367_4790# 8.52e-19
C1205 a_23529_6422# ringtest_0.x4.net6 1.5e-19
C1206 a_12473_23980# muxtest_0.x2.x2.GN3 0.048646f
C1207 ringtest_0.x4.net7 a_24317_4942# 0.084753f
C1208 a_12849_23648# muxtest_0.x2.x2.GN1 6.43e-20
C1209 ringtest_0.x4._21_ a_23837_5878# 0.002821f
C1210 ringtest_0.counter7 ua[2] 2.06e-19
C1211 ringtest_0.x4._11_ ringtest_0.x4._02_ 0.012298f
C1212 ringtest_0.x4._21_ ringtest_0.x4._22_ 2.96e-19
C1213 ringtest_0.x4._17_ a_24317_4942# 1.09e-21
C1214 m2_11882_23495# ui_in[3] 0.130999f
C1215 a_27169_6641# a_26201_5340# 7.7e-20
C1216 a_26749_6422# a_26367_5340# 6.98e-21
C1217 ringtest_0.x4._03_ a_22499_4790# 9.96e-20
C1218 a_22021_4220# VDPWR 0.37664f
C1219 a_21509_4790# ringtest_0.x4._20_ 1.9e-21
C1220 ringtest_0.counter7 ringtest_0.x4.net10 5.8e-20
C1221 a_21951_5878# a_22733_6244# 4.04e-19
C1222 a_22224_6244# a_22139_5878# 0.037333f
C1223 ringtest_0.x4.net8 a_24004_6128# 0.063158f
C1224 a_26640_5156# VDPWR 0.247956f
C1225 ringtest_0.counter3 a_22295_3867# 5.4e-19
C1226 ringtest_0.x4.net4 a_21375_3867# 7.77e-19
C1227 a_21132_8918# a_21049_8598# 2.42e-19
C1228 ringtest_0.x4._12_ a_21780_8964# 0.001666f
C1229 ringtest_0.x4._19_ ringtest_0.x4.net9 4.58e-20
C1230 VDPWR ua[3] 11.3115f
C1231 ringtest_0.x4.net6 ringtest_0.x4._06_ 0.037389f
C1232 a_23879_6940# a_23837_5878# 1.78e-20
C1233 ringtest_0.x4._24_ a_27491_4566# 5.3e-19
C1234 ringtest_0.x4.net6 a_24070_5852# 0.016498f
C1235 ringtest_0.x3.x2.GP2 ringtest_0.counter3 0.148166f
C1236 a_23879_6940# ringtest_0.x4._22_ 7.51e-19
C1237 a_21399_5340# ringtest_0.x4._03_ 1.23e-19
C1238 a_21233_5340# a_22116_4902# 0.001786f
C1239 a_26201_4790# a_26895_3867# 4.75e-20
C1240 a_21840_5308# a_21509_4790# 0.001425f
C1241 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP1 0.051787f
C1242 ringtest_0.x4.net8 a_23963_4790# 8.5e-20
C1243 a_22765_4478# a_22390_4566# 4e-20
C1244 ringtest_0.x4._15_ ringtest_0.x4._08_ 0.030258f
C1245 ringtest_0.x4._11_ a_25593_5156# 0.045045f
C1246 muxtest_0.R3R4 ua[0] 3.1523f
C1247 ui_in[1] ui_in[6] 0.239552f
C1248 a_20492_32319# VDPWR 8.55e-19
C1249 a_21561_9116# a_21780_9142# 0.006169f
C1250 ringtest_0.counter7 ringtest_0.x4.counter[4] 0.007159f
C1251 a_18836_32319# muxtest_0.x1.x3.GN2 8.86e-19
C1252 muxtest_0.x1.x3.GN1 a_19242_32347# 1.22e-20
C1253 a_21675_9686# a_21845_9116# 5.23e-20
C1254 a_20318_32213# muxtest_0.x1.x3.GN3 1.07e-20
C1255 a_21465_9294# a_21852_9416# 0.034054f
C1256 ringtest_0.counter7 a_23399_3867# 2.81e-20
C1257 a_19842_32287# VDPWR 0.261767f
C1258 a_27065_5156# ringtest_0.x4.net11 0.003417f
C1259 ringtest_0.x4._11_ a_22116_4902# 0.004479f
C1260 ringtest_0.x4._19_ ringtest_0.x4.net7 0.552257f
C1261 muxtest_0.x1.x1.nSEL0 a_19290_32287# 0.001174f
C1262 a_22649_6244# a_22795_5334# 1.65e-19
C1263 ringtest_0.x4._15_ a_25336_4902# 4.59e-21
C1264 ringtest_0.x4._11_ a_23993_5654# 5.64e-19
C1265 ringtest_0.x4._16_ a_21672_5334# 1.68e-20
C1266 a_24045_6654# a_24465_6800# 0.036838f
C1267 a_24329_6640# a_24536_6699# 0.260055f
C1268 ringtest_0.x4._17_ ringtest_0.x4._19_ 0.214371f
C1269 a_23949_6654# ringtest_0.x4._05_ 1.85e-19
C1270 ringtest_0.x4._24_ a_27149_5334# 8.56e-19
C1271 a_25761_5058# a_25593_5156# 0.310858f
C1272 a_25168_5156# a_25083_4790# 0.037333f
C1273 ua[0] ui_in[5] 0.483363f
C1274 muxtest_0.R3R4 muxtest_0.x2.x2.GN3 3.9625f
C1275 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x1.nSEL1 0.352716f
C1276 a_21561_8830# VDPWR 0.179712f
C1277 ringtest_0.x4._04_ a_21233_5340# 0.001469f
C1278 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net10 6.99e-20
C1279 ringtest_0.drv_out ui_in[5] 0.391919f
C1280 a_27815_3867# ringtest_0.x4.counter[9] 0.039377f
C1281 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ui_in[4] 1.79e-19
C1282 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x3.x2.GN1 2.09e-20
C1283 ringtest_0.x4._15_ VDPWR 1.68193f
C1284 ringtest_0.x4.clknet_1_0__leaf_clk a_21233_5340# 0.318658f
C1285 a_21675_4790# a_22116_4902# 0.127288f
C1286 a_26808_5308# a_26201_4790# 1.99e-20
C1287 ringtest_0.drv_out ringtest_0.x4.clknet_0_clk 0.00889f
C1288 ui_in[0] ui_in[2] 0.450267f
C1289 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.173286f
C1290 ringtest_0.x4._11_ ringtest_0.x4._04_ 0.257603f
C1291 a_25263_5156# VDPWR 0.00304f
C1292 a_22295_3867# a_23399_3867# 9e-21
C1293 a_25364_5878# a_26627_4246# 1.15e-20
C1294 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._11_ 0.317456f
C1295 a_24536_6699# a_24545_5878# 1.55e-20
C1296 ringtest_0.x4.net7 ringtest_0.x4.net9 0.742565f
C1297 a_22541_5058# VDPWR 0.387929f
C1298 ringtest_0.x4.net3 a_22052_8875# 3.02e-19
C1299 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.ring_out 0.083309f
C1300 ringtest_0.x4.net2 ringtest_0.x4.counter[1] 0.015257f
C1301 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP2 0.100463f
C1302 a_25225_5334# a_25309_5334# 0.008508f
C1303 a_26808_5308# a_26555_5334# 3.39e-19
C1304 a_22052_9116# a_21852_8720# 1.26e-19
C1305 a_21981_9142# a_21845_8816# 5.28e-20
C1306 a_21845_9116# a_22052_8875# 6.88e-20
C1307 ringtest_0.x4._17_ ringtest_0.x4.net9 7.02e-19
C1308 a_24465_6800# a_24699_6200# 1.61e-19
C1309 muxtest_0.x1.x5.GN ui_in[1] 0.141313f
C1310 a_24926_5712# VDPWR 0.001185f
C1311 ringtest_0.x3.x2.GN2 ringtest_0.counter3 0.004367f
C1312 ringtest_0.x4._15_ a_23467_4584# 0.001523f
C1313 ringtest_0.x4.net1 a_21561_8830# 0.030538f
C1314 ringtest_0.x4._15_ ringtest_0.x4._25_ 0.003323f
C1315 ringtest_0.x4.net8 ringtest_0.x4._20_ 0.027217f
C1316 ringtest_0.ring_out a_17405_12123# 1.86e-19
C1317 ringtest_0.x4.net2 a_22052_9116# 1.88e-19
C1318 ringtest_0.ring_out ringtest_0.x3.x2.GN3 0.080584f
C1319 a_21951_5878# ringtest_0.x4._03_ 3.92e-19
C1320 ringtest_0.x4._09_ a_27065_5156# 0.024482f
C1321 a_26201_4790# a_26555_4790# 0.062224f
C1322 ringtest_0.x4._07_ a_24527_5340# 0.029939f
C1323 ringtest_0.x4._22_ a_24968_5308# 0.01767f
C1324 ringtest_0.x4.net5 a_22164_4362# 3.95e-20
C1325 ringtest_0.x4._17_ ringtest_0.x4.net7 0.072785f
C1326 ringtest_0.x4.clknet_1_0__leaf_clk a_21675_4790# 0.021572f
C1327 ringtest_0.counter7 a_26808_4902# 1.4e-19
C1328 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN3 4.01e-20
C1329 ringtest_0.x3.x2.GN4 ringtest_0.counter7 3.94045f
C1330 a_24527_5340# a_25055_3867# 7.09e-22
C1331 ringtest_0.x4._23_ ringtest_0.x4.net10 0.188811f
C1332 ringtest_0.x4.clknet_0_clk ringtest_0.x4._07_ 0.114561f
C1333 ringtest_0.counter3 ringtest_0.x4._02_ 0.001266f
C1334 a_21049_8598# VDPWR 0.226794f
C1335 ringtest_0.x4._20_ a_24729_4790# 0.004564f
C1336 a_22224_6244# a_22097_5334# 0.002298f
C1337 a_26173_4612# VDPWR 0.001618f
C1338 ringtest_0.x4.net10 a_26367_4790# 0.003321f
C1339 a_12849_23648# ua[3] 0.001506f
C1340 a_22224_6244# ringtest_0.x4._16_ 1.81e-20
C1341 ringtest_0.x4.net4 a_21233_5340# 0.007432f
C1342 a_26895_3867# ringtest_0.x4.counter[8] 6.92e-19
C1343 muxtest_0.x1.x4.A a_13025_23980# 3.23e-19
C1344 ringtest_0.x4.clknet_1_1__leaf_clk a_25393_5308# 0.005058f
C1345 ringtest_0.x4.net6 a_21399_5340# 1.26e-19
C1346 ringtest_0.x4._11_ ringtest_0.x4.net4 0.952686f
C1347 ringtest_0.x4.clknet_0_clk a_24264_6788# 1.49e-19
C1348 a_21785_5878# ringtest_0.x4._04_ 0.09532f
C1349 ringtest_0.x4._15_ ringtest_0.x4._21_ 0.054317f
C1350 ringtest_0.x4.clknet_1_0__leaf_clk a_21785_5878# 0.245743f
C1351 a_26627_4246# a_26913_4566# 0.010132f
C1352 muxtest_0.x2.x2.GN1 m2_11882_23495# 0.06935f
C1353 a_22399_9142# ringtest_0.x4.clknet_1_0__leaf_clk 0.012004f
C1354 ringtest_0.x4.net1 a_21049_8598# 0.060735f
C1355 ui_in[3] ua[2] 1.63519f
C1356 a_13501_23906# ui_in[3] 0.220366f
C1357 a_21425_9686# a_21561_8830# 6.59e-20
C1358 ringtest_0.x4.net7 a_26095_6788# 0.00717f
C1359 ringtest_0.x4._21_ a_22541_5058# 1.79e-21
C1360 ringtest_0.x4._17_ a_22817_6146# 1.35e-20
C1361 a_24527_5340# a_26201_5340# 1.33e-19
C1362 a_24968_5308# a_25225_5334# 0.036838f
C1363 a_24361_5340# a_26367_5340# 3.42e-21
C1364 a_21672_5334# a_21587_5334# 0.037333f
C1365 a_21840_5308# a_21798_5712# 4.62e-19
C1366 a_19290_32287# muxtest_0.x1.x3.GN2 0.017048f
C1367 ringtest_0.x4.net9 a_27065_5334# 2.45e-19
C1368 ringtest_0.x4.clknet_1_1__leaf_clk a_26808_4902# 2.7e-19
C1369 ringtest_0.x4.net4 a_21675_4790# 0.019846f
C1370 a_24536_6699# ringtest_0.x4._19_ 0.034076f
C1371 a_13025_23980# muxtest_0.x2.x2.GP2 3.2e-20
C1372 a_23879_6940# ringtest_0.x4._15_ 2.08e-20
C1373 muxtest_0.x2.x2.GP3 ui_in[4] 0.00356f
C1374 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP2 8.45e-19
C1375 ringtest_0.x4._03_ a_23381_4584# 2.93e-20
C1376 a_19794_32347# ui_in[0] 0.001558f
C1377 ringtest_0.x4.net4 a_23899_5654# 7.88e-20
C1378 ringtest_0.x3.x2.GN1 ui_in[4] 0.312198f
C1379 ringtest_0.x4._11_ a_23837_5878# 3.73e-19
C1380 a_15575_12017# ringtest_0.x3.x2.GN2 0.039612f
C1381 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN3 0.012418f
C1382 ringtest_0.x4._11_ ringtest_0.x4._22_ 0.420712f
C1383 a_22373_5156# ringtest_0.x4.net5 0.019334f
C1384 ringtest_0.x4.net3 a_21672_5334# 8.21e-19
C1385 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ui_in[4] 1.03e-20
C1386 rst_n clk 0.031023f
C1387 a_22392_5990# ringtest_0.x4.net8 1.22e-20
C1388 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 5.04e-19
C1389 ringtest_0.x4.net9 a_26627_4246# 0.008597f
C1390 muxtest_0.x1.x3.GP1 muxtest_0.R3R4 4.16645f
C1391 a_21981_8976# ringtest_0.x4._10_ 6.67e-19
C1392 ringtest_0.x4._01_ a_21785_8054# 3.94e-19
C1393 a_24045_6654# a_23770_5308# 7.28e-21
C1394 ringtest_0.x4.net4 a_21785_5878# 0.071607f
C1395 ringtest_0.x4.net9 a_27149_5156# 1.5e-19
C1396 ringtest_0.x4._11_ a_23619_6788# 1.46e-19
C1397 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ui_in[3] 1.18e-19
C1398 a_24336_6544# ringtest_0.x4._16_ 6.29e-20
C1399 ringtest_0.x4._07_ a_25168_5156# 0.008539f
C1400 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.ring_out 0.025177f
C1401 a_24536_6699# ringtest_0.x4.net9 4.56e-19
C1402 ringtest_0.x4._22_ a_25761_5058# 3.11e-19
C1403 a_24883_6800# a_24712_6422# 0.001229f
C1404 ui_in[0] rst_n 0.031023f
C1405 ui_in[4] ui_in[6] 0.178963f
C1406 ringtest_0.x4.clknet_0_clk a_23529_6422# 8e-19
C1407 ringtest_0.x4.net6 a_21951_5878# 0.004467f
C1408 ringtest_0.x4._24_ a_27273_4220# 0.003347f
C1409 a_15575_12017# m2_15612_11606# 0.01297f
C1410 a_26569_6422# a_26749_6422# 0.185422f
C1411 ringtest_0.x4.net6 a_24883_6800# 9.51e-20
C1412 ringtest_0.x4._00_ ringtest_0.x4.clknet_1_0__leaf_clk 0.144154f
C1413 a_15575_12017# ui_in[3] 0.048888f
C1414 ringtest_0.x4._24_ a_26766_4790# 6.57e-19
C1415 ringtest_0.x4._23_ a_26808_4902# 0.005759f
C1416 ringtest_0.x4.net7 a_27149_5156# 3.05e-20
C1417 ringtest_0.x4._05_ a_26569_6422# 6.38e-20
C1418 muxtest_0.x1.x1.nSEL1 VDPWR 0.475048f
C1419 a_24763_6143# a_24715_5334# 1.39e-19
C1420 a_26367_4790# a_26808_4902# 0.118966f
C1421 a_24536_6699# ringtest_0.x4.net7 0.026259f
C1422 ringtest_0.x4._14_ a_22265_5308# 1.02e-20
C1423 ringtest_0.x4.clknet_1_1__leaf_clk a_25083_4790# 0.011819f
C1424 ringtest_0.x4._06_ a_24527_5340# 0.183131f
C1425 ringtest_0.x4.net8 a_26640_5334# 2.79e-19
C1426 ringtest_0.x4._16_ a_24986_5878# 3.12e-19
C1427 ringtest_0.x4._11_ a_25225_5334# 7.12e-21
C1428 ringtest_0.x4._17_ a_24536_6699# 0.032936f
C1429 a_16707_12151# ringtest_0.x3.x2.GN4 3.22e-19
C1430 ringtest_0.x3.x2.GN3 a_17405_12123# 1.07e-20
C1431 a_25975_3867# VDPWR 0.309189f
C1432 a_24004_6128# a_24361_5340# 4.26e-19
C1433 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GN4 8.82e-19
C1434 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP1 1.51569f
C1435 muxtest_0.x2.x1.nSEL1 a_13025_23980# 1.59e-19
C1436 ringtest_0.x4._08_ a_26367_5340# 0.415957f
C1437 ringtest_0.x4.clknet_0_clk ringtest_0.x4._06_ 2.8e-19
C1438 ringtest_0.x4.net5 a_22499_4790# 6.03e-19
C1439 a_24685_6788# VDPWR 0.002269f
C1440 ringtest_0.x4._04_ a_22775_5878# 6.79e-19
C1441 a_21785_5878# a_23837_5878# 9.88e-21
C1442 ringtest_0.x4.clknet_0_clk a_24070_5852# 7.65e-20
C1443 ui_in[1] ui_in[4] 4.85e-19
C1444 ringtest_0.x4.clknet_1_1__leaf_clk a_24715_5334# 0.017223f
C1445 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x3.nselect2 1.41e-19
C1446 ringtest_0.x4._15_ a_24968_5308# 0.03519f
C1447 ringtest_0.x4._22_ a_25345_4612# 0.002279f
C1448 a_21233_5340# a_22021_4220# 3.4e-19
C1449 ringtest_0.x4._01_ a_22695_8304# 0.012244f
C1450 muxtest_0.x1.x5.A ua[3] 4.51865f
C1451 ringtest_0.counter3 ringtest_0.x4.net4 8.11e-19
C1452 a_25393_5308# a_25593_5156# 4.17e-19
C1453 a_24800_5334# a_25083_4790# 0.001307f
C1454 a_26913_4566# a_26721_4246# 6.96e-20
C1455 muxtest_0.x1.x3.GN3 muxtest_0.R4R5 0.123863f
C1456 a_21845_8816# ringtest_0.x4._12_ 0.062549f
C1457 a_16579_11759# VDPWR 0.179803f
C1458 ringtest_0.x4.net8 a_25149_4220# 0.1454f
C1459 ringtest_0.x4._11_ a_22021_4220# 7.66e-19
C1460 a_23770_5308# a_23809_4790# 2.2e-19
C1461 ringtest_0.x4.net9 a_25294_4790# 3.93e-19
C1462 muxtest_0.x1.x5.GN ui_in[4] 2.49e-19
C1463 ringtest_0.x4.net11 a_27489_3702# 0.250513f
C1464 ringtest_0.x4._11_ a_26640_5156# 5.04e-19
C1465 muxtest_0.x1.x3.GN1 muxtest_0.R7R8 4.45989f
C1466 ringtest_0.x3.x2.GN4 ui_in[3] 0.218716f
C1467 a_24329_6640# ringtest_0.x4.net8 0.001356f
C1468 ringtest_0.x4.net2 a_21132_8918# 0.010623f
C1469 a_24968_5308# a_24926_5712# 4.62e-19
C1470 a_22765_5308# a_23151_5334# 0.006406f
C1471 a_24800_5334# a_24715_5334# 0.037333f
C1472 ringtest_0.x4._08_ a_27065_5156# 3.02e-19
C1473 a_26367_5340# VDPWR 0.308687f
C1474 ringtest_0.x4._15_ a_25925_6788# 0.142876f
C1475 ringtest_0.x4._16_ a_23899_5334# 0.008193f
C1476 ringtest_0.x4.net6 a_23381_4584# 1.4e-20
C1477 ringtest_0.drv_out ringtest_0.counter7 2.39e-19
C1478 ringtest_0.x4.net9 a_25351_5712# 3.81e-19
C1479 ringtest_0.x4._24_ a_26201_4790# 0.03301f
C1480 a_19290_32287# a_19666_31955# 3.02e-19
C1481 muxtest_0.x1.x4.A ui_in[3] 0.004014f
C1482 a_24729_4790# a_25149_4220# 0.009169f
C1483 a_24045_6654# ringtest_0.x4.net6 8.38e-19
C1484 a_13025_23980# muxtest_0.x2.x2.GN3 0.004288f
C1485 a_21675_4790# a_22021_4220# 0.010515f
C1486 muxtest_0.x2.x2.GN1 ua[2] 0.430038f
C1487 a_24329_6640# a_24729_4790# 2.6e-21
C1488 ringtest_0.x4._24_ a_26555_5334# 4.8e-19
C1489 ringtest_0.x4.net7 a_25351_5712# 1.38e-19
C1490 ringtest_0.x4.net8 a_24545_5878# 0.009814f
C1491 a_27233_5308# a_27273_4220# 1.35e-20
C1492 ringtest_0.x4._25_ a_26367_5340# 1.11e-19
C1493 ui_in[0] ui_in[6] 0.281408f
C1494 ringtest_0.x3.nselect2 a_16755_12091# 6.01e-20
C1495 a_22765_4478# VDPWR 0.201367f
C1496 a_21951_5878# a_23932_6128# 1.01e-20
C1497 a_21507_9686# VDPWR 0.008578f
C1498 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ui_in[4] 7.73e-20
C1499 a_22392_5990# a_22350_5878# 4.62e-19
C1500 ringtest_0.x4.net8 a_25364_5878# 0.001798f
C1501 ringtest_0.x4.net9 a_26721_4246# 0.003753f
C1502 a_27065_5156# VDPWR 0.210976f
C1503 ringtest_0.x4._15_ a_21233_5340# 8.17e-21
C1504 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.173286f
C1505 a_23949_6654# VDPWR 0.375047f
C1506 muxtest_0.x1.x3.GP2 muxtest_0.R4R5 0.117653f
C1507 ringtest_0.x4._12_ a_22201_8964# 0.002771f
C1508 a_21845_8816# a_22245_8054# 4.04e-19
C1509 ringtest_0.x4.net4 a_23399_3867# 0.003224f
C1510 muxtest_0.x2.x2.GP2 ui_in[3] 6.63e-19
C1511 ringtest_0.x4._11_ ringtest_0.x4._15_ 1.40124f
C1512 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B 0.163894f
C1513 muxtest_0.x1.x3.GN1 muxtest_0.R5R6 0.250509f
C1514 ringtest_0.x4.net6 a_24699_6200# 0.09145f
C1515 a_22265_5308# a_21509_4790# 0.00142f
C1516 a_21672_5334# ringtest_0.x4._03_ 0.001262f
C1517 ringtest_0.x4.net8 a_24551_4790# 5.79e-19
C1518 a_24699_6200# a_24895_4790# 8.41e-19
C1519 a_25364_5878# a_24729_4790# 4.21e-21
C1520 ringtest_0.drv_out ringtest_0.x4.clknet_1_1__leaf_clk 0.008913f
C1521 ringtest_0.drv_out ringtest_0.x3.x2.GP2 4.09557f
C1522 a_21561_9116# a_21845_9116# 0.032244f
C1523 ringtest_0.counter7 a_25055_3867# 2.81e-20
C1524 ringtest_0.x4._22_ ringtest_0.x4.net10 0.074459f
C1525 muxtest_0.x1.x3.GN1 VDPWR 0.915833f
C1526 ringtest_0.x4._11_ a_22541_5058# 0.065594f
C1527 a_21951_5878# ringtest_0.x4.net5 3.57e-21
C1528 ringtest_0.x4.net8 a_24317_4942# 0.236033f
C1529 ringtest_0.x4.net1 a_21507_9686# 0.010028f
C1530 a_22265_5308# a_22765_5308# 0.016344f
C1531 muxtest_0.x1.x1.nSEL0 a_19842_32287# 1.21e-20
C1532 ui_in[0] ui_in[1] 4.44986f
C1533 ringtest_0.x4.net6 a_24479_4790# 1.78e-19
C1534 ringtest_0.x4._15_ a_25761_5058# 7.77e-19
C1535 ringtest_0.x4._16_ a_22097_5334# 1.35e-19
C1536 a_24329_6640# ringtest_0.x4._05_ 0.196756f
C1537 a_24336_6544# a_24465_6800# 0.110715f
C1538 muxtest_0.x1.x3.GN3 ui_in[2] 0.002225f
C1539 a_24004_6128# VDPWR 0.314938f
C1540 a_24729_4790# a_24551_4790# 1.43e-19
C1541 a_21395_6940# a_21840_5308# 3.17e-20
C1542 ringtest_0.x4.net6 a_23809_4790# 0.005791f
C1543 a_24763_6143# ringtest_0.x4._07_ 0.001092f
C1544 a_21852_8720# VDPWR 0.304165f
C1545 muxtest_0.x1.x5.GN ui_in[0] 0.149831f
C1546 a_24317_4942# a_24729_4790# 0.020429f
C1547 ringtest_0.x4._15_ a_23899_5654# 0.005043f
C1548 ringtest_0.x4.net6 a_22795_5334# 0.007899f
C1549 a_22116_4902# a_21948_5156# 0.239923f
C1550 a_24135_3867# ringtest_0.x4.counter[4] 0.110403f
C1551 ringtest_0.x4.net2 VDPWR 2.35179f
C1552 a_21675_4790# a_22541_5058# 0.034054f
C1553 a_23963_4790# VDPWR 2.15e-19
C1554 a_23399_3867# a_24135_3867# 2.31e-20
C1555 ringtest_0.x4._11_ a_26173_4612# 7.08e-19
C1556 a_26749_6422# a_25364_5878# 0.006666f
C1557 muxtest_0.x1.x3.GP3 muxtest_0.R7R8 0.124327f
C1558 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._07_ 0.44529f
C1559 a_23381_4818# VDPWR 0.253456f
C1560 ringtest_0.x4.net3 ringtest_0.x4._01_ 0.006403f
C1561 a_26640_5334# a_26766_5712# 0.005525f
C1562 a_22052_9116# a_21981_8976# 1.77e-19
C1563 ringtest_0.x4.clknet_1_0__leaf_clk a_21465_8830# 0.01132f
C1564 a_23949_6654# ringtest_0.x4._21_ 0.001295f
C1565 ringtest_0.x4._05_ a_25364_5878# 0.003024f
C1566 a_21845_9116# ringtest_0.x4._01_ 6.79e-20
C1567 a_21981_9142# a_22052_8875# 1.77e-19
C1568 ringtest_0.x4._19_ ringtest_0.x4.net8 2.14e-19
C1569 ringtest_0.x4.clknet_1_1__leaf_clk a_25055_3867# 4.13e-21
C1570 a_22181_5334# VDPWR 0.007439f
C1571 ringtest_0.counter7 ringtest_0.x4.counter[5] 0.007023f
C1572 ringtest_0.x4._15_ a_25345_4612# 2.85e-21
C1573 ringtest_0.x4.net1 a_21852_8720# 0.00338f
C1574 muxtest_0.x2.x1.nSEL1 ui_in[3] 0.168511f
C1575 ringtest_0.drv_out ringtest_0.x3.x2.GN2 3.92936f
C1576 a_26201_4790# a_25977_4220# 2.81e-20
C1577 a_21425_9686# a_21507_9686# 0.006406f
C1578 a_21785_5878# a_22541_5058# 3.85e-19
C1579 muxtest_0.x2.x2.GN4 muxtest_0.x2.x2.GP3 3.4436f
C1580 ringtest_0.x4._04_ a_21948_5156# 3.52e-21
C1581 ringtest_0.x4.net8 a_26735_5334# 7.49e-20
C1582 ringtest_0.x4._07_ a_24800_5334# 0.002926f
C1583 ringtest_0.x4.net1 ringtest_0.x4.net2 0.722672f
C1584 a_25421_6641# ringtest_0.x4.net6 0.019537f
C1585 ringtest_0.x4.net3 a_21863_4790# 7.76e-19
C1586 ringtest_0.x4._22_ a_25393_5308# 4.4e-21
C1587 ringtest_0.x4.net5 a_23381_4584# 0.201023f
C1588 muxtest_0.x1.x3.GP2 ui_in[2] 4.34e-19
C1589 ringtest_0.x4.clknet_1_0__leaf_clk a_21948_5156# 0.003461f
C1590 ringtest_0.x4._18_ a_23529_6422# 0.190808f
C1591 a_22399_8976# VDPWR 0.073139f
C1592 a_24800_5334# a_25055_3867# 3e-19
C1593 a_22817_6146# a_22765_5308# 0.004132f
C1594 a_23879_6940# a_23949_6654# 0.022122f
C1595 ringtest_0.x4._20_ a_25336_4902# 6.25e-20
C1596 muxtest_0.R7R8 muxtest_0.R1R2 0.216753f
C1597 a_26375_4612# VDPWR 8.72e-20
C1598 ringtest_0.x4.net10 a_26640_5156# 5.45e-19
C1599 ua[3] ua[2] 8.93455f
C1600 a_13501_23906# ua[3] 0.003273f
C1601 a_24883_6800# a_24527_5340# 1.11e-20
C1602 a_22649_6244# ringtest_0.x4._16_ 0.003542f
C1603 a_15575_12017# a_16027_11759# 0.002207f
C1604 ringtest_0.x4.net8 ringtest_0.x4.net9 0.748324f
C1605 a_24004_6128# ringtest_0.x4._21_ 0.128337f
C1606 a_27815_3867# ringtest_0.x4.counter[8] 0.111116f
C1607 muxtest_0.R4R5 muxtest_0.R3R4 1.39313f
C1608 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN1 1.38e-21
C1609 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ui_in[4] 1.2e-19
C1610 ringtest_0.x4.clknet_1_1__leaf_clk a_26201_5340# 0.285659f
C1611 ringtest_0.x3.x2.GP3 VDPWR 1.79155f
C1612 ringtest_0.x4.net6 a_21672_5334# 6.57e-20
C1613 ringtest_0.x4._13_ ringtest_0.x4.counter[0] 3.39e-20
C1614 ringtest_0.x4.clknet_0_clk a_24883_6800# 0.004448f
C1615 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 5.04e-19
C1616 muxtest_0.x1.x3.GP3 muxtest_0.R5R6 4.11451f
C1617 ringtest_0.x4._20_ VDPWR 0.172559f
C1618 ringtest_0.x4._22_ a_26808_4902# 8.71e-19
C1619 ringtest_0.x4.net3 a_21785_8054# 0.079675f
C1620 muxtest_0.x1.x3.GN2 ua[3] 0.01442f
C1621 ringtest_0.x4.clknet_1_0__leaf_clk a_21780_8964# 0.001172f
C1622 a_27273_4220# a_27491_4566# 0.007234f
C1623 a_22164_4362# a_22295_3867# 0.002548f
C1624 a_26627_4246# a_26721_4246# 0.062574f
C1625 ringtest_0.x4._16_ a_23467_4818# 5.76e-19
C1626 ringtest_0.x4.net7 ringtest_0.x4.net8 1.22349f
C1627 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B 5.04e-19
C1628 a_13675_24012# ui_in[3] 1.4e-19
C1629 a_25364_5878# ringtest_0.x4._09_ 3.55e-20
C1630 ringtest_0.x4.net9 a_24729_4790# 0.006834f
C1631 muxtest_0.x2.x2.GN3 ui_in[3] 0.254283f
C1632 ringtest_0.x4._18_ ringtest_0.x4._06_ 3.12e-20
C1633 ringtest_0.x4.net1 a_22399_8976# 6.38e-20
C1634 muxtest_0.x1.x3.GP3 VDPWR 3.24635f
C1635 muxtest_0.x1.x3.GN3 a_19794_32347# 0.001073f
C1636 ringtest_0.x4._18_ a_24070_5852# 7.58e-19
C1637 muxtest_0.x1.x3.GN2 a_20492_32319# 8.14e-21
C1638 ringtest_0.x4.net7 a_26839_6788# 1.83e-19
C1639 a_23879_6940# a_24004_6128# 1.01e-19
C1640 ringtest_0.x4._17_ ringtest_0.x4.net8 0.172731f
C1641 a_25393_5308# a_25225_5334# 0.310858f
C1642 a_21840_5308# a_22223_5712# 4.67e-20
C1643 a_19842_32287# muxtest_0.x1.x3.GN2 9.62e-20
C1644 ringtest_0.x4.net6 ringtest_0.x4._24_ 0.002355f
C1645 a_21840_5308# VDPWR 0.198342f
C1646 ringtest_0.x4._16_ a_21587_5334# 4.26e-21
C1647 ringtest_0.x4.net2 a_21425_9686# 0.107098f
C1648 ringtest_0.x4.net4 a_21948_5156# 0.004091f
C1649 ringtest_0.x4.clknet_1_1__leaf_clk a_27233_5058# 1.1e-19
C1650 muxtest_0.x1.x1.nSEL1 a_19114_31955# 0.073392f
C1651 ua[2] ua[6] 0.001584f
C1652 ringtest_0.x4._05_ ringtest_0.x4._19_ 0.284135f
C1653 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP2 0.005194f
C1654 ringtest_0.x4.net7 a_24729_4790# 0.003956f
C1655 a_23529_6422# ringtest_0.x4.clknet_1_1__leaf_clk 1.19e-21
C1656 ringtest_0.x4._15_ ringtest_0.x4.net10 0.289356f
C1657 ringtest_0.x4._17_ a_24729_4790# 1.69e-21
C1658 ringtest_0.x3.x2.GP1 ui_in[4] 8.45e-19
C1659 ringtest_0.x4._06_ a_24763_6143# 9.69e-19
C1660 a_16203_12091# ringtest_0.x3.x2.GN2 0.017071f
C1661 a_23809_4790# ringtest_0.x4.net5 5.06e-20
C1662 a_26569_6422# VDPWR 0.205477f
C1663 ringtest_0.x4._23_ a_26201_5340# 0.029216f
C1664 muxtest_0.R1R2 VDPWR 1.61319f
C1665 a_26201_5340# a_26367_4790# 2.64e-19
C1666 ringtest_0.x4.net3 ringtest_0.x4._16_ 6.72e-19
C1667 ringtest_0.x4._11_ a_25975_3867# 2.18e-19
C1668 a_22817_6146# ringtest_0.x4.net8 5.45e-19
C1669 a_26749_6422# ringtest_0.x4.net9 7.48e-22
C1670 a_24329_6640# a_24361_5340# 0.001493f
C1671 ringtest_0.x4.net9 ringtest_0.x4.net11 0.055197f
C1672 ringtest_0.x4._07_ a_25593_5156# 5.62e-20
C1673 ringtest_0.x4._15_ ringtest_0.x4.counter[4] 9.07e-20
C1674 a_24465_6800# ringtest_0.x4._16_ 2.16e-20
C1675 ringtest_0.x3.x2.GP2 m3_17036_9140# 0.004119f
C1676 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._06_ 0.005269f
C1677 ringtest_0.x4._22_ a_25083_4790# 0.012798f
C1678 ringtest_0.x4._05_ ringtest_0.x4.net9 1.93e-19
C1679 ringtest_0.x4.clknet_0_clk a_24045_6654# 0.00222f
C1680 ringtest_0.x4.net6 a_22224_6244# 3.12e-19
C1681 ringtest_0.x4.net2 a_21375_3867# 0.016821f
C1682 ringtest_0.x4._14_ a_21509_4790# 0.008544f
C1683 ringtest_0.x4._21_ ringtest_0.x4._20_ 0.296715f
C1684 ringtest_0.x4._24_ a_27169_6641# 0.006166f
C1685 a_26569_6422# ringtest_0.x4._25_ 0.001476f
C1686 a_25761_5058# a_25975_3867# 2.93e-21
C1687 a_16203_12091# ui_in[3] 0.143958f
C1688 ringtest_0.x4.net7 a_26749_6422# 5.4e-19
C1689 muxtest_0.R3R4 ui_in[2] 2.94e-19
C1690 ringtest_0.x4.net7 ringtest_0.x4.net11 2.47e-20
C1691 ringtest_0.x4._23_ a_27233_5058# 2.3e-19
C1692 a_26367_4790# a_27233_5058# 0.034054f
C1693 a_26808_4902# a_26640_5156# 0.239923f
C1694 ringtest_0.x4._05_ ringtest_0.x4.net7 0.232588f
C1695 ringtest_0.x4._17_ a_26749_6422# 8.24e-19
C1696 ringtest_0.x4._14_ a_22765_5308# 1.74e-20
C1697 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x1.nSEL1 0.352716f
C1698 ringtest_0.x4._06_ a_24800_5334# 3.32e-19
C1699 ringtest_0.x4.net8 a_27065_5334# 1.1e-19
C1700 ringtest_0.x4._11_ a_26367_5340# 2.03e-20
C1701 ringtest_0.x4._17_ ringtest_0.x4._05_ 0.0576f
C1702 a_24699_6200# a_24527_5340# 1.08e-19
C1703 a_27489_3702# VDPWR 0.290806f
C1704 muxtest_0.x2.x1.nSEL1 a_12425_24040# 9.57e-19
C1705 a_22392_5990# VDPWR 0.176029f
C1706 a_11845_23906# a_12019_24012# 0.006584f
C1707 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN1 0.034862f
C1708 ringtest_0.x4._08_ a_26640_5334# 0.030723f
C1709 ui_in[2] ui_in[5] 0.211146f
C1710 a_24287_6422# VDPWR 0.004431f
C1711 ringtest_0.x4._13_ ringtest_0.x4._14_ 0.074354f
C1712 ringtest_0.x4.clknet_0_clk a_24699_6200# 0.034583f
C1713 a_21509_4790# a_22043_5156# 0.002698f
C1714 ringtest_0.x4._15_ a_25393_5308# 0.031321f
C1715 ringtest_0.x4._03_ a_21863_4790# 0.13856f
C1716 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ui_in[4] 1.2e-19
C1717 ringtest_0.x4.counter[0] ringtest_0.x4.counter[1] 0.079742f
C1718 ringtest_0.x4._22_ a_25547_4612# 0.002069f
C1719 uio_in[3] uio_in[2] 0.031023f
C1720 a_21981_8976# a_21395_6940# 1.29e-20
C1721 muxtest_0.x1.x4.A ua[3] 6.48818f
C1722 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 0.173286f
C1723 muxtest_0.x2.nselect2 VDPWR 1.22451f
C1724 a_17231_12017# VDPWR 0.217593f
C1725 a_22052_8875# ringtest_0.x4._12_ 0.032034f
C1726 ringtest_0.x4.net8 a_26627_4246# 4.33e-20
C1727 ringtest_0.x4._11_ a_22765_4478# 0.159397f
C1728 ringtest_0.x4.net9 ringtest_0.x4._09_ 0.571636f
C1729 a_24361_5340# a_24317_4942# 1.28e-19
C1730 ringtest_0.x4._11_ a_27065_5156# 3.81e-21
C1731 muxtest_0.x2.x2.GN1 ua[0] 2.35e-19
C1732 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A 0.17253f
C1733 ringtest_0.x3.x2.GN2 m3_17036_9140# 0.099332f
C1734 muxtest_0.x1.x3.GN1 muxtest_0.x1.x5.A 0.4308f
C1735 a_23770_5308# a_23899_5334# 0.062574f
C1736 a_24536_6699# ringtest_0.x4.net8 5.83e-19
C1737 ringtest_0.x4._11_ a_23949_6654# 8.65e-19
C1738 a_26640_5334# VDPWR 0.246903f
C1739 ringtest_0.x4.clknet_1_1__leaf_clk a_26269_4612# 3.29e-19
C1740 ringtest_0.x4.net6 a_25977_4220# 0.009771f
C1741 a_19666_31955# a_19842_32287# 0.185422f
C1742 a_19114_31955# muxtest_0.x1.x3.GN1 0.012335f
C1743 ringtest_0.x4._15_ a_26808_4902# 0.002208f
C1744 a_25336_4902# a_25149_4220# 3.07e-19
C1745 ringtest_0.x4.net7 ringtest_0.x4._09_ 2.46e-19
C1746 a_24336_6544# ringtest_0.x4.net6 0.001918f
C1747 a_12425_24040# muxtest_0.x2.x2.GN3 5.17e-20
C1748 muxtest_0.x2.x2.GN2 a_12977_24040# 3.11e-20
C1749 a_21948_5156# a_22021_4220# 3.53e-19
C1750 a_22116_4902# a_22164_4362# 5.83e-19
C1751 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN3 0.002859f
C1752 muxtest_0.x2.x2.GP2 ua[3] 0.085048f
C1753 a_18662_32213# ui_in[2] 4.33e-19
C1754 m3_13302_19985# m3_13316_18955# 0.003741f
C1755 ringtest_0.x4.net3 a_21587_5334# 0.003111f
C1756 a_11845_23906# ui_in[4] 0.02803f
C1757 ringtest_0.x4.counter[9] ringtest_0.x4.counter[8] 0.299988f
C1758 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN2 0.154394f
C1759 a_25149_4220# VDPWR 0.405422f
C1760 m2_18699_31802# ui_in[2] 4.4e-19
C1761 a_21465_9294# VDPWR 0.413258f
C1762 a_26735_5156# VDPWR 0.002923f
C1763 ringtest_0.x4._10_ a_21867_8054# 4.63e-20
C1764 a_22649_6244# a_22733_6244# 0.008508f
C1765 ringtest_0.x4.net9 a_27659_4246# 3.29e-19
C1766 a_21785_8054# a_21939_8054# 0.004009f
C1767 ringtest_0.x4._11_ a_24004_6128# 0.043142f
C1768 ringtest_0.x4._19_ a_24361_5340# 9.86e-21
C1769 ringtest_0.x4._08_ a_25364_5878# 0.011527f
C1770 muxtest_0.R7R8 muxtest_0.R6R7 2.27687f
C1771 a_24329_6640# VDPWR 0.427982f
C1772 a_24287_6422# ringtest_0.x4._21_ 1.26e-19
C1773 ringtest_0.x4.net2 a_21233_5340# 3.28e-19
C1774 a_21852_8720# ringtest_0.x4._11_ 4.06e-19
C1775 ringtest_0.x4.net6 a_24986_5878# 0.001357f
C1776 ringtest_0.x4._12_ a_21803_8598# 1.13e-19
C1777 a_22052_8875# a_22245_8054# 2.48e-20
C1778 muxtest_0.x1.x3.GN3 muxtest_0.R2R3 0.27459f
C1779 muxtest_0.x2.x2.GP2 m3_13316_18955# 2.65e-20
C1780 muxtest_0.x1.x3.GN3 ui_in[1] 0.273672f
C1781 ringtest_0.x4.clknet_0_clk a_25421_6641# 0.012442f
C1782 a_21465_8830# a_21561_8830# 0.310858f
C1783 ringtest_0.x4.net6 a_22139_5878# 5.63e-21
C1784 ringtest_0.x4.net2 ringtest_0.x4._11_ 0.001125f
C1785 ringtest_0.x4._11_ a_23963_4790# 0.001879f
C1786 a_25364_5878# a_25336_4902# 2.72e-20
C1787 a_24699_6200# a_25168_5156# 5.18e-21
C1788 a_22052_9116# a_22201_9142# 0.005525f
C1789 a_21981_9142# a_21780_9142# 4.67e-20
C1790 ringtest_0.x4.net11 a_26627_4246# 2.78e-19
C1791 ringtest_0.x4._16_ ringtest_0.x4._03_ 0.005745f
C1792 ringtest_0.x3.x1.nSEL0 m2_15612_11606# 3.43e-19
C1793 ringtest_0.x4._18_ a_21951_5878# 8.49e-20
C1794 a_21561_9116# a_21981_9142# 0.036838f
C1795 a_21852_9416# a_22052_9116# 0.074815f
C1796 ringtest_0.counter7 a_26895_3867# 0.110188f
C1797 a_22224_6244# ringtest_0.x4.net5 1.47e-19
C1798 ringtest_0.x3.x1.nSEL0 ui_in[3] 0.324822f
C1799 ringtest_0.x4._11_ a_23381_4818# 0.163973f
C1800 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN3 1.7e-19
C1801 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN2 0.209954f
C1802 ringtest_0.x4.net1 a_21465_9294# 0.045364f
C1803 ringtest_0.x4._18_ a_24883_6800# 2.19e-20
C1804 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN1 0.002605f
C1805 a_24545_5878# VDPWR 0.011033f
C1806 ringtest_0.x4._06_ a_23993_5654# 6.56e-20
C1807 ringtest_0.x4._13_ a_21509_4790# 6.65e-20
C1808 ringtest_0.x4._15_ a_25083_4790# 7.24e-21
C1809 ringtest_0.x4._11_ a_22181_5334# 7.61e-19
C1810 ringtest_0.x4._16_ a_23770_5308# 0.01721f
C1811 ringtest_0.x4.net9 a_24361_5340# 5.55e-19
C1812 a_24536_6699# ringtest_0.x4._05_ 3.36e-19
C1813 a_24895_4790# a_25677_5156# 3.14e-19
C1814 a_25364_5878# VDPWR 1.34839f
C1815 a_25083_4790# a_25263_5156# 0.001229f
C1816 muxtest_0.x2.x2.GN4 ui_in[4] 0.063283f
C1817 ringtest_0.counter7 ua[1] 5.26868f
C1818 ringtest_0.x4._22_ ringtest_0.x4._07_ 0.503878f
C1819 ringtest_0.x4.net2 a_21675_4790# 3.95e-20
C1820 ringtest_0.drv_out a_25225_5334# 2.32e-21
C1821 muxtest_0.x2.nselect2 a_12849_23648# 1.29e-19
C1822 ringtest_0.x4._14_ ringtest_0.x4.counter[1] 1.03e-21
C1823 a_21981_8976# VDPWR 0.210717f
C1824 ringtest_0.x4.net6 a_23899_5334# 0.044713f
C1825 ringtest_0.x4._15_ a_24715_5334# 0.019231f
C1826 ringtest_0.x4._22_ a_25055_3867# 8.8e-19
C1827 ringtest_0.x4._14_ a_22390_4566# 0.122283f
C1828 a_22116_4902# a_22373_5156# 0.036838f
C1829 a_27065_5334# ringtest_0.x4._09_ 0.001217f
C1830 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ui_in[4] 2.29e-19
C1831 ringtest_0.x4.net7 a_24361_5340# 0.088061f
C1832 a_24135_3867# a_25055_3867# 1.37e-20
C1833 a_21785_5878# a_24004_6128# 1.89e-21
C1834 muxtest_0.R6R7 muxtest_0.R5R6 2.03637f
C1835 ringtest_0.x4._04_ a_24070_5852# 8.65e-21
C1836 a_22399_8976# ringtest_0.x4._11_ 0.001319f
C1837 a_24551_4790# VDPWR 6.66e-20
C1838 ringtest_0.x4.net8 a_26721_4246# 6.89e-20
C1839 muxtest_0.x1.x3.GP2 muxtest_0.R2R3 4.15159f
C1840 ringtest_0.x4._11_ a_26375_4612# 0.001561f
C1841 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A 5.04e-19
C1842 ringtest_0.x4._17_ a_24361_5340# 1.12e-20
C1843 muxtest_0.x1.x3.GP2 ui_in[1] 3.1e-20
C1844 ringtest_0.counter3 a_22765_4478# 8.56e-20
C1845 a_21561_8830# a_21780_8964# 0.006169f
C1846 a_21465_8830# a_21049_8598# 5.03e-19
C1847 muxtest_0.x1.x3.GP3 muxtest_0.x1.x5.A 0.358703f
C1848 a_24317_4942# VDPWR 0.220214f
C1849 muxtest_0.x1.x3.GN4 muxtest_0.R7R8 0.13848f
C1850 muxtest_0.R6R7 VDPWR 1.6078f
C1851 a_26808_5308# a_27191_5712# 4.67e-20
C1852 a_26367_5340# ringtest_0.x4.net10 5.04e-19
C1853 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A 5.04e-19
C1854 ringtest_0.x4.clknet_1_0__leaf_clk a_21845_8816# 0.683552f
C1855 ringtest_0.x4.net4 a_22164_4362# 0.007901f
C1856 a_24329_6640# ringtest_0.x4._21_ 8.19e-20
C1857 a_22399_9142# a_21852_8720# 4.5e-20
C1858 a_23151_5334# VDPWR 0.008519f
C1859 ringtest_0.x4.net2 a_21785_5878# 2.26e-20
C1860 ringtest_0.x4._15_ a_25547_4612# 5.62e-21
C1861 ringtest_0.x4.net1 a_21981_8976# 0.001727f
C1862 ua[3] ua[0] 1.8361f
C1863 ringtest_0.x4._11_ ringtest_0.x4._20_ 0.174111f
C1864 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP2 1.7e-20
C1865 ringtest_0.x4._09_ a_26627_4246# 0.001692f
C1866 ringtest_0.x4.clknet_1_1__leaf_clk a_24883_6800# 3.41e-20
C1867 ringtest_0.x4.net2 a_22399_9142# 1.04e-19
C1868 a_21425_9686# a_21465_9294# 1.32e-19
C1869 ringtest_0.x4._00_ a_21507_9686# 6.18e-19
C1870 ringtest_0.x4._09_ a_27149_5156# 6.12e-19
C1871 ringtest_0.x4._04_ a_22373_5156# 0.001409f
C1872 ringtest_0.x4._07_ a_25225_5334# 0.009837f
C1873 ringtest_0.x4._02_ a_21399_5340# 0.275992f
C1874 a_21233_5340# a_21840_5308# 0.141453f
C1875 ringtest_0.x4._22_ a_26201_5340# 5.82e-21
C1876 ringtest_0.x3.x2.GP2 ua[1] 0.349381f
C1877 ringtest_0.x4.clknet_1_0__leaf_clk a_22373_5156# 6.12e-19
C1878 ringtest_0.counter7 a_26555_4790# 2.77e-20
C1879 muxtest_0.R3R4 muxtest_0.x2.x2.GP3 4.09931f
C1880 ringtest_0.x4._18_ a_24045_6654# 2.33e-19
C1881 a_23349_6422# a_24329_6640# 6.46e-21
C1882 a_22228_8598# VDPWR 0.004407f
C1883 ringtest_0.x4._21_ a_24545_5878# 0.053333f
C1884 a_13675_24012# ua[3] 3.17e-19
C1885 a_16755_12091# ringtest_0.x3.x2.GP2 3.2e-20
C1886 a_23879_6940# a_24329_6640# 0.022305f
C1887 ringtest_0.x4._20_ a_25761_5058# 3.47e-20
C1888 ringtest_0.x4.clknet_1_0__leaf_clk a_21767_5334# 0.001355f
C1889 ringtest_0.x4._11_ a_21840_5308# 0.005658f
C1890 muxtest_0.x2.x2.GN3 ua[3] 0.087947f
C1891 ringtest_0.x4.net10 a_27065_5156# 0.003817f
C1892 a_26913_4566# VDPWR 4.13e-19
C1893 ringtest_0.ring_out VDPWR 4.36398f
C1894 ringtest_0.counter3 m3_17032_8096# 0.119717f
C1895 a_25364_5878# ringtest_0.x4._21_ 3.33e-20
C1896 a_16027_11759# a_16203_12091# 0.185422f
C1897 a_22116_4902# a_22499_4790# 4.67e-20
C1898 a_24135_3867# ringtest_0.x4.counter[5] 4.98e-19
C1899 ringtest_0.x4.clknet_1_1__leaf_clk a_26808_5308# 5.16e-19
C1900 ringtest_0.x4._08_ ringtest_0.x4.net9 0.003243f
C1901 ringtest_0.x4._19_ VDPWR 0.188083f
C1902 ringtest_0.x4.net6 a_22097_5334# 5.09e-19
C1903 ringtest_0.x4.clknet_0_clk a_26007_6788# 5.18e-20
C1904 ringtest_0.x4.net6 ringtest_0.x4._16_ 0.291584f
C1905 muxtest_0.x1.x3.GN4 muxtest_0.R5R6 0.304696f
C1906 ringtest_0.x4._23_ a_26895_3867# 7.52e-20
C1907 muxtest_0.x2.x2.GN3 m3_13316_18955# 0.016026f
C1908 a_27273_4220# a_27303_4246# 0.025037f
C1909 ringtest_0.x4.clknet_1_0__leaf_clk a_22201_8964# 4.64e-19
C1910 ringtest_0.x4._16_ a_24895_4790# 4.88e-21
C1911 ringtest_0.x4.net2 ringtest_0.counter3 0.003151f
C1912 a_23879_6940# a_24545_5878# 2.81e-20
C1913 a_26735_5334# VDPWR 0.002923f
C1914 ringtest_0.counter7 m3_17046_7066# 0.117708f
C1915 a_21840_5308# a_21675_4790# 3.46e-19
C1916 ringtest_0.x4.net9 a_25336_4902# 0.007121f
C1917 a_21399_5340# a_22116_4902# 0.001879f
C1918 ringtest_0.drv_out ringtest_0.x4._15_ 0.005511f
C1919 ringtest_0.x4._00_ a_21852_8720# 4.06e-19
C1920 ringtest_0.counter7 ringtest_0.x4.counter[6] 0.087745f
C1921 ringtest_0.x4.net7 ringtest_0.x4._08_ 1.97e-19
C1922 ringtest_0.x4._21_ a_24317_4942# 0.011629f
C1923 muxtest_0.x1.x3.GN4 VDPWR 1.35388f
C1924 a_25225_5334# a_26201_5340# 1.07e-19
C1925 a_22265_5308# a_22223_5712# 7.84e-20
C1926 a_25393_5308# a_26367_5340# 2.73e-19
C1927 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN2 0.142718f
C1928 ringtest_0.x4._19_ ringtest_0.x4._25_ 9.05e-21
C1929 a_22265_5308# VDPWR 0.418555f
C1930 ringtest_0.x4.net2 ringtest_0.x4._00_ 0.002662f
C1931 a_23529_6422# a_23619_6788# 0.004764f
C1932 muxtest_0.x1.x1.nSEL1 a_19666_31955# 7.84e-19
C1933 ringtest_0.x4.net4 a_22373_5156# 0.022715f
C1934 ringtest_0.x4.clknet_1_1__leaf_clk a_26555_4790# 6.27e-19
C1935 ringtest_0.x4.net7 a_25336_4902# 0.005145f
C1936 ringtest_0.x4.net9 VDPWR 0.934233f
C1937 ringtest_0.x4.net3 ringtest_0.x4._03_ 0.019455f
C1938 a_24045_6654# ringtest_0.x4.clknet_1_1__leaf_clk 1.54e-20
C1939 a_21509_4790# a_22390_4566# 3.11e-19
C1940 ui_in[6] ui_in[5] 6.4498f
C1941 ringtest_0.x3.x2.GN2 ua[1] 0.42933f
C1942 ringtest_0.x4._06_ a_23837_5878# 4.79e-19
C1943 ringtest_0.x4._06_ ringtest_0.x4._22_ 0.004416f
C1944 a_16579_11759# ringtest_0.x3.x2.GN4 6.84e-19
C1945 a_24070_5852# a_23837_5878# 0.005961f
C1946 ringtest_0.x4._04_ a_21399_5340# 0.011144f
C1947 a_16755_12091# ringtest_0.x3.x2.GN2 5.62e-20
C1948 a_21785_5878# a_21840_5308# 0.002941f
C1949 a_21863_4790# ringtest_0.x4.net5 2.02e-19
C1950 a_24699_6200# a_24763_6143# 0.266837f
C1951 ringtest_0.x4._23_ a_26808_5308# 0.006211f
C1952 muxtest_0.R3R4 muxtest_0.R2R3 2.48395f
C1953 ringtest_0.x4.clknet_1_0__leaf_clk a_21399_5340# 0.158653f
C1954 ringtest_0.x4._18_ a_22795_5334# 4.57e-20
C1955 a_26201_5340# a_26640_5156# 1.73e-19
C1956 ringtest_0.x4.net7 VDPWR 1.78561f
C1957 a_26808_5308# a_26367_4790# 2.96e-21
C1958 a_26367_5340# a_26808_4902# 2.96e-21
C1959 ringtest_0.x4._11_ a_22392_5990# 0.032361f
C1960 a_21561_9116# ui_in[5] 2.06e-20
C1961 ringtest_0.x4._15_ ringtest_0.x4._07_ 0.022092f
C1962 ringtest_0.x4.net3 a_21939_8054# 8.45e-20
C1963 a_24336_6544# a_24527_5340# 6.46e-19
C1964 a_27273_4220# ringtest_0.x4.counter[8] 0.001844f
C1965 a_24536_6699# a_24361_5340# 2.08e-22
C1966 a_24329_6640# a_24968_5308# 2.9e-20
C1967 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A 0.173286f
C1968 muxtest_0.x1.x3.GN3 ui_in[4] 7.93e-20
C1969 ringtest_0.x4._17_ VDPWR 2.34858f
C1970 ringtest_0.x4._07_ a_25263_5156# 2.91e-19
C1971 ringtest_0.x3.x2.GP2 m3_17046_7066# 2.65e-20
C1972 ringtest_0.x3.x1.nSEL1 VDPWR 0.646724f
C1973 ringtest_0.x4._19_ ringtest_0.x4._21_ 7.87e-20
C1974 ringtest_0.x4.clknet_0_clk a_24336_6544# 0.025079f
C1975 a_21561_9116# ringtest_0.x4._12_ 1.23e-19
C1976 ringtest_0.x4._00_ a_22399_8976# 0.001531f
C1977 ringtest_0.x4.clknet_1_1__leaf_clk a_24699_6200# 7.2e-19
C1978 a_23963_4790# ringtest_0.x4.counter[4] 4.17e-20
C1979 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y 0.17253f
C1980 ui_in[3] ua[1] 4.1e-22
C1981 ringtest_0.x4.net6 a_22649_6244# 0.021756f
C1982 ringtest_0.x3.x2.GP3 ringtest_0.counter3 4.0653f
C1983 ui_in[1] ui_in[5] 0.187526f
C1984 ringtest_0.x4._09_ a_26721_4246# 2.04e-21
C1985 a_16755_12091# ui_in[3] 0.279858f
C1986 a_22021_4220# a_22164_4362# 0.221119f
C1987 ringtest_0.x4.net8 a_24729_4790# 0.009204f
C1988 ringtest_0.x4.net7 ringtest_0.x4._25_ 3.01e-19
C1989 a_27065_5156# a_27191_4790# 0.006169f
C1990 ringtest_0.x4._23_ a_26555_4790# 0.012973f
C1991 ringtest_0.x4.net4 a_22499_4790# 0.00133f
C1992 a_26808_4902# a_27065_5156# 0.036838f
C1993 a_26367_4790# a_26555_4790# 0.097994f
C1994 a_24329_6640# a_25925_6788# 2.69e-21
C1995 ringtest_0.x4._17_ ringtest_0.x4._25_ 1.89e-19
C1996 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP1 2.55932f
C1997 ringtest_0.x4._06_ a_25225_5334# 9.38e-20
C1998 a_23349_6422# ringtest_0.x4._19_ 0.001413f
C1999 ringtest_0.x4._11_ a_26640_5334# 6.96e-20
C2000 a_23879_6940# ringtest_0.x4._19_ 5.98e-19
C2001 ringtest_0.x4.counter[0] VDPWR 0.656838f
C2002 a_24699_6200# a_24800_5334# 0.001605f
C2003 a_12297_23648# muxtest_0.x2.x2.GN2 0.106178f
C2004 a_22817_6146# VDPWR 0.383645f
C2005 ringtest_0.x4._08_ a_27065_5334# 0.013878f
C2006 ringtest_0.x4.clknet_1_1__leaf_clk a_23809_4790# 2.42e-19
C2007 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VDPWR 0.787508f
C2008 a_26095_6788# VDPWR 0.002069f
C2009 ringtest_0.x4._21_ ringtest_0.x4.net9 0.170283f
C2010 ringtest_0.x4.net4 a_21399_5340# 0.002039f
C2011 ringtest_0.x3.nselect2 ui_in[4] 0.001177f
C2012 ringtest_0.x4.clknet_1_1__leaf_clk a_22795_5334# 7.11e-20
C2013 ringtest_0.x4._15_ a_26201_5340# 0.069151f
C2014 ringtest_0.x3.x1.nSEL0 a_16027_11759# 0.03096f
C2015 ringtest_0.x4.net6 a_21587_5334# 1.35e-20
C2016 ringtest_0.x4._22_ a_26269_4612# 6.12e-20
C2017 ringtest_0.x4._13_ a_22350_5878# 2.65e-20
C2018 a_17405_12123# VDPWR 7.45e-19
C2019 ringtest_0.x4._04_ a_21951_5878# 0.215918f
C2020 ua[2] ua[5] 0.002786f
C2021 a_21785_5878# a_22392_5990# 0.136461f
C2022 ringtest_0.x3.x2.GN3 VDPWR 0.649844f
C2023 muxtest_0.x1.x3.GP1 ua[3] 0.0076f
C2024 ringtest_0.x4._01_ ringtest_0.x4._12_ 0.353697f
C2025 ringtest_0.x4._11_ a_25149_4220# 2.67e-19
C2026 a_25925_6788# a_25364_5878# 0.010774f
C2027 ringtest_0.x4.net7 ringtest_0.x4._21_ 0.326643f
C2028 ringtest_0.x4.clknet_1_0__leaf_clk a_21951_5878# 0.020113f
C2029 ringtest_0.x3.x2.GN4 m3_17032_8096# 7.07e-19
C2030 a_26749_6422# a_26839_6788# 0.004764f
C2031 a_18662_32213# ui_in[1] 0.02803f
C2032 ringtest_0.x4._16_ ringtest_0.x4.net5 0.096932f
C2033 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP3 0.060268f
C2034 muxtest_0.x1.x3.GN1 muxtest_0.x1.x4.A 0.428132f
C2035 ringtest_0.x4._17_ ringtest_0.x4._21_ 0.019243f
C2036 a_23879_6940# ringtest_0.x4.net9 1.97e-19
C2037 ringtest_0.x4._08_ a_27149_5156# 1.22e-19
C2038 ringtest_0.x4._11_ a_24329_6640# 2.33e-19
C2039 a_20318_32213# a_20492_32319# 0.006584f
C2040 a_27065_5334# VDPWR 0.231069f
C2041 ringtest_0.x4._15_ a_22164_4362# 4.86e-20
C2042 ringtest_0.x4.net6 a_27273_4220# 4.97e-21
C2043 m2_18699_31802# ui_in[1] 0.183786f
C2044 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ui_in[3] 1.1e-22
C2045 a_19666_31955# muxtest_0.x1.x3.GN1 7.37e-20
C2046 muxtest_0.x1.x5.GN a_18662_32213# 0.001336f
C2047 ringtest_0.x4.clknet_1_1__leaf_clk a_25421_6641# 0.035969f
C2048 a_23529_6422# ringtest_0.x4._15_ 2e-21
C2049 a_24465_6800# ringtest_0.x4.net6 0.001158f
C2050 a_13501_23906# muxtest_0.R1R2 5.05e-21
C2051 a_23349_6422# ringtest_0.x4.net7 2.88e-19
C2052 a_23879_6940# ringtest_0.x4.net7 0.002812f
C2053 muxtest_0.x1.x5.GN m2_18699_31802# 4e-19
C2054 muxtest_0.x1.x3.GN3 ui_in[0] 0.254198f
C2055 a_19290_32287# ui_in[2] 1.22e-19
C2056 ringtest_0.x4._17_ a_23349_6422# 0.250762f
C2057 a_23879_6940# ringtest_0.x4._17_ 7.15e-19
C2058 ringtest_0.x4.net7 a_25309_5334# 0.001255f
C2059 a_12473_23980# ui_in[4] 0.254026f
C2060 ringtest_0.x4._11_ a_24545_5878# 1.22e-19
C2061 a_22201_9142# VDPWR 0.003202f
C2062 a_26627_4246# VDPWR 0.151674f
C2063 a_21852_9416# VDPWR 0.327097f
C2064 a_27149_5156# VDPWR 0.005027f
C2065 a_22817_6146# ringtest_0.x4._21_ 1.76e-19
C2066 muxtest_0.x1.x3.GN2 muxtest_0.R1R2 0.006936f
C2067 ringtest_0.x4._11_ a_25364_5878# 0.049204f
C2068 ui_in[2] ui_in[3] 0.170107f
C2069 a_24536_6699# VDPWR 0.264477f
C2070 muxtest_0.x1.x5.A muxtest_0.R6R7 4.52052f
C2071 ringtest_0.x4._12_ a_21785_8054# 0.001375f
C2072 ringtest_0.x4._01_ a_22245_8054# 0.014882f
C2073 ringtest_0.x4.net4 a_21951_5878# 0.34974f
C2074 ringtest_0.x4._15_ ringtest_0.x4._06_ 0.139237f
C2075 a_21561_8830# a_21845_8816# 0.030894f
C2076 a_21465_8830# a_21852_8720# 0.034054f
C2077 ringtest_0.x4._15_ a_24070_5852# 6.77e-20
C2078 ringtest_0.x4.net8 ringtest_0.x4._09_ 2.1e-20
C2079 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y 5.04e-19
C2080 a_25149_4220# a_25345_4612# 0.00119f
C2081 a_25593_5156# ringtest_0.x4.counter[6] 2e-19
C2082 ringtest_0.x4._23_ a_26817_4566# 4.18e-19
C2083 ringtest_0.x4._11_ a_24551_4790# 0.001398f
C2084 a_25364_5878# a_25761_5058# 0.001883f
C2085 ringtest_0.x4._18_ a_22224_6244# 5.13e-20
C2086 a_21675_9686# ringtest_0.x4.clknet_1_0__leaf_clk 2.59e-19
C2087 a_21845_9116# a_21981_9142# 0.141453f
C2088 a_21233_5340# a_23151_5334# 4.04e-20
C2089 a_21852_9416# a_21803_9508# 6.32e-19
C2090 ringtest_0.x4.net2 a_21465_8830# 0.004306f
C2091 a_22649_6244# ringtest_0.x4.net5 4.89e-20
C2092 ringtest_0.x4._11_ a_24317_4942# 0.046716f
C2093 a_25421_6641# ringtest_0.x4._23_ 1.03e-19
C2094 a_22111_10993# a_21845_9116# 6.9e-23
C2095 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._24_ 0.041474f
C2096 ringtest_0.x4.net1 a_21852_9416# 0.006588f
C2097 ringtest_0.x4._05_ a_26749_6422# 4.21e-20
C2098 ringtest_0.x4._14_ VDPWR 0.674773f
C2099 ringtest_0.x4.net10 a_27489_3702# 1.3e-21
C2100 ringtest_0.x4._15_ a_23891_4790# 1.25e-19
C2101 ringtest_0.x4.net6 a_26201_4790# 5.6e-22
C2102 a_13025_23980# muxtest_0.x2.x2.GP3 5.21e-19
C2103 ringtest_0.x4._11_ a_23151_5334# 0.00137f
C2104 ringtest_0.x4._16_ a_24527_5340# 9.89e-20
C2105 ringtest_0.x4.net9 a_24968_5308# 2.05e-20
C2106 muxtest_0.x1.x3.GP2 ui_in[0] 4.71e-19
C2107 ringtest_0.x3.x2.GN4 ringtest_0.x3.x2.GP3 3.4436f
C2108 a_22319_6244# VDPWR 0.003715f
C2109 a_25336_4902# a_25294_4790# 4.62e-19
C2110 a_24895_4790# a_26201_4790# 3.23e-19
C2111 ringtest_0.x4._15_ a_22373_5156# 1.6e-20
C2112 muxtest_0.x2.nselect2 a_13501_23906# 9.77e-20
C2113 ringtest_0.x4.clknet_0_clk ringtest_0.x4._16_ 0.019509f
C2114 ringtest_0.x4.net5 a_23467_4818# 2.72e-19
C2115 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VDPWR 0.639974f
C2116 ringtest_0.x4.net6 a_26555_5334# 3.93e-20
C2117 muxtest_0.R7R8 muxtest_0.x2.x2.GN2 1.22e-19
C2118 ringtest_0.x4._22_ a_26895_3867# 1.85e-19
C2119 muxtest_0.R3R4 ui_in[4] 3.8e-21
C2120 a_22392_5990# a_22775_5878# 4.67e-20
C2121 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x2.GN2 3.88e-22
C2122 clk ena 0.031023f
C2123 a_22541_5058# a_22373_5156# 0.310858f
C2124 ringtest_0.x4.net7 a_24968_5308# 0.040813f
C2125 a_25294_4790# VDPWR 9.98e-20
C2126 a_25055_3867# a_25975_3867# 1.37e-20
C2127 a_21785_8054# a_22245_8054# 0.001479f
C2128 a_24883_6800# ringtest_0.x4._22_ 0.001069f
C2129 ringtest_0.x4._12_ a_22695_8304# 0.001754f
C2130 ringtest_0.x4._17_ a_24968_5308# 1.03e-20
C2131 a_22043_5156# VDPWR 0.005794f
C2132 muxtest_0.x1.x3.GP3 muxtest_0.x1.x4.A 0.358376f
C2133 muxtest_0.x1.x3.GN4 muxtest_0.x1.x5.A 0.446595f
C2134 a_26640_5334# ringtest_0.x4.net10 3.33e-19
C2135 a_27233_5308# a_27191_5712# 7.84e-20
C2136 ringtest_0.x4.clknet_1_0__leaf_clk a_22052_8875# 0.037641f
C2137 ringtest_0.x4.net4 a_23381_4584# 0.083888f
C2138 ui_in[4] ui_in[5] 0.285451f
C2139 a_24536_6699# ringtest_0.x4._21_ 0.0043f
C2140 ringtest_0.x4._11_ ringtest_0.x4._19_ 0.032711f
C2141 ringtest_0.x4._15_ a_26269_4612# 0.00403f
C2142 a_19666_31955# muxtest_0.x1.x3.GP3 0.001353f
C2143 ringtest_0.x4._23_ ringtest_0.x4._24_ 0.206353f
C2144 ringtest_0.x4._00_ a_21465_9294# 0.001095f
C2145 a_21425_9686# a_21852_9416# 0.00324f
C2146 a_26749_6422# ringtest_0.x4._09_ 2.51e-21
C2147 ringtest_0.x4._24_ a_26367_4790# 0.03707f
C2148 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ui_in[3] 0.001551f
C2149 ringtest_0.x4.net7 a_25925_6788# 0.168744f
C2150 ringtest_0.x4._09_ ringtest_0.x4.net11 0.071633f
C2151 ringtest_0.x4.net3 ringtest_0.x4.net5 9.15e-21
C2152 ringtest_0.x4._22_ a_26808_5308# 9.3e-20
C2153 ringtest_0.x4._02_ a_21672_5334# 8.22e-19
C2154 a_21233_5340# a_22265_5308# 0.048748f
C2155 ringtest_0.x4._17_ a_25925_6788# 0.139841f
C2156 ringtest_0.x4._04_ a_22795_5334# 0.072162f
C2157 ringtest_0.x4._18_ a_24336_6544# 1.59e-19
C2158 ringtest_0.x4._10_ VDPWR 0.248739f
C2159 ringtest_0.x4.net8 a_24361_5340# 0.036074f
C2160 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP2 0.005192f
C2161 a_23879_6940# a_24536_6699# 0.007109f
C2162 ringtest_0.x4._20_ a_25083_4790# 5.09e-20
C2163 ringtest_0.x4._11_ a_22265_5308# 0.033019f
C2164 a_26721_4246# VDPWR 0.19107f
C2165 muxtest_0.x1.x4.A muxtest_0.R1R2 4.5214f
C2166 muxtest_0.x2.x1.nSEL0 ui_in[4] 0.13767f
C2167 a_22541_5058# a_22499_4790# 7.84e-20
C2168 a_16203_12091# a_16579_11759# 3.02e-19
C2169 ringtest_0.x3.x1.nSEL1 a_15749_12123# 0.00175f
C2170 ringtest_0.x4._11_ ringtest_0.x4.net9 0.233741f
C2171 muxtest_0.x1.x3.GN3 muxtest_0.x2.x2.GN4 8.02e-21
C2172 ringtest_0.x4.clknet_1_1__leaf_clk a_27233_5308# 9.45e-20
C2173 a_12977_24040# VDPWR 0.001496f
C2174 ringtest_0.x4.net6 a_23770_5308# 0.050235f
C2175 ringtest_0.x4.clknet_0_clk a_26201_6788# 6.75e-20
C2176 muxtest_0.x2.x2.GN2 VDPWR 0.601936f
C2177 a_24361_5340# a_24729_4790# 0.012779f
C2178 ringtest_0.x4.net3 a_21007_3867# 0.006292f
C2179 ringtest_0.x4.clknet_1_0__leaf_clk a_21803_8598# 0.002574f
C2180 a_24045_6654# a_23837_5878# 9.42e-20
C2181 a_24336_6544# a_24763_6143# 0.003687f
C2182 ringtest_0.x4._16_ a_25168_5156# 7.37e-22
C2183 a_21509_4790# VDPWR 0.73231f
C2184 ringtest_0.x4._11_ ringtest_0.x4.net7 0.966176f
C2185 ringtest_0.x4.net11 a_27659_4246# 0.004987f
C2186 a_22265_5308# a_21675_4790# 0.00183f
C2187 a_26640_5156# a_26895_3867# 6.36e-19
C2188 ringtest_0.x4.net9 a_25761_5058# 0.115737f
C2189 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A 0.17253f
C2190 ringtest_0.x4.net1 ringtest_0.x4._10_ 0.033245f
C2191 a_25925_6788# a_26095_6788# 0.001675f
C2192 ringtest_0.x4._11_ ringtest_0.x4._17_ 0.113734f
C2193 a_26201_5340# a_26367_5340# 0.970499f
C2194 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GP1 1.17e-19
C2195 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN4 2.26e-20
C2196 ringtest_0.x4.clknet_1_1__leaf_clk a_25977_4220# 3.39e-19
C2197 a_22765_5308# VDPWR 0.250093f
C2198 muxtest_0.x1.x5.GN a_18836_32319# 1.95e-19
C2199 ringtest_0.x4._16_ a_22983_5654# 3.98e-19
C2200 a_23949_6654# a_24264_6788# 7.84e-20
C2201 a_25364_5878# ringtest_0.x4.net10 3.58e-19
C2202 ringtest_0.x4.net7 a_25761_5058# 0.064911f
C2203 a_12297_23648# muxtest_0.x2.x2.GP1 9.92e-19
C2204 ringtest_0.x4._03_ a_22939_4584# 1.17e-19
C2205 a_24336_6544# ringtest_0.x4.clknet_1_1__leaf_clk 0.013843f
C2206 a_21867_8054# VDPWR 1.13e-19
C2207 ringtest_0.x4.net4 a_22795_5334# 0.005199f
C2208 a_24627_6200# a_24545_5878# 2.78e-19
C2209 a_24763_6143# a_24986_5878# 3.74e-19
C2210 ringtest_0.x3.x2.GN2 a_16155_12151# 0.002418f
C2211 a_17231_12017# ringtest_0.x3.x2.GN4 0.134079f
C2212 ringtest_0.x4._13_ VDPWR 0.524307f
C2213 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN2 0.065153f
C2214 ua[3] ua[1] 0.003505f
C2215 a_21785_5878# a_22265_5308# 4.12e-19
C2216 ringtest_0.x4._22_ ringtest_0.x4.counter[6] 9.35e-22
C2217 ringtest_0.x4._04_ a_21672_5334# 3.3e-20
C2218 a_24699_6200# ringtest_0.x4._22_ 0.019192f
C2219 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VDPWR 0.636657f
C2220 ui_in[0] ui_in[5] 0.21609f
C2221 ringtest_0.x4._23_ a_27233_5308# 1.75e-20
C2222 ringtest_0.x4.clknet_1_0__leaf_clk a_21672_5334# 0.032164f
C2223 a_26201_5340# a_27065_5156# 1.29e-19
C2224 a_26640_5334# a_26808_4902# 3.15e-19
C2225 a_26808_5308# a_26640_5156# 3.15e-19
C2226 ringtest_0.x4._18_ a_23899_5334# 3.94e-20
C2227 muxtest_0.x1.x4.A muxtest_0.x2.nselect2 0.01287f
C2228 ringtest_0.x4._16_ a_22486_4246# 0.00427f
C2229 ringtest_0.x4._11_ a_22817_6146# 0.052724f
C2230 a_21845_9116# ui_in[5] 1.25e-19
C2231 ringtest_0.x4.net9 a_25345_4612# 0.001755f
C2232 a_24336_6544# a_24800_5334# 9.47e-20
C2233 ringtest_0.x4._08_ ringtest_0.x4.net8 2.38e-19
C2234 ringtest_0.x4._11_ a_26095_6788# 0.001703f
C2235 muxtest_0.x2.x2.GP3 ui_in[3] 4.18e-19
C2236 ringtest_0.x4.net3 ringtest_0.x4._12_ 0.271994f
C2237 muxtest_0.x1.x3.GN2 muxtest_0.R6R7 4.03742f
C2238 ringtest_0.x4._15_ a_26895_3867# 0.006207f
C2239 ringtest_0.x4.net1 a_21867_8054# 0.00162f
C2240 ringtest_0.x4.clknet_0_clk a_24465_6800# 0.003343f
C2241 a_21845_9116# ringtest_0.x4._12_ 2.52e-19
C2242 ringtest_0.x4._07_ a_23381_4818# 2.73e-21
C2243 ringtest_0.x3.x2.GN1 m2_15612_11606# 0.06935f
C2244 ringtest_0.x4._09_ a_27659_4246# 2.25e-19
C2245 ringtest_0.counter7 ringtest_0.x4.counter[9] 2.14e-19
C2246 ringtest_0.x3.x2.GN1 ui_in[3] 0.021168f
C2247 ringtest_0.drv_out ringtest_0.x3.x2.GP3 0.077808f
C2248 ringtest_0.x4._23_ a_25977_4220# 0.130093f
C2249 ringtest_0.x4.net8 a_25336_4902# 0.00264f
C2250 ringtest_0.x4._17_ a_21785_5878# 1.5e-21
C2251 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A ui_in[3] 1.61e-19
C2252 muxtest_0.x1.x3.GP3 ua[0] 0.17111f
C2253 a_26640_5156# a_26555_4790# 0.037333f
C2254 a_27233_5058# a_27065_5156# 0.310858f
C2255 a_21951_5878# a_22541_5058# 8.13e-20
C2256 ringtest_0.x4.clknet_1_1__leaf_clk a_25677_5156# 1.62e-19
C2257 ringtest_0.x4.net10 a_26913_4566# 0.002966f
C2258 ringtest_0.x4.net6 a_24895_4790# 0.045685f
C2259 a_12849_23648# a_12977_24040# 0.004764f
C2260 a_25364_5878# a_25393_5308# 0.009572f
C2261 a_12849_23648# muxtest_0.x2.x2.GN2 1.63e-19
C2262 ringtest_0.x4.net8 VDPWR 1.74959f
C2263 a_23529_6422# a_23949_6654# 0.017007f
C2264 a_24729_4790# a_25336_4902# 0.141453f
C2265 ui_in[3] ui_in[6] 0.135749f
C2266 a_18662_32213# ui_in[0] 0.048888f
C2267 a_26839_6788# VDPWR 6.35e-19
C2268 ringtest_0.x4.net4 a_21672_5334# 4.27e-19
C2269 ringtest_0.x4.clknet_1_1__leaf_clk a_23899_5334# 0.001857f
C2270 ringtest_0.x3.x1.nSEL0 a_16579_11759# 1.91e-20
C2271 ringtest_0.x4._15_ a_26808_5308# 4.57e-19
C2272 ringtest_0.x4._03_ ringtest_0.x4.net5 3.86e-19
C2273 m2_18699_31802# ui_in[0] 0.130999f
C2274 ringtest_0.x4._22_ a_26817_4566# 1.37e-20
C2275 a_21785_5878# a_22817_6146# 0.048608f
C2276 ringtest_0.x4._04_ a_22224_6244# 0.01404f
C2277 ringtest_0.x4.net10 a_26735_5334# 8.52e-20
C2278 a_24729_4790# VDPWR 0.721729f
C2279 ringtest_0.x4.net3 a_22245_8054# 0.001478f
C2280 muxtest_0.R1R2 ua[0] 2.31469f
C2281 ringtest_0.x4._11_ a_26627_4246# 0.054652f
C2282 a_21845_9116# a_22245_8054# 4.52e-21
C2283 ringtest_0.x4.clknet_1_0__leaf_clk a_22224_6244# 0.002436f
C2284 a_25364_5878# a_26808_4902# 7.13e-20
C2285 ringtest_0.x4._07_ ringtest_0.x4._20_ 1.72e-19
C2286 ringtest_0.x4._18_ ringtest_0.x4._16_ 0.283975f
C2287 ringtest_0.x4._25_ a_26839_6788# 8.17e-20
C2288 a_19290_32287# ui_in[1] 0.254026f
C2289 a_26749_6422# ringtest_0.x4._08_ 0.001905f
C2290 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A 5.04e-19
C2291 a_24968_5308# a_25351_5712# 4.67e-20
C2292 a_21465_9294# a_21465_8830# 0.025128f
C2293 ringtest_0.x4._11_ a_24536_6699# 3.53e-20
C2294 a_23949_6654# a_24070_5852# 0.002561f
C2295 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP1 2.99928f
C2296 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GN4 0.057602f
C2297 a_21798_5712# VDPWR 4.21e-19
C2298 ringtest_0.x4._15_ a_23381_4584# 0.110742f
C2299 a_19242_32347# VDPWR 5.13e-19
C2300 ringtest_0.x4.net9 ringtest_0.x4.net10 0.022804f
C2301 ringtest_0.x4.net6 a_27169_6641# 1.17e-21
C2302 ui_in[1] ui_in[3] 0.006066f
C2303 ui_in[2] ua[3] 0.781024f
C2304 ringtest_0.x4._15_ a_26555_4790# 0.005742f
C2305 a_25593_5156# a_25977_4220# 0.009905f
C2306 muxtest_0.x1.x5.GN a_19290_32287# 3.26e-19
C2307 a_24045_6654# ringtest_0.x4._15_ 1.09e-20
C2308 a_25593_5156# a_25719_4790# 0.006169f
C2309 ringtest_0.x4._14_ a_21233_5340# 0.001276f
C2310 a_22373_5156# a_22765_4478# 0.001309f
C2311 ringtest_0.x4.counter[1] VDPWR 0.336981f
C2312 muxtest_0.R3R4 muxtest_0.x2.x2.GN4 0.269437f
C2313 a_24763_6143# ringtest_0.x4._16_ 0.060109f
C2314 m3_17036_9140# m3_17032_8096# 0.003764f
C2315 ringtest_0.x4.net9 a_24627_6200# 0.004319f
C2316 ringtest_0.x4.net7 ringtest_0.x4.net10 6.54e-19
C2317 a_13025_23980# ui_in[4] 0.127717f
C2318 ringtest_0.x4._11_ ringtest_0.x4._14_ 0.007676f
C2319 muxtest_0.x2.x1.nSEL0 a_11845_23906# 0.081627f
C2320 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.nselect2 0.047548f
C2321 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VDPWR 0.636415f
C2322 a_22390_4566# VDPWR 0.007441f
C2323 ringtest_0.x4._16_ a_22295_3867# 4.24e-19
C2324 a_26749_6422# VDPWR 0.176006f
C2325 a_24004_6128# ringtest_0.x4._06_ 0.111795f
C2326 a_22052_9116# VDPWR 0.285583f
C2327 ringtest_0.x4.net11 VDPWR 0.783893f
C2328 ringtest_0.x4.net8 ringtest_0.x4._21_ 0.333812f
C2329 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A a_16027_11759# 2.51e-19
C2330 ringtest_0.x4._11_ a_22319_6244# 0.00121f
C2331 ringtest_0.counter3 ringtest_0.x4.counter[0] 0.117902f
C2332 a_24070_5852# a_24004_6128# 0.221119f
C2333 a_24329_6640# a_24715_5334# 6.17e-21
C2334 ringtest_0.x4._05_ VDPWR 0.236897f
C2335 ringtest_0.x4._24_ ringtest_0.x4._22_ 0.01067f
C2336 ringtest_0.x4.net4 a_22224_6244# 0.034877f
C2337 ringtest_0.x4._23_ ringtest_0.x4.counter[9] 7.62e-19
C2338 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._16_ 0.001692f
C2339 ringtest_0.x4.net3 a_21591_6128# 0.001185f
C2340 a_21465_8830# a_21981_8976# 1.28e-19
C2341 a_21845_8816# a_21852_8720# 0.969092f
C2342 ringtest_0.x4.net6 a_23932_6128# 0.002624f
C2343 ringtest_0.x4._15_ a_24699_6200# 2.91e-20
C2344 ringtest_0.x4.net3 a_22486_4246# 1.66e-19
C2345 ringtest_0.x4._17_ a_24627_6200# 4.44e-20
C2346 ringtest_0.x4._23_ a_27491_4566# 3.52e-19
C2347 a_25149_4220# a_25547_4612# 0.005781f
C2348 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP2 4.55678f
C2349 ringtest_0.x4.clknet_1_0__leaf_clk a_21780_9142# 0.001704f
C2350 ringtest_0.x4._11_ a_25294_4790# 0.002651f
C2351 ringtest_0.x4._21_ a_24729_4790# 5.62e-21
C2352 ringtest_0.x4._14_ a_21675_4790# 5.98e-19
C2353 ringtest_0.x3.x2.GN3 ringtest_0.counter3 3.89796f
C2354 a_26749_6422# ringtest_0.x4._25_ 0.082413f
C2355 ringtest_0.x4.counter[0] ua[2] 1.11e-19
C2356 a_21852_9416# a_22399_9142# 0.095025f
C2357 ringtest_0.x4.net2 a_21845_8816# 3.07e-19
C2358 a_21845_9116# a_22228_9508# 0.002698f
C2359 a_21561_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.038899f
C2360 ringtest_0.x4._08_ ringtest_0.x4._09_ 0.013938f
C2361 ringtest_0.x4._18_ a_22649_6244# 3.43e-19
C2362 a_23879_6940# ringtest_0.x4.net8 0.001938f
C2363 ringtest_0.x4._11_ a_22043_5156# 6.67e-19
C2364 ringtest_0.ring_out ringtest_0.x3.x2.GN4 0.080391f
C2365 ringtest_0.x4.net1 a_22052_9116# 0.002893f
C2366 ringtest_0.drv_out a_17231_12017# 3.86e-20
C2367 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A ui_in[3] 5.64e-20
C2368 ringtest_0.x4._05_ ringtest_0.x4._25_ 4.6e-21
C2369 ringtest_0.x4.net8 a_25309_5334# 9.28e-20
C2370 ua[2] ua[4] 0.002786f
C2371 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GP3 0.002439f
C2372 ringtest_0.x4._16_ a_24800_5334# 0.00213f
C2373 ringtest_0.x4.net9 a_25393_5308# 0.007609f
C2374 a_25593_5156# a_25677_5156# 0.008508f
C2375 ringtest_0.x4._08_ a_26766_5712# 0.001882f
C2376 a_22350_5878# VDPWR 3.37e-19
C2377 ringtest_0.x4.clknet_0_clk a_23770_5308# 8.98e-21
C2378 ringtest_0.x4._15_ a_23809_4790# 0.080244f
C2379 ringtest_0.x4.net6 ringtest_0.x4.net5 0.003368f
C2380 muxtest_0.x2.nselect2 muxtest_0.x2.x2.GN3 7.39e-21
C2381 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN4 2.26e-20
C2382 ringtest_0.x3.x2.GP2 ui_in[4] 1.37e-19
C2383 ringtest_0.x4.net6 a_24895_5334# 0.001259f
C2384 a_22817_6146# a_22775_5878# 7.84e-20
C2385 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A a_16579_11759# 2.51e-19
C2386 ringtest_0.x3.x1.nSEL1 a_15575_12017# 0.193944f
C2387 a_17377_14114# ui_in[6] 0.040112f
C2388 a_22541_5058# a_23809_4790# 3.71e-21
C2389 ringtest_0.x4.counter[1] ringtest_0.x4.counter[2] 0.070133f
C2390 a_22116_4902# a_21863_4790# 3.39e-19
C2391 ringtest_0.x4.net7 a_25393_5308# 0.08513f
C2392 muxtest_0.x2.x2.GP1 VDPWR 1.85798f
C2393 ringtest_0.x4._10_ ringtest_0.x4._11_ 0.033565f
C2394 ringtest_0.x4._09_ VDPWR 0.254927f
C2395 a_21785_5878# a_22319_6244# 0.002698f
C2396 a_25975_3867# a_26895_3867# 1.37e-20
C2397 ringtest_0.x4._04_ a_22139_5878# 0.126198f
C2398 ringtest_0.x4._11_ a_26721_4246# 0.039972f
C2399 ringtest_0.x4._23_ ringtest_0.x4._16_ 3.32e-22
C2400 a_22795_5334# a_22541_5058# 0.001352f
C2401 ringtest_0.x4._17_ a_25393_5308# 4.35e-22
C2402 a_12297_23648# VDPWR 0.161892f
C2403 ringtest_0.x4.clknet_1_0__leaf_clk a_22139_5878# 0.003123f
C2404 ringtest_0.x4.net9 a_27191_4790# 6.87e-19
C2405 a_21561_8830# a_21803_8598# 0.008508f
C2406 a_21981_8976# a_21780_8964# 4.67e-20
C2407 a_21845_8816# a_22399_8976# 0.057611f
C2408 a_21852_8720# a_22201_8964# 2.36e-19
C2409 a_22074_4790# VDPWR 0.003212f
C2410 ringtest_0.x4.net9 a_26808_4902# 0.022365f
C2411 ringtest_0.x3.x2.GP3 m3_17036_9140# 9.67e-19
C2412 a_23993_5654# a_23899_5334# 1.26e-19
C2413 a_27065_5334# ringtest_0.x4.net10 0.00375f
C2414 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._01_ 0.05158f
C2415 muxtest_0.x1.x3.GP1 muxtest_0.x1.x3.GP3 0.061475f
C2416 muxtest_0.x1.x3.GN4 muxtest_0.x1.x4.A 0.446529f
C2417 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A 0.17253f
C2418 a_12019_24012# ui_in[3] 9.55e-19
C2419 a_21233_5340# a_21509_4790# 0.001876f
C2420 ringtest_0.x4._15_ a_26817_4566# 0.004129f
C2421 a_19666_31955# muxtest_0.x1.x3.GN4 6.84e-19
C2422 ringtest_0.drv_out a_24329_6640# 4.16e-19
C2423 ringtest_0.x4._00_ a_21852_9416# 0.208988f
C2424 ringtest_0.x4._24_ a_26640_5156# 0.010089f
C2425 ringtest_0.x4._11_ a_21509_4790# 0.005486f
C2426 ringtest_0.x4.net3 ringtest_0.counter7 4.2e-20
C2427 ringtest_0.x4.net7 a_26808_4902# 1.23e-19
C2428 ringtest_0.x4.net5 a_22939_4584# 0.002311f
C2429 ringtest_0.x4._02_ a_22097_5334# 3.18e-19
C2430 a_21233_5340# a_22765_5308# 1.05e-19
C2431 ringtest_0.x4.clknet_1_0__leaf_clk a_21863_4790# 0.003207f
C2432 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP2 0.043302f
C2433 ringtest_0.x4._16_ ringtest_0.x4._02_ 3.22e-20
C2434 a_23349_6422# ringtest_0.x4._05_ 4.45e-20
C2435 ringtest_0.x4._18_ a_24465_6800# 7.52e-20
C2436 ringtest_0.x4.net10 a_26627_4246# 0.27342f
C2437 a_23879_6940# ringtest_0.x4._05_ 0.005813f
C2438 ringtest_0.x4._11_ a_22765_5308# 0.001227f
C2439 ringtest_0.x4.net8 a_24968_5308# 0.001066f
C2440 a_18836_32319# ui_in[0] 9.55e-19
C2441 a_27659_4246# VDPWR 0.00908f
C2442 ringtest_0.x4.net10 a_27149_5156# 3.08e-19
C2443 a_16027_11759# a_16155_12151# 0.004764f
C2444 ringtest_0.x3.x2.GN2 ui_in[4] 0.108649f
C2445 ringtest_0.x4._08_ a_24361_5340# 3.42e-20
C2446 a_16027_11759# ringtest_0.x3.x2.GN1 0.012445f
C2447 a_16579_11759# a_16755_12091# 0.185422f
C2448 ringtest_0.x4._13_ a_21233_5340# 3.88e-19
C2449 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VDPWR 0.636415f
C2450 muxtest_0.x1.x3.GP1 muxtest_0.R1R2 2.46e-21
C2451 ringtest_0.x4._11_ a_21867_8054# 1.17e-19
C2452 uio_in[2] uio_in[1] 0.031023f
C2453 ringtest_0.x4.net6 a_24527_5340# 0.048602f
C2454 ringtest_0.x4.clknet_0_clk a_24712_6422# 4.01e-19
C2455 a_21375_3867# ringtest_0.x4.counter[1] 0.1107f
C2456 a_21509_4790# a_21675_4790# 0.970278f
C2457 ringtest_0.x4._07_ a_25149_4220# 9.24e-19
C2458 ringtest_0.x4.net4 a_22139_5878# 0.011292f
C2459 ringtest_0.drv_out a_25364_5878# 1.27e-19
C2460 ringtest_0.x4._22_ a_25977_4220# 0.191159f
C2461 ringtest_0.x4._11_ ringtest_0.x4._13_ 0.217373f
C2462 a_24968_5308# a_24729_4790# 1.62e-19
C2463 a_24527_5340# a_24895_4790# 1.17e-19
C2464 ringtest_0.x4._22_ a_25719_4790# 7.63e-20
C2465 a_24361_5340# a_25336_4902# 3.92e-19
C2466 muxtest_0.x1.x3.GN3 muxtest_0.R3R4 0.377005f
C2467 ringtest_0.x4.clknet_1_0__leaf_clk a_21785_8054# 0.024338f
C2468 a_24329_6640# ringtest_0.x4._07_ 5.99e-19
C2469 ringtest_0.x4.net3 a_22295_3867# 0.001252f
C2470 a_25149_4220# a_25055_3867# 3.27e-19
C2471 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net6 0.087511f
C2472 a_24336_6544# ringtest_0.x4._22_ 8.56e-19
C2473 a_22265_5308# a_21948_5156# 0.005602f
C2474 a_22097_5334# a_22116_4902# 3.73e-19
C2475 a_27233_5058# a_27489_3702# 3.35e-20
C2476 ringtest_0.x4.net9 a_25083_4790# 1.61e-19
C2477 ringtest_0.x4.clknet_0_clk a_24895_4790# 3.43e-21
C2478 ringtest_0.x4._18_ a_22733_6244# 1.72e-19
C2479 m2_15612_11606# ui_in[4] 0.183786f
C2480 ringtest_0.x4._16_ a_22116_4902# 0.005579f
C2481 ui_in[3] ui_in[4] 13.6084f
C2482 a_26367_5340# a_26808_5308# 0.118966f
C2483 a_21399_5340# a_22181_5334# 6.32e-19
C2484 a_26201_5340# a_26640_5334# 0.273138f
C2485 ringtest_0.x4._15_ ringtest_0.x4._24_ 0.032103f
C2486 a_24361_5340# VDPWR 0.419324f
C2487 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A ui_in[3] 9.57e-20
C2488 ringtest_0.x4._16_ a_23993_5654# 3.31e-19
C2489 ringtest_0.x4.net4 a_21863_4790# 4.45e-19
C2490 ringtest_0.x4.net9 a_24715_5334# 1.41e-19
C2491 a_21785_5878# a_21509_4790# 2.82e-20
C2492 ringtest_0.x4.net7 a_25083_4790# 4.68e-19
C2493 a_12849_23648# muxtest_0.x2.x2.GP1 1.21e-20
C2494 a_24465_6800# ringtest_0.x4.clknet_1_1__leaf_clk 1.17e-20
C2495 a_21395_6940# VDPWR 1.51709f
C2496 ringtest_0.x3.x2.GN4 a_17405_12123# 0.001562f
C2497 ringtest_0.counter7 a_26201_4790# 2.09e-20
C2498 ringtest_0.x4._22_ a_24986_5878# 0.006962f
C2499 muxtest_0.x2.x2.GP3 ua[3] 0.084041f
C2500 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GN4 0.071282f
C2501 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP1 2.56189f
C2502 muxtest_0.x1.x1.nSEL1 ui_in[2] 0.164995f
C2503 a_21785_5878# a_22765_5308# 0.002539f
C2504 a_21132_8918# VDPWR 2.08e-19
C2505 ringtest_0.x4._04_ a_22097_5334# 0.001211f
C2506 a_25364_5878# ringtest_0.x4._07_ 0.022424f
C2507 ringtest_0.x4.net7 a_24715_5334# 0.014734f
C2508 ringtest_0.x4._04_ ringtest_0.x4._16_ 0.025302f
C2509 ringtest_0.x4.clknet_1_0__leaf_clk a_22097_5334# 0.004501f
C2510 a_25975_3867# ringtest_0.x4.counter[6] 0.1107f
C2511 a_26367_5340# a_26555_4790# 1.41e-20
C2512 ringtest_0.x4._11_ ringtest_0.x4.net8 0.418201f
C2513 a_21951_5878# a_24004_6128# 1.23e-20
C2514 ringtest_0.x4.net9 a_25547_4612# 6.77e-19
C2515 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._16_ 4.14e-20
C2516 a_21981_9142# ui_in[5] 2.79e-20
C2517 ringtest_0.x4._05_ a_24968_5308# 8.7e-19
C2518 muxtest_0.R7R8 muxtest_0.R5R6 0.318606f
C2519 muxtest_0.x1.x3.GP2 muxtest_0.R3R4 0.170487f
C2520 ringtest_0.x4._13_ a_21785_5878# 0.002226f
C2521 muxtest_0.x2.x2.GP3 m3_13316_18955# 0.006132f
C2522 a_22111_10993# ui_in[5] 0.231636f
C2523 ringtest_0.ring_out ringtest_0.drv_out 2.13841f
C2524 ringtest_0.x4.net1 a_21395_6940# 0.001584f
C2525 muxtest_0.x1.x3.GN1 muxtest_0.R4R5 0.334962f
C2526 muxtest_0.R7R8 VDPWR 3.21675f
C2527 a_21981_9142# ringtest_0.x4._12_ 7.61e-20
C2528 ringtest_0.x3.x2.GP1 ui_in[3] 8.3e-19
C2529 ringtest_0.x4._07_ a_24317_4942# 1.81e-19
C2530 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A 5.04e-19
C2531 ringtest_0.drv_out ringtest_0.x4._19_ 0.013619f
C2532 ringtest_0.x4.net1 a_21132_8918# 0.001512f
C2533 ringtest_0.x4._23_ a_27273_4220# 0.220841f
C2534 ringtest_0.x4._11_ a_24729_4790# 0.029022f
C2535 ringtest_0.x4.net7 a_25547_4612# 0.001525f
C2536 a_22765_4478# a_23381_4584# 0.013543f
C2537 ringtest_0.x4.net8 a_25761_5058# 0.020836f
C2538 a_26808_4902# a_26627_4246# 3.15e-19
C2539 ringtest_0.x4._23_ a_26766_4790# 6.82e-19
C2540 a_19114_31955# a_19242_32347# 0.004764f
C2541 ringtest_0.x4._02_ a_21587_5334# 0.114994f
C2542 a_22224_6244# a_22541_5058# 2.18e-19
C2543 a_26808_4902# a_27149_5156# 9.73e-19
C2544 ringtest_0.x4._05_ a_25925_6788# 1.27e-19
C2545 muxtest_0.x1.x3.GN4 ua[0] 4.10932f
C2546 a_21399_5340# a_21840_5308# 0.127288f
C2547 ringtest_0.x4.clknet_1_1__leaf_clk a_26201_4790# 0.306202f
C2548 ringtest_0.x4.net10 a_26721_4246# 0.007482f
C2549 ringtest_0.x4.net6 a_25168_5156# 6.05e-21
C2550 ringtest_0.x4._11_ a_21798_5712# 4.01e-19
C2551 a_13025_23980# muxtest_0.x2.x2.GN4 0.003699f
C2552 a_25364_5878# a_26201_5340# 0.016172f
C2553 ringtest_0.x4._21_ a_24361_5340# 0.016583f
C2554 muxtest_0.x2.x2.GN1 a_12019_24012# 0.001144f
C2555 a_13501_23906# muxtest_0.x2.x2.GN2 7.58e-21
C2556 a_23529_6422# a_24329_6640# 2.3e-20
C2557 a_23949_6654# a_24045_6654# 0.310858f
C2558 muxtest_0.x2.x2.GN2 ua[2] 0.429379f
C2559 a_24729_4790# a_25761_5058# 0.048748f
C2560 a_24895_4790# a_25168_5156# 0.074022f
C2561 a_19290_32287# ui_in[0] 0.143958f
C2562 ringtest_0.x4._08_ VDPWR 0.45369f
C2563 ringtest_0.x4.net4 a_22097_5334# 0.006897f
C2564 ringtest_0.x4.clknet_1_1__leaf_clk a_26555_5334# 3.58e-19
C2565 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VDPWR 0.636362f
C2566 ringtest_0.x4.net6 a_22983_5654# 0.001315f
C2567 ringtest_0.x4._15_ a_27233_5308# 1.61e-19
C2568 muxtest_0.R2R3 ua[3] 0.017699f
C2569 ringtest_0.x4.net3 ringtest_0.x4._02_ 0.031079f
C2570 ringtest_0.x4.net4 ringtest_0.x4._16_ 0.442589f
C2571 ringtest_0.x4._22_ a_27491_4566# 3.34e-21
C2572 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GN3 1.1e-19
C2573 ringtest_0.drv_out ringtest_0.x4.net9 4.05e-20
C2574 ui_in[0] ui_in[3] 0.001641f
C2575 ringtest_0.counter3 ringtest_0.x4._13_ 0.003357f
C2576 ringtest_0.x4._04_ a_22649_6244# 0.006456f
C2577 a_21785_5878# ringtest_0.x4.net8 9.67e-20
C2578 a_25336_4902# VDPWR 0.183561f
C2579 ringtest_0.x4._18_ a_23770_5308# 0.079699f
C2580 ringtest_0.x4._11_ a_22390_4566# 9.44e-19
C2581 ringtest_0.x4.net8 a_25345_4612# 0.005557f
C2582 a_23879_6940# a_24361_5340# 3.84e-19
C2583 ringtest_0.x4.clknet_1_0__leaf_clk a_22649_6244# 6.75e-21
C2584 a_20492_32319# ui_in[1] 8.84e-19
C2585 ringtest_0.x4._11_ ringtest_0.x4.net11 2.31e-19
C2586 muxtest_0.R5R6 VDPWR 1.61253f
C2587 a_19842_32287# ui_in[1] 0.127717f
C2588 ringtest_0.x4._25_ ringtest_0.x4._08_ 0.208467f
C2589 muxtest_0.x1.x5.GN ua[3] 0.820663f
C2590 a_24329_6640# ringtest_0.x4._06_ 0.002324f
C2591 a_25393_5308# a_25351_5712# 7.84e-20
C2592 ringtest_0.x4._11_ ringtest_0.x4._05_ 0.023537f
C2593 ringtest_0.drv_out ringtest_0.x4.net7 6.87e-19
C2594 ringtest_0.x4.net6 a_21591_6128# 4.71e-21
C2595 a_21561_9116# a_21561_8830# 0.015931f
C2596 ringtest_0.counter7 ringtest_0.x4.counter[8] 0.068429f
C2597 a_24045_6654# a_24004_6128# 0.001715f
C2598 a_22223_5712# VDPWR 0.002609f
C2599 ringtest_0.x4._15_ a_25977_4220# 0.086673f
C2600 ringtest_0.x4._19_ a_24264_6788# 1.38e-19
C2601 ringtest_0.drv_out ringtest_0.x4._17_ 1.68e-19
C2602 muxtest_0.x1.x1.nSEL1 a_19794_32347# 4.08e-19
C2603 muxtest_0.x1.x1.nSEL0 a_19242_32347# 2.51e-19
C2604 ringtest_0.x4._23_ a_26201_4790# 0.029061f
C2605 ringtest_0.x4.net2 a_21675_9686# 0.008042f
C2606 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A ui_in[3] 9.57e-20
C2607 muxtest_0.x1.x5.GN a_19842_32287# 2.26e-19
C2608 a_24336_6544# ringtest_0.x4._15_ 1.53e-20
C2609 a_26201_4790# a_26367_4790# 0.970499f
C2610 ringtest_0.x4.net3 a_22116_4902# 3.22e-20
C2611 ringtest_0.x3.x2.GP3 ua[1] 0.357364f
C2612 a_23381_4818# a_23381_4584# 0.012876f
C2613 a_21675_4790# a_22390_4566# 4.63e-19
C2614 ringtest_0.x4._16_ a_23837_5878# 0.061172f
C2615 ringtest_0.x4._04_ a_21587_5334# 3.27e-21
C2616 muxtest_0.x1.x3.GN1 ui_in[2] 0.054229f
C2617 ringtest_0.x4.net9 ringtest_0.x4._07_ 0.03749f
C2618 ringtest_0.x4._22_ ringtest_0.x4._16_ 0.135659f
C2619 a_16755_12091# ringtest_0.x3.x2.GP3 5.21e-19
C2620 ringtest_0.x4._06_ a_24545_5878# 0.046896f
C2621 m3_17032_8096# m3_17046_7066# 0.003741f
C2622 ringtest_0.x4._23_ a_26555_5334# 0.014354f
C2623 muxtest_0.x2.x2.GN1 ui_in[4] 0.312374f
C2624 a_22795_5334# a_22765_4478# 6.77e-20
C2625 muxtest_0.x2.x1.nSEL0 a_12473_23980# 0.001174f
C2626 ringtest_0.x4.clknet_1_0__leaf_clk a_21587_5334# 0.03291f
C2627 a_26555_5334# a_26367_4790# 1.41e-20
C2628 a_23467_4584# VDPWR 0.002731f
C2629 a_21803_9508# VDPWR 0.005022f
C2630 ringtest_0.x4._25_ VDPWR 0.220602f
C2631 ringtest_0.x4._11_ a_22350_5878# 0.003523f
C2632 a_24004_6128# a_24699_6200# 5.89e-19
C2633 ringtest_0.x4.net1 VDPWR 1.43699f
C2634 ringtest_0.x4.clknet_1_1__leaf_clk a_23770_5308# 0.048773f
C2635 ringtest_0.x4.net7 ringtest_0.x4._07_ 0.047771f
C2636 muxtest_0.x1.x3.GP3 muxtest_0.R4R5 0.346864f
C2637 ringtest_0.x4.net4 a_22649_6244# 0.002624f
C2638 muxtest_0.x1.x3.GP1 muxtest_0.R6R7 0.271251f
C2639 ringtest_0.x4.net3 ringtest_0.x4._04_ 5.28e-22
C2640 a_21852_8720# a_22052_8875# 0.080195f
C2641 a_21785_5878# a_22390_4566# 4.07e-21
C2642 a_21561_8830# ringtest_0.x4._01_ 8.93e-19
C2643 a_21845_8816# a_21981_8976# 0.136009f
C2644 a_26201_5340# a_26735_5334# 0.002698f
C2645 ringtest_0.x4._17_ ringtest_0.x4._07_ 3.97e-20
C2646 ringtest_0.x4._23_ a_27303_4246# 0.113094f
C2647 ringtest_0.x4.net7 a_25055_3867# 0.201574f
C2648 a_25977_4220# a_26173_4612# 0.00119f
C2649 ringtest_0.x4._11_ ringtest_0.x4._09_ 0.004259f
C2650 ringtest_0.x4._14_ a_21948_5156# 9.43e-20
C2651 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net3 0.373279f
C2652 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A 0.17253f
C2653 a_26808_4902# a_26721_4246# 5.71e-20
C2654 a_11845_23906# ui_in[3] 0.048888f
C2655 a_22052_9116# a_22399_9142# 0.037333f
C2656 ringtest_0.x4._06_ a_24317_4942# 2.49e-19
C2657 ringtest_0.x4.net2 a_22052_8875# 3.35e-21
C2658 a_21845_9116# ringtest_0.x4.clknet_1_0__leaf_clk 0.308902f
C2659 ringtest_0.x4.net7 a_24264_6788# 0.001683f
C2660 a_24004_6128# a_23809_4790# 5.65e-20
C2661 ringtest_0.drv_out ringtest_0.x3.x2.GN3 0.243642f
C2662 ringtest_0.x4.net1 a_21803_9508# 8.57e-19
C2663 a_24361_5340# a_24968_5308# 0.136009f
C2664 ringtest_0.x4.net8 ringtest_0.x4.net10 1.02e-19
C2665 ringtest_0.x4.net9 a_26201_5340# 8.34e-19
C2666 a_25593_5156# a_26201_4790# 3.54e-19
C2667 a_23529_6422# ringtest_0.x4._19_ 0.082191f
C2668 ringtest_0.x4._21_ VDPWR 0.483109f
C2669 a_25761_5058# ringtest_0.x4._09_ 0.001669f
C2670 ringtest_0.x4._18_ ringtest_0.x4.net6 0.081404f
C2671 ringtest_0.x4.clknet_0_clk a_24527_5340# 5.94e-19
C2672 ringtest_0.counter7 ringtest_0.x4.net6 6.88e-20
C2673 ringtest_0.x4.counter[2] VDPWR 0.488095f
C2674 a_24045_6654# ringtest_0.x4._20_ 1.76e-19
C2675 ringtest_0.x4.net4 a_21587_5334# 1.97e-19
C2676 a_23809_4790# a_23963_4790# 0.004009f
C2677 ringtest_0.x4._15_ a_23899_5334# 0.046541f
C2678 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VDPWR 0.636314f
C2679 ringtest_0.x4._24_ a_26367_5340# 0.035946f
C2680 muxtest_0.x1.x4.A a_12977_24040# 3.86e-20
C2681 a_16027_11759# ui_in[4] 0.03417f
C2682 a_23381_4818# a_23809_4790# 0.00155f
C2683 a_21675_4790# a_22074_4790# 0.001351f
C2684 a_21948_5156# a_22043_5156# 0.007724f
C2685 ringtest_0.x3.x1.nSEL1 a_16203_12091# 0.041068f
C2686 a_22116_4902# a_22457_5156# 9.73e-19
C2687 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN2 1.03e-20
C2688 ringtest_0.counter3 ringtest_0.x4.counter[1] 0.099026f
C2689 ringtest_0.x4.net7 a_26201_5340# 8.61e-20
C2690 a_22265_5308# a_22164_4362# 6.81e-19
C2691 a_21425_9686# VDPWR 0.25892f
C2692 ringtest_0.x4._16_ a_22021_4220# 0.184103f
C2693 a_21951_5878# a_22392_5990# 0.111047f
C2694 a_23349_6422# VDPWR 0.251829f
C2695 a_12849_23648# VDPWR 0.180589f
C2696 a_21845_8816# a_22228_8598# 0.001632f
C2697 a_21981_8976# a_22201_8964# 4.62e-19
C2698 a_23879_6940# VDPWR 1.2913f
C2699 ringtest_0.x4._23_ ringtest_0.x4.counter[8] 9.18e-19
C2700 a_22052_8875# a_22399_8976# 0.037333f
C2701 a_21852_8720# a_21803_8598# 4.04e-19
C2702 ringtest_0.x4.net9 a_27233_5058# 0.001937f
C2703 ringtest_0.x4.net6 a_24763_6143# 0.027058f
C2704 ringtest_0.x3.x2.GP3 m3_17046_7066# 0.006132f
C2705 ringtest_0.x4._19_ ringtest_0.x4._06_ 7.42e-21
C2706 ringtest_0.x4.net7 ringtest_0.x4.counter[5] 0.002945f
C2707 ringtest_0.x4.net3 ringtest_0.x4.net4 0.0313f
C2708 muxtest_0.x2.x2.GN2 m3_13302_19985# 0.016745f
C2709 muxtest_0.x2.x2.GN4 ui_in[3] 0.218988f
C2710 a_25309_5334# VDPWR 0.004428f
C2711 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP1 0.062377f
C2712 ringtest_0.x4.counter[1] ua[2] 1.11e-19
C2713 muxtest_0.x1.x3.GN2 a_19242_32347# 0.002395f
C2714 a_20318_32213# muxtest_0.x1.x3.GN4 0.134079f
C2715 ringtest_0.x4._24_ a_27065_5156# 0.012283f
C2716 ringtest_0.x4._00_ a_22052_9116# 0.00938f
C2717 ringtest_0.x4.net7 a_27233_5058# 8.32e-20
C2718 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y ui_in[3] 9.57e-20
C2719 ringtest_0.x4.net1 a_21425_9686# 0.224922f
C2720 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4.net6 0.323735f
C2721 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP2 2.14737f
C2722 ringtest_0.ring_out ringtest_0.x3.x1.nSEL0 1.86e-21
C2723 muxtest_0.x1.x3.GP3 ui_in[2] 1.6e-19
C2724 a_23529_6422# ringtest_0.x4.net7 0.002934f
C2725 ringtest_0.x4.clknet_1_1__leaf_clk a_24895_4790# 0.486375f
C2726 ringtest_0.x4.net8 a_25393_5308# 0.084103f
C2727 ringtest_0.x4._11_ a_24361_5340# 1.58e-19
C2728 ringtest_0.x4._17_ a_23529_6422# 0.043588f
C2729 ringtest_0.x4.net10 ringtest_0.x4.net11 0.310558f
C2730 a_21375_3867# VDPWR 0.271691f
C2731 a_16027_11759# ringtest_0.x3.x2.GP1 9.92e-19
C2732 ringtest_0.x4._06_ ringtest_0.x4.net9 0.017291f
C2733 ringtest_0.x4._08_ a_24968_5308# 9.82e-20
C2734 a_16203_12091# ringtest_0.x3.x2.GN3 0.048646f
C2735 a_23809_4790# ringtest_0.x4._20_ 0.237238f
C2736 a_16579_11759# ringtest_0.x3.x2.GN1 6.43e-20
C2737 ua[3] ui_in[4] 1.15229f
C2738 ringtest_0.x4._11_ a_21395_6940# 0.055744f
C2739 a_21509_4790# a_21948_5156# 0.273138f
C2740 ringtest_0.x4._03_ a_22116_4902# 0.006259f
C2741 ringtest_0.x4.net6 a_24800_5334# 0.019975f
C2742 ringtest_0.x4._15_ a_22097_5334# 7.5e-20
C2743 ringtest_0.x4._22_ a_27273_4220# 4.31e-19
C2744 ringtest_0.x4._12_ a_22245_8054# 0.026119f
C2745 muxtest_0.x1.x5.A muxtest_0.R7R8 4.52065f
C2746 a_25393_5308# a_24729_4790# 0.002274f
C2747 a_24527_5340# a_25168_5156# 7.62e-19
C2748 a_24800_5334# a_24895_4790# 8.92e-19
C2749 ringtest_0.x4._15_ ringtest_0.x4._16_ 0.656968f
C2750 a_25977_4220# a_25975_3867# 0.01226f
C2751 ringtest_0.x4.net7 ringtest_0.x4._06_ 0.141876f
C2752 ringtest_0.x4.net7 a_24070_5852# 0.003377f
C2753 ringtest_0.x4.clknet_0_clk a_25168_5156# 4.63e-19
C2754 ringtest_0.x4._18_ a_23932_6128# 0.00112f
C2755 ringtest_0.x4._17_ ringtest_0.x4._06_ 0.001225f
C2756 muxtest_0.x1.x1.nSEL1 ui_in[1] 0.275603f
C2757 ringtest_0.x4._16_ a_22541_5058# 1.37e-19
C2758 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A 5.04e-19
C2759 a_23879_6940# ringtest_0.x4._21_ 0.001038f
C2760 a_26367_5340# a_27233_5308# 0.034054f
C2761 ringtest_0.x4._17_ a_24070_5852# 0.062168f
C2762 a_26808_5308# a_26640_5334# 0.239923f
C2763 a_26201_5340# a_27065_5334# 0.032244f
C2764 a_23770_5308# a_23993_5654# 0.011458f
C2765 a_24968_5308# VDPWR 0.183392f
C2766 a_24329_6640# a_24883_6800# 0.057611f
C2767 a_24045_6654# a_24287_6422# 0.008508f
C2768 ringtest_0.x4.net6 ringtest_0.x4._23_ 0.023006f
C2769 ringtest_0.x4.net4 a_22457_5156# 8.77e-19
C2770 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x5.GN 0.10521f
C2771 muxtest_0.x2.x2.GP1 ua[2] 0.352897f
C2772 a_24895_4790# a_26367_4790# 0.002814f
C2773 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._03_ 0.00668f
C2774 a_18662_32213# m2_18699_31802# 0.01297f
C2775 muxtest_0.x2.x1.nSEL1 a_12977_24040# 4.08e-19
C2776 a_11845_23906# muxtest_0.x2.x2.GN1 0.12869f
C2777 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN2 0.209956f
C2778 ringtest_0.counter7 ringtest_0.x4.net5 6.88e-20
C2779 ringtest_0.x4.net10 ringtest_0.x4._09_ 0.081678f
C2780 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VDPWR 0.636314f
C2781 a_27233_5308# a_27065_5156# 7.04e-19
C2782 a_27065_5334# a_27233_5058# 7.04e-19
C2783 a_25925_6788# VDPWR 0.451929f
C2784 a_22817_6146# ringtest_0.x4._06_ 1.81e-20
C2785 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x1.nSEL1 0.352716f
C2786 a_21395_6940# a_21785_5878# 5.49e-20
C2787 a_21375_3867# ringtest_0.x4.counter[2] 4.98e-19
C2788 a_22817_6146# a_24070_5852# 2.22e-20
C2789 uio_in[7] uio_in[6] 0.031023f
C2790 ringtest_0.x4.net6 ringtest_0.x4._02_ 0.001309f
C2791 muxtest_0.x1.x5.A muxtest_0.R5R6 4.5214f
C2792 ringtest_0.x4._11_ ringtest_0.x4._08_ 1.44e-20
C2793 ringtest_0.x4.clknet_1_0__leaf_clk a_21939_8054# 3.8e-19
C2794 a_15749_12123# VDPWR 9.25e-19
C2795 ringtest_0.x4._22_ a_26201_4790# 4.68e-20
C2796 muxtest_0.x2.x2.GN2 ua[0] 4.0283f
C2797 ringtest_0.x3.x2.GN3 m3_17036_9140# 0.001446f
C2798 a_19794_32347# muxtest_0.x1.x3.GP3 4.39e-19
C2799 muxtest_0.x1.x5.A VDPWR 14.1646f
C2800 ringtest_0.x4.net3 a_22021_4220# 0.002183f
C2801 ringtest_0.x4._15_ a_26201_6788# 0.001194f
C2802 ringtest_0.x4.net7 a_26269_4612# 5.42e-19
C2803 ringtest_0.x4._11_ a_25336_4902# 0.039242f
C2804 ringtest_0.x4._23_ a_27169_6641# 6.47e-19
C2805 a_25925_6788# ringtest_0.x4._25_ 1.87e-19
C2806 ringtest_0.x4.net11 a_27191_4790# 3e-19
C2807 ringtest_0.x4._07_ a_25351_5712# 5.27e-19
C2808 a_19290_32287# muxtest_0.x1.x3.GN3 0.048646f
C2809 ringtest_0.counter7 a_21007_3867# 2.81e-20
C2810 ringtest_0.x4._02_ a_21055_5334# 0.01416f
C2811 a_26749_6422# a_26808_4902# 1.02e-20
C2812 a_21675_9686# a_21465_9294# 3.08e-19
C2813 a_19114_31955# VDPWR 0.164569f
C2814 a_26555_4790# a_26735_5156# 0.001229f
C2815 a_26640_5156# a_26766_4790# 0.005525f
C2816 a_21233_5340# VDPWR 0.680742f
C2817 a_21840_5308# a_21672_5334# 0.239923f
C2818 a_21399_5340# a_22265_5308# 0.034054f
C2819 ringtest_0.x4.net10 a_27659_4246# 0.003077f
C2820 ringtest_0.x4.net4 ringtest_0.x4._03_ 0.031989f
C2821 ringtest_0.ring_out ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.167117f
C2822 muxtest_0.x2.x2.GN3 a_12977_24040# 0.001073f
C2823 ringtest_0.x4.net8 a_24715_5334# 0.005878f
C2824 m2_11882_23495# VDPWR 0.139985f
C2825 muxtest_0.x2.x2.GN2 a_13675_24012# 8.14e-21
C2826 ringtest_0.x4.net6 a_25593_5156# 4.38e-19
C2827 ringtest_0.x4._15_ a_23467_4818# 7.85e-19
C2828 ringtest_0.x4._11_ a_22223_5712# 6.78e-19
C2829 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GN3 0.067465f
C2830 muxtest_0.x2.x2.GN1 muxtest_0.x2.x2.GN4 0.001074f
C2831 a_25364_5878# a_26808_5308# 0.006157f
C2832 a_20492_32319# ui_in[0] 1.77e-19
C2833 a_23949_6654# a_24336_6544# 0.034054f
C2834 a_24045_6654# a_24329_6640# 0.030894f
C2835 ringtest_0.x4._11_ VDPWR 5.08909f
C2836 a_25336_4902# a_25761_5058# 1.28e-19
C2837 a_24729_4790# a_25083_4790# 0.062224f
C2838 a_24895_4790# a_25593_5156# 0.193199f
C2839 a_19842_32287# ui_in[0] 0.279876f
C2840 ringtest_0.x4.net4 a_23770_5308# 1.34e-19
C2841 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN3 4.01e-20
C2842 ringtest_0.x4.clknet_1_1__leaf_clk a_24895_5334# 0.002214f
C2843 ringtest_0.x4._22_ a_27303_4246# 6.52e-20
C2844 a_25975_3867# ringtest_0.x4.counter[9] 2.37e-20
C2845 muxtest_0.R6R7 muxtest_0.R4R5 2.49e-19
C2846 ringtest_0.x4._14_ a_22164_4362# 0.089653f
C2847 a_25761_5058# VDPWR 0.395041f
C2848 ringtest_0.x4.net8 a_25547_4612# 1.72e-20
C2849 ringtest_0.x4._11_ a_23467_4584# 6.46e-19
C2850 a_23879_6940# a_24968_5308# 8.05e-21
C2851 ringtest_0.x4._11_ ringtest_0.x4._25_ 2.54e-20
C2852 muxtest_0.x1.x3.GN1 muxtest_0.R2R3 2.55e-19
C2853 a_21675_4790# VDPWR 0.328278f
C2854 a_25364_5878# a_26555_4790# 1.26e-19
C2855 muxtest_0.x1.x3.GN1 ui_in[1] 0.312176f
C2856 a_24536_6699# ringtest_0.x4._06_ 2.41e-19
C2857 ringtest_0.x4.net3 a_21561_8830# 0.006429f
C2858 a_24968_5308# a_25309_5334# 9.73e-19
C2859 a_24800_5334# a_24895_5334# 0.007724f
C2860 ringtest_0.x4.net1 ringtest_0.x4._11_ 0.002334f
C2861 ringtest_0.x4.clknet_0_clk ringtest_0.x4._18_ 0.002702f
C2862 ringtest_0.x4.net6 ringtest_0.x4._04_ 0.050232f
C2863 a_24336_6544# a_24004_6128# 0.002652f
C2864 a_21561_9116# a_21852_8720# 1.53e-19
C2865 a_24329_6640# a_24699_6200# 0.007926f
C2866 a_21852_9416# a_21845_8816# 3.36e-19
C2867 a_21845_9116# a_21561_8830# 9.64e-20
C2868 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A 0.17253f
C2869 a_23899_5654# VDPWR 5.6e-19
C2870 a_26569_6422# ringtest_0.x4._24_ 0.095435f
C2871 ringtest_0.ring_out ua[1] 4.51997f
C2872 ringtest_0.x4._19_ a_24883_6800# 0.014678f
C2873 ringtest_0.x3.nselect2 ui_in[3] 1.88e-19
C2874 ringtest_0.x4.net2 a_21780_9142# 2.28e-19
C2875 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net6 6.56e-20
C2876 ringtest_0.x4._09_ a_27191_4790# 0.001794f
C2877 ringtest_0.x4.net2 a_21561_9116# 0.019416f
C2878 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN1 0.645006f
C2879 muxtest_0.x1.x1.nSEL0 VDPWR 0.389106f
C2880 ringtest_0.ring_out a_16755_12091# 2.55e-19
C2881 a_26201_4790# a_26640_5156# 0.273138f
C2882 ringtest_0.x4._09_ a_26808_4902# 0.039926f
C2883 a_24465_6800# ringtest_0.x4._15_ 2.35e-21
C2884 a_24763_6143# a_24527_5340# 0.003413f
C2885 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GP3 0.002437f
C2886 a_21785_5878# VDPWR 0.63892f
C2887 muxtest_0.x2.x1.nSEL0 a_13025_23980# 1.21e-20
C2888 a_21951_5878# a_22265_5308# 0.003783f
C2889 a_24045_6654# a_24317_4942# 5.98e-21
C2890 a_24699_6200# a_24545_5878# 0.049785f
C2891 ringtest_0.x4.clknet_0_clk a_24763_6143# 7.62e-19
C2892 ringtest_0.x4.clknet_1_0__leaf_clk a_21055_5334# 1.21e-20
C2893 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP1 1.16e-20
C2894 a_22399_9142# VDPWR 0.077754f
C2895 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VDPWR 0.63819f
C2896 ringtest_0.x4.net9 a_26895_3867# 0.202772f
C2897 muxtest_0.R7R8 ua[2] 4.51509f
C2898 ringtest_0.x4._11_ ringtest_0.x4._21_ 0.059807f
C2899 a_23949_6654# a_23899_5334# 2.76e-21
C2900 ringtest_0.x4.clknet_1_1__leaf_clk a_24527_5340# 0.079788f
C2901 muxtest_0.x2.x2.GP1 m3_13302_19985# 3.25e-21
C2902 muxtest_0.x1.x3.GN4 muxtest_0.R4R5 4.23588f
C2903 ringtest_0.x4.net3 a_21049_8598# 0.042192f
C2904 a_21852_8720# ringtest_0.x4._01_ 0.239739f
C2905 a_22052_8875# a_21981_8976# 0.239923f
C2906 a_26367_5340# a_27149_5334# 6.32e-19
C2907 ringtest_0.x4.clknet_0_clk ringtest_0.x4.clknet_1_1__leaf_clk 0.335671f
C2908 a_25977_4220# a_26375_4612# 0.005781f
C2909 muxtest_0.x1.x3.GN2 muxtest_0.R7R8 0.260757f
C2910 ringtest_0.x4._14_ a_22373_5156# 0.002114f
C2911 a_12473_23980# ui_in[3] 0.143958f
C2912 ringtest_0.x4.net2 ringtest_0.x4._01_ 9.85e-20
C2913 ringtest_0.x4.net6 ringtest_0.x4.net4 0.008308f
C2914 a_21981_9142# ringtest_0.x4.clknet_1_0__leaf_clk 0.050329f
C2915 ringtest_0.x4._11_ a_23349_6422# 0.001422f
C2916 ringtest_0.x4.net7 a_24883_6800# 0.019182f
C2917 ringtest_0.x4._11_ a_23879_6940# 4.59e-19
C2918 ringtest_0.x4._17_ a_21951_5878# 9.29e-21
C2919 ringtest_0.x4.net1 a_22399_9142# 5.53e-20
C2920 a_24527_5340# a_24800_5334# 0.074815f
C2921 a_24361_5340# a_25393_5308# 0.048748f
C2922 a_18662_32213# a_18836_32319# 0.006584f
C2923 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP2 0.043402f
C2924 ringtest_0.x4._17_ a_24883_6800# 0.016586f
C2925 ringtest_0.x4._15_ a_26201_4790# 0.02569f
C2926 ringtest_0.x4._21_ a_23899_5654# 2.03e-19
C2927 ringtest_0.x4.net9 a_26808_5308# 2.66e-21
C2928 ringtest_0.ring_out ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 5.04e-19
C2929 ringtest_0.x4._08_ ringtest_0.x4.net10 0.001321f
C2930 a_24329_6640# a_25421_6641# 5.23e-20
C2931 a_24045_6654# ringtest_0.x4._19_ 0.046625f
C2932 ringtest_0.x4.clknet_0_clk a_24800_5334# 4.59e-20
C2933 ringtest_0.counter3 VDPWR 2.47715f
C2934 a_21509_4790# a_22164_4362# 0.00127f
C2935 ringtest_0.x4._03_ a_22021_4220# 0.112166f
C2936 a_24317_4942# a_24479_4790# 0.004009f
C2937 muxtest_0.x2.x2.GN4 ua[3] 0.085877f
C2938 ringtest_0.x4._15_ a_26555_5334# 0.007874f
C2939 ringtest_0.x4.net8 ringtest_0.x4._07_ 0.001136f
C2940 a_16579_11759# ui_in[4] 0.261734f
C2941 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A ringtest_0.x3.x2.GN3 7.01e-21
C2942 ringtest_0.x4._24_ a_26640_5334# 0.010979f
C2943 ringtest_0.x3.x1.nSEL1 a_16755_12091# 1.59e-19
C2944 a_23809_4790# a_24317_4942# 0.017774f
C2945 a_21948_5156# a_22074_4790# 0.005525f
C2946 a_22116_4902# ringtest_0.x4.net5 0.001073f
C2947 ringtest_0.x4._00_ VDPWR 0.643985f
C2948 a_27489_3702# a_27815_3867# 0.024477f
C2949 ringtest_0.x4.net8 a_25055_3867# 3.76e-19
C2950 ringtest_0.x4._16_ a_22765_4478# 0.01632f
C2951 muxtest_0.x1.x3.GP3 muxtest_0.R2R3 0.115101f
C2952 a_21951_5878# a_22817_6146# 0.034054f
C2953 a_22392_5990# a_22224_6244# 0.239923f
C2954 a_13501_23906# VDPWR 0.218058f
C2955 VDPWR ua[2] 13.246901f
C2956 a_21845_8816# ringtest_0.x4._10_ 0.011255f
C2957 a_21852_8720# a_21785_8054# 1.58e-19
C2958 a_22052_8875# a_22228_8598# 0.007724f
C2959 a_21981_8976# a_21803_8598# 9.73e-19
C2960 ringtest_0.x4._01_ a_22399_8976# 0.121379f
C2961 muxtest_0.x1.x3.GP3 ui_in[1] 0.003199f
C2962 ringtest_0.x4.net6 a_23837_5878# 4.02e-19
C2963 ringtest_0.x4.clknet_0_clk ringtest_0.x4._23_ 2.29e-20
C2964 ringtest_0.x4.net9 a_26555_4790# 0.016338f
C2965 ringtest_0.x4.net6 ringtest_0.x4._22_ 0.641715f
C2966 muxtest_0.x2.x2.GN4 m3_13316_18955# 0.084813f
C2967 muxtest_0.x1.x3.GN2 muxtest_0.R5R6 0.122627f
C2968 a_23949_6654# ringtest_0.x4._16_ 3.45e-20
C2969 ringtest_0.x4._07_ a_24729_4790# 0.112051f
C2970 ringtest_0.x4.net10 VDPWR 1.25953f
C2971 ringtest_0.x4._19_ a_24699_6200# 1.87e-20
C2972 ringtest_0.x4._22_ a_24895_4790# 0.02378f
C2973 ringtest_0.x4.net6 a_24135_3867# 0.195979f
C2974 ringtest_0.x4.net2 a_21785_8054# 0.165774f
C2975 ringtest_0.x4.counter[0] ua[1] 3.21e-19
C2976 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A 5.04e-19
C2977 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GP3 3.82e-20
C2978 ringtest_0.drv_out ringtest_0.x4._05_ 0.0016f
C2979 a_24729_4790# a_25055_3867# 1.63e-21
C2980 muxtest_0.x1.x3.GN2 VDPWR 0.701394f
C2981 ringtest_0.x4.net7 a_23381_4584# 2.04e-20
C2982 ringtest_0.x4._00_ a_21803_9508# 3.7e-19
C2983 ringtest_0.x4._24_ a_26735_5156# 7.21e-19
C2984 ringtest_0.x4._04_ ringtest_0.x4.net5 0.003846f
C2985 ringtest_0.x4.net7 a_26555_4790# 2.26e-19
C2986 ua[1] ua[4] 0.001128f
C2987 ringtest_0.x4.net1 ringtest_0.x4._00_ 0.056053f
C2988 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net5 6.12e-20
C2989 a_24627_6200# VDPWR 0.001263f
C2990 ringtest_0.x4._14_ a_21399_5340# 4.89e-20
C2991 a_24045_6654# ringtest_0.x4.net7 0.037726f
C2992 muxtest_0.x1.x3.GN4 ui_in[2] 5.71e-20
C2993 ringtest_0.x4.counter[4] VDPWR 0.443202f
C2994 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GP1 1.21e-19
C2995 ringtest_0.x4.clknet_1_1__leaf_clk a_25168_5156# 0.042872f
C2996 ringtest_0.x4._06_ a_22765_5308# 1.6e-20
C2997 ringtest_0.x3.x2.GN3 ua[1] 0.429944f
C2998 muxtest_0.R2R3 muxtest_0.R1R2 1.9897f
C2999 ringtest_0.x4.net8 a_26201_5340# 0.001229f
C3000 ringtest_0.x4._11_ a_24968_5308# 7.26e-20
C3001 a_23399_3867# VDPWR 0.316069f
C3002 ringtest_0.x4._17_ a_24045_6654# 0.036473f
C3003 a_16579_11759# ringtest_0.x3.x2.GP1 1.21e-20
C3004 ui_in[3] ui_in[5] 0.141096f
C3005 ringtest_0.x4._08_ a_25393_5308# 9.54e-19
C3006 muxtest_0.x2.x1.nSEL1 a_12297_23648# 0.073392f
C3007 a_16755_12091# ringtest_0.x3.x2.GN3 0.004288f
C3008 muxtest_0.x1.x1.nSEL1 ui_in[0] 0.169954f
C3009 ringtest_0.x4.net9 ringtest_0.x4.counter[6] 3.69e-19
C3010 a_24004_6128# ringtest_0.x4._16_ 0.029136f
C3011 a_24699_6200# ringtest_0.x4.net9 0.170073f
C3012 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VDPWR 0.92605f
C3013 ringtest_0.counter3 ringtest_0.x4.counter[2] 0.16993f
C3014 ringtest_0.x4.net6 a_25225_5334# 8.63e-19
C3015 ringtest_0.x4._15_ a_23770_5308# 0.229149f
C3016 a_21509_4790# a_22373_5156# 0.032244f
C3017 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A ringtest_0.x3.x1.nSEL1 1.23e-19
C3018 ringtest_0.x4._03_ a_22541_5058# 3.08e-19
C3019 a_23899_5334# ringtest_0.x4._20_ 1.05e-19
C3020 a_25225_5334# a_24895_4790# 1.5e-19
C3021 a_25393_5308# a_25336_4902# 6.84e-19
C3022 ringtest_0.x4.net2 ringtest_0.x4._16_ 5.41e-20
C3023 muxtest_0.x2.x2.GP1 ua[0] 0.128232f
C3024 ringtest_0.x4._24_ a_25364_5878# 0.025563f
C3025 a_26627_4246# a_26895_3867# 1.23e-19
C3026 a_15575_12017# VDPWR 0.211635f
C3027 a_22649_6244# a_22765_4478# 3.06e-22
C3028 ringtest_0.x4._16_ a_23963_4790# 5.12e-19
C3029 ringtest_0.x4.net7 ringtest_0.x4.counter[6] 1.8e-19
C3030 ringtest_0.x4._11_ a_25925_6788# 0.087773f
C3031 ringtest_0.x4.net7 a_24699_6200# 6.37e-20
C3032 ringtest_0.x4.net9 a_24479_4790# 8.5e-21
C3033 a_22765_5308# a_22373_5156# 0.006202f
C3034 a_21840_5308# a_21863_4790# 6.87e-19
C3035 a_19666_31955# muxtest_0.R7R8 7.47e-21
C3036 ringtest_0.x4.counter[2] ua[2] 1.11e-19
C3037 ringtest_0.x4._16_ a_23381_4818# 0.113241f
C3038 a_22097_5334# a_22181_5334# 0.008508f
C3039 ringtest_0.x4._17_ a_24699_6200# 7.49e-19
C3040 a_22265_5308# a_22795_5334# 2.84e-19
C3041 a_26808_5308# a_27065_5334# 0.036838f
C3042 a_24361_5340# a_24715_5334# 0.057611f
C3043 muxtest_0.x2.x1.nSEL0 ui_in[3] 0.32698f
C3044 muxtest_0.R7R8 m3_13302_19985# 0.001045f
C3045 a_25393_5308# VDPWR 0.40591f
C3046 a_24465_6800# a_24685_6788# 4.62e-19
C3047 a_24336_6544# a_24287_6422# 4.04e-19
C3048 a_24536_6699# a_24883_6800# 0.037333f
C3049 a_21425_9686# ringtest_0.x4._00_ 0.167554f
C3050 ringtest_0.x4.net4 ringtest_0.x4.net5 0.483177f
C3051 a_25421_6641# ringtest_0.x4._19_ 0.214472f
C3052 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP1 0.001426f
C3053 ringtest_0.x4.net7 a_24479_4790# 1.98e-19
C3054 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.001676f
C3055 a_12297_23648# muxtest_0.x2.x2.GN3 6.68e-19
C3056 ringtest_0.x4.net7 a_23809_4790# 0.003261f
C3057 a_12473_23980# muxtest_0.x2.x2.GN1 1.46e-19
C3058 muxtest_0.R7R8 muxtest_0.x2.x2.GP2 1.13e-20
C3059 a_23932_6128# a_23837_5878# 0.002032f
C3060 ringtest_0.x4._11_ a_21233_5340# 0.00462f
C3061 ringtest_0.x4._17_ a_23809_4790# 1e-20
C3062 a_21951_5878# ringtest_0.x4._14_ 3.24e-22
C3063 a_26749_6422# a_26201_5340# 6.06e-21
C3064 a_27191_4790# VDPWR 3.32e-19
C3065 ringtest_0.x4.net8 ringtest_0.x4._06_ 0.209874f
C3066 ringtest_0.x4.net8 a_24070_5852# 0.028641f
C3067 a_26808_4902# VDPWR 0.183021f
C3068 a_22392_5990# a_22139_5878# 3.39e-19
C3069 ringtest_0.counter3 a_21375_3867# 4.27e-20
C3070 muxtest_0.x1.x4.A muxtest_0.R5R6 1.64e-20
C3071 ringtest_0.x3.x2.GN4 VDPWR 1.23317f
C3072 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.clknet_0_clk 0.004956f
C3073 muxtest_0.x1.x3.GN3 ua[3] 0.014498f
C3074 muxtest_0.x1.x5.GN muxtest_0.x2.nselect2 4.76e-21
C3075 a_25421_6641# ringtest_0.x4.net9 3.61e-20
C3076 ringtest_0.x3.x2.GP1 m3_17032_8096# 3.25e-21
C3077 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._12_ 0.075464f
C3078 ringtest_0.x3.x2.GN3 m3_17046_7066# 0.016026f
C3079 ringtest_0.x4._24_ a_26913_4566# 0.002926f
C3080 ringtest_0.x4._16_ ringtest_0.x4._20_ 0.011071f
C3081 a_21399_5340# a_21509_4790# 0.010101f
C3082 muxtest_0.x1.x4.A VDPWR 15.014299f
C3083 a_21233_5340# a_21675_4790# 2.24e-19
C3084 ringtest_0.x4._22_ ringtest_0.x4.net5 4.26e-20
C3085 a_19794_32347# muxtest_0.x1.x3.GN4 3.22e-19
C3086 muxtest_0.x1.x3.GN3 a_20492_32319# 1.07e-20
C3087 a_22164_4362# a_22390_4566# 0.005961f
C3088 ringtest_0.x4.net8 a_23891_4790# 4.38e-20
C3089 ringtest_0.x4._11_ a_25761_5058# 0.028602f
C3090 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A 0.17253f
C3091 a_21465_9294# a_21780_9142# 7.84e-20
C3092 a_27065_5156# a_27273_4220# 0.003595f
C3093 a_19842_32287# muxtest_0.x1.x3.GN3 0.004289f
C3094 ringtest_0.counter7 a_22295_3867# 2.81e-20
C3095 a_21675_9686# a_21852_9416# 0.001655f
C3096 a_21465_9294# a_21561_9116# 0.310858f
C3097 ringtest_0.x4.net5 a_24135_3867# 0.001724f
C3098 ringtest_0.x4._19_ ringtest_0.x4._24_ 8.27e-21
C3099 a_27233_5058# ringtest_0.x4.net11 0.092457f
C3100 a_19666_31955# VDPWR 0.171399f
C3101 ringtest_0.x4._11_ a_21675_4790# 0.03376f
C3102 ringtest_0.x4.net6 ringtest_0.x4._15_ 0.117386f
C3103 a_25421_6641# ringtest_0.x4.net7 0.030401f
C3104 a_21840_5308# a_22097_5334# 0.036838f
C3105 muxtest_0.x1.x1.nSEL0 a_19114_31955# 0.03096f
C3106 ringtest_0.x4._15_ a_24895_4790# 2.57e-20
C3107 ringtest_0.x4._16_ a_21840_5308# 1.76e-20
C3108 a_23529_6422# ringtest_0.x4._05_ 4.91e-20
C3109 ringtest_0.x4._18_ ringtest_0.x4.clknet_1_1__leaf_clk 3.06e-19
C3110 ringtest_0.x4._17_ a_25421_6641# 0.019971f
C3111 a_24329_6640# a_24336_6544# 0.961627f
C3112 a_23949_6654# a_24465_6800# 1.28e-19
C3113 a_25336_4902# a_25083_4790# 3.39e-19
C3114 ringtest_0.x4._24_ a_26735_5334# 7.21e-19
C3115 ringtest_0.x3.x2.GP2 ringtest_0.counter7 1.13e-20
C3116 ringtest_0.x3.x2.GP3 ui_in[4] 0.003259f
C3117 muxtest_0.x1.x3.GN1 ui_in[0] 0.023343f
C3118 a_21465_8830# VDPWR 0.397883f
C3119 a_23381_4818# a_23467_4818# 0.006584f
C3120 ringtest_0.x4._13_ a_21399_5340# 1.58e-19
C3121 a_21785_5878# a_21233_5340# 0.002682f
C3122 ringtest_0.x4.net6 a_24926_5712# 0.001426f
C3123 a_27489_3702# ringtest_0.x4.counter[9] 0.109832f
C3124 muxtest_0.x2.x2.GP2 VDPWR 1.81003f
C3125 a_26367_5340# a_26201_4790# 2.64e-19
C3126 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A ringtest_0.x3.x1.nSEL1 2.53e-21
C3127 ringtest_0.x4._14_ a_23381_4584# 9.06e-21
C3128 a_26201_5340# ringtest_0.x4._09_ 1.11e-19
C3129 ringtest_0.x4._11_ a_21785_5878# 0.205946f
C3130 a_26721_4246# a_26895_3867# 2.21e-19
C3131 a_25083_4790# VDPWR 0.077706f
C3132 ringtest_0.x4._24_ ringtest_0.x4.net9 0.165357f
C3133 muxtest_0.x1.x3.GP2 ua[3] 0.023177f
C3134 a_25364_5878# a_25977_4220# 4.57e-20
C3135 a_22399_9142# ringtest_0.x4._11_ 2.48e-19
C3136 ringtest_0.x4.clknet_1_0__leaf_clk a_22245_8054# 0.00537f
C3137 a_21948_5156# VDPWR 0.285287f
C3138 ringtest_0.x4.net3 a_21852_8720# 0.005586f
C3139 a_26367_5340# a_26555_5334# 0.097994f
C3140 a_22052_9116# a_21845_8816# 6.88e-20
C3141 a_21852_9416# a_22052_8875# 1.26e-19
C3142 a_21845_9116# a_21852_8720# 3.36e-19
C3143 a_24715_5334# VDPWR 0.084103f
C3144 a_19842_32287# muxtest_0.x1.x3.GP2 2.95e-20
C3145 ringtest_0.x4._15_ a_22939_4584# 1.81e-19
C3146 ringtest_0.x4.net2 ringtest_0.x4.net3 1.28152f
C3147 ringtest_0.x4.net1 a_21465_8830# 0.081622f
C3148 ringtest_0.x4._15_ a_27169_6641# 8.98e-20
C3149 muxtest_0.R7R8 ua[0] 2.33155f
C3150 ringtest_0.x4.net7 ringtest_0.x4._24_ 2.68e-19
C3151 ringtest_0.x4.net2 a_21845_9116# 4.59e-19
C3152 ringtest_0.ring_out ringtest_0.x3.x2.GN1 4.6809f
C3153 a_26201_4790# a_27065_5156# 0.032244f
C3154 a_21951_5878# a_21509_4790# 1.21e-19
C3155 a_21785_5878# a_21675_4790# 3.23e-21
C3156 ringtest_0.x4._09_ a_27233_5058# 0.010518f
C3157 ringtest_0.x4._07_ a_24361_5340# 0.022853f
C3158 ringtest_0.x4._17_ ringtest_0.x4._24_ 0.004444f
C3159 ringtest_0.x4.net5 a_22021_4220# 0.006016f
C3160 ringtest_0.x4._22_ a_24527_5340# 0.015364f
C3161 a_24763_6143# a_24800_5334# 1.41e-19
C3162 ringtest_0.counter7 ringtest_0.x4._23_ 0.004833f
C3163 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A 0.025028f
C3164 ringtest_0.x3.x2.GP1 ringtest_0.x3.x2.GP3 0.001226f
C3165 ringtest_0.x4._04_ a_22983_5654# 0.002919f
C3166 ringtest_0.counter7 a_26367_4790# 5.88e-20
C3167 muxtest_0.R1R2 ui_in[4] 8.73e-20
C3168 muxtest_0.x2.x1.nSEL0 a_12425_24040# 2.51e-19
C3169 a_24361_5340# a_25055_3867# 1.7e-21
C3170 a_21780_8964# VDPWR 1.37e-19
C3171 muxtest_0.x2.x1.nSEL0 muxtest_0.x2.x2.GN1 0.004375f
C3172 a_22224_6244# a_22265_5308# 0.004197f
C3173 a_22392_5990# a_22097_5334# 0.004484f
C3174 a_24336_6544# a_24317_4942# 2.42e-19
C3175 ringtest_0.x4.clknet_0_clk ringtest_0.x4._22_ 0.003156f
C3176 ringtest_0.x4.clknet_1_0__leaf_clk a_22983_5654# 1.8e-20
C3177 muxtest_0.R7R8 muxtest_0.x2.x2.GN3 0.01204f
C3178 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GP3 2.78e-20
C3179 a_22392_5990# ringtest_0.x4._16_ 1.01e-19
C3180 muxtest_0.x1.x4.A a_12849_23648# 1.34e-19
C3181 ringtest_0.ring_out ui_in[6] 0.555069f
C3182 ringtest_0.x4._11_ ringtest_0.counter3 1.13e-19
C3183 uio_in[1] uio_in[0] 0.033505f
C3184 ringtest_0.x4.clknet_1_1__leaf_clk a_24800_5334# 0.033626f
C3185 ringtest_0.x4.clknet_0_clk a_23619_6788# 9.48e-20
C3186 ringtest_0.x4._13_ a_21951_5878# 7.99e-20
C3187 muxtest_0.x2.x1.nSEL1 VDPWR 0.649185f
C3188 ringtest_0.x4.net3 a_22399_8976# 4.27e-20
C3189 a_21981_8976# ringtest_0.x4._01_ 0.00226f
C3190 ringtest_0.x4.clknet_1_0__leaf_clk a_21591_6128# 0.001585f
C3191 a_26627_4246# a_26817_4566# 0.011458f
C3192 ringtest_0.x4._00_ ringtest_0.x4._11_ 0.003231f
C3193 muxtest_0.x1.x3.GN2 muxtest_0.x1.x5.A 0.429373f
C3194 a_27065_5156# a_27303_4246# 3.93e-20
C3195 a_13025_23980# ui_in[3] 0.279858f
C3196 ringtest_0.x4.net1 a_21780_8964# 1.42e-19
C3197 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A 5.04e-19
C3198 ringtest_0.x4.net7 a_26007_6788# 0.003849f
C3199 a_21840_5308# a_21587_5334# 3.39e-19
C3200 a_21399_5340# a_21798_5712# 8.12e-19
C3201 a_24527_5340# a_25225_5334# 0.192206f
C3202 a_24361_5340# a_26201_5340# 0.002059f
C3203 a_21948_5156# ringtest_0.x4.counter[2] 1.99e-20
C3204 a_24968_5308# a_25393_5308# 1.28e-19
C3205 a_19114_31955# muxtest_0.x1.x3.GN2 0.106131f
C3206 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._23_ 0.071442f
C3207 ringtest_0.x4._11_ ringtest_0.x4.net10 0.36244f
C3208 ringtest_0.x4.clknet_1_1__leaf_clk a_26367_4790# 0.031849f
C3209 VDPWR ua[0] 3.15952f
C3210 a_12849_23648# muxtest_0.x2.x2.GP2 3.07e-19
C3211 a_24336_6544# ringtest_0.x4._19_ 0.457296f
C3212 muxtest_0.x1.x3.GP3 ui_in[0] 2.74e-19
C3213 ringtest_0.x4.clknet_0_clk a_25225_5334# 0.013741f
C3214 ringtest_0.x4._15_ ringtest_0.x4.net5 0.016962f
C3215 ringtest_0.x4._03_ a_22765_4478# 1.19e-19
C3216 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP2 2.14737f
C3217 ringtest_0.x4.net4 a_22983_5654# 5.3e-19
C3218 ringtest_0.drv_out VDPWR 16.3479f
C3219 muxtest_0.x2.nselect2 ui_in[4] 0.001201f
C3220 ringtest_0.x4._11_ a_22775_5878# 8.02e-19
C3221 a_15575_12017# a_15749_12123# 0.006584f
C3222 a_17231_12017# ui_in[4] 0.125445f
C3223 ringtest_0.x3.x1.nSEL1 a_16155_12151# 9.57e-19
C3224 ringtest_0.x4._24_ a_27065_5334# 0.013075f
C3225 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GN1 0.034862f
C3226 ringtest_0.x4._11_ a_24627_6200# 4.38e-19
C3227 a_22541_5058# ringtest_0.x4.net5 0.13266f
C3228 ringtest_0.x4._08_ ringtest_0.x4._07_ 9.41e-21
C3229 muxtest_0.R3R4 ua[3] 0.039417f
C3230 ringtest_0.x4._11_ ringtest_0.x4.counter[4] 6.77e-20
C3231 ringtest_0.x4.net8 a_26895_3867# 7.5e-19
C3232 a_13675_24012# VDPWR 8.97e-19
C3233 ringtest_0.x4._18_ a_23993_5654# 6.01e-19
C3234 a_21951_5878# ringtest_0.x4.net8 0.001542f
C3235 muxtest_0.x2.x2.GN3 VDPWR 0.650589f
C3236 a_22392_5990# a_22649_6244# 0.036838f
C3237 a_23879_6940# a_24715_5334# 2.19e-20
C3238 ringtest_0.x4.net9 a_25977_4220# 9.8e-19
C3239 muxtest_0.x1.x3.GN4 muxtest_0.R2R3 0.127088f
C3240 a_23949_6654# a_23770_5308# 8.51e-20
C3241 ringtest_0.x4._01_ a_22228_8598# 5.75e-19
C3242 a_22052_8875# ringtest_0.x4._10_ 2.11e-19
C3243 ringtest_0.x4.net9 a_25719_4790# 0.001933f
C3244 muxtest_0.x1.x3.GN4 ui_in[1] 0.059771f
C3245 ringtest_0.x4.net4 a_22486_4246# 0.003167f
C3246 ringtest_0.x4._07_ a_25336_4902# 0.004454f
C3247 a_24329_6640# ringtest_0.x4._16_ 1.49e-19
C3248 a_24336_6544# ringtest_0.x4.net9 1.52e-20
C3249 ringtest_0.x4._22_ a_25168_5156# 0.002895f
C3250 ringtest_0.x3.x2.GP2 ui_in[3] 5.28e-19
C3251 muxtest_0.R3R4 m3_13316_18955# 1.46e-19
C3252 ringtest_0.x4._24_ a_26627_4246# 0.085832f
C3253 ringtest_0.x4._00_ a_22399_9142# 0.139872f
C3254 ringtest_0.x4._18_ ringtest_0.x4._04_ 0.003255f
C3255 ringtest_0.x4._24_ a_27149_5156# 8.56e-19
C3256 ringtest_0.x4.net7 a_25977_4220# 0.023542f
C3257 muxtest_0.x1.x5.GN muxtest_0.x1.x3.GN4 9.02e-19
C3258 muxtest_0.x1.x1.nSEL1 muxtest_0.x1.x3.GN3 0.012418f
C3259 ringtest_0.x4._23_ a_26367_4790# 0.031117f
C3260 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GN2 0.154394f
C3261 ringtest_0.x4._07_ VDPWR 0.311668f
C3262 a_24336_6544# ringtest_0.x4.net7 0.027472f
C3263 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.001676f
C3264 ringtest_0.x4.clknet_1_1__leaf_clk a_25593_5156# 0.044904f
C3265 ringtest_0.x4._06_ a_24361_5340# 0.091082f
C3266 ringtest_0.x4.net8 a_26808_5308# 8.61e-20
C3267 ringtest_0.x4._16_ a_24545_5878# 0.036674f
C3268 ringtest_0.x4._11_ a_25393_5308# 1.18e-19
C3269 a_25055_3867# VDPWR 0.307891f
C3270 ringtest_0.x4._17_ a_24336_6544# 0.050404f
C3271 a_16155_12151# ringtest_0.x3.x2.GN3 5.17e-20
C3272 ringtest_0.x3.x2.GN2 a_16707_12151# 3.11e-20
C3273 ringtest_0.x4.net2 ringtest_0.x4._03_ 5.34e-20
C3274 muxtest_0.x2.x1.nSEL1 a_12849_23648# 7.84e-19
C3275 ringtest_0.x3.x2.GN1 ringtest_0.x3.x2.GN3 0.002857f
C3276 ringtest_0.x4._08_ a_26201_5340# 0.097891f
C3277 a_25364_5878# ringtest_0.x4._16_ 0.001016f
C3278 a_24264_6788# VDPWR 4.18e-20
C3279 muxtest_0.x2.x1.nSEL0 ua[3] 7.05e-20
C3280 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ui_in[6] 0.108977f
C3281 ringtest_0.x4._03_ a_23381_4818# 2.2e-20
C3282 a_21509_4790# a_23809_4790# 1.62e-21
C3283 ringtest_0.x4._15_ a_24527_5340# 0.027322f
C3284 ringtest_0.x4.net6 a_26367_5340# 1.27e-19
C3285 a_21845_8816# a_21395_6940# 6.92e-20
C3286 a_25225_5334# a_25168_5156# 7.26e-19
C3287 muxtest_0.x1.x4.A muxtest_0.x1.x5.A 2.05508f
C3288 a_27273_4220# a_27489_3702# 1.29e-21
C3289 a_26817_4566# a_26721_4246# 1.26e-19
C3290 muxtest_0.x1.x3.GP1 muxtest_0.R7R8 4.13739f
C3291 ringtest_0.x4.clknet_0_clk ringtest_0.x4._15_ 4.05e-19
C3292 a_21561_8830# ringtest_0.x4._12_ 0.036321f
C3293 a_16203_12091# VDPWR 0.192568f
C3294 ringtest_0.x4.net8 a_23381_4584# 9.57e-20
C3295 ringtest_0.x4._11_ a_27191_4790# 9.67e-22
C3296 ringtest_0.x4.net11 a_26895_3867# 3.2e-20
C3297 ringtest_0.x4.net9 a_25677_5156# 8.89e-19
C3298 ringtest_0.x4._11_ a_26808_4902# 8.51e-19
C3299 ringtest_0.x4.counter[1] ua[1] 3.21e-19
C3300 ringtest_0.x4._16_ a_24317_4942# 1.3e-19
C3301 a_16707_12151# ui_in[3] 0.001558f
C3302 a_22265_5308# a_23899_5334# 2.67e-21
C3303 a_27233_5308# a_27065_5334# 0.310858f
C3304 a_22765_5308# a_22795_5334# 0.025037f
C3305 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._04_ 1.67e-21
C3306 a_24968_5308# a_24715_5334# 3.39e-19
C3307 a_24045_6654# ringtest_0.x4.net8 1.55e-19
C3308 ringtest_0.x3.x2.GN2 ui_in[3] 0.114345f
C3309 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A 0.159172f
C3310 a_26201_5340# VDPWR 0.711087f
C3311 ringtest_0.x4.net6 a_22765_4478# 5.34e-20
C3312 ringtest_0.x4._05_ a_24883_6800# 0.114695f
C3313 ringtest_0.x4._16_ a_23151_5334# 0.010038f
C3314 ringtest_0.x4._18_ ringtest_0.x4.net4 3.06e-19
C3315 a_24465_6800# a_24287_6422# 9.73e-19
C3316 ringtest_0.drv_out a_23879_6940# 0.318051f
C3317 ringtest_0.counter7 ringtest_0.x4.net4 6.88e-20
C3318 ringtest_0.x4.net7 a_25677_5156# 0.002598f
C3319 ringtest_0.x4._23_ a_25593_5156# 0.001187f
C3320 a_25593_5156# a_26367_4790# 2.56e-19
C3321 a_23949_6654# ringtest_0.x4.net6 1.76e-19
C3322 a_24729_4790# a_26555_4790# 4.76e-21
C3323 ringtest_0.x4.counter[5] VDPWR 0.439805f
C3324 a_12849_23648# muxtest_0.x2.x2.GN3 0.104151f
C3325 a_13025_23980# muxtest_0.x2.x2.GN1 3.78e-20
C3326 ringtest_0.x4._21_ ringtest_0.x4._07_ 4.77e-20
C3327 ringtest_0.x4.net7 a_23899_5334# 0.006434f
C3328 a_22224_6244# ringtest_0.x4._14_ 5.19e-22
C3329 ringtest_0.x4.net9 ringtest_0.x4.counter[9] 5.19e-19
C3330 m2_15612_11606# ui_in[3] 0.130999f
C3331 a_26749_6422# a_26808_5308# 2.48e-20
C3332 ringtest_0.x4._25_ a_26201_5340# 1.01e-19
C3333 ringtest_0.x3.nselect2 a_16579_11759# 1.29e-19
C3334 a_22164_4362# VDPWR 0.108683f
C3335 ringtest_0.counter3 ringtest_0.x4.counter[4] 0.07836f
C3336 ringtest_0.x4.net8 ringtest_0.x4.counter[6] 0.079257f
C3337 a_22224_6244# a_22319_6244# 0.007724f
C3338 a_22392_5990# a_22733_6244# 9.73e-19
C3339 ringtest_0.x4.net8 a_24699_6200# 0.003186f
C3340 ringtest_0.x4._17_ a_23899_5334# 9.12e-21
C3341 a_27233_5058# VDPWR 0.459668f
C3342 ringtest_0.counter3 a_23399_3867# 0.110188f
C3343 a_23529_6422# VDPWR 0.182648f
C3344 ringtest_0.x4._12_ a_21049_8598# 0.090947f
C3345 ringtest_0.x4.net4 a_22295_3867# 0.202764f
C3346 muxtest_0.x1.x3.GP1 muxtest_0.R5R6 0.122287f
C3347 ringtest_0.x4._19_ ringtest_0.x4._16_ 0.001191f
C3348 a_23770_5308# ringtest_0.x4._20_ 3.36e-20
C3349 ringtest_0.x4._18_ a_23837_5878# 0.002103f
C3350 ringtest_0.x4.net6 a_24004_6128# 0.074355f
C3351 a_21840_5308# ringtest_0.x4._03_ 0.009555f
C3352 a_21672_5334# a_21509_4790# 4.57e-19
C3353 ringtest_0.counter7 ringtest_0.x4._22_ 1.31e-20
C3354 a_21233_5340# a_21948_5156# 0.001041f
C3355 a_22765_4478# a_22939_4584# 0.006584f
C3356 a_22021_4220# a_22486_4246# 0.005941f
C3357 ringtest_0.x4.net8 a_24479_4790# 0.002158f
C3358 a_25977_4220# a_26627_4246# 0.010893f
C3359 a_21465_9294# ringtest_0.x4.net3 9.98e-20
C3360 ringtest_0.x4._11_ a_25083_4790# 0.016192f
C3361 muxtest_0.x1.x3.GP1 VDPWR 3.2848f
C3362 a_24699_6200# a_24729_4790# 5.07e-21
C3363 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GN3 0.08518f
C3364 a_21465_9294# a_21845_9116# 0.048748f
C3365 a_21561_9116# a_21852_9416# 0.194892f
C3366 ringtest_0.counter7 a_24135_3867# 2.81e-20
C3367 ringtest_0.x4.net9 a_27149_5334# 1.06e-19
C3368 a_20318_32213# VDPWR 0.217349f
C3369 ringtest_0.x4.net8 a_23809_4790# 7.44e-19
C3370 ringtest_0.x4._11_ a_21948_5156# 0.00274f
C3371 ringtest_0.ring_out ui_in[4] 0.016625f
C3372 a_22265_5308# a_22097_5334# 0.310858f
C3373 muxtest_0.x1.x1.nSEL0 a_19666_31955# 1.91e-20
C3374 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A 0.025028f
C3375 ringtest_0.x4._06_ VDPWR 0.273817f
C3376 ringtest_0.x4._16_ a_22265_5308# 7.03e-19
C3377 a_24336_6544# a_24536_6699# 0.074815f
C3378 a_24045_6654# ringtest_0.x4._05_ 9.72e-20
C3379 a_24329_6640# a_24465_6800# 0.136009f
C3380 a_25168_5156# a_25263_5156# 0.007724f
C3381 a_24070_5852# VDPWR 0.084816f
C3382 a_21395_6940# a_21399_5340# 1.82e-21
C3383 ringtest_0.x4.net6 a_23381_4818# 4.93e-21
C3384 ringtest_0.x4.net9 ringtest_0.x4._16_ 0.243936f
C3385 a_24763_6143# ringtest_0.x4._22_ 0.155189f
C3386 a_21845_8816# VDPWR 0.442439f
C3387 ringtest_0.x4._04_ ringtest_0.x4._02_ 1.6e-19
C3388 a_23809_4790# a_24729_4790# 2.37e-21
C3389 ringtest_0.x4._15_ a_22983_5654# 1.54e-19
C3390 ringtest_0.x4.net2 a_21055_5334# 0.002977f
C3391 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._02_ 0.254839f
C3392 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A ui_in[6] 6.29e-19
C3393 a_23399_3867# ringtest_0.x4.counter[4] 0.001146f
C3394 a_26640_5334# a_26201_4790# 1.73e-19
C3395 a_21675_4790# a_21948_5156# 0.081834f
C3396 a_23891_4790# VDPWR 2e-19
C3397 ringtest_0.x4.net7 ringtest_0.x4._16_ 5.07e-19
C3398 a_24465_6800# a_24545_5878# 1.71e-20
C3399 a_22164_4362# ringtest_0.x4.counter[2] 6.46e-19
C3400 a_22373_5156# VDPWR 0.179183f
C3401 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._22_ 0.031888f
C3402 ringtest_0.x3.x1.nSEL0 VDPWR 0.5228f
C3403 ringtest_0.x4.net3 a_21981_8976# 2.06e-19
C3404 ringtest_0.x4._17_ ringtest_0.x4._16_ 0.048058f
C3405 a_26808_5308# a_26766_5712# 4.62e-19
C3406 a_26640_5334# a_26555_5334# 0.037333f
C3407 ringtest_0.x4._05_ a_24699_6200# 3.16e-19
C3408 a_21852_9416# ringtest_0.x4._01_ 8.68e-20
C3409 a_21845_9116# a_21981_8976# 5.28e-20
C3410 ringtest_0.drv_out a_25925_6788# 1.34e-19
C3411 a_22052_9116# a_22052_8875# 0.013851f
C3412 muxtest_0.x2.x1.nSEL1 m2_11882_23495# 0.00815f
C3413 ringtest_0.x3.x2.GN4 ringtest_0.counter3 0.237196f
C3414 a_21767_5334# VDPWR 0.00331f
C3415 muxtest_0.x1.x3.GN1 muxtest_0.x1.x3.GP2 0.068989f
C3416 ringtest_0.x4.net1 a_21845_8816# 0.002755f
C3417 ringtest_0.ring_out ringtest_0.x3.x2.GP1 4.09516f
C3418 ringtest_0.x4.net2 a_21981_9142# 3.46e-19
C3419 a_12977_24040# muxtest_0.x2.x2.GP3 4.39e-19
C3420 a_21785_5878# a_21948_5156# 8.98e-19
C3421 a_22224_6244# a_21509_4790# 5.5e-20
C3422 a_26201_4790# a_26735_5156# 0.002698f
C3423 ringtest_0.x4._09_ a_26555_4790# 0.129132f
C3424 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GP3 0.004298f
C3425 ringtest_0.x4._07_ a_24968_5308# 0.011124f
C3426 ringtest_0.x4.net5 a_22765_4478# 0.081136f
C3427 ringtest_0.x4._22_ a_24800_5334# 0.006172f
C3428 ringtest_0.x4.clknet_1_0__leaf_clk a_22116_4902# 0.001507f
C3429 ringtest_0.x4.net6 ringtest_0.x4._20_ 0.00624f
C3430 muxtest_0.x2.nselect2 muxtest_0.x2.x2.GN4 1.53e-20
C3431 a_23349_6422# a_23529_6422# 0.185422f
C3432 a_22201_8964# VDPWR 0.002269f
C3433 ringtest_0.x4._20_ a_24895_4790# 0.003428f
C3434 a_26269_4612# VDPWR 0.001175f
C3435 ringtest_0.x4.net10 a_26808_4902# 1.26e-19
C3436 ringtest_0.x4._21_ ringtest_0.x4._06_ 0.224771f
C3437 a_13025_23980# ua[3] 9.59e-19
C3438 a_22817_6146# ringtest_0.x4._16_ 0.001048f
C3439 ringtest_0.x4.net4 ringtest_0.x4._02_ 1.19e-19
C3440 ringtest_0.counter7 ua[3] 1.17e-19
C3441 ringtest_0.x3.x1.nSEL1 ui_in[4] 0.272823f
C3442 a_24004_6128# a_23932_6128# 0.005941f
C3443 a_27489_3702# ringtest_0.x4.counter[8] 0.006251f
C3444 a_24070_5852# ringtest_0.x4._21_ 0.114705f
C3445 a_22139_5878# a_22319_6244# 0.001229f
C3446 muxtest_0.x1.x4.A a_13501_23906# 0.001685f
C3447 a_21395_6940# a_21951_5878# 1.63e-19
C3448 ringtest_0.x4.clknet_1_1__leaf_clk a_25225_5334# 0.024694f
C3449 ringtest_0.x4.net6 a_21840_5308# 6.4e-20
C3450 ringtest_0.x4.clknet_0_clk a_24685_6788# 4.62e-19
C3451 ringtest_0.drv_out ringtest_0.x4._11_ 1.2e-19
C3452 ringtest_0.x4._13_ a_22224_6244# 5.02e-20
C3453 ringtest_0.x4._23_ ringtest_0.x4._22_ 0.511385f
C3454 a_22499_4790# VDPWR 3.26e-19
C3455 ringtest_0.x4._22_ a_26367_4790# 3.15e-20
C3456 ringtest_0.x4._24_ ringtest_0.x4.net8 1.23e-20
C3457 a_27065_5334# a_27149_5334# 0.008508f
C3458 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4._04_ 0.005301f
C3459 a_22021_4220# a_22295_3867# 4.71e-19
C3460 a_25364_5878# a_26201_4790# 6.92e-20
C3461 muxtest_0.x1.x3.GN2 muxtest_0.x1.x4.A 0.429199f
C3462 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GP3 5.02073f
C3463 muxtest_0.x2.x2.GN1 ui_in[3] 0.021261f
C3464 a_23879_6940# ringtest_0.x4._06_ 1.96e-20
C3465 ringtest_0.x4.net7 a_26201_6788# 5.71e-19
C3466 ringtest_0.x4._17_ a_22649_6244# 1.03e-20
C3467 a_23879_6940# a_24070_5852# 3.15e-19
C3468 a_21672_5334# a_21798_5712# 0.005525f
C3469 a_24527_5340# a_26367_5340# 0.001861f
C3470 ringtest_0.x4.net6 a_26569_6422# 2.84e-19
C3471 a_19666_31955# muxtest_0.x1.x3.GN2 1.61e-19
C3472 ringtest_0.x4._17_ a_26201_6788# 3.01e-19
C3473 a_21399_5340# VDPWR 0.339296f
C3474 a_25364_5878# a_26555_5334# 9.53e-19
C3475 muxtest_0.x1.x1.nSEL1 a_18662_32213# 0.193944f
C3476 ringtest_0.x4.clknet_1_1__leaf_clk a_26640_5156# 3.02e-19
C3477 ringtest_0.x4.net4 a_22116_4902# 0.007782f
C3478 a_24465_6800# ringtest_0.x4._19_ 0.040707f
C3479 ringtest_0.x4._18_ ringtest_0.x4._15_ 0.045245f
C3480 ringtest_0.x4._05_ a_25421_6641# 0.121098f
C3481 muxtest_0.x2.x2.GP2 ua[2] 0.349855f
C3482 ringtest_0.counter7 ringtest_0.x4._15_ 0.003538f
C3483 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.001676f
C3484 ringtest_0.x4.net2 ringtest_0.x4.net5 7.09e-21
C3485 a_24968_5308# ringtest_0.x4.counter[5] 2.7e-21
C3486 muxtest_0.x1.x3.GN4 ui_in[0] 0.218694f
C3487 muxtest_0.x1.x1.nSEL1 m2_18699_31802# 0.00815f
C3488 ringtest_0.x4.net5 a_23963_4790# 1.04e-20
C3489 ringtest_0.x4._15_ a_27191_5712# 6.51e-20
C3490 a_17405_12123# ui_in[4] 8.84e-19
C3491 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.x2.GP1 1.21e-19
C3492 ringtest_0.x3.x2.GN3 ui_in[4] 0.273713f
C3493 ringtest_0.x4._11_ ringtest_0.x4._07_ 0.161717f
C3494 a_16027_11759# ringtest_0.x3.x2.GN2 0.106178f
C3495 a_21863_4790# a_22043_5156# 0.001229f
C3496 a_23381_4818# ringtest_0.x4.net5 4.5e-19
C3497 muxtest_0.x1.x3.GN3 muxtest_0.R1R2 4.03753f
C3498 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y ui_in[6] 3.49e-19
C3499 a_22817_6146# a_22649_6244# 0.310858f
C3500 muxtest_0.R7R8 muxtest_0.R4R5 0.286971f
C3501 a_22224_6244# ringtest_0.x4.net8 4.11e-20
C3502 uio_in[6] uio_in[5] 0.031023f
C3503 ringtest_0.x4.net9 a_27273_4220# 0.001158f
C3504 ringtest_0.x4._01_ ringtest_0.x4._10_ 0.002197f
C3505 a_24045_6654# a_24361_5340# 1.16e-21
C3506 ringtest_0.x4._15_ a_24763_6143# 1.57e-19
C3507 ringtest_0.x4.net4 ringtest_0.x4._04_ 0.689049f
C3508 ringtest_0.x4.net9 a_26766_4790# 0.002793f
C3509 muxtest_0.x1.x3.GN1 muxtest_0.R3R4 3.99705f
C3510 a_24536_6699# ringtest_0.x4._16_ 1.35e-21
C3511 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VDPWR 0.639695f
C3512 ringtest_0.x4._07_ a_25761_5058# 3.3e-20
C3513 a_24465_6800# ringtest_0.x4.net9 0.004659f
C3514 muxtest_0.x1.x3.GP2 muxtest_0.x1.x3.GP3 0.09552f
C3515 ringtest_0.x4.clknet_1_0__leaf_clk ringtest_0.x4.net4 0.158995f
C3516 ringtest_0.x4._22_ a_25593_5156# 6.29e-19
C3517 ringtest_0.x4.clknet_0_clk a_23949_6654# 0.002548f
C3518 ringtest_0.x4.net6 a_22392_5990# 3.85e-19
C3519 ringtest_0.x4.net2 a_21007_3867# 0.223155f
C3520 ringtest_0.x4._24_ a_26749_6422# 0.197975f
C3521 ringtest_0.x4._24_ ringtest_0.x4.net11 0.002712f
C3522 ringtest_0.x4.net6 a_24287_6422# 1.73e-19
C3523 a_16027_11759# ui_in[3] 0.246189f
C3524 ringtest_0.x4._23_ a_26640_5156# 0.011058f
C3525 a_26808_4902# a_27191_4790# 4.67e-20
C3526 ringtest_0.x4._05_ ringtest_0.x4._24_ 2.08e-20
C3527 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._15_ 0.471647f
C3528 a_26367_4790# a_26640_5156# 0.078545f
C3529 a_24465_6800# ringtest_0.x4.net7 0.035198f
C3530 ringtest_0.x4._14_ a_22097_5334# 2.97e-21
C3531 ringtest_0.x4.clknet_1_1__leaf_clk a_25263_5156# 0.001835f
C3532 ringtest_0.x4._06_ a_24968_5308# 0.001008f
C3533 ringtest_0.x4._16_ ringtest_0.x4._14_ 0.202586f
C3534 ringtest_0.x4.net8 a_27233_5308# 4.93e-20
C3535 ringtest_0.x4._11_ a_26201_5340# 3.54e-20
C3536 a_24699_6200# a_24361_5340# 0.001396f
C3537 ringtest_0.x4._17_ a_24465_6800# 0.016441f
C3538 ringtest_0.x3.x2.GN3 ringtest_0.x3.x2.GP1 0.001426f
C3539 a_26895_3867# VDPWR 0.298665f
C3540 a_21951_5878# VDPWR 0.302152f
C3541 ringtest_0.x4._08_ a_26808_5308# 0.047112f
C3542 ringtest_0.x4.net5 ringtest_0.x4._20_ 8.42e-21
C3543 a_24883_6800# VDPWR 0.084837f
C3544 muxtest_0.x1.x3.GP2 muxtest_0.R1R2 0.153531f
C3545 ringtest_0.x4.clknet_0_clk a_24004_6128# 2.03e-19
C3546 ringtest_0.x4._15_ a_24800_5334# 0.026278f
C3547 a_21509_4790# a_21863_4790# 0.062224f
C3548 muxtest_0.R5R6 muxtest_0.R4R5 2.29244f
C3549 ringtest_0.x4._22_ a_25441_4612# 0.002353f
C3550 a_22052_8875# a_21395_6940# 2.84e-19
C3551 a_21785_8054# ringtest_0.x4._10_ 0.107891f
C3552 ringtest_0.x4._13_ a_22139_5878# 5.97e-20
C3553 VDPWR ua[1] 17.382101f
C3554 ringtest_0.drv_out ringtest_0.counter3 1.91048f
C3555 a_25225_5334# a_25593_5156# 3.78e-19
C3556 a_26555_5334# a_26735_5334# 0.001229f
C3557 a_16755_12091# VDPWR 0.26222f
C3558 a_22224_6244# a_22390_4566# 4.44e-21
C3559 a_21852_8720# ringtest_0.x4._12_ 0.206007f
C3560 ringtest_0.x4.net8 a_25977_4220# 0.004343f
C3561 ringtest_0.x4._11_ a_22164_4362# 1e-19
C3562 muxtest_0.R4R5 VDPWR 1.56678f
C3563 muxtest_0.x1.x3.GP1 muxtest_0.x1.x5.A 0.353808f
C3564 ringtest_0.x4.net9 a_26201_4790# 0.11266f
C3565 ringtest_0.x4.net11 a_27815_3867# 0.003661f
C3566 ringtest_0.x4.net8 a_25719_4790# 5.67e-20
C3567 ringtest_0.x4._11_ a_27233_5058# 5.38e-21
C3568 ua[0] ua[2] 4.5205f
C3569 a_24336_6544# ringtest_0.x4.net8 4.93e-19
C3570 ringtest_0.x4.net2 ringtest_0.x4._12_ 0.10227f
C3571 a_24800_5334# a_24926_5712# 0.005525f
C3572 ringtest_0.x4._11_ a_23529_6422# 0.001495f
C3573 a_19114_31955# muxtest_0.x1.x3.GP1 9.8e-19
C3574 a_26808_5308# VDPWR 0.180852f
C3575 ringtest_0.x4._15_ ringtest_0.x4._23_ 0.683594f
C3576 ringtest_0.x4.net6 a_25149_4220# 0.211407f
C3577 a_24329_6640# a_24712_6422# 0.001632f
C3578 ua[3] ui_in[3] 0.554156f
C3579 ringtest_0.x4._24_ ringtest_0.x4._09_ 0.151845f
C3580 a_18662_32213# muxtest_0.x1.x3.GN1 0.128677f
C3581 ringtest_0.x4._15_ a_26367_4790# 0.036316f
C3582 muxtest_0.R7R8 ui_in[2] 0.054741f
C3583 ringtest_0.x4.net7 a_26201_4790# 0.007864f
C3584 a_24895_4790# a_25149_4220# 0.002313f
C3585 a_24329_6640# ringtest_0.x4.net6 0.001597f
C3586 muxtest_0.x1.x3.GN1 m2_18699_31802# 0.06935f
C3587 a_13501_23906# a_13675_24012# 0.006584f
C3588 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A 0.025028f
C3589 muxtest_0.x2.x2.GN1 a_12425_24040# 1.22e-20
C3590 a_13501_23906# muxtest_0.x2.x2.GN3 1.07e-20
C3591 a_12019_24012# muxtest_0.x2.x2.GN2 8.86e-19
C3592 muxtest_0.x2.x2.GN3 ua[2] 0.429994f
C3593 a_21675_4790# a_22164_4362# 0.010312f
C3594 a_22116_4902# a_22021_4220# 1.66e-20
C3595 a_24329_6640# a_24895_4790# 4.79e-20
C3596 ringtest_0.x4._24_ a_26766_5712# 9.29e-19
C3597 muxtest_0.x1.x4.A muxtest_0.x2.x2.GP2 1.19e-20
C3598 ringtest_0.x4.net8 a_24986_5878# 1.76e-19
C3599 a_27065_5334# a_27273_4220# 9.49e-21
C3600 a_27233_5308# ringtest_0.x4.net11 1.16e-19
C3601 ringtest_0.x3.nselect2 a_17231_12017# 9.77e-20
C3602 ringtest_0.x4._11_ ringtest_0.x4._06_ 0.020042f
C3603 a_23381_4584# VDPWR 0.241858f
C3604 a_21675_9686# VDPWR 0.262771f
C3605 a_22224_6244# a_22350_5878# 0.005525f
C3606 muxtest_0.x1.x3.GN4 muxtest_0.x2.x2.GN4 3.13e-20
C3607 a_21951_5878# ringtest_0.x4._21_ 2.75e-21
C3608 ringtest_0.x4.net9 a_27303_4246# 0.005829f
C3609 a_21785_8054# a_21867_8054# 0.005167f
C3610 ringtest_0.x4._11_ a_24070_5852# 0.002559f
C3611 a_26555_4790# VDPWR 0.077654f
C3612 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ui_in[6] 1.67e-19
C3613 ringtest_0.x4._19_ a_23770_5308# 8.51e-20
C3614 muxtest_0.x1.x3.GP3 muxtest_0.R3R4 0.384927f
C3615 a_24045_6654# VDPWR 0.17352f
C3616 a_21852_8720# a_22245_8054# 0.011211f
C3617 ringtest_0.x4.net6 a_24545_5878# 0.00514f
C3618 ringtest_0.x4._12_ a_22399_8976# 0.023132f
C3619 a_21845_8816# ringtest_0.x4._11_ 9.54e-19
C3620 muxtest_0.x2.x2.GP2 m3_13302_19985# 0.005314f
C3621 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VDPWR 0.637448f
C3622 ringtest_0.x4.net6 a_25364_5878# 0.047825f
C3623 a_22097_5334# a_21509_4790# 0.002525f
C3624 ringtest_0.x4.net2 a_22245_8054# 3.45e-20
C3625 ringtest_0.x4.counter[2] ua[1] 3.21e-19
C3626 a_23381_4584# a_23467_4584# 0.006584f
C3627 a_26627_4246# a_27273_4220# 0.016298f
C3628 ringtest_0.x4._11_ a_23891_4790# 0.002312f
C3629 a_25364_5878# a_24895_4790# 1.98e-20
C3630 ringtest_0.x4._16_ a_21509_4790# 1.96e-20
C3631 ringtest_0.x4.net11 a_25977_4220# 1.29e-21
C3632 a_21233_5340# a_21767_5334# 0.002698f
C3633 a_21465_9294# a_21981_9142# 1.28e-19
C3634 ringtest_0.counter7 a_25975_3867# 8.66e-19
C3635 a_21852_9416# a_21845_9116# 0.966391f
C3636 a_22392_5990# ringtest_0.x4.net5 1.47e-21
C3637 muxtest_0.x1.x1.nSEL0 muxtest_0.x1.x3.GP1 6.21e-20
C3638 ringtest_0.x4._11_ a_22373_5156# 0.045224f
C3639 muxtest_0.x1.x5.GN a_19242_32347# 1.08e-19
C3640 muxtest_0.x2.x2.GP1 muxtest_0.x2.x2.GP3 0.001226f
C3641 muxtest_0.R5R6 ui_in[2] 2.39e-19
C3642 ringtest_0.x4.net1 a_21675_9686# 0.073427f
C3643 a_22265_5308# a_23770_5308# 1e-20
C3644 muxtest_0.x1.x1.nSEL1 a_18836_32319# 0.00175f
C3645 a_23879_6940# a_24883_6800# 8.9e-19
C3646 ringtest_0.x4.net6 a_24551_4790# 7.29e-19
C3647 ringtest_0.x4._15_ a_25593_5156# 1.98e-20
C3648 ringtest_0.x4.net8 a_23899_5334# 2.79e-20
C3649 ringtest_0.x4._11_ a_21767_5334# 3.45e-19
C3650 ringtest_0.x4._16_ a_22765_5308# 0.243866f
C3651 a_24336_6544# ringtest_0.x4._05_ 0.181338f
C3652 a_24536_6699# a_24465_6800# 0.239923f
C3653 ringtest_0.x4.counter[6] VDPWR 0.448598f
C3654 a_24699_6200# VDPWR 0.253923f
C3655 a_21395_6940# a_21672_5334# 7.35e-19
C3656 ringtest_0.x4.net6 a_24317_4942# 0.173962f
C3657 muxtest_0.R3R4 muxtest_0.R1R2 0.184502f
C3658 VDPWR ui_in[2] 4.46272f
C3659 muxtest_0.x2.x2.GN2 ui_in[4] 0.108808f
C3660 ringtest_0.drv_out a_25393_5308# 1.4e-22
C3661 a_22052_8875# VDPWR 0.270616f
C3662 a_24317_4942# a_24895_4790# 0.00145f
C3663 ringtest_0.x4.net9 ringtest_0.x4.counter[8] 2.39e-19
C3664 ringtest_0.x4.net6 a_23151_5334# 7.79e-20
C3665 ringtest_0.x4._15_ a_23993_5654# 0.004604f
C3666 ringtest_0.x4.net8 ringtest_0.x4.counter[9] 1.68e-20
C3667 ringtest_0.x4.net3 ringtest_0.x4._14_ 0.471315f
C3668 a_21675_4790# a_22373_5156# 0.195152f
C3669 a_22116_4902# a_22541_5058# 1.28e-19
C3670 a_27065_5334# a_26201_4790# 1.29e-19
C3671 a_27233_5308# ringtest_0.x4._09_ 5.87e-19
C3672 ringtest_0.x4.net7 a_23770_5308# 0.142058f
C3673 a_22399_8976# a_22245_8054# 6.31e-19
C3674 a_21785_5878# a_24070_5852# 1.55e-21
C3675 a_24479_4790# VDPWR 3.4e-19
C3676 ringtest_0.x4._11_ a_26269_4612# 0.006396f
C3677 ringtest_0.x4.clknet_0_clk a_26569_6422# 2.96e-20
C3678 ringtest_0.x4._17_ a_23770_5308# 1.33e-19
C3679 a_21465_8830# a_21780_8964# 7.84e-20
C3680 a_23809_4790# VDPWR 0.207983f
C3681 muxtest_0.x1.x3.GN3 muxtest_0.R6R7 0.260987f
C3682 a_26201_5340# ringtest_0.x4.net10 4.73e-19
C3683 a_24045_6654# ringtest_0.x4._21_ 9.57e-19
C3684 ringtest_0.x4._15_ ringtest_0.x4._04_ 3.75e-19
C3685 ringtest_0.x4.net4 a_22021_4220# 0.021386f
C3686 a_21981_9142# a_21981_8976# 0.013661f
C3687 ringtest_0.x4.clknet_1_0__leaf_clk a_21561_8830# 0.044938f
C3688 a_22795_5334# VDPWR 0.260656f
C3689 ringtest_0.x4._15_ a_25441_4612# 3.42e-21
C3690 ringtest_0.x4.net1 a_22052_8875# 1.33e-19
C3691 ringtest_0.x4._11_ a_22499_4790# 5.7e-19
C3692 ringtest_0.drv_out ringtest_0.x3.x2.GN4 0.071598f
C3693 ringtest_0.x4._09_ a_25977_4220# 1.89e-19
C3694 a_26201_4790# a_26627_4246# 9.12e-19
C3695 muxtest_0.x1.x4.A ua[0] 4.51511f
C3696 a_21425_9686# a_21675_9686# 0.025037f
C3697 ringtest_0.x4.net8 a_27149_5334# 2.29e-20
C3698 ringtest_0.x4._04_ a_22541_5058# 7.11e-19
C3699 a_21785_5878# a_22373_5156# 0.001131f
C3700 ringtest_0.x4._19_ ringtest_0.x4.net6 0.04173f
C3701 ringtest_0.x4._07_ a_25393_5308# 0.008579f
C3702 ringtest_0.x4.net5 a_25149_4220# 1.18e-20
C3703 ringtest_0.x4._22_ a_25225_5334# 1.1e-21
C3704 a_21233_5340# a_21399_5340# 0.968904f
C3705 ringtest_0.x4.clknet_1_0__leaf_clk a_22541_5058# 1.1e-19
C3706 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.001676f
C3707 ringtest_0.x4._18_ a_23949_6654# 0.006776f
C3708 a_21803_8598# VDPWR 0.004458f
C3709 ringtest_0.x4._20_ a_25168_5156# 9.2e-20
C3710 a_22649_6244# a_22765_5308# 0.001534f
C3711 a_23879_6940# a_24045_6654# 0.017149f
C3712 a_16579_11759# ringtest_0.x3.x2.GP2 3.07e-19
C3713 ringtest_0.x4._11_ a_21399_5340# 0.008371f
C3714 m3_13302_19985# ua[0] 0.003764f
C3715 ringtest_0.x4.net10 a_27233_5058# 0.008159f
C3716 muxtest_0.x2.x2.GN1 ua[3] 4.69116f
C3717 ringtest_0.counter3 m3_17036_9140# 2.1e-20
C3718 ringtest_0.x4.net8 ringtest_0.x4._16_ 0.193029f
C3719 muxtest_0.x1.x4.A a_13675_24012# 2.9e-19
C3720 muxtest_0.x1.x4.A muxtest_0.x2.x2.GN3 8.22e-19
C3721 a_24699_6200# ringtest_0.x4._21_ 0.001146f
C3722 ringtest_0.x4.counter[4] ringtest_0.x4.counter[5] 0.068962f
C3723 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[6] 5.64e-20
C3724 a_25421_6641# VDPWR 0.208917f
C3725 ringtest_0.x4.clknet_1_1__leaf_clk a_26367_5340# 0.026802f
C3726 ringtest_0.x4.net6 a_22265_5308# 6.37e-19
C3727 ringtest_0.x4.clknet_0_clk a_24287_6422# 2.01e-19
C3728 muxtest_0.x2.x2.GP2 ua[0] 4.069f
C3729 ringtest_0.x4._22_ a_26640_5156# 0.004398f
C3730 muxtest_0.x1.x3.GP2 muxtest_0.R6R7 4.11376f
C3731 ringtest_0.x4.net11 ringtest_0.x4.counter[9] 0.066386f
C3732 ringtest_0.x4.net3 ringtest_0.x4._10_ 0.003052f
C3733 a_21587_5334# a_21509_4790# 2.5e-19
C3734 ringtest_0.x4.net6 ringtest_0.x4.net9 0.566537f
C3735 ringtest_0.x4._23_ a_25975_3867# 2.99e-20
C3736 muxtest_0.x2.x2.GN3 m3_13302_19985# 0.087318f
C3737 ringtest_0.x4.clknet_1_0__leaf_clk a_21049_8598# 3.26e-19
C3738 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VDPWR 0.637284f
C3739 ringtest_0.x4._16_ a_24729_4790# 1.25e-20
C3740 ringtest_0.x4.net9 a_24895_4790# 0.017191f
C3741 ringtest_0.counter7 m3_17032_8096# 6.07e-21
C3742 a_21399_5340# a_21675_4790# 6.25e-19
C3743 ringtest_0.x4.net11 a_27491_4566# 0.001149f
C3744 ringtest_0.x4._24_ ringtest_0.x4._08_ 0.423487f
C3745 ringtest_0.x4._15_ ringtest_0.x4.net4 0.003757f
C3746 ringtest_0.x4._00_ a_21845_8816# 8.76e-20
C3747 muxtest_0.x1.x3.GN2 muxtest_0.x1.x3.GP1 4.57902f
C3748 ringtest_0.x4._18_ a_24004_6128# 5.77e-19
C3749 muxtest_0.x1.x3.GN3 muxtest_0.x1.x3.GN4 0.190572f
C3750 a_23879_6940# a_24699_6200# 6.61e-19
C3751 ringtest_0.x4._21_ a_23809_4790# 0.087922f
C3752 a_19794_32347# VDPWR 0.001496f
C3753 a_25393_5308# a_26201_5340# 4.62e-19
C3754 a_25421_6641# ringtest_0.x4._25_ 6.03e-21
C3755 muxtest_0.x1.x3.GN1 a_18836_32319# 0.001144f
C3756 a_20318_32213# muxtest_0.x1.x3.GN2 7.58e-21
C3757 ringtest_0.x4._17_ a_24712_6422# 0.002153f
C3758 a_21672_5334# VDPWR 0.256539f
C3759 ringtest_0.x4.net6 ringtest_0.x4.net7 0.905861f
C3760 ringtest_0.x4.net4 a_22541_5058# 0.020834f
C3761 muxtest_0.x1.x1.nSEL1 a_19290_32287# 0.041068f
C3762 ringtest_0.x4.clknet_1_1__leaf_clk a_27065_5156# 2.2e-19
C3763 muxtest_0.x2.x2.GN3 muxtest_0.x2.x2.GP2 2.65608f
C3764 ringtest_0.ring_out ringtest_0.x3.nselect2 0.006614f
C3765 ringtest_0.x4.net7 a_24895_4790# 0.030766f
C3766 ringtest_0.x4.net3 a_21509_4790# 0.005671f
C3767 ringtest_0.x4._17_ ringtest_0.x4.net6 0.277113f
C3768 a_23949_6654# ringtest_0.x4.clknet_1_1__leaf_clk 1.77e-20
C3769 ringtest_0.x4.net2 ringtest_0.counter7 6.88e-20
C3770 muxtest_0.R7R8 muxtest_0.x2.x2.GP3 0.17349f
C3771 ringtest_0.x4._17_ a_24895_4790# 6.74e-21
C3772 a_16579_11759# a_16707_12151# 0.004764f
C3773 a_21785_5878# a_21399_5340# 1.36e-19
C3774 a_21951_5878# a_21233_5340# 9.16e-19
C3775 a_16579_11759# ringtest_0.x3.x2.GN2 1.63e-19
C3776 ringtest_0.x4._18_ a_23381_4818# 1.7e-19
C3777 a_22097_5334# a_22390_4566# 3.78e-21
C3778 ringtest_0.x4._23_ a_26367_5340# 0.031087f
C3779 ringtest_0.x4._24_ VDPWR 0.670774f
C3780 a_26201_5340# a_26808_4902# 1.99e-20
C3781 a_26367_5340# a_26367_4790# 0.027195f
C3782 a_22649_6244# ringtest_0.x4.net8 3.5e-19
C3783 ringtest_0.x4._16_ a_22390_4566# 3.76e-19
C3784 ringtest_0.x4._11_ a_21951_5878# 0.082924f
C3785 muxtest_0.x1.x5.A muxtest_0.R4R5 4.5151f
C3786 ringtest_0.x4.net3 a_21867_8054# 1.25e-19
C3787 a_24336_6544# a_24361_5340# 1.6e-20
C3788 a_24329_6640# a_24527_5340# 3.93e-19
C3789 ringtest_0.x4._15_ a_23837_5878# 9.44e-19
C3790 ringtest_0.x4._15_ ringtest_0.x4._22_ 0.422897f
C3791 ringtest_0.x4._11_ a_24883_6800# 7.39e-21
C3792 ringtest_0.x4._05_ ringtest_0.x4._16_ 0.001611f
C3793 ringtest_0.x4._07_ a_25083_4790# 0.128255f
C3794 ringtest_0.x3.x2.GP2 m3_17032_8096# 0.005314f
C3795 ringtest_0.x4.net3 ringtest_0.x4._13_ 0.031667f
C3796 ringtest_0.x4.clknet_0_clk a_24329_6640# 0.043419f
C3797 a_23891_4790# ringtest_0.x4.counter[4] 4.37e-20
C3798 a_21465_9294# ringtest_0.x4._12_ 6.08e-20
C3799 ringtest_0.x4.clknet_1_1__leaf_clk a_24004_6128# 0.007927f
C3800 muxtest_0.x1.x3.GN4 muxtest_0.x1.x3.GP2 0.059353f
C3801 ringtest_0.x4.net6 a_22817_6146# 0.129987f
C3802 ringtest_0.x4._14_ ringtest_0.x4._03_ 0.071143f
C3803 ringtest_0.x4._24_ ringtest_0.x4._25_ 0.095329f
C3804 a_25593_5156# a_25975_3867# 3.85e-20
C3805 a_25083_4790# a_25055_3867# 7.39e-20
C3806 ringtest_0.x4._09_ a_27491_4566# 0.002954f
C3807 a_16579_11759# ui_in[3] 0.086353f
C3808 ringtest_0.x4.net7 a_27169_6641# 2.85e-19
C3809 a_27233_5058# a_27191_4790# 7.84e-20
C3810 ringtest_0.x4._23_ a_27065_5156# 0.006274f
C3811 a_26367_4790# a_27065_5156# 0.194892f
C3812 a_26808_4902# a_27233_5058# 1.28e-19
C3813 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A ui_in[4] 2.42e-19
C3814 ringtest_0.x4._06_ a_25393_5308# 1.75e-19
C3815 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A 0.025028f
C3816 a_23879_6940# a_25421_6641# 1.59e-19
C3817 a_24699_6200# a_24968_5308# 1e-18
C3818 a_27815_3867# VDPWR 0.270825f
C3819 ringtest_0.x3.x2.GP3 ringtest_0.counter7 0.165274f
C3820 muxtest_0.x2.x1.nSEL1 muxtest_0.x2.x2.GN3 0.012418f
C3821 a_11845_23906# muxtest_0.x2.x2.GN2 0.039612f
C3822 a_22224_6244# VDPWR 0.253899f
C3823 ringtest_0.x4.clknet_1_1__leaf_clk a_23381_4818# 2.67e-20
C3824 ringtest_0.x4._08_ a_27233_5308# 0.004928f
C3825 a_27149_5334# ringtest_0.x4._09_ 1.2e-19
C3826 a_22350_5878# ringtest_0.x4._16_ 2.63e-21
C3827 a_26007_6788# VDPWR 0.001434f
C3828 ringtest_0.x4.clknet_0_clk a_25364_5878# 0.316676f
C3829 ringtest_0.x3.x1.nSEL1 ringtest_0.x3.nselect2 0.047548f
C3830 muxtest_0.x2.x2.GP3 VDPWR 1.78328f
C3831 ringtest_0.x4._15_ a_25225_5334# 0.0351f
C3832 ringtest_0.x3.x1.nSEL0 a_15575_12017# 0.081627f
C3833 ringtest_0.x4._22_ a_26173_4612# 0.001961f
C3834 muxtest_0.R7R8 muxtest_0.R2R3 0.215077f
C3835 ringtest_0.x4._01_ a_21395_6940# 3.77e-19
C3836 muxtest_0.R7R8 ui_in[1] 4.98e-22
C3837 a_21785_5878# a_21951_5878# 0.966818f
C3838 a_16155_12151# VDPWR 2.96e-19
C3839 ringtest_0.x3.x2.GN1 VDPWR 1.47002f
C3840 a_21981_8976# ringtest_0.x4._12_ 0.039032f
C3841 ringtest_0.x4._11_ a_23381_4584# 0.002917f
C3842 a_22265_5308# ringtest_0.x4.net5 6.71e-21
C3843 muxtest_0.x2.x2.GN3 ua[0] 0.214839f
C3844 muxtest_0.x1.x3.GP1 muxtest_0.x1.x4.A 0.354981f
C3845 ringtest_0.x3.x2.GN4 m3_17036_9140# 7.17e-19
C3846 ringtest_0.x4._11_ a_26555_4790# 2.79e-20
C3847 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VDPWR 0.637855f
C3848 ringtest_0.x3.x2.GN2 m3_17032_8096# 0.016745f
C3849 a_24361_5340# a_23899_5334# 1.44e-19
C3850 a_24465_6800# ringtest_0.x4.net8 0.00192f
C3851 muxtest_0.x1.x5.GN muxtest_0.R7R8 0.558172f
C3852 ringtest_0.x4._17_ a_23932_6128# 0.002503f
C3853 ringtest_0.x4._11_ a_24045_6654# 1.82e-19
C3854 a_27233_5308# VDPWR 0.486506f
C3855 a_19666_31955# muxtest_0.x1.x3.GP1 1.19e-20
C3856 ringtest_0.x4.clknet_1_1__leaf_clk a_26375_4612# 5.67e-20
C3857 a_24536_6699# a_24712_6422# 0.007724f
C3858 ringtest_0.x4.net6 a_26627_4246# 5.59e-20
C3859 ringtest_0.x4._15_ a_22021_4220# 3.5e-20
C3860 ringtest_0.x4._15_ a_26640_5156# 0.001788f
C3861 a_19290_32287# muxtest_0.x1.x3.GN1 1.45e-19
C3862 a_25168_5156# a_25149_4220# 1.83e-19
C3863 muxtest_0.x1.x5.A ui_in[2] 5.67943f
C3864 VDPWR ui_in[6] 1.09983f
C3865 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B ringtest_0.x3.nselect2 2.88e-20
C3866 a_12977_24040# muxtest_0.x2.x2.GN4 3.22e-19
C3867 muxtest_0.x2.x2.GN3 a_13675_24012# 1.07e-20
C3868 a_25336_4902# a_25719_4790# 4.67e-20
C3869 a_24536_6699# ringtest_0.x4.net6 6.81e-19
C3870 muxtest_0.x2.x2.GN2 muxtest_0.x2.x2.GN4 8.84e-19
C3871 ringtest_0.x3.x2.GP2 ringtest_0.x3.x2.GP3 0.031766f
C3872 muxtest_0.x2.x2.GP1 ui_in[4] 0.001143f
C3873 a_21948_5156# a_22164_4362# 0.003601f
C3874 ua[3] ua[6] 0.008019f
C3875 ringtest_0.x4.clknet_1_1__leaf_clk ringtest_0.x4._20_ 0.0051f
C3876 a_24329_6640# a_25168_5156# 7.91e-22
C3877 a_19114_31955# ui_in[2] 8.66e-20
C3878 a_12297_23648# ui_in[4] 0.03417f
C3879 ringtest_0.x3.x1.nSEL0 ringtest_0.x3.x2.GN4 2.26e-20
C3880 ringtest_0.x3.nselect2 ringtest_0.x3.x2.GN3 7.39e-21
C3881 a_21780_9142# VDPWR 1.77e-19
C3882 a_25977_4220# VDPWR 0.418373f
C3883 a_21561_9116# VDPWR 0.189203f
C3884 ringtest_0.x4._11_ ringtest_0.x4.counter[6] 0.002692f
C3885 a_21785_8054# a_21395_6940# 5.68e-19
C3886 ringtest_0.x4._10_ a_21939_8054# 5.49e-20
C3887 a_25719_4790# VDPWR 1.93e-19
C3888 ringtest_0.x4._11_ a_24699_6200# 0.042839f
C3889 uio_in[0] ui_in[7] 0.031023f
C3890 ringtest_0.x4._19_ a_24527_5340# 4.93e-21
C3891 a_21509_4790# ringtest_0.x4._03_ 0.095111f
C3892 a_24336_6544# VDPWR 0.310723f
C3893 ringtest_0.x4.net2 ringtest_0.x4._02_ 0.035742f
C3894 ringtest_0.x4.net3 ringtest_0.x4.counter[1] 0.103986f
C3895 muxtest_0.x1.x3.GN4 muxtest_0.R3R4 0.237766f
C3896 muxtest_0.R2R3 VDPWR 1.6072f
C3897 ringtest_0.x4.clknet_0_clk ringtest_0.x4._19_ 0.038005f
C3898 ringtest_0.x4._04_ a_22765_4478# 1.25e-20
C3899 a_21465_8830# a_21845_8816# 0.048748f
C3900 VDPWR ui_in[1] 2.66846f
C3901 ringtest_0.x4.net3 a_22390_4566# 9.94e-20
C3902 ringtest_0.counter3 ua[1] 4.52195f
C3903 muxtest_0.x1.x5.GN muxtest_0.R5R6 7.03e-21
C3904 ringtest_0.x4._23_ a_26375_4612# 1.08e-20
C3905 ringtest_0.x4.net8 a_26201_4790# 3.27e-19
C3906 a_25761_5058# ringtest_0.x4.counter[6] 4.54e-21
C3907 ringtest_0.x4._11_ a_24479_4790# 0.001677f
C3908 a_21981_9142# a_22201_9142# 4.62e-19
C3909 ringtest_0.x4.net11 a_27273_4220# 0.088145f
C3910 a_21845_9116# a_22052_9116# 0.273138f
C3911 a_21561_9116# a_21803_9508# 0.008508f
C3912 a_21233_5340# a_22795_5334# 2.77e-19
C3913 ringtest_0.x4._18_ a_22392_5990# 1.41e-19
C3914 ringtest_0.counter7 a_27489_3702# 3.7e-19
C3915 a_21852_9416# a_21981_9142# 0.110715f
C3916 ringtest_0.x4.net1 a_21780_9142# 2.14e-19
C3917 ringtest_0.x4._11_ a_23809_4790# 0.222369f
C3918 ringtest_0.x4._14_ a_21055_5334# 6.31e-19
C3919 muxtest_0.x1.x5.GN VDPWR 3.74211f
C3920 ringtest_0.x4.net1 a_21561_9116# 0.017118f
C3921 ringtest_0.x4.clknet_1_1__leaf_clk a_26569_6422# 7.87e-19
C3922 a_22111_10993# a_21852_9416# 4.65e-23
C3923 ringtest_0.x4.net10 a_26895_3867# 2.65e-20
C3924 ringtest_0.x4._06_ a_24715_5334# 0.114717f
C3925 a_24986_5878# VDPWR 1.76e-19
C3926 ringtest_0.x4.net8 a_26555_5334# 1.28e-19
C3927 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A ui_in[4] 8.27e-22
C3928 ringtest_0.x4._11_ a_22795_5334# 2.49e-20
C3929 a_12849_23648# muxtest_0.x2.x2.GP3 0.00144f
C3930 ringtest_0.x4._16_ a_24361_5340# 1.57e-19
C3931 a_24465_6800# ringtest_0.x4._05_ 0.001005f
C3932 ringtest_0.x4.net9 a_24527_5340# 0.002182f
C3933 a_24729_4790# a_26201_4790# 0.003146f
C3934 a_22139_5878# VDPWR 0.093135f
C3935 a_16707_12151# ringtest_0.x3.x2.GP3 4.39e-19
C3936 a_25336_4902# a_25677_5156# 9.73e-19
C3937 ua[2] ua[1] 1.12657f
C3938 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A 0.001676f
C3939 ringtest_0.x4._15_ a_22541_5058# 2.99e-20
C3940 ringtest_0.x3.x2.GN2 ringtest_0.x3.x2.GP3 0.004296f
C3941 muxtest_0.x2.nselect2 a_13025_23980# 6.01e-20
C3942 muxtest_0.x1.x1.nSEL0 ui_in[2] 0.131256f
C3943 ringtest_0.x4._01_ VDPWR 0.464547f
C3944 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net9 0.132797f
C3945 ringtest_0.x4._07_ a_25055_3867# 7.51e-19
C3946 ringtest_0.x4._15_ a_24926_5712# 0.002542f
C3947 ringtest_0.x4._22_ a_25975_3867# 2.78e-19
C3948 ringtest_0.x4._14_ a_22939_4584# 5.76e-19
C3949 ringtest_0.x4.net7 a_24527_5340# 0.456298f
C3950 a_21007_3867# ringtest_0.x4.counter[0] 0.109791f
C3951 ringtest_0.x4._04_ a_24004_6128# 3.15e-21
C3952 a_25677_5156# VDPWR 0.004404f
C3953 ringtest_0.x4._17_ a_24527_5340# 1.22e-20
C3954 a_21863_4790# VDPWR 0.079882f
C3955 muxtest_0.x1.x3.GN2 muxtest_0.R4R5 0.116214f
C3956 ringtest_0.x4.clknet_0_clk ringtest_0.x4.net7 0.043959f
C3957 a_26808_5308# ringtest_0.x4.net10 2.56e-19
C3958 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VDPWR 0.637064f
C3959 ringtest_0.x4.net4 a_22765_4478# 0.130038f
C3960 ringtest_0.x3.x2.GP3 ui_in[3] 2.82e-19
C3961 ringtest_0.x4.clknet_1_0__leaf_clk a_21852_8720# 0.083453f
C3962 a_24336_6544# ringtest_0.x4._21_ 0.001538f
C3963 ringtest_0.x4.counter[4] ua[1] 3.21e-19
C3964 ringtest_0.x4._11_ a_25421_6641# 0.004334f
C3965 a_23899_5334# VDPWR 0.205163f
C3966 ringtest_0.x4.net2 ringtest_0.x4._04_ 4.09e-22
C3967 ringtest_0.x4.clknet_0_clk ringtest_0.x4._17_ 0.029087f
C3968 ringtest_0.x4._15_ a_26173_4612# 0.006963f
C3969 ringtest_0.x4.net6 a_26721_4246# 7.2e-20
C3970 ua[4] VSS 0.139799f
C3971 ua[5] VSS 0.141076f
C3972 ua[6] VSS 0.141964f
C3973 ua[7] VSS 0.146962f
C3974 ena VSS 0.072324f
C3975 clk VSS 0.044814f
C3976 rst_n VSS 0.044814f
C3977 ui_in[7] VSS 0.044814f
C3978 uio_in[0] VSS 0.047326f
C3979 uio_in[1] VSS 0.048926f
C3980 uio_in[2] VSS 0.044814f
C3981 uio_in[3] VSS 0.044814f
C3982 uio_in[4] VSS 0.044814f
C3983 uio_in[5] VSS 0.044814f
C3984 uio_in[6] VSS 0.044814f
C3985 uio_in[7] VSS 0.075838f
C3986 ua[1] VSS 28.486887f
C3987 ui_in[5] VSS 18.12969f
C3988 ui_in[6] VSS 24.902954f
C3989 ua[2] VSS 34.46381f
C3990 ua[0] VSS 51.530293f
C3991 ui_in[4] VSS 32.182537f
C3992 ui_in[3] VSS 33.128075f
C3993 ua[3] VSS 54.146942f
C3994 ui_in[2] VSS 26.529623f
C3995 ui_in[1] VSS 10.570298f
C3996 ui_in[0] VSS 10.700917f
C3997 VDPWR VSS 0.629686p
C3998 m3_17046_7066# VSS 0.075151f $ **FLOATING
C3999 m3_17032_8096# VSS 0.073094f $ **FLOATING
C4000 m3_17036_9140# VSS 0.148749f $ **FLOATING
C4001 m3_13316_18955# VSS 0.066786f $ **FLOATING
C4002 m3_13302_19985# VSS 0.064102f $ **FLOATING
C4003 m2_15612_11606# VSS 0.070212f $ **FLOATING
C4004 m2_11882_23495# VSS 0.065655f $ **FLOATING
C4005 m2_18699_31802# VSS 0.065655f $ **FLOATING
C4006 ringtest_0.x4.counter[8] VSS 0.584764f
C4007 ringtest_0.x4.counter[9] VSS 0.886603f
C4008 ringtest_0.x4.counter[6] VSS 0.659065f
C4009 ringtest_0.x4.counter[5] VSS 0.636147f
C4010 ringtest_0.x4.counter[4] VSS 0.790245f
C4011 ringtest_0.x4.counter[2] VSS 0.6063f
C4012 ringtest_0.x4.counter[1] VSS 0.590824f
C4013 ringtest_0.x4.counter[0] VSS 0.938192f
C4014 a_27815_3867# VSS 0.269591f
C4015 a_27489_3702# VSS 0.256771f
C4016 a_26895_3867# VSS 0.29547f
C4017 a_25975_3867# VSS 0.269288f
C4018 a_25055_3867# VSS 0.277656f
C4019 a_24135_3867# VSS 0.327843f
C4020 a_23399_3867# VSS 0.269041f
C4021 a_22295_3867# VSS 0.275662f
C4022 a_21375_3867# VSS 0.316839f
C4023 a_21007_3867# VSS 0.251452f
C4024 a_27659_4246# VSS 4.27e-19
C4025 a_27303_4246# VSS 0.004592f
C4026 a_26721_4246# VSS 0.018483f
C4027 a_27491_4566# VSS 0.00589f
C4028 a_26913_4566# VSS 0.009736f
C4029 a_26817_4566# VSS 0.006433f
C4030 a_26375_4612# VSS 0.001527f
C4031 a_26269_4612# VSS 0.003564f
C4032 a_26173_4612# VSS 0.003656f
C4033 a_25547_4612# VSS 0.003203f
C4034 a_25441_4612# VSS 0.005457f
C4035 a_25345_4612# VSS 0.005167f
C4036 a_22486_4246# VSS 5.31e-19
C4037 a_23467_4584# VSS 0.004685f
C4038 a_22939_4584# VSS 0.007506f
C4039 a_22390_4566# VSS 0.179568f
C4040 a_27273_4220# VSS 0.362051f
C4041 a_26627_4246# VSS 0.339432f
C4042 a_25977_4220# VSS 0.256933f
C4043 a_25149_4220# VSS 0.289797f
C4044 a_23381_4584# VSS 0.253144f
C4045 a_22765_4478# VSS 0.281913f
C4046 a_22164_4362# VSS 0.205675f
C4047 a_22021_4220# VSS 0.201965f
C4048 a_27191_4790# VSS 0.004798f
C4049 ringtest_0.x4.net11 VSS 0.751523f
C4050 a_26766_4790# VSS 0.009249f
C4051 a_27149_5156# VSS 3.75e-19
C4052 a_25719_4790# VSS 0.004081f
C4053 a_26735_5156# VSS 0.002645f
C4054 a_26555_4790# VSS 0.063295f
C4055 a_27065_5156# VSS 0.268999f
C4056 a_27233_5058# VSS 0.379334f
C4057 a_26640_5156# VSS 0.227962f
C4058 a_26808_4902# VSS 0.257432f
C4059 a_26367_4790# VSS 0.333607f
C4060 ringtest_0.x4._09_ VSS 0.53373f
C4061 a_26201_4790# VSS 0.49567f
C4062 a_25294_4790# VSS 0.008648f
C4063 a_25677_5156# VSS 2.5e-19
C4064 a_24551_4790# VSS 7.4e-19
C4065 a_24479_4790# VSS 0.00237f
C4066 a_23963_4790# VSS 0.002571f
C4067 a_23891_4790# VSS 7.07e-19
C4068 a_25263_5156# VSS 7.5e-19
C4069 a_25083_4790# VSS 0.062171f
C4070 a_25593_5156# VSS 0.274347f
C4071 a_25761_5058# VSS 0.355731f
C4072 a_25168_5156# VSS 0.21761f
C4073 a_25336_4902# VSS 0.278138f
C4074 a_24895_4790# VSS 0.322796f
C4075 a_24729_4790# VSS 0.48451f
C4076 a_23467_4818# VSS 0.004685f
C4077 ringtest_0.x4._20_ VSS 0.296242f
C4078 a_22499_4790# VSS 0.004654f
C4079 ringtest_0.x4.net5 VSS 1.49846f
C4080 a_22074_4790# VSS 0.007478f
C4081 a_22457_5156# VSS 3.28e-19
C4082 a_21863_4790# VSS 0.067973f
C4083 a_24317_4942# VSS 0.231129f
C4084 a_23809_4790# VSS 0.250882f
C4085 a_23381_4818# VSS 0.250336f
C4086 a_22373_5156# VSS 0.28936f
C4087 a_22541_5058# VSS 0.404768f
C4088 a_21948_5156# VSS 0.210208f
C4089 a_22116_4902# VSS 0.255122f
C4090 a_21675_4790# VSS 0.414612f
C4091 ringtest_0.x4._03_ VSS 0.568022f
C4092 a_21509_4790# VSS 0.556893f
C4093 a_27149_5334# VSS 7.44e-19
C4094 a_26735_5334# VSS 0.002645f
C4095 ringtest_0.x4.net10 VSS 1.55164f
C4096 a_27191_5712# VSS 0.00478f
C4097 a_25309_5334# VSS 0.002002f
C4098 a_26766_5712# VSS 0.010952f
C4099 a_26555_5334# VSS 0.068133f
C4100 a_25351_5712# VSS 0.005844f
C4101 a_23899_5334# VSS 0.01364f
C4102 a_23151_5334# VSS 9.17e-19
C4103 a_22795_5334# VSS 0.025384f
C4104 a_22181_5334# VSS 4.07e-19
C4105 a_21767_5334# VSS 3.97e-19
C4106 a_24926_5712# VSS 0.006742f
C4107 a_24715_5334# VSS 0.060578f
C4108 a_23993_5654# VSS 0.006535f
C4109 a_23899_5654# VSS 0.007251f
C4110 a_22983_5654# VSS 0.006594f
C4111 a_22223_5712# VSS 0.004473f
C4112 a_21055_5334# VSS 2.59e-19
C4113 a_21798_5712# VSS 0.007899f
C4114 a_21587_5334# VSS 0.080556f
C4115 a_27065_5334# VSS 0.271f
C4116 a_27233_5308# VSS 0.369643f
C4117 a_26640_5334# VSS 0.236761f
C4118 a_26808_5308# VSS 0.26375f
C4119 a_26367_5340# VSS 0.339249f
C4120 a_26201_5340# VSS 0.527463f
C4121 a_25225_5334# VSS 0.287672f
C4122 a_25393_5308# VSS 0.390363f
C4123 a_24800_5334# VSS 0.199335f
C4124 a_24968_5308# VSS 0.244436f
C4125 a_24527_5340# VSS 0.30834f
C4126 a_24361_5340# VSS 0.476837f
C4127 a_23770_5308# VSS 0.3495f
C4128 a_22765_5308# VSS 0.426063f
C4129 a_22097_5334# VSS 0.278482f
C4130 a_22265_5308# VSS 0.362892f
C4131 a_21672_5334# VSS 0.210395f
C4132 a_21840_5308# VSS 0.26005f
C4133 a_21399_5340# VSS 0.408899f
C4134 ringtest_0.x4._02_ VSS 0.380851f
C4135 a_21233_5340# VSS 0.547022f
C4136 ringtest_0.x4._14_ VSS 1.22018f
C4137 a_24986_5878# VSS 0.00398f
C4138 a_24545_5878# VSS 0.153731f
C4139 ringtest_0.x4._07_ VSS 0.455737f
C4140 a_23837_5878# VSS 0.202457f
C4141 a_22775_5878# VSS 0.00681f
C4142 ringtest_0.x4._16_ VSS 2.056043f
C4143 ringtest_0.x4._22_ VSS 1.53821f
C4144 a_24627_6200# VSS 4.54e-20
C4145 a_24763_6143# VSS 0.188859f
C4146 ringtest_0.x4.net9 VSS 1.94148f
C4147 ringtest_0.x4._06_ VSS 0.345483f
C4148 ringtest_0.x4._21_ VSS 0.479535f
C4149 a_23932_6128# VSS 5.66e-19
C4150 a_22350_5878# VSS 0.006923f
C4151 a_22733_6244# VSS 0.002478f
C4152 a_22319_6244# VSS 2.95e-19
C4153 a_22139_5878# VSS 0.062642f
C4154 a_25364_5878# VSS 2.06251f
C4155 a_24699_6200# VSS 0.164646f
C4156 a_24004_6128# VSS 0.20664f
C4157 a_24070_5852# VSS 0.228407f
C4158 ringtest_0.x4.net8 VSS 1.74106f
C4159 a_22649_6244# VSS 0.330474f
C4160 a_22817_6146# VSS 0.422968f
C4161 a_22224_6244# VSS 0.217913f
C4162 a_22392_5990# VSS 0.26464f
C4163 a_21951_5878# VSS 0.380288f
C4164 ringtest_0.x4._04_ VSS 0.637317f
C4165 a_21785_5878# VSS 0.555262f
C4166 a_21591_6128# VSS 0.005123f
C4167 ringtest_0.x4._13_ VSS 1.12775f
C4168 ringtest_0.x4.net4 VSS 1.27471f
C4169 ringtest_0.x4._08_ VSS 0.709311f
C4170 a_26839_6788# VSS 0.008414f
C4171 a_26201_6788# VSS 0.003851f
C4172 a_26095_6788# VSS 0.003674f
C4173 a_26007_6788# VSS 0.001688f
C4174 a_24287_6422# VSS 7.93e-19
C4175 a_24883_6800# VSS 0.060771f
C4176 a_24685_6788# VSS 0.006624f
C4177 a_24264_6788# VSS 0.005504f
C4178 a_23619_6788# VSS 0.005146f
C4179 ringtest_0.x4._25_ VSS 0.365803f
C4180 a_27169_6641# VSS 0.272731f
C4181 a_26749_6422# VSS 0.26247f
C4182 ringtest_0.x4._24_ VSS 0.681525f
C4183 a_26569_6422# VSS 0.271803f
C4184 ringtest_0.x4._23_ VSS 0.94177f
C4185 a_25925_6788# VSS 0.263758f
C4186 ringtest_0.x4._15_ VSS 3.49608f
C4187 ringtest_0.x4.net7 VSS 2.68462f
C4188 ringtest_0.x4.net6 VSS 3.121006f
C4189 ringtest_0.x4._19_ VSS 0.323337f
C4190 a_25421_6641# VSS 0.252712f
C4191 ringtest_0.x4.clknet_1_1__leaf_clk VSS 3.376462f
C4192 ringtest_0.x4._05_ VSS 0.317001f
C4193 a_24465_6800# VSS 0.240387f
C4194 a_24536_6699# VSS 0.197853f
C4195 a_24336_6544# VSS 0.302006f
C4196 a_24329_6640# VSS 0.464687f
C4197 a_24045_6654# VSS 0.281097f
C4198 a_23949_6654# VSS 0.378482f
C4199 a_23529_6422# VSS 0.233246f
C4200 ringtest_0.x4._18_ VSS 0.453422f
C4201 a_23349_6422# VSS 0.254342f
C4202 ringtest_0.x4._17_ VSS 0.620105f
C4203 ringtest_0.counter7 VSS 17.348873f
C4204 a_23879_6940# VSS 2.26754f
C4205 ringtest_0.x4.clknet_0_clk VSS 4.126871f
C4206 a_21395_6940# VSS 2.26943f
C4207 a_21939_8054# VSS 0.002324f
C4208 a_21867_8054# VSS 0.001217f
C4209 a_22695_8304# VSS 0.005104f
C4210 ringtest_0.counter3 VSS 14.330247f
C4211 ringtest_0.x4._11_ VSS 5.567417f
C4212 a_22245_8054# VSS 0.294759f
C4213 ringtest_0.x4._10_ VSS 0.338654f
C4214 a_21785_8054# VSS 0.248451f
C4215 a_21803_8598# VSS 2.93e-19
C4216 a_22399_8976# VSS 0.062869f
C4217 a_22201_8964# VSS 0.006624f
C4218 a_21049_8598# VSS 0.014348f
C4219 a_21780_8964# VSS 0.004174f
C4220 ringtest_0.x4._12_ VSS 1.24358f
C4221 a_21132_8918# VSS 0.00439f
C4222 ringtest_0.x4._01_ VSS 0.392316f
C4223 a_21981_8976# VSS 0.237918f
C4224 a_22052_8875# VSS 0.194948f
C4225 a_21852_8720# VSS 0.308329f
C4226 a_21845_8816# VSS 0.548694f
C4227 a_21561_8830# VSS 0.278058f
C4228 a_21465_8830# VSS 0.389128f
C4229 ringtest_0.x4.net3 VSS 2.243398f
C4230 a_22201_9142# VSS 0.007478f
C4231 a_21780_9142# VSS 0.004654f
C4232 ringtest_0.x4.clknet_1_0__leaf_clk VSS 3.939619f
C4233 a_22399_9142# VSS 0.069066f
C4234 a_21803_9508# VSS 3.83e-19
C4235 a_21981_9142# VSS 0.264294f
C4236 a_22052_9116# VSS 0.210441f
C4237 a_21845_9116# VSS 0.577647f
C4238 a_21852_9416# VSS 0.335522f
C4239 a_21561_9116# VSS 0.285682f
C4240 a_21465_9294# VSS 0.411301f
C4241 a_21675_9686# VSS 0.008029f
C4242 a_21507_9686# VSS 0.006974f
C4243 ringtest_0.x4._00_ VSS 0.734028f
C4244 a_21675_10006# VSS 0.006039f
C4245 a_21425_9686# VSS 0.39001f
C4246 ringtest_0.x4.net2 VSS 3.435971f
C4247 ringtest_0.x4.net1 VSS 1.77359f
C4248 a_22111_10993# VSS 0.292622f
C4249 ringtest_0.x3.x2.GP3 VSS 1.64575f
C4250 ringtest_0.x3.x2.GP2 VSS 5.54164f
C4251 ringtest_0.x3.x2.GP1 VSS 4.63625f
C4252 a_17405_12123# VSS 0.006782f
C4253 ringtest_0.x3.x2.GN4 VSS 3.79271f
C4254 a_16707_12151# VSS 0.007327f
C4255 ringtest_0.x3.x2.GN3 VSS 3.64172f
C4256 a_16155_12151# VSS 0.004704f
C4257 ringtest_0.x3.x2.GN2 VSS 3.91967f
C4258 a_15749_12123# VSS 0.006793f
C4259 ringtest_0.x3.x2.GN1 VSS 4.84443f
C4260 a_17231_12017# VSS 0.3167f
C4261 a_16755_12091# VSS 0.251626f
C4262 a_16579_11759# VSS 0.236732f
C4263 a_16203_12091# VSS 0.236633f
C4264 a_16027_11759# VSS 0.222621f
C4265 a_15575_12017# VSS 0.270062f
C4266 ringtest_0.x3.nselect2 VSS 0.455447f
C4267 ringtest_0.x3.x1.nSEL1 VSS 0.740163f
C4268 ringtest_0.x3.x1.nSEL0 VSS 0.685116f
C4269 ringtest_0.x1.sky130_fd_sc_hd__inv_2_11.A VSS 0.505562f
C4270 ringtest_0.x1.sky130_fd_sc_hd__inv_2_12.A VSS 0.498424f
C4271 ringtest_0.x1.sky130_fd_sc_hd__inv_2_13.A VSS 0.498285f
C4272 ringtest_0.x1.sky130_fd_sc_hd__inv_2_14.A VSS 0.499488f
C4273 ringtest_0.x1.sky130_fd_sc_hd__inv_2_15.A VSS 0.500758f
C4274 ringtest_0.x1.sky130_fd_sc_hd__inv_2_16.A VSS 0.50136f
C4275 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.A VSS 0.501617f
C4276 ringtest_0.x1.sky130_fd_sc_hd__inv_2_17.Y VSS 0.52312f
C4277 ringtest_0.drv_out VSS 29.21638f
C4278 a_17377_14114# VSS 0.332619f
C4279 ringtest_0.ring_out VSS 16.284393f
C4280 ringtest_0.x1.sky130_fd_sc_hd__nand2_2_0.B VSS 0.632983f
C4281 ringtest_0.x1.sky130_fd_sc_hd__inv_2_9.A VSS 0.508122f
C4282 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.Y VSS 0.498331f
C4283 ringtest_0.x1.sky130_fd_sc_hd__inv_2_7.A VSS 0.498331f
C4284 ringtest_0.x1.sky130_fd_sc_hd__inv_2_6.A VSS 0.498339f
C4285 ringtest_0.x1.sky130_fd_sc_hd__inv_2_5.A VSS 0.498632f
C4286 ringtest_0.x1.sky130_fd_sc_hd__inv_2_4.A VSS 0.498682f
C4287 ringtest_0.x1.sky130_fd_sc_hd__inv_2_3.A VSS 0.498707f
C4288 ringtest_0.x1.sky130_fd_sc_hd__inv_2_2.A VSS 0.507755f
C4289 ringtest_0.x1.sky130_fd_sc_hd__inv_2_8.Y VSS 0.971227f
C4290 muxtest_0.x2.x2.GP3 VSS 1.68554f
C4291 muxtest_0.x2.x2.GP2 VSS 5.5641f
C4292 muxtest_0.x2.x2.GP1 VSS 4.625069f
C4293 muxtest_0.R1R2 VSS 6.645506f
C4294 a_13675_24012# VSS 0.006439f
C4295 muxtest_0.x2.x2.GN4 VSS 3.796f
C4296 a_12977_24040# VSS 0.006801f
C4297 muxtest_0.x2.x2.GN3 VSS 3.65554f
C4298 a_12425_24040# VSS 0.004461f
C4299 muxtest_0.x2.x2.GN2 VSS 3.88834f
C4300 a_12019_24012# VSS 0.006505f
C4301 muxtest_0.x2.x2.GN1 VSS 4.79625f
C4302 a_13501_23906# VSS 0.306555f
C4303 a_13025_23980# VSS 0.249538f
C4304 a_12849_23648# VSS 0.232764f
C4305 a_12473_23980# VSS 0.23458f
C4306 a_12297_23648# VSS 0.220868f
C4307 a_11845_23906# VSS 0.267622f
C4308 muxtest_0.x2.nselect2 VSS 0.451665f
C4309 muxtest_0.x2.x1.nSEL1 VSS 0.686441f
C4310 muxtest_0.x2.x1.nSEL0 VSS 0.647345f
C4311 muxtest_0.R2R3 VSS 7.982832f
C4312 muxtest_0.R3R4 VSS 15.859409f
C4313 muxtest_0.R4R5 VSS 7.656276f
C4314 muxtest_0.R5R6 VSS 7.957228f
C4315 muxtest_0.R6R7 VSS 7.795067f
C4316 muxtest_0.R7R8 VSS 29.82938f
C4317 muxtest_0.x1.x5.A VSS 13.867701f
C4318 muxtest_0.x1.x4.A VSS 16.1317f
C4319 muxtest_0.x1.x3.GP3 VSS 3.18231f
C4320 muxtest_0.x1.x3.GP2 VSS 10.304811f
C4321 muxtest_0.x1.x3.GP1 VSS 10.781407f
C4322 a_20492_32319# VSS 0.006616f
C4323 muxtest_0.x1.x3.GN4 VSS 7.04004f
C4324 a_19794_32347# VSS 0.006984f
C4325 muxtest_0.x1.x3.GN3 VSS 6.77674f
C4326 a_19242_32347# VSS 0.004523f
C4327 muxtest_0.x1.x3.GN2 VSS 7.175951f
C4328 a_18836_32319# VSS 0.006515f
C4329 muxtest_0.x1.x3.GN1 VSS 8.91731f
C4330 a_20318_32213# VSS 0.311491f
C4331 a_19842_32287# VSS 0.24978f
C4332 a_19666_31955# VSS 0.233122f
C4333 a_19290_32287# VSS 0.234813f
C4334 a_19114_31955# VSS 0.221018f
C4335 a_18662_32213# VSS 0.267639f
C4336 muxtest_0.x1.x5.GN VSS 5.73587f
C4337 muxtest_0.x1.x1.nSEL1 VSS 0.683011f
C4338 muxtest_0.x1.x1.nSEL0 VSS 0.650421f
C4339 ui_in[5].t1 VSS 0.002404f
C4340 ui_in[5].t0 VSS 0.003855f
C4341 ui_in[5].n0 VSS 0.007767f
C4342 ui_in[5].n1 VSS 0.003276f
C4343 ui_in[5].n2 VSS 0.31852f
C4344 ui_in[5].n3 VSS 3.27959f
C4345 ui_in[6].t0 VSS 0.002431f
C4346 ui_in[6].t2 VSS 0.001432f
C4347 ui_in[6].n0 VSS 0.003276f
C4348 ui_in[6].t1 VSS 0.002431f
C4349 ui_in[6].t3 VSS 0.001432f
C4350 ui_in[6].n1 VSS 0.003276f
C4351 ui_in[6].n2 VSS 0.001614f
C4352 ui_in[6].n3 VSS 0.214753f
C4353 muxtest_0.R2R3.t4 VSS 0.626391f
C4354 muxtest_0.R2R3.t5 VSS 0.443113f
C4355 muxtest_0.R2R3.n0 VSS 3.43546f
C4356 muxtest_0.R2R3.t1 VSS 0.347912f
C4357 muxtest_0.R2R3.t2 VSS 0.638083f
C4358 muxtest_0.R2R3.n1 VSS 3.5698f
C4359 muxtest_0.R2R3.n2 VSS 0.568983f
C4360 muxtest_0.R2R3.n3 VSS 0.116677f
C4361 muxtest_0.R2R3.t0 VSS 0.210663f
C4362 muxtest_0.R2R3.t3 VSS 0.170342f
C4363 muxtest_0.R2R3.n4 VSS 3.38019f
C4364 muxtest_0.R4R5.t1 VSS 0.627578f
C4365 muxtest_0.R4R5.t2 VSS 0.443953f
C4366 muxtest_0.R4R5.n0 VSS 3.44197f
C4367 muxtest_0.R4R5.t4 VSS 0.348571f
C4368 muxtest_0.R4R5.t5 VSS 0.639293f
C4369 muxtest_0.R4R5.n1 VSS 3.57657f
C4370 muxtest_0.R4R5.n2 VSS 0.570061f
C4371 muxtest_0.R4R5.n3 VSS 0.119407f
C4372 muxtest_0.R4R5.t0 VSS 0.212944f
C4373 muxtest_0.R4R5.t3 VSS 0.170665f
C4374 muxtest_0.R4R5.n4 VSS 3.47489f
C4375 muxtest_0.x2.x2.x4.GP VSS 2.57727f
C4376 muxtest_0.x2.x1.gpo3 VSS 1.20603f
C4377 muxtest_0.x2.x2.GP4.t3 VSS 0.012374f
C4378 muxtest_0.x2.x2.GP4.t2 VSS 0.012374f
C4379 muxtest_0.x2.x2.GP4.n0 VSS 0.027184f
C4380 muxtest_0.x2.x1.x14.Y VSS 0.076955f
C4381 muxtest_0.x2.x2.GP4.n1 VSS 0.01052f
C4382 muxtest_0.x2.x2.GP4.t5 VSS 0.626223f
C4383 muxtest_0.x2.x2.GP4.t4 VSS 0.643686f
C4384 muxtest_0.x2.x2.GP4.n2 VSS 2.28835f
C4385 muxtest_0.x2.x2.GP4.n3 VSS 0.048401f
C4386 muxtest_0.x2.x2.GP4.t1 VSS 0.019037f
C4387 muxtest_0.x2.x2.GP4.t0 VSS 0.019037f
C4388 muxtest_0.x2.x2.GP4.n4 VSS 0.043773f
C4389 muxtest_0.x2.x2.GP4.n5 VSS 0.088779f
C4390 ringtest_0.x3.x2.GP2.t3 VSS 0.016198f
C4391 ringtest_0.x3.x2.GP2.t2 VSS 0.016198f
C4392 ringtest_0.x3.x2.GP2.n0 VSS 0.035585f
C4393 ringtest_0.x3.x2.GP2.n1 VSS 0.023f
C4394 ringtest_0.x3.x2.GP2.t5 VSS 0.819754f
C4395 ringtest_0.x3.x2.GP2.t4 VSS 0.842614f
C4396 ringtest_0.x3.x2.GP2.n2 VSS 2.98946f
C4397 ringtest_0.x3.x2.GP2.t1 VSS 0.02492f
C4398 ringtest_0.x3.x2.GP2.t0 VSS 0.02492f
C4399 ringtest_0.x3.x2.GP2.n3 VSS 0.051391f
C4400 ringtest_0.x3.x2.GP2.n4 VSS 0.120168f
C4401 ringtest_0.x3.x2.GP2.n5 VSS 0.027176f
C4402 ringtest_0.ring_out.t13 VSS 0.143976f
C4403 ringtest_0.ring_out.t12 VSS 0.066482f
C4404 ringtest_0.ring_out.n0 VSS 1.43742f
C4405 ringtest_0.ring_out.t1 VSS 0.011895f
C4406 ringtest_0.ring_out.t0 VSS 0.011895f
C4407 ringtest_0.ring_out.n1 VSS 0.036116f
C4408 ringtest_0.ring_out.t6 VSS 0.011895f
C4409 ringtest_0.ring_out.t7 VSS 0.011895f
C4410 ringtest_0.ring_out.n2 VSS 0.026441f
C4411 ringtest_0.ring_out.n3 VSS 0.119642f
C4412 ringtest_0.ring_out.t8 VSS 0.007732f
C4413 ringtest_0.ring_out.t9 VSS 0.007732f
C4414 ringtest_0.ring_out.n4 VSS 0.017154f
C4415 ringtest_0.ring_out.n5 VSS 0.032249f
C4416 ringtest_0.ring_out.n6 VSS 0.009203f
C4417 ringtest_0.ring_out.t14 VSS 0.010903f
C4418 ringtest_0.ring_out.t10 VSS 0.018503f
C4419 ringtest_0.ring_out.t15 VSS 0.010903f
C4420 ringtest_0.ring_out.t11 VSS 0.018503f
C4421 ringtest_0.ring_out.n7 VSS 0.031045f
C4422 ringtest_0.ring_out.n8 VSS 0.04596f
C4423 ringtest_0.ring_out.n9 VSS 0.181049f
C4424 ringtest_0.ring_out.n10 VSS 0.421446f
C4425 ringtest_0.ring_out.t4 VSS 0.673389f
C4426 ringtest_0.ring_out.t5 VSS 0.47636f
C4427 ringtest_0.ring_out.n11 VSS 3.69323f
C4428 ringtest_0.ring_out.t2 VSS 0.374016f
C4429 ringtest_0.ring_out.t3 VSS 0.685959f
C4430 ringtest_0.ring_out.n12 VSS 3.83764f
C4431 ringtest_0.ring_out.n13 VSS 0.611674f
C4432 ringtest_0.x3.x2.GP1.t3 VSS 0.012908f
C4433 ringtest_0.x3.x2.GP1.t2 VSS 0.012908f
C4434 ringtest_0.x3.x2.GP1.n0 VSS 0.028358f
C4435 ringtest_0.x3.x2.GP1.n1 VSS 0.018329f
C4436 ringtest_0.x3.x2.GP1.t4 VSS 0.653268f
C4437 ringtest_0.x3.x2.GP1.t5 VSS 0.671486f
C4438 ringtest_0.x3.x2.GP1.n2 VSS 2.37213f
C4439 ringtest_0.x3.x2.GP1.t1 VSS 0.019859f
C4440 ringtest_0.x3.x2.GP1.t0 VSS 0.019859f
C4441 ringtest_0.x3.x2.GP1.n3 VSS 0.04092f
C4442 ringtest_0.x3.x2.GP1.n4 VSS 0.100085f
C4443 ringtest_0.x3.x2.GP1.n5 VSS 0.021877f
C4444 ui_in[3].t3 VSS 0.007328f
C4445 ui_in[3].t12 VSS 0.004318f
C4446 ui_in[3].t18 VSS 0.007328f
C4447 ui_in[3].t2 VSS 0.004318f
C4448 ui_in[3].n0 VSS 0.012295f
C4449 ui_in[3].n1 VSS 0.018171f
C4450 ui_in[3].n2 VSS 0.00571f
C4451 ui_in[3].t6 VSS 0.003609f
C4452 ui_in[3].t10 VSS 0.005242f
C4453 ui_in[3].n3 VSS 0.012487f
C4454 ui_in[3].n4 VSS 0.006935f
C4455 ui_in[3].t9 VSS 0.004274f
C4456 ui_in[3].t19 VSS 0.006294f
C4457 ui_in[3].n5 VSS 0.01487f
C4458 ui_in[3].n6 VSS 0.003088f
C4459 ui_in[3].n7 VSS 0.001204f
C4460 ui_in[3].n8 VSS 0.109977f
C4461 ui_in[3].t17 VSS 0.007151f
C4462 ui_in[3].t15 VSS 0.003391f
C4463 ui_in[3].n9 VSS 0.025678f
C4464 ui_in[3].n10 VSS 0.004976f
C4465 ui_in[3].n11 VSS 0.126174f
C4466 ui_in[3].n12 VSS 0.081988f
C4467 ui_in[3].t8 VSS 0.007328f
C4468 ui_in[3].t16 VSS 0.004318f
C4469 ui_in[3].t5 VSS 0.007328f
C4470 ui_in[3].t13 VSS 0.004318f
C4471 ui_in[3].n13 VSS 0.012295f
C4472 ui_in[3].n14 VSS 0.018171f
C4473 ui_in[3].n15 VSS 0.00571f
C4474 ui_in[3].t7 VSS 0.003609f
C4475 ui_in[3].t11 VSS 0.005242f
C4476 ui_in[3].n16 VSS 0.012487f
C4477 ui_in[3].n17 VSS 0.006935f
C4478 ui_in[3].t14 VSS 0.004274f
C4479 ui_in[3].t0 VSS 0.006294f
C4480 ui_in[3].n18 VSS 0.01487f
C4481 ui_in[3].n19 VSS 0.003088f
C4482 ui_in[3].n20 VSS 0.001204f
C4483 ui_in[3].n21 VSS 0.109977f
C4484 ui_in[3].t4 VSS 0.007151f
C4485 ui_in[3].t1 VSS 0.003391f
C4486 ui_in[3].n22 VSS 0.025678f
C4487 ui_in[3].n23 VSS 0.004976f
C4488 ui_in[3].n24 VSS 0.126174f
C4489 ui_in[3].n25 VSS 0.081988f
C4490 ui_in[3].n26 VSS 9.89241f
C4491 muxtest_0.R7R8.t8 VSS 0.570638f
C4492 muxtest_0.R7R8.t7 VSS 0.403673f
C4493 muxtest_0.R7R8.n0 VSS 3.12968f
C4494 muxtest_0.R7R8.t5 VSS 0.316945f
C4495 muxtest_0.R7R8.t6 VSS 0.58129f
C4496 muxtest_0.R7R8.n1 VSS 3.25206f
C4497 muxtest_0.R7R8.n2 VSS 0.51834f
C4498 muxtest_0.R7R8.n3 VSS 0.107649f
C4499 muxtest_0.R7R8.t9 VSS 0.157299f
C4500 muxtest_0.R7R8.t2 VSS 0.858788f
C4501 muxtest_0.R7R8.n4 VSS 1.55412f
C4502 muxtest_0.R7R8.t0 VSS 0.570638f
C4503 muxtest_0.R7R8.t1 VSS 0.403673f
C4504 muxtest_0.R7R8.n5 VSS 3.12968f
C4505 muxtest_0.R7R8.t3 VSS 0.316945f
C4506 muxtest_0.R7R8.t4 VSS 0.58129f
C4507 muxtest_0.R7R8.n6 VSS 3.25206f
C4508 muxtest_0.R7R8.n7 VSS 0.51834f
C4509 muxtest_0.R7R8.n8 VSS 0.108573f
C4510 muxtest_0.R7R8.n9 VSS 9.50513f
C4511 ua[0].t0 VSS 0.319126f
C4512 ua[0].t1 VSS 0.225752f
C4513 ua[0].n0 VSS 1.75026f
C4514 ua[0].t8 VSS 0.17725f
C4515 ua[0].t7 VSS 0.325083f
C4516 ua[0].n1 VSS 1.8187f
C4517 ua[0].n2 VSS 0.289879f
C4518 ua[0].n3 VSS 0.060719f
C4519 ua[0].t2 VSS 0.086784f
C4520 ua[0].n4 VSS 1.50131f
C4521 ua[0].n5 VSS 11.5833f
C4522 ua[0].t6 VSS 0.319126f
C4523 ua[0].t5 VSS 0.225752f
C4524 ua[0].n6 VSS 1.75026f
C4525 ua[0].t4 VSS 0.17725f
C4526 ua[0].t3 VSS 0.325083f
C4527 ua[0].n7 VSS 1.8187f
C4528 ua[0].n8 VSS 0.289879f
C4529 ua[0].n9 VSS 0.059443f
C4530 muxtest_0.R6R7.t3 VSS 0.693928f
C4531 muxtest_0.R6R7.t2 VSS 0.490889f
C4532 muxtest_0.R6R7.n0 VSS 3.80587f
C4533 muxtest_0.R6R7.t0 VSS 0.385423f
C4534 muxtest_0.R6R7.t1 VSS 0.706881f
C4535 muxtest_0.R6R7.n1 VSS 3.95469f
C4536 muxtest_0.R6R7.n2 VSS 0.63033f
C4537 muxtest_0.R6R7.n3 VSS 0.129257f
C4538 muxtest_0.R6R7.t4 VSS 0.920517f
C4539 muxtest_0.R6R7.t5 VSS 0.188708f
C4540 muxtest_0.R6R7.n4 VSS 2.80583f
C4541 muxtest_0.R6R7.n5 VSS 1.24461f
C4542 muxtest_0.x2.x2.GP2.t2 VSS 0.016198f
C4543 muxtest_0.x2.x2.GP2.t3 VSS 0.016198f
C4544 muxtest_0.x2.x2.GP2.n0 VSS 0.035585f
C4545 muxtest_0.x2.x2.GP2.n1 VSS 0.023f
C4546 muxtest_0.x2.x2.GP2.t5 VSS 0.819754f
C4547 muxtest_0.x2.x2.GP2.t4 VSS 0.842614f
C4548 muxtest_0.x2.x2.GP2.n2 VSS 2.98946f
C4549 muxtest_0.x2.x2.GP2.t1 VSS 0.02492f
C4550 muxtest_0.x2.x2.GP2.t0 VSS 0.02492f
C4551 muxtest_0.x2.x2.GP2.n3 VSS 0.051391f
C4552 muxtest_0.x2.x2.GP2.n4 VSS 0.120168f
C4553 muxtest_0.x2.x2.GP2.n5 VSS 0.027176f
C4554 ringtest_0.x4._16_.t1 VSS 0.046376f
C4555 ringtest_0.x4._16_.n0 VSS 0.026397f
C4556 ringtest_0.x4._16_.t7 VSS 0.021164f
C4557 ringtest_0.x4._16_.t2 VSS 0.017507f
C4558 ringtest_0.x4._16_.n1 VSS 0.047954f
C4559 ringtest_0.x4._16_.n2 VSS 0.154756f
C4560 ringtest_0.x4._16_.t9 VSS 0.020065f
C4561 ringtest_0.x4._16_.t3 VSS 0.031953f
C4562 ringtest_0.x4._16_.n3 VSS 0.045672f
C4563 ringtest_0.x4._16_.n4 VSS 0.0375f
C4564 ringtest_0.x4._16_.t4 VSS 0.020065f
C4565 ringtest_0.x4._16_.t8 VSS 0.031953f
C4566 ringtest_0.x4._16_.n5 VSS 0.058943f
C4567 ringtest_0.x4._16_.n6 VSS 0.063595f
C4568 ringtest_0.x4._16_.n7 VSS 0.426096f
C4569 ringtest_0.x4._16_.t5 VSS 0.012893f
C4570 ringtest_0.x4._16_.t6 VSS 0.013824f
C4571 ringtest_0.x4._16_.n8 VSS 0.03796f
C4572 ringtest_0.x4._16_.n9 VSS 0.022428f
C4573 ringtest_0.x4._16_.n10 VSS 0.327394f
C4574 ringtest_0.x4._16_.n11 VSS 0.020414f
C4575 ringtest_0.x4._16_.t0 VSS 0.119992f
C4576 ringtest_0.x4._16_.n12 VSS 0.021583f
C4577 ringtest_0.x4._16_.n13 VSS 0.021194f
C4578 muxtest_0.R5R6.t1 VSS 0.695132f
C4579 muxtest_0.R5R6.t2 VSS 0.491742f
C4580 muxtest_0.R5R6.n0 VSS 3.81248f
C4581 muxtest_0.R5R6.t5 VSS 0.386092f
C4582 muxtest_0.R5R6.t4 VSS 0.708108f
C4583 muxtest_0.R5R6.n1 VSS 3.96156f
C4584 muxtest_0.R5R6.n2 VSS 0.631424f
C4585 muxtest_0.R5R6.n3 VSS 0.129973f
C4586 muxtest_0.R5R6.t3 VSS 0.191095f
C4587 muxtest_0.R5R6.t0 VSS 1.13104f
C4588 muxtest_0.R5R6.n4 VSS 2.8297f
C4589 muxtest_0.x1.x3.GP2.t2 VSS 0.018287f
C4590 muxtest_0.x1.x3.GP2.t3 VSS 0.018287f
C4591 muxtest_0.x1.x3.GP2.n0 VSS 0.040174f
C4592 muxtest_0.x1.x3.GP2.n1 VSS 0.025967f
C4593 muxtest_0.x1.x3.GP2.t6 VSS 0.925483f
C4594 muxtest_0.x1.x3.GP2.t7 VSS 0.951291f
C4595 muxtest_0.x1.x3.GP2.n2 VSS 3.37503f
C4596 muxtest_0.x1.x3.GP2.t5 VSS 0.925483f
C4597 muxtest_0.x1.x3.GP2.t4 VSS 0.951291f
C4598 muxtest_0.x1.x3.GP2.n3 VSS 3.37503f
C4599 muxtest_0.x1.x3.GP2.n4 VSS 1.97357f
C4600 muxtest_0.x1.x3.GP2.t0 VSS 0.028134f
C4601 muxtest_0.x1.x3.GP2.t1 VSS 0.028134f
C4602 muxtest_0.x1.x3.GP2.n5 VSS 0.058019f
C4603 muxtest_0.x1.x3.GP2.n6 VSS 0.132927f
C4604 muxtest_0.x1.x3.GP2.n7 VSS 0.030681f
C4605 ringtest_0.counter3.t0 VSS 0.033829f
C4606 ringtest_0.counter3.n0 VSS 0.005886f
C4607 ringtest_0.counter3.t1 VSS 0.023398f
C4608 ringtest_0.counter3.n1 VSS 0.028682f
C4609 ringtest_0.counter3.n2 VSS 0.036901f
C4610 ringtest_0.counter3.n3 VSS 0.371589f
C4611 ringtest_0.counter3.t3 VSS 0.740343f
C4612 ringtest_0.counter3.t2 VSS 0.523724f
C4613 ringtest_0.counter3.n4 VSS 4.06044f
C4614 ringtest_0.counter3.t4 VSS 0.410954f
C4615 ringtest_0.counter3.t5 VSS 0.761665f
C4616 ringtest_0.counter3.n5 VSS 4.29752f
C4617 ringtest_0.counter3.n6 VSS 0.672491f
C4618 ringtest_0.x4.clknet_1_0__leaf_clk.t38 VSS 0.022262f
C4619 ringtest_0.x4.clknet_1_0__leaf_clk.t41 VSS 0.014894f
C4620 ringtest_0.x4.clknet_1_0__leaf_clk.n0 VSS 0.04068f
C4621 ringtest_0.x4.clknet_1_0__leaf_clk.n1 VSS 0.107083f
C4622 ringtest_0.x4.clknet_1_0__leaf_clk.t37 VSS 0.014894f
C4623 ringtest_0.x4.clknet_1_0__leaf_clk.t32 VSS 0.022262f
C4624 ringtest_0.x4.clknet_1_0__leaf_clk.n2 VSS 0.041145f
C4625 ringtest_0.x4.clknet_1_0__leaf_clk.n3 VSS 0.437523f
C4626 ringtest_0.x4.clknet_1_0__leaf_clk.t14 VSS 0.014222f
C4627 ringtest_0.x4.clknet_1_0__leaf_clk.t0 VSS 0.014222f
C4628 ringtest_0.x4.clknet_1_0__leaf_clk.n4 VSS 0.029978f
C4629 ringtest_0.x4.clknet_1_0__leaf_clk.t11 VSS 0.014222f
C4630 ringtest_0.x4.clknet_1_0__leaf_clk.t13 VSS 0.014222f
C4631 ringtest_0.x4.clknet_1_0__leaf_clk.n5 VSS 0.029589f
C4632 ringtest_0.x4.clknet_1_0__leaf_clk.t24 VSS 0.005973f
C4633 ringtest_0.x4.clknet_1_0__leaf_clk.t27 VSS 0.005973f
C4634 ringtest_0.x4.clknet_1_0__leaf_clk.n6 VSS 0.021211f
C4635 ringtest_0.x4.clknet_1_0__leaf_clk.t29 VSS 0.005973f
C4636 ringtest_0.x4.clknet_1_0__leaf_clk.t31 VSS 0.005973f
C4637 ringtest_0.x4.clknet_1_0__leaf_clk.n7 VSS 0.013636f
C4638 ringtest_0.x4.clknet_1_0__leaf_clk.n8 VSS 0.086164f
C4639 ringtest_0.x4.clknet_1_0__leaf_clk.t26 VSS 0.005973f
C4640 ringtest_0.x4.clknet_1_0__leaf_clk.t28 VSS 0.005973f
C4641 ringtest_0.x4.clknet_1_0__leaf_clk.n9 VSS 0.013636f
C4642 ringtest_0.x4.clknet_1_0__leaf_clk.n10 VSS 0.051791f
C4643 ringtest_0.x4.clknet_1_0__leaf_clk.t30 VSS 0.005973f
C4644 ringtest_0.x4.clknet_1_0__leaf_clk.t25 VSS 0.005973f
C4645 ringtest_0.x4.clknet_1_0__leaf_clk.n11 VSS 0.013644f
C4646 ringtest_0.x4.clknet_1_0__leaf_clk.n12 VSS 0.053424f
C4647 ringtest_0.x4.clknet_1_0__leaf_clk.t17 VSS 0.005973f
C4648 ringtest_0.x4.clknet_1_0__leaf_clk.t20 VSS 0.005973f
C4649 ringtest_0.x4.clknet_1_0__leaf_clk.n13 VSS 0.013636f
C4650 ringtest_0.x4.clknet_1_0__leaf_clk.n14 VSS 0.051791f
C4651 ringtest_0.x4.clknet_1_0__leaf_clk.t22 VSS 0.005973f
C4652 ringtest_0.x4.clknet_1_0__leaf_clk.t23 VSS 0.005973f
C4653 ringtest_0.x4.clknet_1_0__leaf_clk.n15 VSS 0.013636f
C4654 ringtest_0.x4.clknet_1_0__leaf_clk.n16 VSS 0.05205f
C4655 ringtest_0.x4.clknet_1_0__leaf_clk.t19 VSS 0.005973f
C4656 ringtest_0.x4.clknet_1_0__leaf_clk.t21 VSS 0.005973f
C4657 ringtest_0.x4.clknet_1_0__leaf_clk.n17 VSS 0.013636f
C4658 ringtest_0.x4.clknet_1_0__leaf_clk.n18 VSS 0.04471f
C4659 ringtest_0.x4.clknet_1_0__leaf_clk.t16 VSS 0.005973f
C4660 ringtest_0.x4.clknet_1_0__leaf_clk.t18 VSS 0.005973f
C4661 ringtest_0.x4.clknet_1_0__leaf_clk.n19 VSS 0.013163f
C4662 ringtest_0.x4.clknet_1_0__leaf_clk.n20 VSS 0.043256f
C4663 ringtest_0.x4.clknet_1_0__leaf_clk.n21 VSS 0.09308f
C4664 ringtest_0.x4.clknet_1_0__leaf_clk.n22 VSS 0.067594f
C4665 ringtest_0.x4.clknet_1_0__leaf_clk.t3 VSS 0.014222f
C4666 ringtest_0.x4.clknet_1_0__leaf_clk.t6 VSS 0.014222f
C4667 ringtest_0.x4.clknet_1_0__leaf_clk.n23 VSS 0.036128f
C4668 ringtest_0.x4.clknet_1_0__leaf_clk.t8 VSS 0.014222f
C4669 ringtest_0.x4.clknet_1_0__leaf_clk.t10 VSS 0.014222f
C4670 ringtest_0.x4.clknet_1_0__leaf_clk.n24 VSS 0.029978f
C4671 ringtest_0.x4.clknet_1_0__leaf_clk.n25 VSS 0.136621f
C4672 ringtest_0.x4.clknet_1_0__leaf_clk.t5 VSS 0.014222f
C4673 ringtest_0.x4.clknet_1_0__leaf_clk.t7 VSS 0.014222f
C4674 ringtest_0.x4.clknet_1_0__leaf_clk.n26 VSS 0.029978f
C4675 ringtest_0.x4.clknet_1_0__leaf_clk.n27 VSS 0.0787f
C4676 ringtest_0.x4.clknet_1_0__leaf_clk.t9 VSS 0.014222f
C4677 ringtest_0.x4.clknet_1_0__leaf_clk.t4 VSS 0.014222f
C4678 ringtest_0.x4.clknet_1_0__leaf_clk.n28 VSS 0.029978f
C4679 ringtest_0.x4.clknet_1_0__leaf_clk.n29 VSS 0.078334f
C4680 ringtest_0.x4.clknet_1_0__leaf_clk.t12 VSS 0.014222f
C4681 ringtest_0.x4.clknet_1_0__leaf_clk.t15 VSS 0.014222f
C4682 ringtest_0.x4.clknet_1_0__leaf_clk.n30 VSS 0.029978f
C4683 ringtest_0.x4.clknet_1_0__leaf_clk.n31 VSS 0.078334f
C4684 ringtest_0.x4.clknet_1_0__leaf_clk.n32 VSS 0.04742f
C4685 ringtest_0.x4.clknet_1_0__leaf_clk.t1 VSS 0.014222f
C4686 ringtest_0.x4.clknet_1_0__leaf_clk.t2 VSS 0.014222f
C4687 ringtest_0.x4.clknet_1_0__leaf_clk.n33 VSS 0.028445f
C4688 ringtest_0.x4.clknet_1_0__leaf_clk.n34 VSS 0.022411f
C4689 ringtest_0.x4.clknet_1_0__leaf_clk.n35 VSS 0.171468f
C4690 ringtest_0.x4.clknet_1_0__leaf_clk.t39 VSS 0.014894f
C4691 ringtest_0.x4.clknet_1_0__leaf_clk.t36 VSS 0.022262f
C4692 ringtest_0.x4.clknet_1_0__leaf_clk.n36 VSS 0.040782f
C4693 ringtest_0.x4.clknet_1_0__leaf_clk.n37 VSS 0.024896f
C4694 ringtest_0.x4.clknet_1_0__leaf_clk.t33 VSS 0.022262f
C4695 ringtest_0.x4.clknet_1_0__leaf_clk.t40 VSS 0.014894f
C4696 ringtest_0.x4.clknet_1_0__leaf_clk.n38 VSS 0.040732f
C4697 ringtest_0.x4.clknet_1_0__leaf_clk.n39 VSS 0.086433f
C4698 ringtest_0.x4.clknet_1_0__leaf_clk.n40 VSS 0.225449f
C4699 ringtest_0.x4.clknet_1_0__leaf_clk.t35 VSS 0.022262f
C4700 ringtest_0.x4.clknet_1_0__leaf_clk.t34 VSS 0.014894f
C4701 ringtest_0.x4.clknet_1_0__leaf_clk.n41 VSS 0.04068f
C4702 ringtest_0.x4.clknet_1_0__leaf_clk.n42 VSS 0.027948f
C4703 ringtest_0.x4.clknet_1_0__leaf_clk.n43 VSS 0.145937f
C4704 ua[1].t4 VSS 0.322568f
C4705 ua[1].n0 VSS 0.401178f
C4706 ua[1].t1 VSS 0.24977f
C4707 ua[1].t5 VSS 0.33145f
C4708 ua[1].n1 VSS 1.6726f
C4709 ua[1].n2 VSS 0.565936f
C4710 ua[1].t2 VSS 0.244855f
C4711 ua[1].n3 VSS 0.365612f
C4712 ua[1].n4 VSS 0.509787f
C4713 ua[1].t3 VSS 0.322568f
C4714 ua[1].n5 VSS 0.401178f
C4715 ua[1].t12 VSS 0.24977f
C4716 ua[1].t11 VSS 0.33145f
C4717 ua[1].n6 VSS 1.6726f
C4718 ua[1].n7 VSS 0.565936f
C4719 ua[1].t13 VSS 0.244855f
C4720 ua[1].n8 VSS 0.365612f
C4721 ua[1].n9 VSS 0.495416f
C4722 ua[1].n10 VSS 0.270615f
C4723 ua[1].t0 VSS 0.322568f
C4724 ua[1].n11 VSS 0.401178f
C4725 ua[1].t10 VSS 0.24977f
C4726 ua[1].t6 VSS 0.33145f
C4727 ua[1].n12 VSS 1.6726f
C4728 ua[1].n13 VSS 0.565936f
C4729 ua[1].t9 VSS 0.244855f
C4730 ua[1].n14 VSS 0.365612f
C4731 ua[1].n15 VSS 0.495991f
C4732 ua[1].n16 VSS 0.268745f
C4733 ua[1].n17 VSS 0.801201f
C4734 ua[1].t8 VSS 0.322568f
C4735 ua[1].n18 VSS 0.401178f
C4736 ua[1].t14 VSS 0.24977f
C4737 ua[1].t7 VSS 0.33145f
C4738 ua[1].n19 VSS 1.6726f
C4739 ua[1].n20 VSS 0.565936f
C4740 ua[1].t15 VSS 0.244855f
C4741 ua[1].n21 VSS 0.365612f
C4742 ua[1].n22 VSS 0.500412f
C4743 ua[1].n23 VSS 0.264233f
C4744 ua[1].n24 VSS 0.382993f
C4745 ua[1].n25 VSS 7.827061f
C4746 ringtest_0.counter7.t2 VSS 0.031678f
C4747 ringtest_0.counter7.n0 VSS 0.005512f
C4748 ringtest_0.counter7.t3 VSS 0.021911f
C4749 ringtest_0.counter7.n1 VSS 0.026858f
C4750 ringtest_0.counter7.n2 VSS 0.039564f
C4751 ringtest_0.counter7.n3 VSS 0.38767f
C4752 ringtest_0.counter7.t4 VSS 0.693272f
C4753 ringtest_0.counter7.t5 VSS 0.490426f
C4754 ringtest_0.counter7.n4 VSS 3.80227f
C4755 ringtest_0.counter7.t0 VSS 0.385059f
C4756 ringtest_0.counter7.t1 VSS 0.706213f
C4757 ringtest_0.counter7.n5 VSS 3.95096f
C4758 ringtest_0.counter7.n6 VSS 0.629734f
C4759 ringtest_0.x3.x2.x4.GP VSS 2.5438f
C4760 ringtest_0.x3.x1.gpo3 VSS 1.19037f
C4761 ringtest_0.x3.x2.GP4.t3 VSS 0.012213f
C4762 ringtest_0.x3.x2.GP4.t2 VSS 0.012213f
C4763 ringtest_0.x3.x2.GP4.n0 VSS 0.026831f
C4764 ringtest_0.x3.x1.x14.Y VSS 0.075955f
C4765 ringtest_0.x3.x2.GP4.n1 VSS 0.010383f
C4766 ringtest_0.x3.x2.GP4.t4 VSS 0.618091f
C4767 ringtest_0.x3.x2.GP4.t5 VSS 0.635327f
C4768 ringtest_0.x3.x2.GP4.n2 VSS 2.25863f
C4769 ringtest_0.x3.x2.GP4.n3 VSS 0.047772f
C4770 ringtest_0.x3.x2.GP4.t1 VSS 0.01879f
C4771 ringtest_0.x3.x2.GP4.t0 VSS 0.01879f
C4772 ringtest_0.x3.x2.GP4.n4 VSS 0.043205f
C4773 ringtest_0.x3.x2.GP4.n5 VSS 0.087626f
C4774 ui_in[2].t7 VSS 0.320078f
C4775 ui_in[2].t1 VSS 0.312355f
C4776 ui_in[2].n0 VSS 1.40142f
C4777 ui_in[2].n1 VSS 0.46615f
C4778 ui_in[2].t6 VSS 0.375993f
C4779 ui_in[2].t0 VSS 0.386477f
C4780 ui_in[2].n2 VSS 1.40813f
C4781 ui_in[2].n3 VSS 0.945344f
C4782 ui_in[2].n4 VSS 2.4766f
C4783 ui_in[2].t3 VSS 0.01778f
C4784 ui_in[2].t5 VSS 0.010478f
C4785 ui_in[2].t2 VSS 0.01778f
C4786 ui_in[2].t4 VSS 0.010478f
C4787 ui_in[2].n5 VSS 0.029832f
C4788 ui_in[2].n6 VSS 0.044104f
C4789 ui_in[2].n7 VSS 0.043804f
C4790 ui_in[2].n8 VSS 0.708274f
C4791 ringtest_0.x4.net3.t0 VSS 0.067779f
C4792 ringtest_0.x4.net3.t2 VSS 0.019614f
C4793 ringtest_0.x4.net3.t7 VSS 0.031428f
C4794 ringtest_0.x4.net3.n0 VSS 0.061838f
C4795 ringtest_0.x4.net3.n1 VSS 0.008618f
C4796 ringtest_0.x4.net3.n2 VSS 0.005246f
C4797 ringtest_0.x4.net3.t6 VSS 0.029572f
C4798 ringtest_0.x4.net3.t5 VSS 0.018443f
C4799 ringtest_0.x4.net3.n3 VSS 0.059457f
C4800 ringtest_0.x4.net3.n4 VSS 0.019056f
C4801 ringtest_0.x4.net3.t4 VSS 0.030361f
C4802 ringtest_0.x4.net3.t3 VSS 0.055573f
C4803 ringtest_0.x4.net3.n5 VSS 0.744487f
C4804 ringtest_0.x4.net3.n6 VSS 0.124162f
C4805 ringtest_0.x4.net3.n7 VSS 0.092279f
C4806 ringtest_0.x4.net3.t1 VSS 0.037792f
C4807 ringtest_0.x4.net3.n8 VSS 0.040884f
C4808 ringtest_0.drv_out.t0 VSS 0.589631f
C4809 ringtest_0.drv_out.t17 VSS 0.41711f
C4810 ringtest_0.drv_out.n0 VSS 3.23385f
C4811 ringtest_0.drv_out.t19 VSS 0.327495f
C4812 ringtest_0.drv_out.t18 VSS 0.600638f
C4813 ringtest_0.drv_out.n1 VSS 3.36031f
C4814 ringtest_0.drv_out.n2 VSS 0.535592f
C4815 ringtest_0.drv_out.n3 VSS 0.10983f
C4816 ringtest_0.drv_out.t21 VSS 0.015218f
C4817 ringtest_0.drv_out.t25 VSS 0.007117f
C4818 ringtest_0.drv_out.t20 VSS 0.015218f
C4819 ringtest_0.drv_out.t24 VSS 0.007117f
C4820 ringtest_0.drv_out.t23 VSS 0.015218f
C4821 ringtest_0.drv_out.t27 VSS 0.007117f
C4822 ringtest_0.drv_out.t22 VSS 0.015218f
C4823 ringtest_0.drv_out.t26 VSS 0.007117f
C4824 ringtest_0.drv_out.n4 VSS 0.034741f
C4825 ringtest_0.drv_out.n5 VSS 0.045758f
C4826 ringtest_0.drv_out.n6 VSS 0.045758f
C4827 ringtest_0.drv_out.n7 VSS 0.055575f
C4828 ringtest_0.drv_out.n8 VSS 0.0154f
C4829 ringtest_0.drv_out.n9 VSS 0.345763f
C4830 ringtest_0.drv_out.n10 VSS 0.761878f
C4831 ringtest_0.drv_out.n11 VSS 5.52133f
C4832 ringtest_0.drv_out.t7 VSS 0.114568f
C4833 ringtest_0.drv_out.t2 VSS 0.114568f
C4834 ringtest_0.drv_out.n12 VSS 0.27282f
C4835 ringtest_0.drv_out.t4 VSS 0.114568f
C4836 ringtest_0.drv_out.t6 VSS 0.114568f
C4837 ringtest_0.drv_out.n13 VSS 0.27282f
C4838 ringtest_0.drv_out.t3 VSS 0.114568f
C4839 ringtest_0.drv_out.t5 VSS 0.114568f
C4840 ringtest_0.drv_out.n14 VSS 0.27282f
C4841 ringtest_0.drv_out.t8 VSS 0.114568f
C4842 ringtest_0.drv_out.t1 VSS 0.114568f
C4843 ringtest_0.drv_out.n15 VSS 0.27282f
C4844 ringtest_0.drv_out.n16 VSS 4.30752f
C4845 ringtest_0.drv_out.t12 VSS 0.038189f
C4846 ringtest_0.drv_out.t14 VSS 0.038189f
C4847 ringtest_0.drv_out.n17 VSS 0.093f
C4848 ringtest_0.drv_out.t13 VSS 0.038189f
C4849 ringtest_0.drv_out.t15 VSS 0.038189f
C4850 ringtest_0.drv_out.n18 VSS 0.093f
C4851 ringtest_0.drv_out.t9 VSS 0.038189f
C4852 ringtest_0.drv_out.t10 VSS 0.038189f
C4853 ringtest_0.drv_out.n19 VSS 0.093f
C4854 ringtest_0.drv_out.t16 VSS 0.038189f
C4855 ringtest_0.drv_out.t11 VSS 0.038189f
C4856 ringtest_0.drv_out.n20 VSS 0.093f
C4857 ringtest_0.drv_out.n21 VSS 1.98913f
C4858 ringtest_0.drv_out.n22 VSS 2.13865f
C4859 a_19289_13081.t12 VSS 0.136375f
C4860 a_19289_13081.t2 VSS 0.13635f
C4861 a_19289_13081.n0 VSS 0.157675f
C4862 a_19289_13081.t13 VSS 0.13635f
C4863 a_19289_13081.n1 VSS 0.086028f
C4864 a_19289_13081.t7 VSS 0.13635f
C4865 a_19289_13081.n2 VSS 0.160734f
C4866 a_19289_13081.t4 VSS 0.049796f
C4867 a_19289_13081.t15 VSS 0.049764f
C4868 a_19289_13081.n3 VSS 0.09498f
C4869 a_19289_13081.t5 VSS 0.049764f
C4870 a_19289_13081.n4 VSS 0.055718f
C4871 a_19289_13081.t11 VSS 0.049764f
C4872 a_19289_13081.n5 VSS 0.086134f
C4873 a_19289_13081.t0 VSS 0.098833f
C4874 a_19289_13081.n6 VSS 0.831842f
C4875 a_19289_13081.t6 VSS 0.049771f
C4876 a_19289_13081.t9 VSS 0.13635f
C4877 a_19289_13081.n7 VSS 0.503671f
C4878 a_19289_13081.t16 VSS 0.049764f
C4879 a_19289_13081.n8 VSS 0.212248f
C4880 a_19289_13081.t17 VSS 0.13635f
C4881 a_19289_13081.n9 VSS 0.242932f
C4882 a_19289_13081.t8 VSS 0.049764f
C4883 a_19289_13081.n10 VSS 0.212248f
C4884 a_19289_13081.t10 VSS 0.13635f
C4885 a_19289_13081.n11 VSS 0.242932f
C4886 a_19289_13081.t3 VSS 0.049764f
C4887 a_19289_13081.n12 VSS 0.212248f
C4888 a_19289_13081.t14 VSS 0.13635f
C4889 a_19289_13081.n13 VSS 0.494157f
C4890 a_19289_13081.n14 VSS 1.47337f
C4891 a_19289_13081.n15 VSS 2.33573f
C4892 a_19289_13081.t1 VSS 0.309542f
C4893 muxtest_0.R1R2.t3 VSS 0.625209f
C4894 muxtest_0.R1R2.t2 VSS 0.442278f
C4895 muxtest_0.R1R2.n0 VSS 3.42898f
C4896 muxtest_0.R1R2.t4 VSS 0.347255f
C4897 muxtest_0.R1R2.t5 VSS 0.63688f
C4898 muxtest_0.R1R2.n1 VSS 3.56307f
C4899 muxtest_0.R1R2.n2 VSS 0.56791f
C4900 muxtest_0.R1R2.n3 VSS 0.116899f
C4901 muxtest_0.R1R2.t0 VSS 0.97499f
C4902 muxtest_0.R1R2.t1 VSS 0.169683f
C4903 muxtest_0.R1R2.n4 VSS 2.37063f
C4904 muxtest_0.R1R2.n5 VSS 1.09366f
C4905 ui_in[4].t4 VSS 0.008164f
C4906 ui_in[4].t10 VSS 0.004811f
C4907 ui_in[4].t6 VSS 0.008164f
C4908 ui_in[4].t16 VSS 0.004811f
C4909 ui_in[4].n0 VSS 0.013698f
C4910 ui_in[4].n1 VSS 0.020239f
C4911 ui_in[4].n2 VSS 0.012348f
C4912 ui_in[4].t19 VSS 0.007967f
C4913 ui_in[4].t13 VSS 0.003778f
C4914 ui_in[4].n3 VSS 0.028608f
C4915 ui_in[4].n4 VSS 0.005547f
C4916 ui_in[4].n5 VSS 0.004735f
C4917 ui_in[4].t7 VSS 0.003955f
C4918 ui_in[4].t12 VSS 0.005756f
C4919 ui_in[4].n6 VSS 0.016725f
C4920 ui_in[4].n7 VSS 0.003853f
C4921 ui_in[4].n8 VSS 0.027592f
C4922 ui_in[4].n9 VSS 0.099963f
C4923 ui_in[4].t5 VSS 0.004762f
C4924 ui_in[4].t0 VSS 0.007012f
C4925 ui_in[4].n10 VSS 0.016567f
C4926 ui_in[4].n11 VSS 0.002158f
C4927 ui_in[4].n12 VSS 0.024381f
C4928 ui_in[4].n13 VSS 0.115377f
C4929 ui_in[4].n14 VSS 0.150704f
C4930 ui_in[4].n15 VSS 0.034799f
C4931 ui_in[4].t15 VSS 0.008164f
C4932 ui_in[4].t2 VSS 0.004811f
C4933 ui_in[4].t9 VSS 0.008164f
C4934 ui_in[4].t18 VSS 0.004811f
C4935 ui_in[4].n16 VSS 0.013698f
C4936 ui_in[4].n17 VSS 0.020239f
C4937 ui_in[4].n18 VSS 0.012348f
C4938 ui_in[4].t1 VSS 0.007967f
C4939 ui_in[4].t17 VSS 0.003778f
C4940 ui_in[4].n19 VSS 0.028608f
C4941 ui_in[4].n20 VSS 0.005547f
C4942 ui_in[4].n21 VSS 0.004735f
C4943 ui_in[4].t11 VSS 0.003955f
C4944 ui_in[4].t14 VSS 0.005756f
C4945 ui_in[4].n22 VSS 0.016725f
C4946 ui_in[4].n23 VSS 0.003853f
C4947 ui_in[4].n24 VSS 0.027592f
C4948 ui_in[4].n25 VSS 0.099963f
C4949 ui_in[4].t8 VSS 0.004762f
C4950 ui_in[4].t3 VSS 0.007012f
C4951 ui_in[4].n26 VSS 0.016567f
C4952 ui_in[4].n27 VSS 0.002158f
C4953 ui_in[4].n28 VSS 0.024381f
C4954 ui_in[4].n29 VSS 0.115377f
C4955 ui_in[4].n30 VSS 0.150704f
C4956 ui_in[4].n31 VSS 11.8341f
C4957 muxtest_0.R3R4.t9 VSS 0.65338f
C4958 muxtest_0.R3R4.t8 VSS 0.462206f
C4959 muxtest_0.R3R4.n0 VSS 3.58349f
C4960 muxtest_0.R3R4.t5 VSS 0.362902f
C4961 muxtest_0.R3R4.t4 VSS 0.665576f
C4962 muxtest_0.R3R4.n1 VSS 3.72361f
C4963 muxtest_0.R3R4.n2 VSS 0.593498f
C4964 muxtest_0.R3R4.n3 VSS 0.123258f
C4965 muxtest_0.R3R4.t2 VSS 1.02738f
C4966 muxtest_0.R3R4.t3 VSS 0.177328f
C4967 muxtest_0.R3R4.n4 VSS 2.29699f
C4968 muxtest_0.R3R4.t1 VSS 0.65338f
C4969 muxtest_0.R3R4.t0 VSS 0.462206f
C4970 muxtest_0.R3R4.n5 VSS 3.58349f
C4971 muxtest_0.R3R4.t6 VSS 0.362902f
C4972 muxtest_0.R3R4.t7 VSS 0.665576f
C4973 muxtest_0.R3R4.n6 VSS 3.72361f
C4974 muxtest_0.R3R4.n7 VSS 0.593498f
C4975 muxtest_0.R3R4.n8 VSS 0.122166f
C4976 muxtest_0.R3R4.n9 VSS 0.05979f
C4977 muxtest_0.R3R4.n10 VSS 6.98972f
C4978 muxtest_0.R3R4.n11 VSS 7.31123f
C4979 muxtest_0.R3R4.n12 VSS 1.03011f
C4980 ui_in[0].t6 VSS 0.006125f
C4981 ui_in[0].t0 VSS 0.003609f
C4982 ui_in[0].t8 VSS 0.006125f
C4983 ui_in[0].t3 VSS 0.003609f
C4984 ui_in[0].n0 VSS 0.010276f
C4985 ui_in[0].n1 VSS 0.015187f
C4986 ui_in[0].n2 VSS 0.004773f
C4987 ui_in[0].t9 VSS 0.003016f
C4988 ui_in[0].t5 VSS 0.004381f
C4989 ui_in[0].n3 VSS 0.010436f
C4990 ui_in[0].n4 VSS 0.005796f
C4991 ui_in[0].t1 VSS 0.003572f
C4992 ui_in[0].t7 VSS 0.00526f
C4993 ui_in[0].n5 VSS 0.012428f
C4994 ui_in[0].n6 VSS 0.002581f
C4995 ui_in[0].n7 VSS 0.001006f
C4996 ui_in[0].n8 VSS 0.091917f
C4997 ui_in[0].t4 VSS 0.005977f
C4998 ui_in[0].t2 VSS 0.002834f
C4999 ui_in[0].n9 VSS 0.021461f
C5000 ui_in[0].n10 VSS 0.004159f
C5001 ui_in[0].n11 VSS 0.105454f
C5002 ui_in[0].n12 VSS 0.068524f
C5003 ui_in[0].n13 VSS 2.54475f
C5004 ringtest_0.x4._11_.t1 VSS 0.025225f
C5005 ringtest_0.x4._11_.t0 VSS 0.025225f
C5006 ringtest_0.x4._11_.n0 VSS 0.052677f
C5007 ringtest_0.x4._11_.t12 VSS 0.042009f
C5008 ringtest_0.x4._11_.t9 VSS 0.026026f
C5009 ringtest_0.x4._11_.n1 VSS 0.085106f
C5010 ringtest_0.x4._11_.n2 VSS 0.023941f
C5011 ringtest_0.x4._11_.t7 VSS 0.026693f
C5012 ringtest_0.x4._11_.t13 VSS 0.042509f
C5013 ringtest_0.x4._11_.n3 VSS 0.057921f
C5014 ringtest_0.x4._11_.n4 VSS 0.032385f
C5015 ringtest_0.x4._11_.t17 VSS 0.023291f
C5016 ringtest_0.x4._11_.t5 VSS 0.034186f
C5017 ringtest_0.x4._11_.n5 VSS 0.06887f
C5018 ringtest_0.x4._11_.n6 VSS 0.034225f
C5019 ringtest_0.x4._11_.n7 VSS 0.488008f
C5020 ringtest_0.x4._11_.t21 VSS 0.026693f
C5021 ringtest_0.x4._11_.t10 VSS 0.042509f
C5022 ringtest_0.x4._11_.n8 VSS 0.057923f
C5023 ringtest_0.x4._11_.n9 VSS 0.132067f
C5024 ringtest_0.x4._11_.n10 VSS 0.755195f
C5025 ringtest_0.x4._11_.t11 VSS 0.020809f
C5026 ringtest_0.x4._11_.t18 VSS 0.017218f
C5027 ringtest_0.x4._11_.n11 VSS 0.090942f
C5028 ringtest_0.x4._11_.n12 VSS 0.043352f
C5029 ringtest_0.x4._11_.n13 VSS 0.147952f
C5030 ringtest_0.x4._11_.t14 VSS 0.027662f
C5031 ringtest_0.x4._11_.t4 VSS 0.01901f
C5032 ringtest_0.x4._11_.n14 VSS 0.080385f
C5033 ringtest_0.x4._11_.n15 VSS 0.011211f
C5034 ringtest_0.x4._11_.n16 VSS 0.03692f
C5035 ringtest_0.x4._11_.n17 VSS 0.154085f
C5036 ringtest_0.x4._11_.t15 VSS 0.019326f
C5037 ringtest_0.x4._11_.t19 VSS 0.028069f
C5038 ringtest_0.x4._11_.n18 VSS 0.066826f
C5039 ringtest_0.x4._11_.n19 VSS 0.141997f
C5040 ringtest_0.x4._11_.n20 VSS 0.485842f
C5041 ringtest_0.x4._11_.t8 VSS 0.04177f
C5042 ringtest_0.x4._11_.t16 VSS 0.026083f
C5043 ringtest_0.x4._11_.n21 VSS 0.079052f
C5044 ringtest_0.x4._11_.n22 VSS 0.023129f
C5045 ringtest_0.x4._11_.n23 VSS 0.351737f
C5046 ringtest_0.x4._11_.t20 VSS 0.023291f
C5047 ringtest_0.x4._11_.t6 VSS 0.034186f
C5048 ringtest_0.x4._11_.n24 VSS 0.06887f
C5049 ringtest_0.x4._11_.n25 VSS 0.014294f
C5050 ringtest_0.x4._11_.n26 VSS 0.484067f
C5051 ringtest_0.x4._11_.n27 VSS 1.17395f
C5052 ringtest_0.x4._11_.n28 VSS 0.348867f
C5053 ringtest_0.x4._11_.n29 VSS 0.0216f
C5054 ringtest_0.x4._11_.t2 VSS 0.010594f
C5055 ringtest_0.x4._11_.t3 VSS 0.010594f
C5056 ringtest_0.x4._11_.n30 VSS 0.026112f
C5057 muxtest_0.x1.x3.x4.GP VSS 2.932f
C5058 muxtest_0.x1.x2.x4.GP VSS 2.29581f
C5059 muxtest_0.x1.x1.gpo3 VSS 1.43031f
C5060 muxtest_0.x1.x3.GP4.t3 VSS 0.01297f
C5061 muxtest_0.x1.x3.GP4.t2 VSS 0.01297f
C5062 muxtest_0.x1.x3.GP4.n0 VSS 0.028494f
C5063 muxtest_0.x1.x1.x14.Y VSS 0.080663f
C5064 muxtest_0.x1.x3.GP4.n1 VSS 0.011026f
C5065 muxtest_0.x1.x3.GP4.t6 VSS 0.656398f
C5066 muxtest_0.x1.x3.GP4.t7 VSS 0.674702f
C5067 muxtest_0.x1.x3.GP4.n2 VSS 2.39862f
C5068 muxtest_0.x1.x3.GP4.t4 VSS 0.656398f
C5069 muxtest_0.x1.x3.GP4.t5 VSS 0.674702f
C5070 muxtest_0.x1.x3.GP4.n3 VSS 2.39862f
C5071 muxtest_0.x1.x3.GP4.n4 VSS 2.8073f
C5072 muxtest_0.x1.x3.GP4.n5 VSS 0.050183f
C5073 muxtest_0.x1.x3.GP4.t0 VSS 0.019954f
C5074 muxtest_0.x1.x3.GP4.t1 VSS 0.019954f
C5075 muxtest_0.x1.x3.GP4.n6 VSS 0.045883f
C5076 muxtest_0.x1.x3.GP4.n7 VSS 0.093057f
C5077 muxtest_0.x1.x3.GP1.t3 VSS 0.018021f
C5078 muxtest_0.x1.x3.GP1.t2 VSS 0.018021f
C5079 muxtest_0.x1.x3.GP1.n0 VSS 0.039591f
C5080 muxtest_0.x1.x3.GP1.n1 VSS 0.02559f
C5081 muxtest_0.x1.x3.GP1.t7 VSS 0.912037f
C5082 muxtest_0.x1.x3.GP1.t6 VSS 0.937471f
C5083 muxtest_0.x1.x3.GP1.n2 VSS 3.31176f
C5084 muxtest_0.x1.x3.GP1.t5 VSS 0.912037f
C5085 muxtest_0.x1.x3.GP1.t4 VSS 0.937471f
C5086 muxtest_0.x1.x3.GP1.n3 VSS 3.31176f
C5087 muxtest_0.x1.x3.GP1.n4 VSS 1.73806f
C5088 muxtest_0.x1.x3.GP1.t0 VSS 0.027725f
C5089 muxtest_0.x1.x3.GP1.t1 VSS 0.027725f
C5090 muxtest_0.x1.x3.GP1.n5 VSS 0.057129f
C5091 muxtest_0.x1.x3.GP1.n6 VSS 0.132634f
C5092 muxtest_0.x1.x3.GP1.n7 VSS 0.030542f
C5093 ui_in[1].t2 VSS 0.013664f
C5094 ui_in[1].t6 VSS 0.008052f
C5095 ui_in[1].t0 VSS 0.013664f
C5096 ui_in[1].t5 VSS 0.008052f
C5097 ui_in[1].n0 VSS 0.022926f
C5098 ui_in[1].n1 VSS 0.033873f
C5099 ui_in[1].n2 VSS 0.020666f
C5100 ui_in[1].t1 VSS 0.013334f
C5101 ui_in[1].t4 VSS 0.006323f
C5102 ui_in[1].n3 VSS 0.047881f
C5103 ui_in[1].n4 VSS 0.009284f
C5104 ui_in[1].n5 VSS 0.007925f
C5105 ui_in[1].t3 VSS 0.00662f
C5106 ui_in[1].t7 VSS 0.009633f
C5107 ui_in[1].n6 VSS 0.027992f
C5108 ui_in[1].n7 VSS 0.006448f
C5109 ui_in[1].n8 VSS 0.04618f
C5110 ui_in[1].n9 VSS 0.167305f
C5111 ui_in[1].t9 VSS 0.007969f
C5112 ui_in[1].t8 VSS 0.011736f
C5113 ui_in[1].n10 VSS 0.027728f
C5114 ui_in[1].n11 VSS 0.003611f
C5115 ui_in[1].n12 VSS 0.040805f
C5116 ui_in[1].n13 VSS 0.193102f
C5117 ui_in[1].n14 VSS 0.252228f
C5118 ui_in[1].n15 VSS 0.051098f
C5119 ui_in[1].n16 VSS 5.24829f
C5120 ringtest_0.x4.clknet_1_1__leaf_clk.t29 VSS 0.005541f
C5121 ringtest_0.x4.clknet_1_1__leaf_clk.t30 VSS 0.005541f
C5122 ringtest_0.x4.clknet_1_1__leaf_clk.n0 VSS 0.019676f
C5123 ringtest_0.x4.clknet_1_1__leaf_clk.t31 VSS 0.005541f
C5124 ringtest_0.x4.clknet_1_1__leaf_clk.t28 VSS 0.005541f
C5125 ringtest_0.x4.clknet_1_1__leaf_clk.n1 VSS 0.01265f
C5126 ringtest_0.x4.clknet_1_1__leaf_clk.n2 VSS 0.07993f
C5127 ringtest_0.x4.clknet_1_1__leaf_clk.t27 VSS 0.005541f
C5128 ringtest_0.x4.clknet_1_1__leaf_clk.t26 VSS 0.005541f
C5129 ringtest_0.x4.clknet_1_1__leaf_clk.n3 VSS 0.01265f
C5130 ringtest_0.x4.clknet_1_1__leaf_clk.n4 VSS 0.048044f
C5131 ringtest_0.x4.clknet_1_1__leaf_clk.t22 VSS 0.005541f
C5132 ringtest_0.x4.clknet_1_1__leaf_clk.t24 VSS 0.005541f
C5133 ringtest_0.x4.clknet_1_1__leaf_clk.n5 VSS 0.012657f
C5134 ringtest_0.x4.clknet_1_1__leaf_clk.n6 VSS 0.049559f
C5135 ringtest_0.x4.clknet_1_1__leaf_clk.t18 VSS 0.005541f
C5136 ringtest_0.x4.clknet_1_1__leaf_clk.t20 VSS 0.005541f
C5137 ringtest_0.x4.clknet_1_1__leaf_clk.n7 VSS 0.01265f
C5138 ringtest_0.x4.clknet_1_1__leaf_clk.n8 VSS 0.048044f
C5139 ringtest_0.x4.clknet_1_1__leaf_clk.t21 VSS 0.005541f
C5140 ringtest_0.x4.clknet_1_1__leaf_clk.t23 VSS 0.005541f
C5141 ringtest_0.x4.clknet_1_1__leaf_clk.n9 VSS 0.011247f
C5142 ringtest_0.x4.clknet_1_1__leaf_clk.t37 VSS 0.013817f
C5143 ringtest_0.x4.clknet_1_1__leaf_clk.t32 VSS 0.020651f
C5144 ringtest_0.x4.clknet_1_1__leaf_clk.n10 VSS 0.038168f
C5145 ringtest_0.x4.clknet_1_1__leaf_clk.t41 VSS 0.020651f
C5146 ringtest_0.x4.clknet_1_1__leaf_clk.t35 VSS 0.013817f
C5147 ringtest_0.x4.clknet_1_1__leaf_clk.n11 VSS 0.037785f
C5148 ringtest_0.x4.clknet_1_1__leaf_clk.n12 VSS 0.039947f
C5149 ringtest_0.x4.clknet_1_1__leaf_clk.t38 VSS 0.013817f
C5150 ringtest_0.x4.clknet_1_1__leaf_clk.t34 VSS 0.020651f
C5151 ringtest_0.x4.clknet_1_1__leaf_clk.n13 VSS 0.038168f
C5152 ringtest_0.x4.clknet_1_1__leaf_clk.n14 VSS 0.30833f
C5153 ringtest_0.x4.clknet_1_1__leaf_clk.t33 VSS 0.020651f
C5154 ringtest_0.x4.clknet_1_1__leaf_clk.t40 VSS 0.013817f
C5155 ringtest_0.x4.clknet_1_1__leaf_clk.n15 VSS 0.037785f
C5156 ringtest_0.x4.clknet_1_1__leaf_clk.n16 VSS 0.030886f
C5157 ringtest_0.x4.clknet_1_1__leaf_clk.n17 VSS 0.118422f
C5158 ringtest_0.x4.clknet_1_1__leaf_clk.t39 VSS 0.013817f
C5159 ringtest_0.x4.clknet_1_1__leaf_clk.t36 VSS 0.020651f
C5160 ringtest_0.x4.clknet_1_1__leaf_clk.n18 VSS 0.037832f
C5161 ringtest_0.x4.clknet_1_1__leaf_clk.n19 VSS 0.022005f
C5162 ringtest_0.x4.clknet_1_1__leaf_clk.n20 VSS 0.128874f
C5163 ringtest_0.x4.clknet_1_1__leaf_clk.n21 VSS 0.280206f
C5164 ringtest_0.x4.clknet_1_1__leaf_clk.n22 VSS 0.023331f
C5165 ringtest_0.x4.clknet_1_1__leaf_clk.n23 VSS 0.030986f
C5166 ringtest_0.x4.clknet_1_1__leaf_clk.t17 VSS 0.005541f
C5167 ringtest_0.x4.clknet_1_1__leaf_clk.t25 VSS 0.005541f
C5168 ringtest_0.x4.clknet_1_1__leaf_clk.n24 VSS 0.01265f
C5169 ringtest_0.x4.clknet_1_1__leaf_clk.n25 VSS 0.041476f
C5170 ringtest_0.x4.clknet_1_1__leaf_clk.t9 VSS 0.013193f
C5171 ringtest_0.x4.clknet_1_1__leaf_clk.t6 VSS 0.013193f
C5172 ringtest_0.x4.clknet_1_1__leaf_clk.n26 VSS 0.027449f
C5173 ringtest_0.x4.clknet_1_1__leaf_clk.t3 VSS 0.013193f
C5174 ringtest_0.x4.clknet_1_1__leaf_clk.t4 VSS 0.013193f
C5175 ringtest_0.x4.clknet_1_1__leaf_clk.n27 VSS 0.033515f
C5176 ringtest_0.x4.clknet_1_1__leaf_clk.t5 VSS 0.013193f
C5177 ringtest_0.x4.clknet_1_1__leaf_clk.t2 VSS 0.013193f
C5178 ringtest_0.x4.clknet_1_1__leaf_clk.n28 VSS 0.02781f
C5179 ringtest_0.x4.clknet_1_1__leaf_clk.n29 VSS 0.126738f
C5180 ringtest_0.x4.clknet_1_1__leaf_clk.t1 VSS 0.013193f
C5181 ringtest_0.x4.clknet_1_1__leaf_clk.t0 VSS 0.013193f
C5182 ringtest_0.x4.clknet_1_1__leaf_clk.n30 VSS 0.02781f
C5183 ringtest_0.x4.clknet_1_1__leaf_clk.n31 VSS 0.073006f
C5184 ringtest_0.x4.clknet_1_1__leaf_clk.t12 VSS 0.013193f
C5185 ringtest_0.x4.clknet_1_1__leaf_clk.t14 VSS 0.013193f
C5186 ringtest_0.x4.clknet_1_1__leaf_clk.n32 VSS 0.02781f
C5187 ringtest_0.x4.clknet_1_1__leaf_clk.n33 VSS 0.072667f
C5188 ringtest_0.x4.clknet_1_1__leaf_clk.t8 VSS 0.013193f
C5189 ringtest_0.x4.clknet_1_1__leaf_clk.t10 VSS 0.013193f
C5190 ringtest_0.x4.clknet_1_1__leaf_clk.n34 VSS 0.02781f
C5191 ringtest_0.x4.clknet_1_1__leaf_clk.n35 VSS 0.072667f
C5192 ringtest_0.x4.clknet_1_1__leaf_clk.t11 VSS 0.013193f
C5193 ringtest_0.x4.clknet_1_1__leaf_clk.t13 VSS 0.013193f
C5194 ringtest_0.x4.clknet_1_1__leaf_clk.n36 VSS 0.02781f
C5195 ringtest_0.x4.clknet_1_1__leaf_clk.n37 VSS 0.073006f
C5196 ringtest_0.x4.clknet_1_1__leaf_clk.t7 VSS 0.013193f
C5197 ringtest_0.x4.clknet_1_1__leaf_clk.t15 VSS 0.013193f
C5198 ringtest_0.x4.clknet_1_1__leaf_clk.n38 VSS 0.02781f
C5199 ringtest_0.x4.clknet_1_1__leaf_clk.n39 VSS 0.062704f
C5200 ringtest_0.x4.clknet_1_1__leaf_clk.n40 VSS 0.086346f
C5201 ringtest_0.x4.clknet_1_1__leaf_clk.n41 VSS 0.040127f
C5202 ringtest_0.x4.clknet_1_1__leaf_clk.t19 VSS 0.005541f
C5203 ringtest_0.x4.clknet_1_1__leaf_clk.t16 VSS 0.005541f
C5204 ringtest_0.x4.clknet_1_1__leaf_clk.n42 VSS 0.012211f
C5205 ringtest_0.x4.net6.t8 VSS 0.022834f
C5206 ringtest_0.x4.net6.t4 VSS 0.03372f
C5207 ringtest_0.x4.net6.n0 VSS 0.093952f
C5208 ringtest_0.x4.net6.t2 VSS 0.039666f
C5209 ringtest_0.x4.net6.t12 VSS 0.024738f
C5210 ringtest_0.x4.net6.n1 VSS 0.079752f
C5211 ringtest_0.x4.net6.n2 VSS 0.121996f
C5212 ringtest_0.x4.net6.t6 VSS 0.022834f
C5213 ringtest_0.x4.net6.t13 VSS 0.03372f
C5214 ringtest_0.x4.net6.n3 VSS 0.093952f
C5215 ringtest_0.x4.net6.n4 VSS 0.409696f
C5216 ringtest_0.x4.net6.t10 VSS 0.021035f
C5217 ringtest_0.x4.net6.t3 VSS 0.017406f
C5218 ringtest_0.x4.net6.n5 VSS 0.091932f
C5219 ringtest_0.x4.net6.n6 VSS 0.078947f
C5220 ringtest_0.x4.net6.n7 VSS 0.280597f
C5221 ringtest_0.x4.net6.t11 VSS 0.026984f
C5222 ringtest_0.x4.net6.t5 VSS 0.042972f
C5223 ringtest_0.x4.net6.n8 VSS 0.058552f
C5224 ringtest_0.x4.net6.n9 VSS 0.143174f
C5225 ringtest_0.x4.net6.n10 VSS 0.757332f
C5226 ringtest_0.x4.net6.n11 VSS 0.718043f
C5227 ringtest_0.x4.net6.t9 VSS 0.023374f
C5228 ringtest_0.x4.net6.t14 VSS 0.039666f
C5229 ringtest_0.x4.net6.n12 VSS 0.050658f
C5230 ringtest_0.x4.net6.t15 VSS 0.023374f
C5231 ringtest_0.x4.net6.t7 VSS 0.039666f
C5232 ringtest_0.x4.net6.n13 VSS 0.056268f
C5233 ringtest_0.x4.net6.n14 VSS 0.026662f
C5234 ringtest_0.x4.net6.n15 VSS 0.104019f
C5235 ringtest_0.x4.net6.n16 VSS 0.481924f
C5236 ringtest_0.x4.net6.t0 VSS 0.090914f
C5237 ringtest_0.x4.net6.n17 VSS 0.124778f
C5238 ringtest_0.x4.net6.t1 VSS 0.049897f
C5239 ringtest_0.x4.net6.n18 VSS 0.063008f
C5240 ringtest_0.x4.clknet_0_clk.t18 VSS 0.004717f
C5241 ringtest_0.x4.clknet_0_clk.t31 VSS 0.004717f
C5242 ringtest_0.x4.clknet_0_clk.n0 VSS 0.016749f
C5243 ringtest_0.x4.clknet_0_clk.t20 VSS 0.004717f
C5244 ringtest_0.x4.clknet_0_clk.t22 VSS 0.004717f
C5245 ringtest_0.x4.clknet_0_clk.n1 VSS 0.010767f
C5246 ringtest_0.x4.clknet_0_clk.n2 VSS 0.068037f
C5247 ringtest_0.x4.clknet_0_clk.t24 VSS 0.004717f
C5248 ringtest_0.x4.clknet_0_clk.t26 VSS 0.004717f
C5249 ringtest_0.x4.clknet_0_clk.n3 VSS 0.010767f
C5250 ringtest_0.x4.clknet_0_clk.n4 VSS 0.040895f
C5251 ringtest_0.x4.clknet_0_clk.t21 VSS 0.004717f
C5252 ringtest_0.x4.clknet_0_clk.t23 VSS 0.004717f
C5253 ringtest_0.x4.clknet_0_clk.n5 VSS 0.010774f
C5254 ringtest_0.x4.clknet_0_clk.n6 VSS 0.042184f
C5255 ringtest_0.x4.clknet_0_clk.t25 VSS 0.004717f
C5256 ringtest_0.x4.clknet_0_clk.t27 VSS 0.004717f
C5257 ringtest_0.x4.clknet_0_clk.n7 VSS 0.010767f
C5258 ringtest_0.x4.clknet_0_clk.n8 VSS 0.040895f
C5259 ringtest_0.x4.clknet_0_clk.t16 VSS 0.004717f
C5260 ringtest_0.x4.clknet_0_clk.t29 VSS 0.004717f
C5261 ringtest_0.x4.clknet_0_clk.n9 VSS 0.009573f
C5262 ringtest_0.x4.clknet_0_clk.t39 VSS 0.015823f
C5263 ringtest_0.x4.clknet_0_clk.t47 VSS 0.0074f
C5264 ringtest_0.x4.clknet_0_clk.t40 VSS 0.015823f
C5265 ringtest_0.x4.clknet_0_clk.t32 VSS 0.0074f
C5266 ringtest_0.x4.clknet_0_clk.t37 VSS 0.015823f
C5267 ringtest_0.x4.clknet_0_clk.t44 VSS 0.0074f
C5268 ringtest_0.x4.clknet_0_clk.t41 VSS 0.015823f
C5269 ringtest_0.x4.clknet_0_clk.t33 VSS 0.0074f
C5270 ringtest_0.x4.clknet_0_clk.n10 VSS 0.036121f
C5271 ringtest_0.x4.clknet_0_clk.n11 VSS 0.047576f
C5272 ringtest_0.x4.clknet_0_clk.n12 VSS 0.047576f
C5273 ringtest_0.x4.clknet_0_clk.n13 VSS 0.057784f
C5274 ringtest_0.x4.clknet_0_clk.n14 VSS 0.075138f
C5275 ringtest_0.x4.clknet_0_clk.t46 VSS 0.015823f
C5276 ringtest_0.x4.clknet_0_clk.t38 VSS 0.0074f
C5277 ringtest_0.x4.clknet_0_clk.t43 VSS 0.015823f
C5278 ringtest_0.x4.clknet_0_clk.t35 VSS 0.0074f
C5279 ringtest_0.x4.clknet_0_clk.t42 VSS 0.015823f
C5280 ringtest_0.x4.clknet_0_clk.t34 VSS 0.0074f
C5281 ringtest_0.x4.clknet_0_clk.t45 VSS 0.015823f
C5282 ringtest_0.x4.clknet_0_clk.t36 VSS 0.0074f
C5283 ringtest_0.x4.clknet_0_clk.n15 VSS 0.036121f
C5284 ringtest_0.x4.clknet_0_clk.n16 VSS 0.047576f
C5285 ringtest_0.x4.clknet_0_clk.n17 VSS 0.047576f
C5286 ringtest_0.x4.clknet_0_clk.n18 VSS 0.057941f
C5287 ringtest_0.x4.clknet_0_clk.n19 VSS 0.038186f
C5288 ringtest_0.x4.clknet_0_clk.n20 VSS 0.145873f
C5289 ringtest_0.x4.clknet_0_clk.n21 VSS 0.015919f
C5290 ringtest_0.x4.clknet_0_clk.n22 VSS 0.026375f
C5291 ringtest_0.x4.clknet_0_clk.t30 VSS 0.004717f
C5292 ringtest_0.x4.clknet_0_clk.t28 VSS 0.004717f
C5293 ringtest_0.x4.clknet_0_clk.n23 VSS 0.010767f
C5294 ringtest_0.x4.clknet_0_clk.n24 VSS 0.035304f
C5295 ringtest_0.x4.clknet_0_clk.t10 VSS 0.01123f
C5296 ringtest_0.x4.clknet_0_clk.t12 VSS 0.01123f
C5297 ringtest_0.x4.clknet_0_clk.n25 VSS 0.023364f
C5298 ringtest_0.x4.clknet_0_clk.t7 VSS 0.01123f
C5299 ringtest_0.x4.clknet_0_clk.t5 VSS 0.01123f
C5300 ringtest_0.x4.clknet_0_clk.n26 VSS 0.023672f
C5301 ringtest_0.x4.clknet_0_clk.t9 VSS 0.01123f
C5302 ringtest_0.x4.clknet_0_clk.t6 VSS 0.01123f
C5303 ringtest_0.x4.clknet_0_clk.n27 VSS 0.023672f
C5304 ringtest_0.x4.clknet_0_clk.t2 VSS 0.01123f
C5305 ringtest_0.x4.clknet_0_clk.t4 VSS 0.01123f
C5306 ringtest_0.x4.clknet_0_clk.n28 VSS 0.023672f
C5307 ringtest_0.x4.clknet_0_clk.t14 VSS 0.01123f
C5308 ringtest_0.x4.clknet_0_clk.t0 VSS 0.01123f
C5309 ringtest_0.x4.clknet_0_clk.n29 VSS 0.023672f
C5310 ringtest_0.x4.clknet_0_clk.t1 VSS 0.01123f
C5311 ringtest_0.x4.clknet_0_clk.t3 VSS 0.01123f
C5312 ringtest_0.x4.clknet_0_clk.n30 VSS 0.023672f
C5313 ringtest_0.x4.clknet_0_clk.t11 VSS 0.01123f
C5314 ringtest_0.x4.clknet_0_clk.t8 VSS 0.01123f
C5315 ringtest_0.x4.clknet_0_clk.n31 VSS 0.028528f
C5316 ringtest_0.x4.clknet_0_clk.t13 VSS 0.01123f
C5317 ringtest_0.x4.clknet_0_clk.t15 VSS 0.01123f
C5318 ringtest_0.x4.clknet_0_clk.n32 VSS 0.023672f
C5319 ringtest_0.x4.clknet_0_clk.n33 VSS 0.107879f
C5320 ringtest_0.x4.clknet_0_clk.n34 VSS 0.062143f
C5321 ringtest_0.x4.clknet_0_clk.n35 VSS 0.061854f
C5322 ringtest_0.x4.clknet_0_clk.n36 VSS 0.061854f
C5323 ringtest_0.x4.clknet_0_clk.n37 VSS 0.062143f
C5324 ringtest_0.x4.clknet_0_clk.n38 VSS 0.053374f
C5325 ringtest_0.x4.clknet_0_clk.n39 VSS 0.073498f
C5326 ringtest_0.x4.clknet_0_clk.n40 VSS 0.034156f
C5327 ringtest_0.x4.clknet_0_clk.t17 VSS 0.004717f
C5328 ringtest_0.x4.clknet_0_clk.t19 VSS 0.004717f
C5329 ringtest_0.x4.clknet_0_clk.n41 VSS 0.010394f
C5330 ua[2].t0 VSS 0.247385f
C5331 ua[2].n0 VSS 0.307673f
C5332 ua[2].t6 VSS 0.191554f
C5333 ua[2].t1 VSS 0.254197f
C5334 ua[2].n1 VSS 1.28275f
C5335 ua[2].n2 VSS 0.434029f
C5336 ua[2].t7 VSS 0.187785f
C5337 ua[2].n3 VSS 0.280396f
C5338 ua[2].n4 VSS 0.390968f
C5339 ua[2].t15 VSS 0.247385f
C5340 ua[2].n5 VSS 0.307673f
C5341 ua[2].t13 VSS 0.191554f
C5342 ua[2].t14 VSS 0.254197f
C5343 ua[2].n6 VSS 1.28275f
C5344 ua[2].n7 VSS 0.434029f
C5345 ua[2].t12 VSS 0.187785f
C5346 ua[2].n8 VSS 0.280396f
C5347 ua[2].n9 VSS 0.385643f
C5348 ua[2].n10 VSS 0.201153f
C5349 ua[2].n11 VSS 0.0295f
C5350 ua[2].n12 VSS 0.068599f
C5351 ua[2].n13 VSS 0.274656f
C5352 ua[2].t4 VSS 0.247385f
C5353 ua[2].n14 VSS 0.307673f
C5354 ua[2].t11 VSS 0.191554f
C5355 ua[2].t5 VSS 0.254197f
C5356 ua[2].n15 VSS 1.28275f
C5357 ua[2].n16 VSS 0.434029f
C5358 ua[2].t10 VSS 0.187785f
C5359 ua[2].n17 VSS 0.280396f
C5360 ua[2].n18 VSS 0.380387f
C5361 ua[2].n19 VSS 0.206106f
C5362 ua[2].n20 VSS 0.522334f
C5363 ua[2].t3 VSS 0.247385f
C5364 ua[2].n21 VSS 0.307673f
C5365 ua[2].t8 VSS 0.191554f
C5366 ua[2].t2 VSS 0.254197f
C5367 ua[2].n22 VSS 1.28275f
C5368 ua[2].n23 VSS 0.434029f
C5369 ua[2].t9 VSS 0.187785f
C5370 ua[2].n24 VSS 0.280396f
C5371 ua[2].n25 VSS 0.383777f
C5372 ua[2].n26 VSS 0.202647f
C5373 ua[2].n27 VSS 0.509311f
C5374 ua[2].n28 VSS 9.99833f
C5375 ua[3].t1 VSS 0.195583f
C5376 ua[3].n0 VSS 0.292041f
C5377 ua[3].t11 VSS 0.199509f
C5378 ua[3].t5 VSS 0.264753f
C5379 ua[3].n1 VSS 1.33602f
C5380 ua[3].n2 VSS 0.452054f
C5381 ua[3].t4 VSS 0.257658f
C5382 ua[3].n3 VSS 0.32045f
C5383 ua[3].n4 VSS 0.405279f
C5384 ua[3].t2 VSS 0.195583f
C5385 ua[3].n5 VSS 0.292041f
C5386 ua[3].t3 VSS 0.199509f
C5387 ua[3].t0 VSS 0.264753f
C5388 ua[3].n6 VSS 1.33602f
C5389 ua[3].n7 VSS 0.452054f
C5390 ua[3].t10 VSS 0.257658f
C5391 ua[3].n8 VSS 0.32045f
C5392 ua[3].n9 VSS 0.407204f
C5393 ua[3].t9 VSS 0.370241f
C5394 ua[3].t8 VSS 0.261912f
C5395 ua[3].n10 VSS 2.0306f
C5396 ua[3].t6 VSS 0.205641f
C5397 ua[3].t7 VSS 0.377153f
C5398 ua[3].n11 VSS 2.11001f
C5399 ua[3].n12 VSS 0.336309f
C5400 ua[3].n13 VSS 0.069845f
C5401 ua[3].n14 VSS 0.028001f
C5402 ua[3].n15 VSS 1.71586f
C5403 ua[3].n16 VSS 0.514233f
C5404 ua[3].n17 VSS 0.337655f
C5405 muxtest_0.x2.x2.GP1.t3 VSS 0.012908f
C5406 muxtest_0.x2.x2.GP1.t2 VSS 0.012908f
C5407 muxtest_0.x2.x2.GP1.n0 VSS 0.028358f
C5408 muxtest_0.x2.x2.GP1.n1 VSS 0.018329f
C5409 muxtest_0.x2.x2.GP1.t5 VSS 0.653268f
C5410 muxtest_0.x2.x2.GP1.t4 VSS 0.671486f
C5411 muxtest_0.x2.x2.GP1.n2 VSS 2.37213f
C5412 muxtest_0.x2.x2.GP1.t1 VSS 0.019859f
C5413 muxtest_0.x2.x2.GP1.t0 VSS 0.019859f
C5414 muxtest_0.x2.x2.GP1.n3 VSS 0.04092f
C5415 muxtest_0.x2.x2.GP1.n4 VSS 0.100085f
C5416 muxtest_0.x2.x2.GP1.n5 VSS 0.021877f
C5417 VDPWR.n0 VSS 0.003685f
C5418 VDPWR.t591 VSS 0.007576f
C5419 VDPWR.n1 VSS 0.008433f
C5420 VDPWR.t419 VSS 7.99e-19
C5421 VDPWR.t40 VSS 0.001213f
C5422 VDPWR.n2 VSS 0.002095f
C5423 VDPWR.t589 VSS 0.007579f
C5424 VDPWR.t612 VSS 0.007436f
C5425 VDPWR.n3 VSS 0.007083f
C5426 VDPWR.n4 VSS 0.003685f
C5427 VDPWR.n5 VSS 0.003336f
C5428 VDPWR.t458 VSS 0.001094f
C5429 VDPWR.n6 VSS 0.003106f
C5430 VDPWR.t198 VSS 0.004499f
C5431 VDPWR.n7 VSS 0.004141f
C5432 VDPWR.n8 VSS 0.003696f
C5433 VDPWR.t610 VSS 0.007579f
C5434 VDPWR.n9 VSS 6.09e-19
C5435 VDPWR.t684 VSS 0.003185f
C5436 VDPWR.t1067 VSS 0.005265f
C5437 VDPWR.n10 VSS 0.00519f
C5438 VDPWR.n11 VSS 0.00622f
C5439 VDPWR.t1217 VSS 0.021971f
C5440 VDPWR.n12 VSS 0.019873f
C5441 VDPWR.t451 VSS 5.96e-19
C5442 VDPWR.t42 VSS 0.001598f
C5443 VDPWR.n13 VSS 0.007294f
C5444 VDPWR.n14 VSS 0.003852f
C5445 VDPWR.t1068 VSS 0.005265f
C5446 VDPWR.n15 VSS 0.014377f
C5447 VDPWR.n16 VSS 0.011359f
C5448 VDPWR.n17 VSS 0.014754f
C5449 VDPWR.n18 VSS 0.008519f
C5450 VDPWR.n19 VSS 0.00622f
C5451 VDPWR.n20 VSS 0.004665f
C5452 VDPWR.n21 VSS 0.005655f
C5453 VDPWR.n22 VSS 0.00641f
C5454 VDPWR.n23 VSS 0.014463f
C5455 VDPWR.t697 VSS 0.014949f
C5456 VDPWR.n24 VSS 7.78e-19
C5457 VDPWR.n25 VSS 0.004665f
C5458 VDPWR.n26 VSS 0.001437f
C5459 VDPWR.t648 VSS 7.99e-19
C5460 VDPWR.t632 VSS 0.001213f
C5461 VDPWR.n27 VSS 0.002095f
C5462 VDPWR.n28 VSS 0.006187f
C5463 VDPWR.n29 VSS 0.003685f
C5464 VDPWR.t1282 VSS 0.021971f
C5465 VDPWR.n30 VSS 0.005477f
C5466 VDPWR.n31 VSS 0.003685f
C5467 VDPWR.t144 VSS 5.96e-19
C5468 VDPWR.t55 VSS 0.001598f
C5469 VDPWR.n32 VSS 0.007294f
C5470 VDPWR.t1268 VSS 0.021971f
C5471 VDPWR.t16 VSS 0.003219f
C5472 VDPWR.n33 VSS 0.010195f
C5473 VDPWR.n34 VSS 0.005646f
C5474 VDPWR.n35 VSS 0.003098f
C5475 VDPWR.t934 VSS 0.005265f
C5476 VDPWR.n36 VSS 0.00519f
C5477 VDPWR.n37 VSS 0.019873f
C5478 VDPWR.n38 VSS 0.008519f
C5479 VDPWR.n39 VSS 0.014754f
C5480 VDPWR.t15 VSS 0.030097f
C5481 VDPWR.t54 VSS 0.0291f
C5482 VDPWR.t933 VSS 0.021526f
C5483 VDPWR.t143 VSS 0.030894f
C5484 VDPWR.t776 VSS 0.030097f
C5485 VDPWR.t19 VSS 0.034282f
C5486 VDPWR.t631 VSS 0.024914f
C5487 VDPWR.t647 VSS 0.013354f
C5488 VDPWR.t145 VSS 0.006179f
C5489 VDPWR.t147 VSS 0.021726f
C5490 VDPWR.n40 VSS 0.02835f
C5491 VDPWR.t148 VSS 0.007539f
C5492 VDPWR.n41 VSS 0.00213f
C5493 VDPWR.n42 VSS 0.002535f
C5494 VDPWR.n43 VSS 0.01966f
C5495 VDPWR.n44 VSS 0.005779f
C5496 VDPWR.t935 VSS 0.005265f
C5497 VDPWR.n45 VSS 0.009272f
C5498 VDPWR.n46 VSS 0.011359f
C5499 VDPWR.n47 VSS 0.003854f
C5500 VDPWR.n48 VSS 0.030698f
C5501 VDPWR.n49 VSS 0.041758f
C5502 VDPWR.t1117 VSS 0.005265f
C5503 VDPWR.n50 VSS 0.010295f
C5504 VDPWR.n51 VSS 0.019873f
C5505 VDPWR.n52 VSS 0.012246f
C5506 VDPWR.t707 VSS 0.007576f
C5507 VDPWR.n53 VSS 0.008852f
C5508 VDPWR.n54 VSS 0.003685f
C5509 VDPWR.n55 VSS 0.001604f
C5510 VDPWR.n56 VSS 0.001604f
C5511 VDPWR.n57 VSS 0.108279f
C5512 VDPWR.t974 VSS 0.005265f
C5513 VDPWR.n58 VSS 0.00519f
C5514 VDPWR.n59 VSS 0.00622f
C5515 VDPWR.t1215 VSS 0.021971f
C5516 VDPWR.n60 VSS 0.019873f
C5517 VDPWR.n61 VSS 0.003852f
C5518 VDPWR.t975 VSS 0.005265f
C5519 VDPWR.n62 VSS 0.014377f
C5520 VDPWR.n63 VSS 0.015796f
C5521 VDPWR.n64 VSS 0.012246f
C5522 VDPWR.n65 VSS 0.00622f
C5523 VDPWR.n66 VSS 0.004665f
C5524 VDPWR.n67 VSS 0.00592f
C5525 VDPWR.t425 VSS 0.007579f
C5526 VDPWR.n68 VSS 0.009801f
C5527 VDPWR.n69 VSS 0.003685f
C5528 VDPWR.n70 VSS 0.00622f
C5529 VDPWR.n71 VSS 0.004665f
C5530 VDPWR.t462 VSS 0.007576f
C5531 VDPWR.n72 VSS 0.008948f
C5532 VDPWR.t18 VSS 0.007579f
C5533 VDPWR.n73 VSS 0.009682f
C5534 VDPWR.n74 VSS 0.003685f
C5535 VDPWR.n75 VSS 0.00622f
C5536 VDPWR.n76 VSS 0.004665f
C5537 VDPWR.t263 VSS 0.007576f
C5538 VDPWR.n77 VSS 0.008948f
C5539 VDPWR.t704 VSS 0.007579f
C5540 VDPWR.n78 VSS 0.009682f
C5541 VDPWR.n79 VSS 0.001604f
C5542 VDPWR.n80 VSS 0.00622f
C5543 VDPWR.n81 VSS 0.004665f
C5544 VDPWR.n82 VSS 0.002366f
C5545 VDPWR.t1116 VSS 0.06771f
C5546 VDPWR.t973 VSS 0.041598f
C5547 VDPWR.t424 VSS 0.017069f
C5548 VDPWR.t461 VSS 0.023625f
C5549 VDPWR.t17 VSS 0.017069f
C5550 VDPWR.t262 VSS 0.023625f
C5551 VDPWR.t703 VSS 0.017069f
C5552 VDPWR.t706 VSS 0.025547f
C5553 VDPWR.n83 VSS 0.027965f
C5554 VDPWR.n84 VSS 0.012927f
C5555 VDPWR.n85 VSS 0.005779f
C5556 VDPWR.t1118 VSS 0.005265f
C5557 VDPWR.n86 VSS 0.009272f
C5558 VDPWR.n87 VSS 0.015796f
C5559 VDPWR.n88 VSS 0.003144f
C5560 VDPWR.n89 VSS 0.028569f
C5561 VDPWR.n90 VSS 0.027702f
C5562 VDPWR.n91 VSS 6.42e-19
C5563 VDPWR.t146 VSS 0.007539f
C5564 VDPWR.n92 VSS 0.014062f
C5565 VDPWR.t778 VSS 0.007576f
C5566 VDPWR.n93 VSS 0.008828f
C5567 VDPWR.t20 VSS 0.002496f
C5568 VDPWR.t698 VSS 0.006635f
C5569 VDPWR.n94 VSS 0.003764f
C5570 VDPWR.t777 VSS 0.007438f
C5571 VDPWR.n95 VSS 0.007848f
C5572 VDPWR.n96 VSS 0.010094f
C5573 VDPWR.n97 VSS 0.001329f
C5574 VDPWR.n98 VSS 0.00622f
C5575 VDPWR.n99 VSS 0.003685f
C5576 VDPWR.n100 VSS 0.00213f
C5577 VDPWR.n101 VSS 0.002366f
C5578 VDPWR.n102 VSS 0.012967f
C5579 VDPWR.n103 VSS 0.034728f
C5580 VDPWR.t418 VSS 0.006577f
C5581 VDPWR.t590 VSS 0.017141f
C5582 VDPWR.t588 VSS 0.019134f
C5583 VDPWR.t39 VSS 0.013354f
C5584 VDPWR.t457 VSS 0.024914f
C5585 VDPWR.t611 VSS 0.03508f
C5586 VDPWR.t609 VSS 0.017141f
C5587 VDPWR.t197 VSS 0.013354f
C5588 VDPWR.t450 VSS 0.030894f
C5589 VDPWR.t1066 VSS 0.021526f
C5590 VDPWR.t41 VSS 0.0291f
C5591 VDPWR.t683 VSS 0.030097f
C5592 VDPWR.n104 VSS 0.020496f
C5593 VDPWR.n105 VSS 0.005954f
C5594 VDPWR.n106 VSS 0.004079f
C5595 VDPWR.n107 VSS 0.009795f
C5596 VDPWR.n108 VSS 0.002848f
C5597 VDPWR.n109 VSS 0.00622f
C5598 VDPWR.n110 VSS 0.004665f
C5599 VDPWR.n111 VSS 0.002773f
C5600 VDPWR.n112 VSS 0.009427f
C5601 VDPWR.n113 VSS 0.006495f
C5602 VDPWR.n114 VSS 0.004293f
C5603 VDPWR.n115 VSS 0.012141f
C5604 VDPWR.n116 VSS 0.077221f
C5605 VDPWR.n117 VSS 4.2675f
C5606 VDPWR.n118 VSS 0.516647f
C5607 VDPWR.t614 VSS 0.007576f
C5608 VDPWR.n119 VSS 0.008852f
C5609 VDPWR.t171 VSS 0.007579f
C5610 VDPWR.n120 VSS 0.009538f
C5611 VDPWR.n121 VSS 0.02527f
C5612 VDPWR.t173 VSS 0.007576f
C5613 VDPWR.t782 VSS 0.007579f
C5614 VDPWR.n122 VSS 0.011536f
C5615 VDPWR.t784 VSS 0.007576f
C5616 VDPWR.n123 VSS 0.008948f
C5617 VDPWR.t767 VSS 0.007579f
C5618 VDPWR.t769 VSS 0.007576f
C5619 VDPWR.n124 VSS 0.008948f
C5620 VDPWR.t324 VSS 0.007579f
C5621 VDPWR.t322 VSS 0.007576f
C5622 VDPWR.n125 VSS 0.008948f
C5623 VDPWR.t326 VSS 0.007579f
C5624 VDPWR.t328 VSS 0.007576f
C5625 VDPWR.n126 VSS 0.008948f
C5626 VDPWR.n127 VSS 0.015292f
C5627 VDPWR.n128 VSS 0.014125f
C5628 VDPWR.t357 VSS 0.007576f
C5629 VDPWR.n129 VSS 0.008948f
C5630 VDPWR.n130 VSS 0.001604f
C5631 VDPWR.n131 VSS 0.001604f
C5632 VDPWR.n132 VSS 0.001604f
C5633 VDPWR.n133 VSS 0.001604f
C5634 VDPWR.n134 VSS 0.024235f
C5635 VDPWR.t180 VSS 0.007576f
C5636 VDPWR.n135 VSS 0.008852f
C5637 VDPWR.n136 VSS 0.012476f
C5638 VDPWR.n137 VSS 0.009071f
C5639 VDPWR.n138 VSS 0.013996f
C5640 VDPWR.t252 VSS 0.007584f
C5641 VDPWR.t652 VSS 0.001902f
C5642 VDPWR.t254 VSS 0.001902f
C5643 VDPWR.n139 VSS 0.004082f
C5644 VDPWR.n140 VSS 0.005585f
C5645 VDPWR.t650 VSS 0.007372f
C5646 VDPWR.n141 VSS 0.010484f
C5647 VDPWR.n142 VSS 0.050368f
C5648 VDPWR.n143 VSS 0.001808f
C5649 VDPWR.n144 VSS 0.010569f
C5650 VDPWR.n145 VSS 0.012476f
C5651 VDPWR.t649 VSS 0.043859f
C5652 VDPWR.t651 VSS 0.018991f
C5653 VDPWR.t253 VSS 0.018991f
C5654 VDPWR.t251 VSS 0.01673f
C5655 VDPWR.n146 VSS 0.022426f
C5656 VDPWR.n147 VSS 0.024235f
C5657 VDPWR.n148 VSS 0.012476f
C5658 VDPWR.n149 VSS 0.009071f
C5659 VDPWR.n150 VSS 0.009071f
C5660 VDPWR.n151 VSS 0.014125f
C5661 VDPWR.n152 VSS 0.001604f
C5662 VDPWR.n153 VSS 0.001604f
C5663 VDPWR.n154 VSS 0.001604f
C5664 VDPWR.t359 VSS 0.007579f
C5665 VDPWR.n155 VSS 0.009682f
C5666 VDPWR.n156 VSS 0.014125f
C5667 VDPWR.n157 VSS 0.023845f
C5668 VDPWR.n158 VSS 0.017884f
C5669 VDPWR.t361 VSS 0.007576f
C5670 VDPWR.n159 VSS 0.008948f
C5671 VDPWR.t136 VSS 0.007579f
C5672 VDPWR.n160 VSS 0.009682f
C5673 VDPWR.n161 VSS 0.014125f
C5674 VDPWR.n162 VSS 0.023845f
C5675 VDPWR.n163 VSS 0.017884f
C5676 VDPWR.t138 VSS 0.007576f
C5677 VDPWR.n164 VSS 0.008948f
C5678 VDPWR.t583 VSS 0.007579f
C5679 VDPWR.n165 VSS 0.009682f
C5680 VDPWR.n166 VSS 0.014125f
C5681 VDPWR.n167 VSS 0.023845f
C5682 VDPWR.n168 VSS 0.017884f
C5683 VDPWR.t585 VSS 0.007576f
C5684 VDPWR.n169 VSS 0.008948f
C5685 VDPWR.t178 VSS 0.007579f
C5686 VDPWR.n170 VSS 0.009682f
C5687 VDPWR.n171 VSS 0.001604f
C5688 VDPWR.n172 VSS 0.023845f
C5689 VDPWR.n173 VSS 0.017884f
C5690 VDPWR.n174 VSS 0.009071f
C5691 VDPWR.n175 VSS 0.01262f
C5692 VDPWR.n176 VSS 0.029887f
C5693 VDPWR.t179 VSS 0.025547f
C5694 VDPWR.t177 VSS 0.016704f
C5695 VDPWR.t584 VSS 0.023625f
C5696 VDPWR.t582 VSS 0.017069f
C5697 VDPWR.t137 VSS 0.023625f
C5698 VDPWR.t135 VSS 0.017069f
C5699 VDPWR.t360 VSS 0.023625f
C5700 VDPWR.t358 VSS 0.017069f
C5701 VDPWR.t356 VSS 0.023625f
C5702 VDPWR.t354 VSS 0.017069f
C5703 VDPWR.t519 VSS 0.023625f
C5704 VDPWR.t517 VSS 0.017069f
C5705 VDPWR.t216 VSS 0.023625f
C5706 VDPWR.t218 VSS 0.017069f
C5707 VDPWR.t214 VSS 0.023625f
C5708 VDPWR.t212 VSS 0.017069f
C5709 VDPWR.t619 VSS 0.023625f
C5710 VDPWR.t617 VSS 0.017069f
C5711 VDPWR.n177 VSS 0.009071f
C5712 VDPWR.n178 VSS 0.027524f
C5713 VDPWR.t618 VSS 0.007579f
C5714 VDPWR.n179 VSS 0.009538f
C5715 VDPWR.n180 VSS 0.014125f
C5716 VDPWR.n181 VSS 0.023845f
C5717 VDPWR.n182 VSS 0.017884f
C5718 VDPWR.t620 VSS 0.007576f
C5719 VDPWR.n183 VSS 0.008948f
C5720 VDPWR.t213 VSS 0.007579f
C5721 VDPWR.n184 VSS 0.009682f
C5722 VDPWR.n185 VSS 0.014125f
C5723 VDPWR.n186 VSS 0.023845f
C5724 VDPWR.n187 VSS 0.017884f
C5725 VDPWR.t215 VSS 0.007576f
C5726 VDPWR.n188 VSS 0.008948f
C5727 VDPWR.t219 VSS 0.007579f
C5728 VDPWR.n189 VSS 0.009682f
C5729 VDPWR.n190 VSS 0.014125f
C5730 VDPWR.n191 VSS 0.023845f
C5731 VDPWR.n192 VSS 0.017884f
C5732 VDPWR.t217 VSS 0.007576f
C5733 VDPWR.n193 VSS 0.008948f
C5734 VDPWR.t518 VSS 0.007579f
C5735 VDPWR.n194 VSS 0.009682f
C5736 VDPWR.n195 VSS 0.014125f
C5737 VDPWR.n196 VSS 0.023845f
C5738 VDPWR.n197 VSS 0.017884f
C5739 VDPWR.t520 VSS 0.007576f
C5740 VDPWR.n198 VSS 0.008948f
C5741 VDPWR.t355 VSS 0.007579f
C5742 VDPWR.n199 VSS 0.009682f
C5743 VDPWR.n200 VSS 0.001604f
C5744 VDPWR.n201 VSS 0.014514f
C5745 VDPWR.n202 VSS 1.71998f
C5746 VDPWR.n203 VSS 1.7218f
C5747 VDPWR.t530 VSS 0.007579f
C5748 VDPWR.t528 VSS 0.007576f
C5749 VDPWR.n204 VSS 0.008948f
C5750 VDPWR.t551 VSS 0.007579f
C5751 VDPWR.t549 VSS 0.007576f
C5752 VDPWR.n205 VSS 0.008948f
C5753 VDPWR.t553 VSS 0.007579f
C5754 VDPWR.t555 VSS 0.007576f
C5755 VDPWR.n206 VSS 0.008948f
C5756 VDPWR.t616 VSS 0.007579f
C5757 VDPWR.n207 VSS 0.02527f
C5758 VDPWR.n208 VSS 0.030581f
C5759 VDPWR.n209 VSS 0.001604f
C5760 VDPWR.n210 VSS 0.009682f
C5761 VDPWR.n211 VSS 0.011536f
C5762 VDPWR.n212 VSS 0.02527f
C5763 VDPWR.n213 VSS 0.030581f
C5764 VDPWR.n214 VSS 0.001604f
C5765 VDPWR.n215 VSS 0.009682f
C5766 VDPWR.n216 VSS 0.011536f
C5767 VDPWR.n217 VSS 0.02527f
C5768 VDPWR.n218 VSS 0.030581f
C5769 VDPWR.n219 VSS 0.001604f
C5770 VDPWR.n220 VSS 0.009682f
C5771 VDPWR.n221 VSS 0.011536f
C5772 VDPWR.n222 VSS 0.02527f
C5773 VDPWR.n223 VSS 0.030581f
C5774 VDPWR.n224 VSS 0.001604f
C5775 VDPWR.n225 VSS 0.009682f
C5776 VDPWR.n226 VSS 0.011536f
C5777 VDPWR.n227 VSS 0.02527f
C5778 VDPWR.n228 VSS 0.020509f
C5779 VDPWR.n229 VSS 0.001604f
C5780 VDPWR.n230 VSS 0.009682f
C5781 VDPWR.n231 VSS 0.011536f
C5782 VDPWR.n232 VSS 0.02527f
C5783 VDPWR.n233 VSS 0.030581f
C5784 VDPWR.n234 VSS 0.001604f
C5785 VDPWR.n235 VSS 0.009682f
C5786 VDPWR.n236 VSS 0.011536f
C5787 VDPWR.n237 VSS 0.02527f
C5788 VDPWR.n238 VSS 0.030581f
C5789 VDPWR.n239 VSS 0.001604f
C5790 VDPWR.n240 VSS 0.009682f
C5791 VDPWR.n241 VSS 0.011536f
C5792 VDPWR.n242 VSS 0.02527f
C5793 VDPWR.n243 VSS 0.030581f
C5794 VDPWR.n244 VSS 0.001604f
C5795 VDPWR.n245 VSS 0.009682f
C5796 VDPWR.n246 VSS 0.008948f
C5797 VDPWR.n247 VSS 0.001604f
C5798 VDPWR.n248 VSS 0.030581f
C5799 VDPWR.n249 VSS 0.011536f
C5800 VDPWR.n250 VSS 0.032879f
C5801 VDPWR.t170 VSS 0.013225f
C5802 VDPWR.t172 VSS 0.027468f
C5803 VDPWR.t781 VSS 0.013225f
C5804 VDPWR.t783 VSS 0.027468f
C5805 VDPWR.t766 VSS 0.013225f
C5806 VDPWR.t768 VSS 0.027468f
C5807 VDPWR.t323 VSS 0.013225f
C5808 VDPWR.t321 VSS 0.027468f
C5809 VDPWR.t325 VSS 0.013225f
C5810 VDPWR.t327 VSS 0.027468f
C5811 VDPWR.t529 VSS 0.013225f
C5812 VDPWR.t527 VSS 0.027468f
C5813 VDPWR.t550 VSS 0.013225f
C5814 VDPWR.t548 VSS 0.027468f
C5815 VDPWR.t552 VSS 0.013225f
C5816 VDPWR.t554 VSS 0.027468f
C5817 VDPWR.t615 VSS 0.013225f
C5818 VDPWR.t613 VSS 0.038494f
C5819 VDPWR.n251 VSS 0.037336f
C5820 VDPWR.n252 VSS 0.012818f
C5821 VDPWR.n253 VSS 14.456599f
C5822 VDPWR.n254 VSS 0.061316f
C5823 VDPWR.n255 VSS 0.111329f
C5824 VDPWR.n256 VSS 2.79006f
C5825 VDPWR.n257 VSS 0.003685f
C5826 VDPWR.t132 VSS 0.007576f
C5827 VDPWR.n258 VSS 0.008433f
C5828 VDPWR.t104 VSS 7.99e-19
C5829 VDPWR.t686 VSS 0.001213f
C5830 VDPWR.n259 VSS 0.002095f
C5831 VDPWR.t134 VSS 0.007579f
C5832 VDPWR.t343 VSS 0.007436f
C5833 VDPWR.n260 VSS 0.007083f
C5834 VDPWR.n261 VSS 0.003685f
C5835 VDPWR.n262 VSS 0.003336f
C5836 VDPWR.t108 VSS 0.001094f
C5837 VDPWR.n263 VSS 0.003106f
C5838 VDPWR.t341 VSS 0.004499f
C5839 VDPWR.n264 VSS 0.004141f
C5840 VDPWR.n265 VSS 0.003696f
C5841 VDPWR.t345 VSS 0.007579f
C5842 VDPWR.n266 VSS 6.09e-19
C5843 VDPWR.t38 VSS 0.003185f
C5844 VDPWR.t945 VSS 0.005265f
C5845 VDPWR.n267 VSS 0.00519f
C5846 VDPWR.n268 VSS 0.00622f
C5847 VDPWR.t1228 VSS 0.021971f
C5848 VDPWR.n269 VSS 0.019873f
C5849 VDPWR.t119 VSS 5.96e-19
C5850 VDPWR.t347 VSS 0.001598f
C5851 VDPWR.n270 VSS 0.007294f
C5852 VDPWR.n271 VSS 0.003852f
C5853 VDPWR.t946 VSS 0.005265f
C5854 VDPWR.n272 VSS 0.014377f
C5855 VDPWR.n273 VSS 0.011359f
C5856 VDPWR.n274 VSS 0.014754f
C5857 VDPWR.n275 VSS 0.008519f
C5858 VDPWR.n276 VSS 0.00622f
C5859 VDPWR.n277 VSS 0.004665f
C5860 VDPWR.n278 VSS 0.005655f
C5861 VDPWR.n279 VSS 0.00641f
C5862 VDPWR.n280 VSS 0.014463f
C5863 VDPWR.t567 VSS 0.014949f
C5864 VDPWR.n281 VSS 7.78e-19
C5865 VDPWR.n282 VSS 0.004665f
C5866 VDPWR.n283 VSS 0.001437f
C5867 VDPWR.t628 VSS 7.99e-19
C5868 VDPWR.t239 VSS 0.001213f
C5869 VDPWR.n284 VSS 0.002095f
C5870 VDPWR.n285 VSS 0.006187f
C5871 VDPWR.n286 VSS 0.003685f
C5872 VDPWR.t1201 VSS 0.021971f
C5873 VDPWR.n287 VSS 0.005477f
C5874 VDPWR.n288 VSS 0.003685f
C5875 VDPWR.t624 VSS 5.96e-19
C5876 VDPWR.t110 VSS 0.001598f
C5877 VDPWR.n289 VSS 0.007294f
C5878 VDPWR.t1200 VSS 0.021971f
C5879 VDPWR.t102 VSS 0.003219f
C5880 VDPWR.n290 VSS 0.010195f
C5881 VDPWR.n291 VSS 0.005646f
C5882 VDPWR.n292 VSS 0.003098f
C5883 VDPWR.t1005 VSS 0.005265f
C5884 VDPWR.n293 VSS 0.00519f
C5885 VDPWR.n294 VSS 0.019873f
C5886 VDPWR.n295 VSS 0.008519f
C5887 VDPWR.n296 VSS 0.014754f
C5888 VDPWR.t101 VSS 0.030097f
C5889 VDPWR.t109 VSS 0.0291f
C5890 VDPWR.t1004 VSS 0.021526f
C5891 VDPWR.t623 VSS 0.030894f
C5892 VDPWR.t758 VSS 0.030097f
C5893 VDPWR.t434 VSS 0.034282f
C5894 VDPWR.t238 VSS 0.024914f
C5895 VDPWR.t627 VSS 0.013354f
C5896 VDPWR.t774 VSS 0.006179f
C5897 VDPWR.t772 VSS 0.021726f
C5898 VDPWR.n297 VSS 0.02835f
C5899 VDPWR.t773 VSS 0.007539f
C5900 VDPWR.n298 VSS 0.00213f
C5901 VDPWR.n299 VSS 0.002535f
C5902 VDPWR.n300 VSS 0.01966f
C5903 VDPWR.n301 VSS 0.005779f
C5904 VDPWR.t1006 VSS 0.005265f
C5905 VDPWR.n302 VSS 0.009272f
C5906 VDPWR.n303 VSS 0.011359f
C5907 VDPWR.n304 VSS 0.003854f
C5908 VDPWR.n305 VSS 0.030698f
C5909 VDPWR.n306 VSS 0.041758f
C5910 VDPWR.t1002 VSS 0.005265f
C5911 VDPWR.n307 VSS 0.010295f
C5912 VDPWR.n308 VSS 0.019873f
C5913 VDPWR.n309 VSS 0.012246f
C5914 VDPWR.t752 VSS 0.007576f
C5915 VDPWR.n310 VSS 0.008852f
C5916 VDPWR.n311 VSS 0.003685f
C5917 VDPWR.n312 VSS 0.001604f
C5918 VDPWR.n313 VSS 0.001604f
C5919 VDPWR.n314 VSS 0.108279f
C5920 VDPWR.t841 VSS 0.005265f
C5921 VDPWR.n315 VSS 0.00519f
C5922 VDPWR.n316 VSS 0.00622f
C5923 VDPWR.t1263 VSS 0.021971f
C5924 VDPWR.n317 VSS 0.019873f
C5925 VDPWR.t842 VSS 0.005265f
C5926 VDPWR.n318 VSS 0.003852f
C5927 VDPWR.n319 VSS 0.014377f
C5928 VDPWR.n320 VSS 0.015796f
C5929 VDPWR.n321 VSS 0.012246f
C5930 VDPWR.n322 VSS 0.00622f
C5931 VDPWR.n323 VSS 0.004665f
C5932 VDPWR.n324 VSS 0.00592f
C5933 VDPWR.t626 VSS 0.007579f
C5934 VDPWR.n325 VSS 0.009801f
C5935 VDPWR.n326 VSS 0.003685f
C5936 VDPWR.n327 VSS 0.00622f
C5937 VDPWR.n328 VSS 0.004665f
C5938 VDPWR.t630 VSS 0.007576f
C5939 VDPWR.n329 VSS 0.008948f
C5940 VDPWR.t433 VSS 0.007579f
C5941 VDPWR.n330 VSS 0.009682f
C5942 VDPWR.n331 VSS 0.003685f
C5943 VDPWR.n332 VSS 0.00622f
C5944 VDPWR.n333 VSS 0.004665f
C5945 VDPWR.t351 VSS 0.007576f
C5946 VDPWR.n334 VSS 0.008948f
C5947 VDPWR.t754 VSS 0.007579f
C5948 VDPWR.n335 VSS 0.009682f
C5949 VDPWR.n336 VSS 0.001604f
C5950 VDPWR.n337 VSS 0.00622f
C5951 VDPWR.n338 VSS 0.004665f
C5952 VDPWR.n339 VSS 0.002366f
C5953 VDPWR.t1001 VSS 0.06771f
C5954 VDPWR.t840 VSS 0.041598f
C5955 VDPWR.t625 VSS 0.017069f
C5956 VDPWR.t629 VSS 0.023625f
C5957 VDPWR.t432 VSS 0.017069f
C5958 VDPWR.t350 VSS 0.023625f
C5959 VDPWR.t753 VSS 0.017069f
C5960 VDPWR.t751 VSS 0.025547f
C5961 VDPWR.n340 VSS 0.027965f
C5962 VDPWR.n341 VSS 0.012927f
C5963 VDPWR.n342 VSS 0.005779f
C5964 VDPWR.t1003 VSS 0.005265f
C5965 VDPWR.n343 VSS 0.009272f
C5966 VDPWR.n344 VSS 0.015796f
C5967 VDPWR.n345 VSS 0.003144f
C5968 VDPWR.n346 VSS 0.028569f
C5969 VDPWR.n347 VSS 0.027702f
C5970 VDPWR.n348 VSS 6.42e-19
C5971 VDPWR.t775 VSS 0.007539f
C5972 VDPWR.n349 VSS 0.014062f
C5973 VDPWR.t757 VSS 0.007576f
C5974 VDPWR.n350 VSS 0.008828f
C5975 VDPWR.t435 VSS 0.002496f
C5976 VDPWR.t568 VSS 0.006635f
C5977 VDPWR.n351 VSS 0.003764f
C5978 VDPWR.t759 VSS 0.007438f
C5979 VDPWR.n352 VSS 0.007848f
C5980 VDPWR.n353 VSS 0.010094f
C5981 VDPWR.n354 VSS 0.001329f
C5982 VDPWR.n355 VSS 0.00622f
C5983 VDPWR.n356 VSS 0.003685f
C5984 VDPWR.n357 VSS 0.00213f
C5985 VDPWR.n358 VSS 0.002366f
C5986 VDPWR.n359 VSS 0.012967f
C5987 VDPWR.n360 VSS 0.034728f
C5988 VDPWR.t103 VSS 0.006577f
C5989 VDPWR.t131 VSS 0.017141f
C5990 VDPWR.t133 VSS 0.019134f
C5991 VDPWR.t685 VSS 0.013354f
C5992 VDPWR.t107 VSS 0.024914f
C5993 VDPWR.t342 VSS 0.03508f
C5994 VDPWR.t344 VSS 0.017141f
C5995 VDPWR.t340 VSS 0.013354f
C5996 VDPWR.t118 VSS 0.030894f
C5997 VDPWR.t944 VSS 0.021526f
C5998 VDPWR.t346 VSS 0.0291f
C5999 VDPWR.t37 VSS 0.030097f
C6000 VDPWR.n361 VSS 0.020496f
C6001 VDPWR.n362 VSS 0.005954f
C6002 VDPWR.n363 VSS 0.004079f
C6003 VDPWR.n364 VSS 0.009795f
C6004 VDPWR.n365 VSS 0.002848f
C6005 VDPWR.n366 VSS 0.00622f
C6006 VDPWR.n367 VSS 0.004665f
C6007 VDPWR.n368 VSS 0.002773f
C6008 VDPWR.n369 VSS 0.009427f
C6009 VDPWR.n370 VSS 0.006495f
C6010 VDPWR.n371 VSS 0.004293f
C6011 VDPWR.n372 VSS 0.012141f
C6012 VDPWR.n373 VSS 0.094729f
C6013 VDPWR.n374 VSS 0.062411f
C6014 VDPWR.n375 VSS 0.121043f
C6015 VDPWR.n376 VSS 0.336123f
C6016 VDPWR.n377 VSS 0.120947f
C6017 VDPWR.n378 VSS 0.059393f
C6018 VDPWR.n379 VSS 0.080969f
C6019 VDPWR.n380 VSS 0.059303f
C6020 VDPWR.n381 VSS 0.491964f
C6021 VDPWR.t362 VSS 0.654139f
C6022 VDPWR.n384 VSS 0.491964f
C6023 VDPWR.n385 VSS 0.058532f
C6024 VDPWR.n386 VSS 0.038385f
C6025 VDPWR.n387 VSS 0.077333f
C6026 VDPWR.n388 VSS 0.040191f
C6027 VDPWR.n389 VSS 0.120947f
C6028 VDPWR.n390 VSS 0.059393f
C6029 VDPWR.n391 VSS 0.080969f
C6030 VDPWR.n392 VSS 0.059303f
C6031 VDPWR.n393 VSS 0.491964f
C6032 VDPWR.t547 VSS 0.654139f
C6033 VDPWR.n396 VSS 0.491964f
C6034 VDPWR.n397 VSS 0.058532f
C6035 VDPWR.n398 VSS 0.038385f
C6036 VDPWR.n399 VSS 0.077333f
C6037 VDPWR.n400 VSS 0.075451f
C6038 VDPWR.n401 VSS 0.180684f
C6039 VDPWR.n402 VSS 0.077737f
C6040 VDPWR.n403 VSS 0.037257f
C6041 VDPWR.n404 VSS 0.120941f
C6042 VDPWR.n405 VSS 0.058602f
C6043 VDPWR.n406 VSS 0.058602f
C6044 VDPWR.n407 VSS 0.058411f
C6045 VDPWR.n408 VSS 0.080977f
C6046 VDPWR.n409 VSS 0.261065f
C6047 VDPWR.t662 VSS 0.376779f
C6048 VDPWR.n410 VSS 0.363781f
C6049 VDPWR.t661 VSS 0.376779f
C6050 VDPWR.n411 VSS 0.261065f
C6051 VDPWR.n412 VSS 2.27e-19
C6052 VDPWR.n413 VSS 0.027354f
C6053 VDPWR.n414 VSS 0.037257f
C6054 VDPWR.n415 VSS 0.080977f
C6055 VDPWR.n416 VSS 0.261065f
C6056 VDPWR.n417 VSS 2.51e-19
C6057 VDPWR.n418 VSS 0.261065f
C6058 VDPWR.t466 VSS 0.376779f
C6059 VDPWR.t467 VSS 0.376779f
C6060 VDPWR.n419 VSS 0.058411f
C6061 VDPWR.n420 VSS 0.058602f
C6062 VDPWR.n421 VSS 0.363781f
C6063 VDPWR.n422 VSS 0.058602f
C6064 VDPWR.n423 VSS 0.120941f
C6065 VDPWR.n424 VSS 0.064054f
C6066 VDPWR.n425 VSS 0.019206f
C6067 VDPWR.n426 VSS 0.031115f
C6068 VDPWR.n427 VSS 0.077293f
C6069 VDPWR.n428 VSS 0.089305f
C6070 VDPWR.n429 VSS 0.037221f
C6071 VDPWR.n430 VSS 0.120941f
C6072 VDPWR.n431 VSS 0.004701f
C6073 VDPWR.n432 VSS 0.058602f
C6074 VDPWR.n433 VSS 0.058602f
C6075 VDPWR.n434 VSS 0.058411f
C6076 VDPWR.n435 VSS 0.080977f
C6077 VDPWR.n436 VSS 0.261065f
C6078 VDPWR.t711 VSS 0.376779f
C6079 VDPWR.n437 VSS 0.363781f
C6080 VDPWR.t714 VSS 0.376779f
C6081 VDPWR.n438 VSS 0.261065f
C6082 VDPWR.n439 VSS 0.002139f
C6083 VDPWR.n440 VSS 0.064116f
C6084 VDPWR.n441 VSS 0.019206f
C6085 VDPWR.n442 VSS 0.030814f
C6086 VDPWR.n443 VSS 0.071389f
C6087 VDPWR.n444 VSS 0.086966f
C6088 VDPWR.n445 VSS 0.037101f
C6089 VDPWR.n446 VSS 0.120941f
C6090 VDPWR.n447 VSS 0.004709f
C6091 VDPWR.n448 VSS 0.058602f
C6092 VDPWR.n449 VSS 0.058602f
C6093 VDPWR.n450 VSS 0.058411f
C6094 VDPWR.n451 VSS 0.080977f
C6095 VDPWR.n452 VSS 0.261065f
C6096 VDPWR.t247 VSS 0.376779f
C6097 VDPWR.n453 VSS 0.363781f
C6098 VDPWR.t248 VSS 0.376779f
C6099 VDPWR.n454 VSS 0.261065f
C6100 VDPWR.n455 VSS 0.002259f
C6101 VDPWR.n456 VSS 0.064116f
C6102 VDPWR.n457 VSS 0.019206f
C6103 VDPWR.n458 VSS 0.030814f
C6104 VDPWR.n459 VSS 0.068877f
C6105 VDPWR.n460 VSS 0.07947f
C6106 VDPWR.n461 VSS 0.006609f
C6107 VDPWR.n462 VSS 0.064079f
C6108 VDPWR.n463 VSS 0.019206f
C6109 VDPWR.n464 VSS 0.031091f
C6110 VDPWR.n465 VSS 0.068139f
C6111 VDPWR.n466 VSS 0.091071f
C6112 VDPWR.n467 VSS 0.037257f
C6113 VDPWR.n468 VSS 0.120941f
C6114 VDPWR.n469 VSS 0.058602f
C6115 VDPWR.n470 VSS 0.058602f
C6116 VDPWR.n471 VSS 0.058411f
C6117 VDPWR.n472 VSS 0.080977f
C6118 VDPWR.n473 VSS 0.261065f
C6119 VDPWR.t464 VSS 0.376779f
C6120 VDPWR.n474 VSS 0.363781f
C6121 VDPWR.t465 VSS 0.376779f
C6122 VDPWR.n475 VSS 0.261065f
C6123 VDPWR.n476 VSS 2.51e-19
C6124 VDPWR.n477 VSS 0.006628f
C6125 VDPWR.n478 VSS 0.064054f
C6126 VDPWR.n479 VSS 0.019206f
C6127 VDPWR.n480 VSS 0.031115f
C6128 VDPWR.n481 VSS 0.046281f
C6129 VDPWR.n482 VSS 0.112591f
C6130 VDPWR.n483 VSS 0.037221f
C6131 VDPWR.n484 VSS 0.120941f
C6132 VDPWR.n485 VSS 0.004701f
C6133 VDPWR.n486 VSS 0.058602f
C6134 VDPWR.n487 VSS 0.058602f
C6135 VDPWR.n488 VSS 0.058411f
C6136 VDPWR.n489 VSS 0.080977f
C6137 VDPWR.n490 VSS 0.261065f
C6138 VDPWR.t713 VSS 0.376779f
C6139 VDPWR.n491 VSS 0.363781f
C6140 VDPWR.t712 VSS 0.376779f
C6141 VDPWR.n492 VSS 0.261065f
C6142 VDPWR.n493 VSS 0.002139f
C6143 VDPWR.n494 VSS 0.064116f
C6144 VDPWR.n495 VSS 0.019206f
C6145 VDPWR.n496 VSS 0.030814f
C6146 VDPWR.n497 VSS 0.071389f
C6147 VDPWR.n498 VSS 0.086966f
C6148 VDPWR.n499 VSS 0.037101f
C6149 VDPWR.n500 VSS 0.120941f
C6150 VDPWR.n501 VSS 0.004709f
C6151 VDPWR.n502 VSS 0.058602f
C6152 VDPWR.n503 VSS 0.058602f
C6153 VDPWR.n504 VSS 0.058411f
C6154 VDPWR.n505 VSS 0.080977f
C6155 VDPWR.n506 VSS 0.261065f
C6156 VDPWR.t246 VSS 0.376779f
C6157 VDPWR.n507 VSS 0.363781f
C6158 VDPWR.t49 VSS 0.376779f
C6159 VDPWR.n508 VSS 0.261065f
C6160 VDPWR.n509 VSS 0.002259f
C6161 VDPWR.n510 VSS 0.064116f
C6162 VDPWR.n511 VSS 0.019206f
C6163 VDPWR.n512 VSS 0.030814f
C6164 VDPWR.n513 VSS 0.068509f
C6165 VDPWR.n514 VSS 0.090982f
C6166 VDPWR.n515 VSS 0.037257f
C6167 VDPWR.n516 VSS 0.120941f
C6168 VDPWR.n517 VSS 0.058602f
C6169 VDPWR.n518 VSS 0.058602f
C6170 VDPWR.n519 VSS 0.058411f
C6171 VDPWR.n520 VSS 0.080977f
C6172 VDPWR.n521 VSS 0.261065f
C6173 VDPWR.t660 VSS 0.376779f
C6174 VDPWR.n522 VSS 0.363781f
C6175 VDPWR.t659 VSS 0.376779f
C6176 VDPWR.n523 VSS 0.261065f
C6177 VDPWR.n524 VSS 2.27e-19
C6178 VDPWR.n525 VSS 0.006609f
C6179 VDPWR.n526 VSS 0.064079f
C6180 VDPWR.n527 VSS 0.019206f
C6181 VDPWR.n528 VSS 0.031091f
C6182 VDPWR.n529 VSS 0.114673f
C6183 VDPWR.n530 VSS 0.429043f
C6184 VDPWR.n531 VSS 1.08249f
C6185 VDPWR.t708 VSS 0.002958f
C6186 VDPWR.t1202 VSS 0.001743f
C6187 VDPWR.t699 VSS 0.002958f
C6188 VDPWR.t1193 VSS 0.001743f
C6189 VDPWR.n532 VSS 0.004963f
C6190 VDPWR.n533 VSS 0.007338f
C6191 VDPWR.n534 VSS 0.007288f
C6192 VDPWR.n535 VSS 0.002975f
C6193 VDPWR.n536 VSS 0.387509f
C6194 VDPWR.n537 VSS 0.003685f
C6195 VDPWR.t534 VSS 0.007576f
C6196 VDPWR.n538 VSS 0.008433f
C6197 VDPWR.t417 VSS 7.99e-19
C6198 VDPWR.t106 VSS 0.001213f
C6199 VDPWR.n539 VSS 0.002095f
C6200 VDPWR.t532 VSS 0.007579f
C6201 VDPWR.t658 VSS 0.007436f
C6202 VDPWR.n540 VSS 0.007083f
C6203 VDPWR.n541 VSS 0.003685f
C6204 VDPWR.n542 VSS 0.003336f
C6205 VDPWR.t57 VSS 0.001094f
C6206 VDPWR.n543 VSS 0.003106f
C6207 VDPWR.t738 VSS 0.004499f
C6208 VDPWR.n544 VSS 0.004141f
C6209 VDPWR.n545 VSS 0.003696f
C6210 VDPWR.t656 VSS 0.007579f
C6211 VDPWR.n546 VSS 6.09e-19
C6212 VDPWR.t274 VSS 0.003185f
C6213 VDPWR.t1087 VSS 0.005265f
C6214 VDPWR.n547 VSS 0.00519f
C6215 VDPWR.n548 VSS 0.00622f
C6216 VDPWR.t1207 VSS 0.021971f
C6217 VDPWR.n549 VSS 0.019873f
C6218 VDPWR.t516 VSS 5.96e-19
C6219 VDPWR.t117 VSS 0.001598f
C6220 VDPWR.n550 VSS 0.007294f
C6221 VDPWR.n551 VSS 0.003852f
C6222 VDPWR.t1088 VSS 0.005265f
C6223 VDPWR.n552 VSS 0.014377f
C6224 VDPWR.n553 VSS 0.011359f
C6225 VDPWR.n554 VSS 0.014754f
C6226 VDPWR.n555 VSS 0.008519f
C6227 VDPWR.n556 VSS 0.00622f
C6228 VDPWR.n557 VSS 0.004665f
C6229 VDPWR.n558 VSS 0.005655f
C6230 VDPWR.n559 VSS 0.00641f
C6231 VDPWR.n560 VSS 0.014463f
C6232 VDPWR.t723 VSS 0.014949f
C6233 VDPWR.n561 VSS 7.78e-19
C6234 VDPWR.n562 VSS 0.004665f
C6235 VDPWR.n563 VSS 0.001437f
C6236 VDPWR.t53 VSS 7.99e-19
C6237 VDPWR.t227 VSS 0.001213f
C6238 VDPWR.n564 VSS 0.002095f
C6239 VDPWR.n565 VSS 0.006187f
C6240 VDPWR.n566 VSS 0.003685f
C6241 VDPWR.t1261 VSS 0.021971f
C6242 VDPWR.n567 VSS 0.005477f
C6243 VDPWR.n568 VSS 0.003685f
C6244 VDPWR.t36 VSS 5.96e-19
C6245 VDPWR.t427 VSS 0.001598f
C6246 VDPWR.n569 VSS 0.007294f
C6247 VDPWR.t1214 VSS 0.021971f
C6248 VDPWR.t265 VSS 0.003219f
C6249 VDPWR.n570 VSS 0.010195f
C6250 VDPWR.n571 VSS 0.005646f
C6251 VDPWR.n572 VSS 0.003098f
C6252 VDPWR.t1073 VSS 0.005265f
C6253 VDPWR.n573 VSS 0.00519f
C6254 VDPWR.n574 VSS 0.019873f
C6255 VDPWR.n575 VSS 0.008519f
C6256 VDPWR.n576 VSS 0.014754f
C6257 VDPWR.t264 VSS 0.030097f
C6258 VDPWR.t426 VSS 0.0291f
C6259 VDPWR.t1072 VSS 0.021526f
C6260 VDPWR.t35 VSS 0.030894f
C6261 VDPWR.t429 VSS 0.030097f
C6262 VDPWR.t266 VSS 0.034282f
C6263 VDPWR.t226 VSS 0.024914f
C6264 VDPWR.t52 VSS 0.013354f
C6265 VDPWR.t228 VSS 0.006179f
C6266 VDPWR.t230 VSS 0.021726f
C6267 VDPWR.n577 VSS 0.02835f
C6268 VDPWR.t231 VSS 0.007539f
C6269 VDPWR.n578 VSS 0.00213f
C6270 VDPWR.n579 VSS 0.002535f
C6271 VDPWR.n580 VSS 0.01966f
C6272 VDPWR.n581 VSS 0.005779f
C6273 VDPWR.t1074 VSS 0.005265f
C6274 VDPWR.n582 VSS 0.009272f
C6275 VDPWR.n583 VSS 0.011359f
C6276 VDPWR.n584 VSS 0.003854f
C6277 VDPWR.n585 VSS 0.030698f
C6278 VDPWR.n586 VSS 0.041758f
C6279 VDPWR.t1105 VSS 0.005265f
C6280 VDPWR.n587 VSS 0.010295f
C6281 VDPWR.n588 VSS 0.019873f
C6282 VDPWR.n589 VSS 0.012246f
C6283 VDPWR.t701 VSS 0.007576f
C6284 VDPWR.n590 VSS 0.008852f
C6285 VDPWR.n591 VSS 0.003685f
C6286 VDPWR.n592 VSS 0.001604f
C6287 VDPWR.n593 VSS 0.001604f
C6288 VDPWR.n594 VSS 0.108279f
C6289 VDPWR.t922 VSS 0.005265f
C6290 VDPWR.n595 VSS 0.00519f
C6291 VDPWR.n596 VSS 0.00622f
C6292 VDPWR.t1205 VSS 0.021971f
C6293 VDPWR.n597 VSS 0.019873f
C6294 VDPWR.n598 VSS 0.003852f
C6295 VDPWR.t923 VSS 0.005265f
C6296 VDPWR.n599 VSS 0.014377f
C6297 VDPWR.n600 VSS 0.015796f
C6298 VDPWR.n601 VSS 0.012246f
C6299 VDPWR.n602 VSS 0.00622f
C6300 VDPWR.n603 VSS 0.004665f
C6301 VDPWR.n604 VSS 0.00592f
C6302 VDPWR.t460 VSS 0.007579f
C6303 VDPWR.n605 VSS 0.009801f
C6304 VDPWR.n606 VSS 0.003685f
C6305 VDPWR.n607 VSS 0.00622f
C6306 VDPWR.n608 VSS 0.004665f
C6307 VDPWR.t51 VSS 0.007576f
C6308 VDPWR.n609 VSS 0.008948f
C6309 VDPWR.t421 VSS 0.007579f
C6310 VDPWR.n610 VSS 0.009682f
C6311 VDPWR.n611 VSS 0.003685f
C6312 VDPWR.n612 VSS 0.00622f
C6313 VDPWR.n613 VSS 0.004665f
C6314 VDPWR.t423 VSS 0.007576f
C6315 VDPWR.n614 VSS 0.008948f
C6316 VDPWR.t710 VSS 0.007579f
C6317 VDPWR.n615 VSS 0.009682f
C6318 VDPWR.n616 VSS 0.001604f
C6319 VDPWR.n617 VSS 0.00622f
C6320 VDPWR.n618 VSS 0.004665f
C6321 VDPWR.n619 VSS 0.002366f
C6322 VDPWR.t1104 VSS 0.06771f
C6323 VDPWR.t921 VSS 0.041598f
C6324 VDPWR.t459 VSS 0.017069f
C6325 VDPWR.t50 VSS 0.023625f
C6326 VDPWR.t420 VSS 0.017069f
C6327 VDPWR.t422 VSS 0.023625f
C6328 VDPWR.t709 VSS 0.017069f
C6329 VDPWR.t700 VSS 0.025547f
C6330 VDPWR.n620 VSS 0.027965f
C6331 VDPWR.n621 VSS 0.012927f
C6332 VDPWR.n622 VSS 0.005779f
C6333 VDPWR.t1106 VSS 0.005265f
C6334 VDPWR.n623 VSS 0.009272f
C6335 VDPWR.n624 VSS 0.015796f
C6336 VDPWR.n625 VSS 0.003144f
C6337 VDPWR.n626 VSS 0.028569f
C6338 VDPWR.n627 VSS 0.027702f
C6339 VDPWR.n628 VSS 6.42e-19
C6340 VDPWR.t229 VSS 0.007539f
C6341 VDPWR.n629 VSS 0.014062f
C6342 VDPWR.t428 VSS 0.007576f
C6343 VDPWR.n630 VSS 0.008828f
C6344 VDPWR.t267 VSS 0.002496f
C6345 VDPWR.t724 VSS 0.006635f
C6346 VDPWR.n631 VSS 0.003764f
C6347 VDPWR.t430 VSS 0.007438f
C6348 VDPWR.n632 VSS 0.007848f
C6349 VDPWR.n633 VSS 0.010094f
C6350 VDPWR.n634 VSS 0.001329f
C6351 VDPWR.n635 VSS 0.00622f
C6352 VDPWR.n636 VSS 0.003685f
C6353 VDPWR.n637 VSS 0.00213f
C6354 VDPWR.n638 VSS 0.002366f
C6355 VDPWR.n639 VSS 0.012967f
C6356 VDPWR.n640 VSS 0.034728f
C6357 VDPWR.t416 VSS 0.006577f
C6358 VDPWR.t533 VSS 0.017141f
C6359 VDPWR.t531 VSS 0.019134f
C6360 VDPWR.t105 VSS 0.013354f
C6361 VDPWR.t56 VSS 0.024914f
C6362 VDPWR.t657 VSS 0.03508f
C6363 VDPWR.t655 VSS 0.017141f
C6364 VDPWR.t737 VSS 0.013354f
C6365 VDPWR.t515 VSS 0.030894f
C6366 VDPWR.t1086 VSS 0.021526f
C6367 VDPWR.t116 VSS 0.0291f
C6368 VDPWR.t273 VSS 0.030097f
C6369 VDPWR.n641 VSS 0.020496f
C6370 VDPWR.n642 VSS 0.005954f
C6371 VDPWR.n643 VSS 0.004079f
C6372 VDPWR.n644 VSS 0.009795f
C6373 VDPWR.n645 VSS 0.002848f
C6374 VDPWR.n646 VSS 0.00622f
C6375 VDPWR.n647 VSS 0.004665f
C6376 VDPWR.n648 VSS 0.002773f
C6377 VDPWR.n649 VSS 0.009427f
C6378 VDPWR.n650 VSS 0.006495f
C6379 VDPWR.n651 VSS 0.004293f
C6380 VDPWR.n652 VSS 0.012141f
C6381 VDPWR.n653 VSS 0.077221f
C6382 VDPWR.n654 VSS 0.039488f
C6383 VDPWR.n655 VSS 0.124227f
C6384 VDPWR.n656 VSS 0.027354f
C6385 VDPWR.n657 VSS 0.037257f
C6386 VDPWR.n658 VSS 0.080977f
C6387 VDPWR.n659 VSS 0.261065f
C6388 VDPWR.n660 VSS 2.51e-19
C6389 VDPWR.n661 VSS 0.261065f
C6390 VDPWR.t5 VSS 0.376779f
C6391 VDPWR.t4 VSS 0.376779f
C6392 VDPWR.n662 VSS 0.058411f
C6393 VDPWR.n663 VSS 0.058602f
C6394 VDPWR.n664 VSS 0.363781f
C6395 VDPWR.n665 VSS 0.058602f
C6396 VDPWR.n666 VSS 0.120941f
C6397 VDPWR.n667 VSS 0.064054f
C6398 VDPWR.n668 VSS 0.019206f
C6399 VDPWR.n669 VSS 0.031115f
C6400 VDPWR.n670 VSS 0.077293f
C6401 VDPWR.n671 VSS 0.089305f
C6402 VDPWR.n672 VSS 0.037221f
C6403 VDPWR.n673 VSS 0.120941f
C6404 VDPWR.n674 VSS 0.004701f
C6405 VDPWR.n675 VSS 0.058602f
C6406 VDPWR.n676 VSS 0.058602f
C6407 VDPWR.n677 VSS 0.058411f
C6408 VDPWR.n678 VSS 0.080977f
C6409 VDPWR.n679 VSS 0.261065f
C6410 VDPWR.t75 VSS 0.376779f
C6411 VDPWR.n680 VSS 0.363781f
C6412 VDPWR.t76 VSS 0.376779f
C6413 VDPWR.n681 VSS 0.261065f
C6414 VDPWR.n682 VSS 0.002139f
C6415 VDPWR.n683 VSS 0.064116f
C6416 VDPWR.n684 VSS 0.019206f
C6417 VDPWR.n685 VSS 0.030814f
C6418 VDPWR.n686 VSS 0.071389f
C6419 VDPWR.n687 VSS 0.086966f
C6420 VDPWR.n688 VSS 0.037101f
C6421 VDPWR.n689 VSS 0.120941f
C6422 VDPWR.n690 VSS 0.004709f
C6423 VDPWR.n691 VSS 0.058602f
C6424 VDPWR.n692 VSS 0.058602f
C6425 VDPWR.n693 VSS 0.058411f
C6426 VDPWR.n694 VSS 0.080977f
C6427 VDPWR.n695 VSS 0.261065f
C6428 VDPWR.t111 VSS 0.376779f
C6429 VDPWR.n696 VSS 0.363781f
C6430 VDPWR.t94 VSS 0.376779f
C6431 VDPWR.n697 VSS 0.261065f
C6432 VDPWR.n698 VSS 0.002259f
C6433 VDPWR.n699 VSS 0.064116f
C6434 VDPWR.n700 VSS 0.019206f
C6435 VDPWR.n701 VSS 0.030814f
C6436 VDPWR.n702 VSS 0.068509f
C6437 VDPWR.n703 VSS 0.090904f
C6438 VDPWR.n704 VSS 0.037257f
C6439 VDPWR.n705 VSS 0.120941f
C6440 VDPWR.n706 VSS 0.058602f
C6441 VDPWR.n707 VSS 0.058602f
C6442 VDPWR.n708 VSS 0.058411f
C6443 VDPWR.n709 VSS 0.080977f
C6444 VDPWR.n710 VSS 0.261065f
C6445 VDPWR.t536 VSS 0.376779f
C6446 VDPWR.n711 VSS 0.363781f
C6447 VDPWR.t535 VSS 0.376779f
C6448 VDPWR.n712 VSS 0.261065f
C6449 VDPWR.n713 VSS 2.27e-19
C6450 VDPWR.n714 VSS 0.006609f
C6451 VDPWR.n715 VSS 0.064079f
C6452 VDPWR.n716 VSS 0.019206f
C6453 VDPWR.n717 VSS 0.031091f
C6454 VDPWR.n718 VSS 0.062837f
C6455 VDPWR.n719 VSS 0.378608f
C6456 VDPWR.n720 VSS 5.63728f
C6457 VDPWR.t175 VSS 0.126772f
C6458 VDPWR.t44 VSS 0.078772f
C6459 VDPWR.t483 VSS 0.020918f
C6460 VDPWR.t716 VSS 0.020918f
C6461 VDPWR.n721 VSS 0.050136f
C6462 VDPWR.n722 VSS 0.447486f
C6463 VDPWR.t48 VSS 0.078753f
C6464 VDPWR.t485 VSS 0.020918f
C6465 VDPWR.t481 VSS 0.020918f
C6466 VDPWR.n723 VSS 0.050136f
C6467 VDPWR.n724 VSS 0.437151f
C6468 VDPWR.t469 VSS 0.020918f
C6469 VDPWR.t46 VSS 0.020918f
C6470 VDPWR.n725 VSS 0.050136f
C6471 VDPWR.n726 VSS 0.167913f
C6472 VDPWR.n727 VSS 0.068395f
C6473 VDPWR.n728 VSS 0.024369f
C6474 VDPWR.n729 VSS 0.037597f
C6475 VDPWR.n730 VSS 0.037597f
C6476 VDPWR.n731 VSS 0.037597f
C6477 VDPWR.n732 VSS 0.036475f
C6478 VDPWR.n733 VSS 0.230589f
C6479 VDPWR.t43 VSS 0.221262f
C6480 VDPWR.t482 VSS 0.151317f
C6481 VDPWR.t715 VSS 0.151317f
C6482 VDPWR.t468 VSS 0.113488f
C6483 VDPWR.n734 VSS 0.075658f
C6484 VDPWR.t45 VSS 0.113488f
C6485 VDPWR.t484 VSS 0.151317f
C6486 VDPWR.t480 VSS 0.151317f
C6487 VDPWR.t47 VSS 0.221262f
C6488 VDPWR.n735 VSS 0.230589f
C6489 VDPWR.n736 VSS 0.036464f
C6490 VDPWR.n737 VSS 0.024368f
C6491 VDPWR.n738 VSS 0.319602f
C6492 VDPWR.n739 VSS 0.015428f
C6493 VDPWR.n740 VSS 0.029611f
C6494 VDPWR.n741 VSS 0.029611f
C6495 VDPWR.t174 VSS 0.285184f
C6496 VDPWR.n742 VSS 0.028847f
C6497 VDPWR.n744 VSS 0.218999f
C6498 VDPWR.n745 VSS 0.029611f
C6499 VDPWR.n747 VSS 0.218999f
C6500 VDPWR.n748 VSS 0.028833f
C6501 VDPWR.n749 VSS 0.015424f
C6502 VDPWR.n750 VSS 0.180441f
C6503 VDPWR.n751 VSS 0.335772f
C6504 VDPWR.n752 VSS 0.491355f
C6505 VDPWR.n753 VSS 1.00522f
C6506 VDPWR.n754 VSS 1.15962f
C6507 VDPWR.n755 VSS 4.50177f
C6508 VDPWR.n756 VSS 3.34127f
C6509 VDPWR.n757 VSS 1.35096f
C6510 VDPWR.n758 VSS 0.170679f
C6511 VDPWR.n759 VSS 0.037257f
C6512 VDPWR.n760 VSS 0.120941f
C6513 VDPWR.n761 VSS 0.058602f
C6514 VDPWR.n762 VSS 0.058602f
C6515 VDPWR.n763 VSS 0.058411f
C6516 VDPWR.n764 VSS 0.080977f
C6517 VDPWR.n765 VSS 0.261065f
C6518 VDPWR.t602 VSS 0.376779f
C6519 VDPWR.n766 VSS 0.363781f
C6520 VDPWR.t176 VSS 0.376779f
C6521 VDPWR.n767 VSS 0.261065f
C6522 VDPWR.n768 VSS 2.27e-19
C6523 VDPWR.n769 VSS 0.367889f
C6524 VDPWR.n770 VSS 0.013567f
C6525 VDPWR.n771 VSS 0.003227f
C6526 VDPWR.n772 VSS 0.001668f
C6527 VDPWR.n773 VSS 0.001668f
C6528 VDPWR.n774 VSS 0.248273f
C6529 VDPWR.n775 VSS 0.231572f
C6530 VDPWR.n776 VSS 0.297449f
C6531 VDPWR.n777 VSS 0.13021f
C6532 VDPWR.n778 VSS 0.12621f
C6533 VDPWR.n779 VSS 0.001668f
C6534 VDPWR.n780 VSS 0.003227f
C6535 VDPWR.n781 VSS 0.003227f
C6536 VDPWR.n782 VSS 0.002085f
C6537 VDPWR.n783 VSS 0.002164f
C6538 VDPWR.n784 VSS 5.79e-19
C6539 VDPWR.t636 VSS 0.003189f
C6540 VDPWR.n785 VSS 0.00651f
C6541 VDPWR.n786 VSS 0.002366f
C6542 VDPWR.t936 VSS 0.055011f
C6543 VDPWR.t260 VSS 0.030495f
C6544 VDPWR.t442 VSS 0.023719f
C6545 VDPWR.t947 VSS 0.030894f
C6546 VDPWR.t1160 VSS 0.036276f
C6547 VDPWR.t477 VSS 0.023719f
C6548 VDPWR.t912 VSS 0.030894f
C6549 VDPWR.t876 VSS 0.033286f
C6550 VDPWR.t679 VSS 0.035478f
C6551 VDPWR.t717 VSS 0.024117f
C6552 VDPWR.t329 VSS 0.043451f
C6553 VDPWR.t279 VSS 0.01754f
C6554 VDPWR.t639 VSS 0.011162f
C6555 VDPWR.t691 VSS 0.018337f
C6556 VDPWR.t749 VSS 0.0584f
C6557 VDPWR.t689 VSS 0.063582f
C6558 VDPWR.t1032 VSS 0.021526f
C6559 VDPWR.t645 VSS 0.0291f
C6560 VDPWR.t633 VSS 0.030097f
C6561 VDPWR.n787 VSS 0.040309f
C6562 VDPWR.t1033 VSS 0.005265f
C6563 VDPWR.n788 VSS 0.009272f
C6564 VDPWR.t634 VSS 0.003189f
C6565 VDPWR.t1198 VSS 0.038955f
C6566 VDPWR.n789 VSS 0.012601f
C6567 VDPWR.n790 VSS 0.004665f
C6568 VDPWR.t690 VSS 5.96e-19
C6569 VDPWR.t646 VSS 0.001598f
C6570 VDPWR.n791 VSS 0.007294f
C6571 VDPWR.n792 VSS 0.014754f
C6572 VDPWR.t750 VSS 0.007935f
C6573 VDPWR.n793 VSS 0.017811f
C6574 VDPWR.t1034 VSS 0.005265f
C6575 VDPWR.n794 VSS 0.005101f
C6576 VDPWR.t640 VSS 0.001614f
C6577 VDPWR.t330 VSS 0.001614f
C6578 VDPWR.n795 VSS 0.003509f
C6579 VDPWR.n796 VSS 0.008256f
C6580 VDPWR.n797 VSS 0.002164f
C6581 VDPWR.n798 VSS 0.002085f
C6582 VDPWR.n799 VSS 0.001668f
C6583 VDPWR.n800 VSS 0.003227f
C6584 VDPWR.n801 VSS 0.002085f
C6585 VDPWR.n802 VSS 0.003115f
C6586 VDPWR.t280 VSS 0.007746f
C6587 VDPWR.n803 VSS 0.005712f
C6588 VDPWR.n804 VSS 0.001832f
C6589 VDPWR.n805 VSS 0.001555f
C6590 VDPWR.n806 VSS 0.001555f
C6591 VDPWR.n807 VSS 8.79e-19
C6592 VDPWR.n808 VSS 0.001689f
C6593 VDPWR.t718 VSS 0.001449f
C6594 VDPWR.t680 VSS 0.002395f
C6595 VDPWR.n809 VSS 0.00662f
C6596 VDPWR.n810 VSS 0.00858f
C6597 VDPWR.t1259 VSS 0.030953f
C6598 VDPWR.n811 VSS 0.016328f
C6599 VDPWR.n812 VSS 0.003685f
C6600 VDPWR.t913 VSS 0.005308f
C6601 VDPWR.t1265 VSS 0.011265f
C6602 VDPWR.n814 VSS 0.028883f
C6603 VDPWR.t914 VSS 0.005308f
C6604 VDPWR.n815 VSS 0.014284f
C6605 VDPWR.t948 VSS 0.005302f
C6606 VDPWR.n816 VSS 0.002464f
C6607 VDPWR.t1245 VSS 0.040015f
C6608 VDPWR.n817 VSS 0.068285f
C6609 VDPWR.n818 VSS 0.021111f
C6610 VDPWR.t443 VSS 0.001614f
C6611 VDPWR.t261 VSS 0.001614f
C6612 VDPWR.n819 VSS 0.003509f
C6613 VDPWR.n820 VSS 0.02258f
C6614 VDPWR.n821 VSS 7.78e-19
C6615 VDPWR.n822 VSS 0.002085f
C6616 VDPWR.n823 VSS 0.00311f
C6617 VDPWR.t949 VSS 0.005265f
C6618 VDPWR.n824 VSS 0.009272f
C6619 VDPWR.n825 VSS 0.005779f
C6620 VDPWR.t937 VSS 0.005308f
C6621 VDPWR.t1248 VSS 0.011265f
C6622 VDPWR.n827 VSS 0.028883f
C6623 VDPWR.t938 VSS 0.005308f
C6624 VDPWR.n828 VSS 0.015733f
C6625 VDPWR.n829 VSS 0.002164f
C6626 VDPWR.t1061 VSS 0.005308f
C6627 VDPWR.t1185 VSS 0.011265f
C6628 VDPWR.n831 VSS 0.028883f
C6629 VDPWR.t1062 VSS 0.005308f
C6630 VDPWR.n832 VSS 0.015733f
C6631 VDPWR.n833 VSS 0.002085f
C6632 VDPWR.n834 VSS 0.002231f
C6633 VDPWR.n835 VSS 0.003047f
C6634 VDPWR.n836 VSS 0.001454f
C6635 VDPWR.n837 VSS 0.013261f
C6636 VDPWR.n838 VSS 0.002164f
C6637 VDPWR.n839 VSS 0.001555f
C6638 VDPWR.n840 VSS 0.002085f
C6639 VDPWR.n841 VSS 0.003227f
C6640 VDPWR.n842 VSS 0.003115f
C6641 VDPWR.n843 VSS 0.005443f
C6642 VDPWR.n844 VSS 0.00213f
C6643 VDPWR.n845 VSS 0.016328f
C6644 VDPWR.n846 VSS 0.0134f
C6645 VDPWR.n847 VSS 0.002366f
C6646 VDPWR.n848 VSS 0.005827f
C6647 VDPWR.t478 VSS 0.001614f
C6648 VDPWR.t1161 VSS 0.001614f
C6649 VDPWR.n849 VSS 0.00353f
C6650 VDPWR.n850 VSS 0.020862f
C6651 VDPWR.n851 VSS 0.00213f
C6652 VDPWR.n852 VSS 0.00213f
C6653 VDPWR.n853 VSS 0.005018f
C6654 VDPWR.t878 VSS 0.005349f
C6655 VDPWR.n854 VSS 0.007928f
C6656 VDPWR.n855 VSS 0.01998f
C6657 VDPWR.n856 VSS 0.021356f
C6658 VDPWR.n857 VSS 0.00622f
C6659 VDPWR.n858 VSS 0.004665f
C6660 VDPWR.n859 VSS 0.002535f
C6661 VDPWR.n860 VSS 0.042017f
C6662 VDPWR.t877 VSS 0.005265f
C6663 VDPWR.n861 VSS 0.009272f
C6664 VDPWR.n862 VSS 0.002988f
C6665 VDPWR.n863 VSS 0.002164f
C6666 VDPWR.n864 VSS 0.001555f
C6667 VDPWR.n865 VSS 0.002085f
C6668 VDPWR.n866 VSS 0.001668f
C6669 VDPWR.n867 VSS 0.245208f
C6670 VDPWR.n868 VSS 0.003595f
C6671 VDPWR.n869 VSS 0.003719f
C6672 VDPWR.n870 VSS 0.003115f
C6673 VDPWR.n871 VSS 0.001668f
C6674 VDPWR.n872 VSS 0.002164f
C6675 VDPWR.n873 VSS 0.002164f
C6676 VDPWR.n874 VSS 0.003257f
C6677 VDPWR.n875 VSS 0.003115f
C6678 VDPWR.t98 VSS 0.001426f
C6679 VDPWR.t100 VSS 0.002942f
C6680 VDPWR.n876 VSS 0.00599f
C6681 VDPWR.n877 VSS 0.001976f
C6682 VDPWR.t194 VSS 0.002994f
C6683 VDPWR.n878 VSS 0.004665f
C6684 VDPWR.t113 VSS 0.001902f
C6685 VDPWR.t320 VSS 0.001902f
C6686 VDPWR.n879 VSS 0.004259f
C6687 VDPWR.n880 VSS 0.005483f
C6688 VDPWR.n881 VSS 0.004665f
C6689 VDPWR.t722 VSS 0.006676f
C6690 VDPWR.n882 VSS 0.012783f
C6691 VDPWR.t449 VSS 0.001902f
C6692 VDPWR.t730 VSS 0.001902f
C6693 VDPWR.n883 VSS 0.004139f
C6694 VDPWR.n884 VSS 0.002164f
C6695 VDPWR.n885 VSS 0.002085f
C6696 VDPWR.n886 VSS 0.003719f
C6697 VDPWR.n887 VSS 0.245208f
C6698 VDPWR.n888 VSS 0.003719f
C6699 VDPWR.n889 VSS 0.002912f
C6700 VDPWR.n890 VSS 0.001668f
C6701 VDPWR.n891 VSS 0.001668f
C6702 VDPWR.n892 VSS 0.002085f
C6703 VDPWR.n893 VSS 0.00311f
C6704 VDPWR.t1270 VSS 0.021971f
C6705 VDPWR.t28 VSS 0.001598f
C6706 VDPWR.t256 VSS 5.96e-19
C6707 VDPWR.n894 VSS 0.007294f
C6708 VDPWR.n895 VSS 0.001703f
C6709 VDPWR.n896 VSS 0.008296f
C6710 VDPWR.t32 VSS 0.002465f
C6711 VDPWR.t696 VSS 0.002395f
C6712 VDPWR.n897 VSS 0.005711f
C6713 VDPWR.t728 VSS 0.002324f
C6714 VDPWR.t502 VSS 0.002324f
C6715 VDPWR.n898 VSS 0.004738f
C6716 VDPWR.n899 VSS 0.00622f
C6717 VDPWR.t150 VSS 0.001183f
C6718 VDPWR.t158 VSS -0.001244f
C6719 VDPWR.n900 VSS 0.007903f
C6720 VDPWR.n901 VSS 0.00182f
C6721 VDPWR.n902 VSS 0.00622f
C6722 VDPWR.t80 VSS 0.001183f
C6723 VDPWR.t66 VSS -0.001244f
C6724 VDPWR.n903 VSS 0.007903f
C6725 VDPWR.t414 VSS 0.001217f
C6726 VDPWR.t542 VSS 0.001217f
C6727 VDPWR.n904 VSS 0.002534f
C6728 VDPWR.t581 VSS 0.002921f
C6729 VDPWR.n905 VSS 0.005646f
C6730 VDPWR.n906 VSS 0.001589f
C6731 VDPWR.t575 VSS 7.99e-19
C6732 VDPWR.t665 VSS 7.99e-19
C6733 VDPWR.n907 VSS 0.001849f
C6734 VDPWR.t560 VSS 0.001217f
C6735 VDPWR.t644 VSS 0.001217f
C6736 VDPWR.n908 VSS 0.002534f
C6737 VDPWR.n909 VSS 0.007542f
C6738 VDPWR.n910 VSS 0.002231f
C6739 VDPWR.n911 VSS 0.002085f
C6740 VDPWR.n912 VSS 0.003719f
C6741 VDPWR.n913 VSS 0.245208f
C6742 VDPWR.n914 VSS 0.189315f
C6743 VDPWR.n915 VSS 0.003719f
C6744 VDPWR.n916 VSS 0.003115f
C6745 VDPWR.n917 VSS 0.001668f
C6746 VDPWR.n918 VSS 0.005882f
C6747 VDPWR.t544 VSS 0.002933f
C6748 VDPWR.t573 VSS 0.001426f
C6749 VDPWR.t233 VSS 0.002942f
C6750 VDPWR.n919 VSS 0.00599f
C6751 VDPWR.n920 VSS 0.002203f
C6752 VDPWR.n921 VSS 0.00622f
C6753 VDPWR.t349 VSS 0.001426f
C6754 VDPWR.t339 VSS 0.002942f
C6755 VDPWR.n922 VSS 0.00599f
C6756 VDPWR.t188 VSS 0.002968f
C6757 VDPWR.n923 VSS 0.002107f
C6758 VDPWR.n924 VSS 0.004665f
C6759 VDPWR.t335 VSS 0.002968f
C6760 VDPWR.t901 VSS 0.005308f
C6761 VDPWR.t1267 VSS 0.011265f
C6762 VDPWR.n926 VSS 0.028883f
C6763 VDPWR.t902 VSS 0.005308f
C6764 VDPWR.n927 VSS 0.015733f
C6765 VDPWR.t337 VSS 0.001902f
C6766 VDPWR.t142 VSS 0.001902f
C6767 VDPWR.n928 VSS 0.004275f
C6768 VDPWR.n929 VSS 0.015248f
C6769 VDPWR.n930 VSS 0.002164f
C6770 VDPWR.n931 VSS 0.002085f
C6771 VDPWR.n932 VSS 0.003719f
C6772 VDPWR.n933 VSS 0.245208f
C6773 VDPWR.n934 VSS 0.12621f
C6774 VDPWR.n935 VSS 0.003719f
C6775 VDPWR.n936 VSS 0.003115f
C6776 VDPWR.n937 VSS 0.001668f
C6777 VDPWR.n938 VSS 0.001425f
C6778 VDPWR.t331 VSS 0.001217f
C6779 VDPWR.t571 VSS 0.001217f
C6780 VDPWR.n939 VSS 0.002534f
C6781 VDPWR.n940 VSS 0.00622f
C6782 VDPWR.n941 VSS 0.002203f
C6783 VDPWR.n942 VSS 0.00622f
C6784 VDPWR.t456 VSS 0.001426f
C6785 VDPWR.t192 VSS 0.002942f
C6786 VDPWR.n943 VSS 0.00599f
C6787 VDPWR.t271 VSS 0.001426f
C6788 VDPWR.t272 VSS 0.002942f
C6789 VDPWR.n944 VSS 0.00599f
C6790 VDPWR.n945 VSS 0.002203f
C6791 VDPWR.n946 VSS 0.003178f
C6792 VDPWR.t125 VSS 0.001902f
C6793 VDPWR.t333 VSS 0.001902f
C6794 VDPWR.n947 VSS 0.004259f
C6795 VDPWR.t827 VSS 0.001902f
C6796 VDPWR.t366 VSS 0.001902f
C6797 VDPWR.n948 VSS 0.004259f
C6798 VDPWR.n949 VSS 0.009864f
C6799 VDPWR.n950 VSS 0.00311f
C6800 VDPWR.n951 VSS 0.002236f
C6801 VDPWR.n952 VSS 0.001668f
C6802 VDPWR.n953 VSS 0.003719f
C6803 VDPWR.n954 VSS 0.245208f
C6804 VDPWR.n955 VSS 0.003595f
C6805 VDPWR.n956 VSS 0.003719f
C6806 VDPWR.n957 VSS 0.007619f
C6807 VDPWR.n958 VSS 0.001668f
C6808 VDPWR.n959 VSS 0.00311f
C6809 VDPWR.n960 VSS 0.016932f
C6810 VDPWR.n961 VSS 0.016932f
C6811 VDPWR.t1030 VSS 0.005308f
C6812 VDPWR.t1218 VSS 0.011265f
C6813 VDPWR.n963 VSS 0.028883f
C6814 VDPWR.t1031 VSS 0.005308f
C6815 VDPWR.n964 VSS 0.015733f
C6816 VDPWR.t1127 VSS 0.005308f
C6817 VDPWR.t1277 VSS 0.011265f
C6818 VDPWR.n966 VSS 0.028883f
C6819 VDPWR.t1128 VSS 0.005308f
C6820 VDPWR.n967 VSS 0.015733f
C6821 VDPWR.n968 VSS 0.013309f
C6822 VDPWR.n969 VSS 0.004061f
C6823 VDPWR.n970 VSS 0.002366f
C6824 VDPWR.n971 VSS 0.001509f
C6825 VDPWR.n972 VSS 0.018606f
C6826 VDPWR.t993 VSS 0.005265f
C6827 VDPWR.n973 VSS 0.031863f
C6828 VDPWR.t1231 VSS 0.030423f
C6829 VDPWR.n974 VSS 0.020527f
C6830 VDPWR.n975 VSS 0.008799f
C6831 VDPWR.t992 VSS 0.005265f
C6832 VDPWR.n976 VSS 0.004111f
C6833 VDPWR.n977 VSS 0.004318f
C6834 VDPWR.n978 VSS 0.0024f
C6835 VDPWR.n979 VSS 0.005282f
C6836 VDPWR.n980 VSS 0.002085f
C6837 VDPWR.n981 VSS 0.003719f
C6838 VDPWR.n982 VSS 0.001668f
C6839 VDPWR.t1204 VSS 0.039717f
C6840 VDPWR.t977 VSS 0.005265f
C6841 VDPWR.n983 VSS 0.071594f
C6842 VDPWR.n984 VSS 0.020892f
C6843 VDPWR.t9 VSS 0.001614f
C6844 VDPWR.t599 VSS 0.001614f
C6845 VDPWR.n985 VSS 0.003509f
C6846 VDPWR.t978 VSS 0.005265f
C6847 VDPWR.n986 VSS 0.009272f
C6848 VDPWR.n987 VSS 0.004665f
C6849 VDPWR.t397 VSS 0.006962f
C6850 VDPWR.n988 VSS 0.003471f
C6851 VDPWR.n989 VSS 0.00622f
C6852 VDPWR.t391 VSS 0.001972f
C6853 VDPWR.t393 VSS 0.001972f
C6854 VDPWR.n990 VSS 0.004109f
C6855 VDPWR.t522 VSS 0.001213f
C6856 VDPWR.t823 VSS 7.99e-19
C6857 VDPWR.n991 VSS 0.002095f
C6858 VDPWR.n992 VSS 0.004913f
C6859 VDPWR.t409 VSS 0.001972f
C6860 VDPWR.t401 VSS 0.001972f
C6861 VDPWR.n993 VSS 0.004099f
C6862 VDPWR.t405 VSS 0.001972f
C6863 VDPWR.t395 VSS 0.001972f
C6864 VDPWR.n994 VSS 0.004108f
C6865 VDPWR.n995 VSS 0.007693f
C6866 VDPWR.n996 VSS 0.00622f
C6867 VDPWR.n997 VSS 0.0048f
C6868 VDPWR.t765 VSS 0.003028f
C6869 VDPWR.t34 VSS 0.004145f
C6870 VDPWR.n998 VSS 0.010723f
C6871 VDPWR.t399 VSS 0.001902f
C6872 VDPWR.t403 VSS 0.001972f
C6873 VDPWR.n999 VSS 0.004f
C6874 VDPWR.t407 VSS 0.001972f
C6875 VDPWR.t381 VSS 0.001972f
C6876 VDPWR.n1000 VSS 0.004071f
C6877 VDPWR.n1001 VSS 0.00612f
C6878 VDPWR.n1002 VSS 0.003115f
C6879 VDPWR.n1003 VSS 0.002366f
C6880 VDPWR.n1004 VSS 0.003257f
C6881 VDPWR.n1005 VSS 0.002085f
C6882 VDPWR.n1006 VSS 0.001668f
C6883 VDPWR.n1007 VSS 0.002085f
C6884 VDPWR.n1008 VSS 0.002164f
C6885 VDPWR.t726 VSS 0.002895f
C6886 VDPWR.t379 VSS 0.001972f
C6887 VDPWR.t389 VSS 0.001972f
C6888 VDPWR.n1009 VSS 0.004071f
C6889 VDPWR.t489 VSS 0.001094f
C6890 VDPWR.t669 VSS 0.001094f
C6891 VDPWR.n1010 VSS 0.002291f
C6892 VDPWR.n1011 VSS 0.00706f
C6893 VDPWR.n1012 VSS 0.00311f
C6894 VDPWR.n1013 VSS 0.002164f
C6895 VDPWR.n1014 VSS 0.00133f
C6896 VDPWR.n1015 VSS 0.001651f
C6897 VDPWR.n1016 VSS 0.006255f
C6898 VDPWR.n1017 VSS 0.004382f
C6899 VDPWR.n1018 VSS 0.002366f
C6900 VDPWR.t383 VSS 0.001972f
C6901 VDPWR.t385 VSS 0.001972f
C6902 VDPWR.n1019 VSS 0.004071f
C6903 VDPWR.n1020 VSS 0.006317f
C6904 VDPWR.t1029 VSS 0.054613f
C6905 VDPWR.t991 VSS 0.078929f
C6906 VDPWR.t976 VSS 0.049231f
C6907 VDPWR.t8 VSS 0.023719f
C6908 VDPWR.t598 VSS 0.030495f
C6909 VDPWR.t6 VSS 0.028104f
C6910 VDPWR.t396 VSS 0.020729f
C6911 VDPWR.t390 VSS 0.031891f
C6912 VDPWR.t677 VSS 0.017141f
C6913 VDPWR.t392 VSS 0.01754f
C6914 VDPWR.t521 VSS 0.017141f
C6915 VDPWR.t408 VSS 0.019134f
C6916 VDPWR.t400 VSS 0.01754f
C6917 VDPWR.t822 VSS 0.013354f
C6918 VDPWR.t404 VSS 0.020928f
C6919 VDPWR.t394 VSS 0.020729f
C6920 VDPWR.t764 VSS 0.017141f
C6921 VDPWR.t398 VSS 0.030495f
C6922 VDPWR.t402 VSS 0.019533f
C6923 VDPWR.t33 VSS 0.017141f
C6924 VDPWR.t406 VSS 0.017141f
C6925 VDPWR.t488 VSS 0.017141f
C6926 VDPWR.t380 VSS 0.020729f
C6927 VDPWR.t668 VSS 0.017141f
C6928 VDPWR.t378 VSS 0.019932f
C6929 VDPWR.t725 VSS 0.017141f
C6930 VDPWR.t388 VSS 0.012955f
C6931 VDPWR.t382 VSS 0.014949f
C6932 VDPWR.n1021 VSS 0.005779f
C6933 VDPWR.n1022 VSS 0.002164f
C6934 VDPWR.n1023 VSS 0.002085f
C6935 VDPWR.n1024 VSS 0.003719f
C6936 VDPWR.n1025 VSS 0.001668f
C6937 VDPWR.n1026 VSS 0.002164f
C6938 VDPWR.n1027 VSS 0.00311f
C6939 VDPWR.t1236 VSS 0.021971f
C6940 VDPWR.n1028 VSS 0.007544f
C6941 VDPWR.t78 VSS 0.008077f
C6942 VDPWR.n1029 VSS 0.011929f
C6943 VDPWR.n1030 VSS 0.00622f
C6944 VDPWR.t604 VSS 0.001902f
C6945 VDPWR.t223 VSS 0.001902f
C6946 VDPWR.n1031 VSS 0.004259f
C6947 VDPWR.t225 VSS 0.002994f
C6948 VDPWR.n1032 VSS 0.00677f
C6949 VDPWR.n1033 VSS 0.005646f
C6950 VDPWR.n1034 VSS 0.001161f
C6951 VDPWR.n1035 VSS 0.003115f
C6952 VDPWR.n1036 VSS 0.002918f
C6953 VDPWR.n1037 VSS 0.003043f
C6954 VDPWR.n1038 VSS 0.001668f
C6955 VDPWR.n1039 VSS 0.003626f
C6956 VDPWR.n1040 VSS 0.003227f
C6957 VDPWR.n1041 VSS 0.003115f
C6958 VDPWR.t720 VSS 0.001213f
C6959 VDPWR.t601 VSS -7.69e-19
C6960 VDPWR.n1042 VSS 0.007741f
C6961 VDPWR.n1043 VSS 0.005961f
C6962 VDPWR.t771 VSS 0.002933f
C6963 VDPWR.n1044 VSS 0.001425f
C6964 VDPWR.n1045 VSS 0.001216f
C6965 VDPWR.t387 VSS 0.001972f
C6966 VDPWR.t496 VSS 0.001972f
C6967 VDPWR.n1046 VSS 0.004306f
C6968 VDPWR.n1047 VSS 0.007138f
C6969 VDPWR.n1048 VSS 0.001799f
C6970 VDPWR.n1049 VSS 0.004665f
C6971 VDPWR.n1050 VSS 0.003955f
C6972 VDPWR.n1051 VSS 0.00213f
C6973 VDPWR.n1052 VSS 0.001281f
C6974 VDPWR.t202 VSS 0.001614f
C6975 VDPWR.t269 VSS 0.001614f
C6976 VDPWR.n1053 VSS 0.003585f
C6977 VDPWR.t740 VSS 0.001972f
C6978 VDPWR.t744 VSS 0.001972f
C6979 VDPWR.n1054 VSS 0.004301f
C6980 VDPWR.n1055 VSS 0.015277f
C6981 VDPWR.n1056 VSS 0.005646f
C6982 VDPWR.n1057 VSS 0.004665f
C6983 VDPWR.n1058 VSS 0.00213f
C6984 VDPWR.t742 VSS 0.007366f
C6985 VDPWR.n1059 VSS 0.009322f
C6986 VDPWR.t538 VSS 0.001217f
C6987 VDPWR.t236 VSS 0.001217f
C6988 VDPWR.n1060 VSS 0.002534f
C6989 VDPWR.n1061 VSS 0.006799f
C6990 VDPWR.n1062 VSS 0.002164f
C6991 VDPWR.n1063 VSS 0.005612f
C6992 VDPWR.n1064 VSS 0.005882f
C6993 VDPWR.n1065 VSS 0.006044f
C6994 VDPWR.t593 VSS 0.002319f
C6995 VDPWR.t365 VSS 0.002808f
C6996 VDPWR.n1066 VSS 0.006664f
C6997 VDPWR.n1067 VSS 0.004035f
C6998 VDPWR.n1068 VSS 0.001798f
C6999 VDPWR.n1069 VSS 0.002164f
C7000 VDPWR.n1070 VSS 0.002164f
C7001 VDPWR.n1071 VSS 0.00311f
C7002 VDPWR.n1072 VSS 0.002085f
C7003 VDPWR.n1073 VSS 0.002085f
C7004 VDPWR.n1074 VSS 0.001668f
C7005 VDPWR.n1075 VSS 0.003719f
C7006 VDPWR.n1077 VSS 0.003719f
C7007 VDPWR.n1078 VSS 0.003626f
C7008 VDPWR.n1079 VSS 0.003227f
C7009 VDPWR.n1080 VSS 0.002085f
C7010 VDPWR.n1081 VSS 0.002231f
C7011 VDPWR.n1082 VSS 0.002164f
C7012 VDPWR.n1083 VSS 0.002138f
C7013 VDPWR.t447 VSS 0.002942f
C7014 VDPWR.t780 VSS 0.001426f
C7015 VDPWR.n1084 VSS 0.00599f
C7016 VDPWR.t734 VSS 0.003026f
C7017 VDPWR.n1085 VSS 0.008534f
C7018 VDPWR.n1086 VSS 0.004594f
C7019 VDPWR.n1087 VSS 0.001688f
C7020 VDPWR.n1088 VSS 0.004124f
C7021 VDPWR.n1089 VSS 0.004665f
C7022 VDPWR.n1090 VSS 0.00213f
C7023 VDPWR.n1091 VSS 0.001976f
C7024 VDPWR.t732 VSS 0.001449f
C7025 VDPWR.t411 VSS 0.002395f
C7026 VDPWR.n1092 VSS 0.006638f
C7027 VDPWR.n1093 VSS 0.008136f
C7028 VDPWR.n1094 VSS 8.26e-19
C7029 VDPWR.n1095 VSS 0.00622f
C7030 VDPWR.n1096 VSS 0.00622f
C7031 VDPWR.n1097 VSS 0.00622f
C7032 VDPWR.t570 VSS 0.007766f
C7033 VDPWR.n1098 VSS 0.007356f
C7034 VDPWR.n1099 VSS 0.005459f
C7035 VDPWR.n1100 VSS 0.001197f
C7036 VDPWR.n1101 VSS 0.001245f
C7037 VDPWR.n1102 VSS 0.004665f
C7038 VDPWR.n1103 VSS 0.00311f
C7039 VDPWR.n1104 VSS 0.001151f
C7040 VDPWR.t200 VSS 0.004499f
C7041 VDPWR.t694 VSS 0.001094f
C7042 VDPWR.n1105 VSS 0.003115f
C7043 VDPWR.n1106 VSS 0.004141f
C7044 VDPWR.n1107 VSS 0.00284f
C7045 VDPWR.n1108 VSS 0.003175f
C7046 VDPWR.n1109 VSS 0.002366f
C7047 VDPWR.n1110 VSS 0.002366f
C7048 VDPWR.n1111 VSS 0.002085f
C7049 VDPWR.n1112 VSS 0.003595f
C7050 VDPWR.n1113 VSS 0.003257f
C7051 VDPWR.n1114 VSS 0.002912f
C7052 VDPWR.n1115 VSS 0.002299f
C7053 VDPWR.n1116 VSS 0.003911f
C7054 VDPWR.t907 VSS 0.005265f
C7055 VDPWR.n1117 VSS 0.00519f
C7056 VDPWR.n1118 VSS 0.019873f
C7057 VDPWR.n1119 VSS 0.012246f
C7058 VDPWR.t96 VSS 0.001213f
C7059 VDPWR.t820 VSS 7.99e-19
C7060 VDPWR.n1120 VSS 0.00207f
C7061 VDPWR.t908 VSS 0.005265f
C7062 VDPWR.n1121 VSS 0.009095f
C7063 VDPWR.n1122 VSS 0.011757f
C7064 VDPWR.n1123 VSS 0.008342f
C7065 VDPWR.n1124 VSS 0.002164f
C7066 VDPWR.n1125 VSS 0.00311f
C7067 VDPWR.n1126 VSS 0.002085f
C7068 VDPWR.n1127 VSS 0.001668f
C7069 VDPWR.n1128 VSS 0.003719f
C7070 VDPWR.n1129 VSS 0.003595f
C7071 VDPWR.n1130 VSS 0.003257f
C7072 VDPWR.n1131 VSS 5.79e-19
C7073 VDPWR.n1132 VSS 0.002366f
C7074 VDPWR.n1133 VSS 0.003194f
C7075 VDPWR.n1134 VSS 0.00622f
C7076 VDPWR.t91 VSS 0.001902f
C7077 VDPWR.t566 VSS 0.001902f
C7078 VDPWR.n1135 VSS 0.004259f
C7079 VDPWR.t1120 VSS 0.005792f
C7080 VDPWR.n1136 VSS 9.21e-19
C7081 VDPWR.n1137 VSS 0.008045f
C7082 VDPWR.t93 VSS 0.002968f
C7083 VDPWR.t1178 VSS 0.076721f
C7084 VDPWR.n1138 VSS 0.035835f
C7085 VDPWR.n1139 VSS 0.00622f
C7086 VDPWR.t70 VSS 0.001426f
C7087 VDPWR.t72 VSS 0.002942f
C7088 VDPWR.n1140 VSS 0.00599f
C7089 VDPWR.n1141 VSS 0.007472f
C7090 VDPWR.n1142 VSS 0.004936f
C7091 VDPWR.n1143 VSS 0.007585f
C7092 VDPWR.n1144 VSS 0.003115f
C7093 VDPWR.n1145 VSS 0.002231f
C7094 VDPWR.n1146 VSS 0.003257f
C7095 VDPWR.n1147 VSS 0.002085f
C7096 VDPWR.n1148 VSS 0.001668f
C7097 VDPWR.n1149 VSS 0.002085f
C7098 VDPWR.n1150 VSS 0.00622f
C7099 VDPWR.t579 VSS 0.00291f
C7100 VDPWR.t1121 VSS 0.005792f
C7101 VDPWR.n1151 VSS 0.0045f
C7102 VDPWR.n1152 VSS 0.002164f
C7103 VDPWR.n1153 VSS 0.00311f
C7104 VDPWR.n1154 VSS 0.001589f
C7105 VDPWR.n1155 VSS 9.74e-19
C7106 VDPWR.n1156 VSS 0.005891f
C7107 VDPWR.t562 VSS 0.001217f
C7108 VDPWR.t59 VSS 0.001217f
C7109 VDPWR.n1157 VSS 0.002507f
C7110 VDPWR.n1158 VSS 0.004176f
C7111 VDPWR.n1159 VSS 0.003651f
C7112 VDPWR.t1187 VSS 0.076721f
C7113 VDPWR.t638 VSS 0.007445f
C7114 VDPWR.n1160 VSS 0.012566f
C7115 VDPWR.n1161 VSS 0.035579f
C7116 VDPWR.t868 VSS 0.005265f
C7117 VDPWR.n1162 VSS 0.012091f
C7118 VDPWR.n1163 VSS 0.00622f
C7119 VDPWR.t1247 VSS 0.030953f
C7120 VDPWR.n1164 VSS 0.021249f
C7121 VDPWR.n1165 VSS 7.78e-19
C7122 VDPWR.n1166 VSS 0.002085f
C7123 VDPWR.n1167 VSS 0.248273f
C7124 VDPWR.n1168 VSS 0.003595f
C7125 VDPWR.n1169 VSS 0.003257f
C7126 VDPWR.n1170 VSS 0.003719f
C7127 VDPWR.n1171 VSS 0.002085f
C7128 VDPWR.n1172 VSS 0.002164f
C7129 VDPWR.n1173 VSS 0.007742f
C7130 VDPWR.t989 VSS 0.005308f
C7131 VDPWR.t1234 VSS 0.011265f
C7132 VDPWR.n1175 VSS 0.028883f
C7133 VDPWR.t990 VSS 0.005308f
C7134 VDPWR.n1176 VSS 0.015733f
C7135 VDPWR.n1177 VSS 0.00622f
C7136 VDPWR.t1284 VSS 0.021971f
C7137 VDPWR.n1178 VSS 0.004233f
C7138 VDPWR.n1179 VSS 0.00622f
C7139 VDPWR.t288 VSS 0.001972f
C7140 VDPWR.t310 VSS 0.001972f
C7141 VDPWR.n1180 VSS 0.004071f
C7142 VDPWR.t1230 VSS 0.076721f
C7143 VDPWR.n1181 VSS 0.035825f
C7144 VDPWR.n1182 VSS 0.00622f
C7145 VDPWR.t318 VSS 0.001972f
C7146 VDPWR.t290 VSS 0.001972f
C7147 VDPWR.n1183 VSS 0.004071f
C7148 VDPWR.t995 VSS 0.005792f
C7149 VDPWR.n1184 VSS 0.004533f
C7150 VDPWR.n1185 VSS 0.00254f
C7151 VDPWR.t296 VSS 0.001972f
C7152 VDPWR.t312 VSS 0.001902f
C7153 VDPWR.n1186 VSS 0.004012f
C7154 VDPWR.t1037 VSS 0.005792f
C7155 VDPWR.n1187 VSS 0.004533f
C7156 VDPWR.n1188 VSS 0.002164f
C7157 VDPWR.n1189 VSS 0.001668f
C7158 VDPWR.n1190 VSS 0.003719f
C7159 VDPWR.n1191 VSS 0.245208f
C7160 VDPWR.n1193 VSS 0.003719f
C7161 VDPWR.n1194 VSS 0.003115f
C7162 VDPWR.n1195 VSS 0.001668f
C7163 VDPWR.t308 VSS 0.001972f
C7164 VDPWR.t298 VSS 0.001972f
C7165 VDPWR.n1196 VSS 0.004071f
C7166 VDPWR.n1197 VSS 0.009136f
C7167 VDPWR.n1198 VSS 0.00622f
C7168 VDPWR.t300 VSS 0.001972f
C7169 VDPWR.t304 VSS 0.001972f
C7170 VDPWR.n1199 VSS 0.004071f
C7171 VDPWR.n1200 VSS 0.004726f
C7172 VDPWR.n1201 VSS 0.00622f
C7173 VDPWR.t500 VSS 0.001972f
C7174 VDPWR.t498 VSS 0.001972f
C7175 VDPWR.n1202 VSS 0.004238f
C7176 VDPWR.t1036 VSS 0.005792f
C7177 VDPWR.n1203 VSS 0.004372f
C7178 VDPWR.t1143 VSS 0.005792f
C7179 VDPWR.n1204 VSS 0.0045f
C7180 VDPWR.t988 VSS 0.055011f
C7181 VDPWR.t1101 VSS 0.089892f
C7182 VDPWR.t313 VSS 0.073348f
C7183 VDPWR.t994 VSS 0.017141f
C7184 VDPWR.t309 VSS 0.019932f
C7185 VDPWR.t287 VSS 0.034282f
C7186 VDPWR.t315 VSS 0.034282f
C7187 VDPWR.t291 VSS 0.034282f
C7188 VDPWR.t289 VSS 0.034282f
C7189 VDPWR.t317 VSS 0.034282f
C7190 VDPWR.t311 VSS 0.027306f
C7191 VDPWR.t295 VSS 0.023918f
C7192 VDPWR.t305 VSS 0.034282f
C7193 VDPWR.t301 VSS 0.034282f
C7194 VDPWR.t297 VSS 0.034282f
C7195 VDPWR.t307 VSS 0.034282f
C7196 VDPWR.t303 VSS 0.028901f
C7197 VDPWR.t1035 VSS 0.017141f
C7198 VDPWR.t299 VSS 0.022523f
C7199 VDPWR.t293 VSS 0.034282f
C7200 VDPWR.t491 VSS 0.034282f
C7201 VDPWR.t497 VSS 0.034282f
C7202 VDPWR.t499 VSS 0.034282f
C7203 VDPWR.t493 VSS 0.023519f
C7204 VDPWR.n1205 VSS 0.039521f
C7205 VDPWR.t1134 VSS 0.005265f
C7206 VDPWR.n1206 VSS 0.012091f
C7207 VDPWR.n1207 VSS 0.00311f
C7208 VDPWR.n1208 VSS 0.002085f
C7209 VDPWR.n1209 VSS 0.003719f
C7210 VDPWR.n1210 VSS 0.245208f
C7211 VDPWR.n1211 VSS 0.003719f
C7212 VDPWR.n1212 VSS 0.002912f
C7213 VDPWR.n1213 VSS 0.001668f
C7214 VDPWR.n1214 VSS 0.001668f
C7215 VDPWR.n1215 VSS 0.002085f
C7216 VDPWR.n1216 VSS 0.00311f
C7217 VDPWR.t1273 VSS 0.021971f
C7218 VDPWR.n1217 VSS 0.007471f
C7219 VDPWR.n1218 VSS 0.00622f
C7220 VDPWR.t812 VSS 0.006928f
C7221 VDPWR.t1173 VSS 0.076721f
C7222 VDPWR.t798 VSS 0.001972f
C7223 VDPWR.t808 VSS 0.001972f
C7224 VDPWR.n1219 VSS 0.004071f
C7225 VDPWR.n1220 VSS 0.009034f
C7226 VDPWR.n1221 VSS 0.005646f
C7227 VDPWR.t800 VSS 0.001972f
C7228 VDPWR.t802 VSS 0.001972f
C7229 VDPWR.n1222 VSS 0.004071f
C7230 VDPWR.t839 VSS 0.005792f
C7231 VDPWR.n1223 VSS 0.003974f
C7232 VDPWR.n1224 VSS 0.00622f
C7233 VDPWR.t788 VSS 0.001972f
C7234 VDPWR.t792 VSS 0.001902f
C7235 VDPWR.n1225 VSS 0.004f
C7236 VDPWR.n1226 VSS 0.006272f
C7237 VDPWR.n1227 VSS 0.002164f
C7238 VDPWR.n1228 VSS 0.002085f
C7239 VDPWR.n1229 VSS 0.003719f
C7240 VDPWR.n1230 VSS 0.245208f
C7241 VDPWR.n1231 VSS 0.003719f
C7242 VDPWR.n1232 VSS 0.003115f
C7243 VDPWR.n1233 VSS 0.001668f
C7244 VDPWR.n1234 VSS 0.002164f
C7245 VDPWR.n1235 VSS 0.002231f
C7246 VDPWR.n1236 VSS 0.001668f
C7247 VDPWR.n1237 VSS 0.002085f
C7248 VDPWR.n1238 VSS 0.003043f
C7249 VDPWR.t818 VSS 0.001972f
C7250 VDPWR.t790 VSS 0.001972f
C7251 VDPWR.n1239 VSS 0.004071f
C7252 VDPWR.t1283 VSS 0.076721f
C7253 VDPWR.t804 VSS 0.001972f
C7254 VDPWR.t814 VSS 0.001972f
C7255 VDPWR.n1240 VSS 0.004071f
C7256 VDPWR.n1241 VSS 0.009136f
C7257 VDPWR.n1242 VSS 0.00622f
C7258 VDPWR.t474 VSS 0.001972f
C7259 VDPWR.t810 VSS 0.001972f
C7260 VDPWR.n1243 VSS 0.004228f
C7261 VDPWR.n1244 VSS 0.006119f
C7262 VDPWR.t472 VSS 0.007287f
C7263 VDPWR.n1245 VSS 0.007275f
C7264 VDPWR.n1246 VSS 0.006165f
C7265 VDPWR.t1240 VSS 0.0218f
C7266 VDPWR.n1247 VSS 0.010829f
C7267 VDPWR.n1248 VSS 0.004163f
C7268 VDPWR.t968 VSS 0.005265f
C7269 VDPWR.n1249 VSS 0.002806f
C7270 VDPWR.t930 VSS 0.06996f
C7271 VDPWR.t1083 VSS 0.058599f
C7272 VDPWR.t961 VSS 0.097466f
C7273 VDPWR.t897 VSS 0.067568f
C7274 VDPWR.t1045 VSS 0.115803f
C7275 VDPWR.t1109 VSS 0.104242f
C7276 VDPWR.t1132 VSS 0.067568f
C7277 VDPWR.t1141 VSS 0.042853f
C7278 VDPWR.t811 VSS 0.051623f
C7279 VDPWR.t807 VSS 0.034282f
C7280 VDPWR.t797 VSS 0.034282f
C7281 VDPWR.t801 VSS 0.034282f
C7282 VDPWR.t799 VSS 0.023719f
C7283 VDPWR.t805 VSS 0.027705f
C7284 VDPWR.t795 VSS 0.034282f
C7285 VDPWR.t791 VSS 0.034083f
C7286 VDPWR.t787 VSS 0.034083f
C7287 VDPWR.t815 VSS 0.034282f
C7288 VDPWR.t793 VSS 0.025313f
C7289 VDPWR.t837 VSS 0.017141f
C7290 VDPWR.t789 VSS 0.02611f
C7291 VDPWR.t817 VSS 0.034282f
C7292 VDPWR.t813 VSS 0.034282f
C7293 VDPWR.t803 VSS 0.034282f
C7294 VDPWR.t809 VSS 0.034282f
C7295 VDPWR.t473 VSS 0.034282f
C7296 VDPWR.t475 VSS 0.021127f
C7297 VDPWR.t62 VSS 0.030296f
C7298 VDPWR.t471 VSS 0.017739f
C7299 VDPWR.t967 VSS 0.006378f
C7300 VDPWR.n1250 VSS 0.039521f
C7301 VDPWR.n1251 VSS 0.018083f
C7302 VDPWR.n1252 VSS 0.003115f
C7303 VDPWR.n1253 VSS 0.013477f
C7304 VDPWR.n1254 VSS 0.002164f
C7305 VDPWR.n1255 VSS 0.001668f
C7306 VDPWR.n1256 VSS 0.003719f
C7307 VDPWR.n1257 VSS 0.245208f
C7308 VDPWR.n1258 VSS 0.003595f
C7309 VDPWR.n1259 VSS 0.003719f
C7310 VDPWR.n1260 VSS 0.003115f
C7311 VDPWR.n1261 VSS 0.001668f
C7312 VDPWR.n1262 VSS 0.002164f
C7313 VDPWR.n1263 VSS 0.002164f
C7314 VDPWR.n1264 VSS 0.003257f
C7315 VDPWR.n1265 VSS 0.003115f
C7316 VDPWR.t1224 VSS 0.076721f
C7317 VDPWR.n1266 VSS 0.013477f
C7318 VDPWR.n1267 VSS 0.005646f
C7319 VDPWR.t984 VSS 0.005792f
C7320 VDPWR.n1268 VSS 0.007319f
C7321 VDPWR.n1269 VSS 0.00622f
C7322 VDPWR.n1270 VSS 0.009235f
C7323 VDPWR.n1271 VSS 0.00622f
C7324 VDPWR.t1210 VSS 0.076721f
C7325 VDPWR.n1272 VSS 0.042898f
C7326 VDPWR.n1273 VSS 0.003043f
C7327 VDPWR.n1274 VSS 0.002085f
C7328 VDPWR.n1275 VSS 0.003719f
C7329 VDPWR.n1276 VSS 0.251293f
C7330 VDPWR.n1277 VSS 0.003595f
C7331 VDPWR.n1278 VSS 0.003719f
C7332 VDPWR.n1279 VSS 0.002777f
C7333 VDPWR.n1280 VSS 0.001668f
C7334 VDPWR.n1281 VSS 0.00311f
C7335 VDPWR.t1199 VSS 0.038277f
C7336 VDPWR.n1282 VSS 0.028878f
C7337 VDPWR.t986 VSS 0.005792f
C7338 VDPWR.t1123 VSS 0.005265f
C7339 VDPWR.n1283 VSS 0.012671f
C7340 VDPWR.t1095 VSS 0.005308f
C7341 VDPWR.t1221 VSS 0.011265f
C7342 VDPWR.n1285 VSS 0.028883f
C7343 VDPWR.t1096 VSS 0.005308f
C7344 VDPWR.n1286 VSS 0.015733f
C7345 VDPWR.t942 VSS 0.005308f
C7346 VDPWR.t1266 VSS 0.011265f
C7347 VDPWR.n1288 VSS 0.028883f
C7348 VDPWR.t943 VSS 0.005308f
C7349 VDPWR.n1289 VSS 0.015733f
C7350 VDPWR.n1290 VSS 0.012962f
C7351 VDPWR.t925 VSS 0.005308f
C7352 VDPWR.t1227 VSS 0.011265f
C7353 VDPWR.n1292 VSS 0.028883f
C7354 VDPWR.t926 VSS 0.005308f
C7355 VDPWR.n1293 VSS 0.015733f
C7356 VDPWR.n1294 VSS 0.004061f
C7357 VDPWR.n1295 VSS 0.005237f
C7358 VDPWR.t1107 VSS 0.005308f
C7359 VDPWR.t1197 VSS 0.011265f
C7360 VDPWR.n1297 VSS 0.028883f
C7361 VDPWR.t1108 VSS 0.005308f
C7362 VDPWR.n1298 VSS 0.015733f
C7363 VDPWR.n1299 VSS 0.014221f
C7364 VDPWR.n1300 VSS 0.003497f
C7365 VDPWR.n1301 VSS 0.004059f
C7366 VDPWR.n1302 VSS 0.004665f
C7367 VDPWR.n1303 VSS 0.003719f
C7368 VDPWR.n1304 VSS 0.016116f
C7369 VDPWR.n1305 VSS 0.027133f
C7370 VDPWR.t1246 VSS 0.076721f
C7371 VDPWR.n1306 VSS 0.042898f
C7372 VDPWR.n1307 VSS 0.00622f
C7373 VDPWR.t1124 VSS 0.005265f
C7374 VDPWR.n1308 VSS 0.012091f
C7375 VDPWR.t874 VSS 0.005792f
C7376 VDPWR.n1309 VSS 0.007319f
C7377 VDPWR.n1310 VSS 0.00622f
C7378 VDPWR.t1286 VSS 0.078173f
C7379 VDPWR.n1311 VSS 0.036257f
C7380 VDPWR.n1312 VSS 0.00622f
C7381 VDPWR.n1313 VSS 0.010328f
C7382 VDPWR.n1314 VSS 0.002164f
C7383 VDPWR.n1315 VSS 0.002085f
C7384 VDPWR.n1316 VSS 0.001668f
C7385 VDPWR.n1317 VSS 0.001668f
C7386 VDPWR.n1318 VSS 0.002085f
C7387 VDPWR.n1319 VSS 0.002164f
C7388 VDPWR.t1260 VSS 0.076721f
C7389 VDPWR.n1320 VSS 0.038654f
C7390 VDPWR.n1321 VSS 0.009888f
C7391 VDPWR.n1322 VSS 0.002907f
C7392 VDPWR.n1323 VSS 0.002085f
C7393 VDPWR.n1324 VSS 0.002366f
C7394 VDPWR.n1325 VSS 0.00311f
C7395 VDPWR.n1326 VSS 0.002164f
C7396 VDPWR.n1327 VSS 0.013477f
C7397 VDPWR.n1328 VSS 0.013038f
C7398 VDPWR.t875 VSS 0.005792f
C7399 VDPWR.n1329 VSS 0.007319f
C7400 VDPWR.t941 VSS 0.06996f
C7401 VDPWR.t924 VSS 0.076737f
C7402 VDPWR.t1122 VSS 0.115803f
C7403 VDPWR.t985 VSS 0.067568f
C7404 VDPWR.t873 VSS 0.115803f
C7405 VDPWR.t955 VSS 0.104242f
C7406 VDPWR.n1330 VSS 0.039521f
C7407 VDPWR.n1331 VSS 0.006604f
C7408 VDPWR.n1332 VSS 0.00449f
C7409 VDPWR.t1158 VSS 0.00581f
C7410 VDPWR.t1016 VSS 0.005792f
C7411 VDPWR.n1333 VSS 0.007319f
C7412 VDPWR.n1334 VSS 0.00622f
C7413 VDPWR.t1175 VSS 0.076721f
C7414 VDPWR.t1235 VSS 0.076721f
C7415 VDPWR.n1335 VSS 0.038654f
C7416 VDPWR.n1336 VSS 0.002164f
C7417 VDPWR.n1337 VSS 0.002085f
C7418 VDPWR.n1338 VSS 0.003719f
C7419 VDPWR.n1339 VSS 0.248927f
C7420 VDPWR.n1340 VSS 0.003719f
C7421 VDPWR.n1341 VSS 0.002085f
C7422 VDPWR.n1342 VSS 0.002164f
C7423 VDPWR.n1343 VSS 0.00622f
C7424 VDPWR.n1344 VSS 0.009888f
C7425 VDPWR.n1345 VSS 0.00311f
C7426 VDPWR.n1346 VSS 0.002231f
C7427 VDPWR.n1347 VSS 0.001668f
C7428 VDPWR.n1348 VSS 0.001668f
C7429 VDPWR.n1349 VSS 0.002085f
C7430 VDPWR.n1350 VSS 0.003043f
C7431 VDPWR.n1351 VSS 0.002164f
C7432 VDPWR.n1352 VSS 0.013477f
C7433 VDPWR.n1353 VSS 0.013477f
C7434 VDPWR.t1017 VSS 0.005811f
C7435 VDPWR.n1354 VSS 0.011885f
C7436 VDPWR.t1056 VSS 0.00581f
C7437 VDPWR.t980 VSS 0.005792f
C7438 VDPWR.n1355 VSS 0.007319f
C7439 VDPWR.n1356 VSS 0.00622f
C7440 VDPWR.t1223 VSS 0.076721f
C7441 VDPWR.t1177 VSS 0.076721f
C7442 VDPWR.n1357 VSS 0.038654f
C7443 VDPWR.n1358 VSS 0.00622f
C7444 VDPWR.n1359 VSS 0.013477f
C7445 VDPWR.n1360 VSS 0.002366f
C7446 VDPWR.n1361 VSS 0.002085f
C7447 VDPWR.n1362 VSS 0.003719f
C7448 VDPWR.n1363 VSS 0.250504f
C7449 VDPWR.n1364 VSS 0.003719f
C7450 VDPWR.n1365 VSS 0.002085f
C7451 VDPWR.n1366 VSS 0.002164f
C7452 VDPWR.t1129 VSS 0.036674f
C7453 VDPWR.t1157 VSS 0.115803f
C7454 VDPWR.t1015 VSS 0.104242f
C7455 VDPWR.t1055 VSS 0.115803f
C7456 VDPWR.t979 VSS 0.104242f
C7457 VDPWR.t1007 VSS 0.055011f
C7458 VDPWR.t1018 VSS 0.073747f
C7459 VDPWR.t209 VSS 0.014949f
C7460 VDPWR.t0 VSS 0.016743f
C7461 VDPWR.t444 VSS 0.016743f
C7462 VDPWR.t607 VSS 0.016743f
C7463 VDPWR.t440 VSS 0.033087f
C7464 VDPWR.t205 VSS 0.025512f
C7465 VDPWR.t2 VSS 0.031492f
C7466 VDPWR.t370 VSS 0.028701f
C7467 VDPWR.t10 VSS 0.016743f
C7468 VDPWR.t526 VSS 0.02611f
C7469 VDPWR.t371 VSS 0.029897f
C7470 VDPWR.t755 VSS 0.046839f
C7471 VDPWR.t525 VSS 0.039465f
C7472 VDPWR.t369 VSS 0.035877f
C7473 VDPWR.t281 VSS 0.03488f
C7474 VDPWR.t858 VSS 0.037471f
C7475 VDPWR.t523 VSS 0.036276f
C7476 VDPWR.t244 VSS 0.022921f
C7477 VDPWR.t1149 VSS 0.055011f
C7478 VDPWR.n1367 VSS 0.039919f
C7479 VDPWR.n1368 VSS 0.002164f
C7480 VDPWR.n1369 VSS 0.001668f
C7481 VDPWR.n1370 VSS 0.001668f
C7482 VDPWR.n1371 VSS 0.002085f
C7483 VDPWR.n1372 VSS 0.00311f
C7484 VDPWR.n1373 VSS 0.00311f
C7485 VDPWR.n1374 VSS 0.002164f
C7486 VDPWR.n1375 VSS 0.013038f
C7487 VDPWR.t1057 VSS 0.005792f
C7488 VDPWR.n1376 VSS 0.007319f
C7489 VDPWR.n1377 VSS 0.006356f
C7490 VDPWR.t981 VSS 0.005814f
C7491 VDPWR.n1378 VSS 0.003868f
C7492 VDPWR.t1181 VSS 0.02239f
C7493 VDPWR.t1150 VSS 0.005265f
C7494 VDPWR.n1379 VSS 0.008287f
C7495 VDPWR.n1380 VSS 0.00847f
C7496 VDPWR.t1151 VSS 0.00534f
C7497 VDPWR.n1381 VSS 0.037596f
C7498 VDPWR.n1382 VSS 0.013535f
C7499 VDPWR.t859 VSS 0.00581f
C7500 VDPWR.n1383 VSS 0.017249f
C7501 VDPWR.t1219 VSS 0.076721f
C7502 VDPWR.t245 VSS 0.001217f
C7503 VDPWR.t524 VSS 0.001217f
C7504 VDPWR.n1384 VSS 0.002507f
C7505 VDPWR.n1385 VSS 0.007542f
C7506 VDPWR.n1386 VSS 0.00622f
C7507 VDPWR.t282 VSS 0.002909f
C7508 VDPWR.n1387 VSS 0.00752f
C7509 VDPWR.n1388 VSS 0.00784f
C7510 VDPWR.n1389 VSS 0.002164f
C7511 VDPWR.n1390 VSS 0.002085f
C7512 VDPWR.n1391 VSS 0.003719f
C7513 VDPWR.n1392 VSS 0.256026f
C7514 VDPWR.n1393 VSS 0.003719f
C7515 VDPWR.n1394 VSS 0.002085f
C7516 VDPWR.n1395 VSS 0.00622f
C7517 VDPWR.t860 VSS 0.005792f
C7518 VDPWR.n1396 VSS 0.002412f
C7519 VDPWR.n1397 VSS 0.003043f
C7520 VDPWR.n1398 VSS 0.001668f
C7521 VDPWR.n1399 VSS 0.001668f
C7522 VDPWR.n1400 VSS 0.002085f
C7523 VDPWR.n1401 VSS 0.002231f
C7524 VDPWR.t756 VSS 0.002942f
C7525 VDPWR.t372 VSS 0.001426f
C7526 VDPWR.n1402 VSS 0.00599f
C7527 VDPWR.n1403 VSS 0.007216f
C7528 VDPWR.n1404 VSS 0.006008f
C7529 VDPWR.n1405 VSS 0.002164f
C7530 VDPWR.n1406 VSS 0.00311f
C7531 VDPWR.n1407 VSS 0.001589f
C7532 VDPWR.n1408 VSS 0.003253f
C7533 VDPWR.t206 VSS 0.006676f
C7534 VDPWR.n1409 VSS 0.00357f
C7535 VDPWR.n1410 VSS 0.00622f
C7536 VDPWR.t3 VSS 0.002994f
C7537 VDPWR.t441 VSS 0.001902f
C7538 VDPWR.t445 VSS 0.001902f
C7539 VDPWR.n1411 VSS 0.004125f
C7540 VDPWR.t608 VSS 0.001902f
C7541 VDPWR.t1 VSS 0.001902f
C7542 VDPWR.n1412 VSS 0.004259f
C7543 VDPWR.n1413 VSS 0.002203f
C7544 VDPWR.t1152 VSS 0.005265f
C7545 VDPWR.t1166 VSS 0.022165f
C7546 VDPWR.n1415 VSS 0.038508f
C7547 VDPWR.t1153 VSS 0.005265f
C7548 VDPWR.n1416 VSS 0.022096f
C7549 VDPWR.n1417 VSS 7.78e-19
C7550 VDPWR.n1418 VSS 0.008248f
C7551 VDPWR.t1019 VSS 0.005265f
C7552 VDPWR.t1237 VSS 0.022165f
C7553 VDPWR.n1420 VSS 0.038508f
C7554 VDPWR.t1020 VSS 0.005265f
C7555 VDPWR.n1421 VSS 0.022096f
C7556 VDPWR.t1147 VSS 0.005308f
C7557 VDPWR.t1220 VSS 0.011265f
C7558 VDPWR.n1423 VSS 0.028883f
C7559 VDPWR.t1148 VSS 0.005308f
C7560 VDPWR.n1424 VSS 0.015733f
C7561 VDPWR.n1425 VSS 0.002164f
C7562 VDPWR.n1426 VSS 0.002164f
C7563 VDPWR.t1008 VSS 0.005308f
C7564 VDPWR.t1242 VSS 0.011265f
C7565 VDPWR.n1428 VSS 0.028883f
C7566 VDPWR.t1009 VSS 0.005308f
C7567 VDPWR.n1429 VSS 0.015733f
C7568 VDPWR.n1430 VSS 0.002231f
C7569 VDPWR.n1431 VSS 0.002085f
C7570 VDPWR.n1432 VSS 0.003595f
C7571 VDPWR.n1433 VSS 0.003257f
C7572 VDPWR.n1434 VSS 0.003719f
C7573 VDPWR.n1435 VSS 0.002085f
C7574 VDPWR.n1436 VSS 0.002164f
C7575 VDPWR.n1437 VSS 0.004785f
C7576 VDPWR.t856 VSS 0.005308f
C7577 VDPWR.t1257 VSS 0.011265f
C7578 VDPWR.n1439 VSS 0.028883f
C7579 VDPWR.t857 VSS 0.005308f
C7580 VDPWR.n1440 VSS 0.015733f
C7581 VDPWR.n1441 VSS 0.00622f
C7582 VDPWR.n1442 VSS 0.013477f
C7583 VDPWR.n1443 VSS 0.00622f
C7584 VDPWR.t1195 VSS 0.076721f
C7585 VDPWR.t1170 VSS 0.076721f
C7586 VDPWR.n1444 VSS 0.07057f
C7587 VDPWR.n1445 VSS 0.00622f
C7588 VDPWR.t865 VSS 0.005792f
C7589 VDPWR.t1013 VSS 0.005792f
C7590 VDPWR.n1446 VSS 0.007899f
C7591 VDPWR.t1060 VSS 0.005792f
C7592 VDPWR.n1447 VSS 0.0045f
C7593 VDPWR.n1448 VSS 0.00311f
C7594 VDPWR.n1449 VSS 0.002085f
C7595 VDPWR.n1450 VSS 0.003719f
C7596 VDPWR.n1451 VSS 0.001668f
C7597 VDPWR.n1452 VSS 0.002468f
C7598 VDPWR.t68 VSS 0.001614f
C7599 VDPWR.t204 VSS 0.001614f
C7600 VDPWR.n1453 VSS 0.003509f
C7601 VDPWR.n1454 VSS 0.009456f
C7602 VDPWR.n1455 VSS 0.00622f
C7603 VDPWR.n1456 VSS 0.016116f
C7604 VDPWR.n1457 VSS 0.00622f
C7605 VDPWR.t1171 VSS 0.038955f
C7606 VDPWR.t1059 VSS 0.005792f
C7607 VDPWR.n1458 VSS 0.004169f
C7608 VDPWR.n1459 VSS 0.023406f
C7609 VDPWR.n1460 VSS 0.002164f
C7610 VDPWR.n1461 VSS 0.002085f
C7611 VDPWR.n1462 VSS 0.003719f
C7612 VDPWR.n1463 VSS 0.001668f
C7613 VDPWR.n1464 VSS 0.002164f
C7614 VDPWR.n1465 VSS 0.00311f
C7615 VDPWR.n1466 VSS 0.013477f
C7616 VDPWR.n1467 VSS 0.00622f
C7617 VDPWR.t1191 VSS 0.076721f
C7618 VDPWR.t1168 VSS 0.076721f
C7619 VDPWR.n1468 VSS 0.07057f
C7620 VDPWR.n1469 VSS 0.00622f
C7621 VDPWR.t871 VSS 0.005792f
C7622 VDPWR.t1027 VSS 0.005792f
C7623 VDPWR.n1470 VSS 0.007899f
C7624 VDPWR.t972 VSS 0.005792f
C7625 VDPWR.t1115 VSS 0.005792f
C7626 VDPWR.n1471 VSS 0.007899f
C7627 VDPWR.n1472 VSS 0.004124f
C7628 VDPWR.n1473 VSS 0.013477f
C7629 VDPWR.n1474 VSS 0.002231f
C7630 VDPWR.n1475 VSS 0.002085f
C7631 VDPWR.n1476 VSS 0.003719f
C7632 VDPWR.n1477 VSS 0.001668f
C7633 VDPWR.n1478 VSS 0.002164f
C7634 VDPWR.n1479 VSS 0.00622f
C7635 VDPWR.t1281 VSS 0.076721f
C7636 VDPWR.t1252 VSS 0.076721f
C7637 VDPWR.n1480 VSS 0.013477f
C7638 VDPWR.n1481 VSS 0.004665f
C7639 VDPWR.t892 VSS 0.005308f
C7640 VDPWR.t1244 VSS 0.011265f
C7641 VDPWR.n1483 VSS 0.028883f
C7642 VDPWR.t893 VSS 0.005308f
C7643 VDPWR.n1484 VSS 0.015733f
C7644 VDPWR.t1080 VSS 0.005809f
C7645 VDPWR.n1485 VSS 0.017223f
C7646 VDPWR.t1026 VSS 0.005792f
C7647 VDPWR.n1486 VSS 0.007319f
C7648 VDPWR.n1487 VSS 0.002164f
C7649 VDPWR.n1488 VSS 0.002085f
C7650 VDPWR.n1489 VSS 0.003719f
C7651 VDPWR.n1490 VSS 0.003719f
C7652 VDPWR.n1491 VSS 0.003115f
C7653 VDPWR.n1492 VSS 0.001668f
C7654 VDPWR.n1493 VSS 0.002164f
C7655 VDPWR.n1494 VSS 0.00311f
C7656 VDPWR.t1213 VSS 0.076721f
C7657 VDPWR.n1495 VSS 0.013477f
C7658 VDPWR.n1496 VSS 0.005646f
C7659 VDPWR.t1192 VSS 0.078173f
C7660 VDPWR.t929 VSS 0.005792f
C7661 VDPWR.n1497 VSS 0.007319f
C7662 VDPWR.n1498 VSS 0.00622f
C7663 VDPWR.n1499 VSS 0.009235f
C7664 VDPWR.n1500 VSS 0.00622f
C7665 VDPWR.t1272 VSS 0.076721f
C7666 VDPWR.n1501 VSS 0.042898f
C7667 VDPWR.n1502 VSS 0.003043f
C7668 VDPWR.n1503 VSS 0.002085f
C7669 VDPWR.n1504 VSS 0.003719f
C7670 VDPWR.n1505 VSS 0.001668f
C7671 VDPWR.n1506 VSS 0.002164f
C7672 VDPWR.t1239 VSS 0.038277f
C7673 VDPWR.n1507 VSS 0.028878f
C7674 VDPWR.t928 VSS 0.005792f
C7675 VDPWR.t910 VSS 0.005265f
C7676 VDPWR.n1508 VSS 0.012671f
C7677 VDPWR.t862 VSS 0.005308f
C7678 VDPWR.t1258 VSS 0.011265f
C7679 VDPWR.n1510 VSS 0.028883f
C7680 VDPWR.t863 VSS 0.005308f
C7681 VDPWR.n1511 VSS 0.015733f
C7682 VDPWR.t1051 VSS 0.005308f
C7683 VDPWR.t1225 VSS 0.011265f
C7684 VDPWR.n1513 VSS 0.028883f
C7685 VDPWR.t1052 VSS 0.005308f
C7686 VDPWR.n1514 VSS 0.015733f
C7687 VDPWR.n1515 VSS 0.012962f
C7688 VDPWR.t835 VSS 0.005308f
C7689 VDPWR.t1262 VSS 0.011265f
C7690 VDPWR.n1517 VSS 0.028883f
C7691 VDPWR.t836 VSS 0.005308f
C7692 VDPWR.n1518 VSS 0.015733f
C7693 VDPWR.n1519 VSS 0.004061f
C7694 VDPWR.n1520 VSS 0.005237f
C7695 VDPWR.t1038 VSS 0.005308f
C7696 VDPWR.t1233 VSS 0.011265f
C7697 VDPWR.n1522 VSS 0.028883f
C7698 VDPWR.t1039 VSS 0.005308f
C7699 VDPWR.n1523 VSS 0.015733f
C7700 VDPWR.n1524 VSS 0.014221f
C7701 VDPWR.n1525 VSS 0.003497f
C7702 VDPWR.n1526 VSS 0.004059f
C7703 VDPWR.n1527 VSS 0.004665f
C7704 VDPWR.n1528 VSS 0.002502f
C7705 VDPWR.n1529 VSS 0.002085f
C7706 VDPWR.n1530 VSS 0.003595f
C7707 VDPWR.n1531 VSS 0.003257f
C7708 VDPWR.n1532 VSS 0.002777f
C7709 VDPWR.n1533 VSS 0.003719f
C7710 VDPWR.n1534 VSS 0.016116f
C7711 VDPWR.n1535 VSS 0.027133f
C7712 VDPWR.n1536 VSS 0.016116f
C7713 VDPWR.n1537 VSS 0.016832f
C7714 VDPWR.n1538 VSS 0.002164f
C7715 VDPWR.n1539 VSS 0.00311f
C7716 VDPWR.n1540 VSS 0.002085f
C7717 VDPWR.n1541 VSS 0.001668f
C7718 VDPWR.n1542 VSS 0.003719f
C7719 VDPWR.n1543 VSS 0.003595f
C7720 VDPWR.n1544 VSS 0.003257f
C7721 VDPWR.n1545 VSS 0.002236f
C7722 VDPWR.n1546 VSS 0.003178f
C7723 VDPWR.n1547 VSS 0.016116f
C7724 VDPWR.n1548 VSS 0.021966f
C7725 VDPWR.t911 VSS 0.005265f
C7726 VDPWR.n1549 VSS 0.012091f
C7727 VDPWR.n1550 VSS 0.021249f
C7728 VDPWR.n1551 VSS 0.00622f
C7729 VDPWR.n1552 VSS 0.003685f
C7730 VDPWR.n1553 VSS 0.004665f
C7731 VDPWR.n1554 VSS 0.005928f
C7732 VDPWR.t1025 VSS 0.005792f
C7733 VDPWR.n1555 VSS 0.007319f
C7734 VDPWR.n1556 VSS 0.013038f
C7735 VDPWR.n1557 VSS 0.013038f
C7736 VDPWR.n1558 VSS 0.00622f
C7737 VDPWR.n1559 VSS 0.003685f
C7738 VDPWR.n1560 VSS 0.00339f
C7739 VDPWR.n1561 VSS 0.036257f
C7740 VDPWR.n1562 VSS 0.003026f
C7741 VDPWR.t1079 VSS 0.005792f
C7742 VDPWR.n1563 VSS 0.007319f
C7743 VDPWR.n1564 VSS 0.013038f
C7744 VDPWR.n1565 VSS 0.00622f
C7745 VDPWR.n1566 VSS 0.00622f
C7746 VDPWR.n1567 VSS 0.0048f
C7747 VDPWR.n1568 VSS 0.010328f
C7748 VDPWR.n1569 VSS 0.038654f
C7749 VDPWR.n1570 VSS 0.009888f
C7750 VDPWR.n1571 VSS 0.013038f
C7751 VDPWR.n1572 VSS 0.013477f
C7752 VDPWR.n1573 VSS 0.002164f
C7753 VDPWR.n1574 VSS 0.001668f
C7754 VDPWR.n1575 VSS 0.002085f
C7755 VDPWR.n1576 VSS 0.002366f
C7756 VDPWR.n1577 VSS 0.002907f
C7757 VDPWR.n1578 VSS 0.002085f
C7758 VDPWR.n1579 VSS 0.003257f
C7759 VDPWR.n1580 VSS 0.003595f
C7760 VDPWR.n1581 VSS 0.256026f
C7761 VDPWR.n1582 VSS 0.003595f
C7762 VDPWR.n1583 VSS 0.003257f
C7763 VDPWR.n1584 VSS 0.003115f
C7764 VDPWR.n1585 VSS 0.002671f
C7765 VDPWR.n1586 VSS 0.006356f
C7766 VDPWR.t861 VSS 0.06996f
C7767 VDPWR.t834 VSS 0.076737f
C7768 VDPWR.t909 VSS 0.115803f
C7769 VDPWR.t927 VSS 0.067568f
C7770 VDPWR.t1024 VSS 0.115803f
C7771 VDPWR.t1078 VSS 0.104242f
C7772 VDPWR.t855 VSS 0.055011f
C7773 VDPWR.t864 VSS 0.220045f
C7774 VDPWR.t203 VSS 0.030495f
C7775 VDPWR.t67 VSS 0.023719f
C7776 VDPWR.t1058 VSS 0.067568f
C7777 VDPWR.t1089 VSS 0.097266f
C7778 VDPWR.n1587 VSS 0.043147f
C7779 VDPWR.t870 VSS 0.220045f
C7780 VDPWR.t970 VSS 0.220045f
C7781 VDPWR.t891 VSS 0.0584f
C7782 VDPWR.n1588 VSS 0.054868f
C7783 VDPWR.n1589 VSS 0.016847f
C7784 VDPWR.n1590 VSS 0.003347f
C7785 VDPWR.n1591 VSS 0.005232f
C7786 VDPWR.n1592 VSS 0.010931f
C7787 VDPWR.n1593 VSS 0.004675f
C7788 VDPWR.t971 VSS 0.005792f
C7789 VDPWR.t1114 VSS 0.005792f
C7790 VDPWR.n1594 VSS 0.007899f
C7791 VDPWR.n1595 VSS 0.013038f
C7792 VDPWR.n1596 VSS 0.00622f
C7793 VDPWR.n1597 VSS 0.00622f
C7794 VDPWR.n1598 VSS 0.00622f
C7795 VDPWR.n1599 VSS 0.010328f
C7796 VDPWR.n1600 VSS 0.07057f
C7797 VDPWR.n1601 VSS 0.009888f
C7798 VDPWR.n1602 VSS 0.013477f
C7799 VDPWR.n1603 VSS 0.013477f
C7800 VDPWR.n1604 VSS 0.005882f
C7801 VDPWR.n1605 VSS 0.003115f
C7802 VDPWR.n1606 VSS 0.003595f
C7803 VDPWR.n1607 VSS 0.003257f
C7804 VDPWR.n1608 VSS 0.002085f
C7805 VDPWR.n1609 VSS 0.00311f
C7806 VDPWR.n1610 VSS 0.002164f
C7807 VDPWR.n1611 VSS 0.003043f
C7808 VDPWR.n1612 VSS 0.002085f
C7809 VDPWR.n1613 VSS 0.001668f
C7810 VDPWR.n1614 VSS 0.003719f
C7811 VDPWR.n1615 VSS 0.003595f
C7812 VDPWR.n1616 VSS 0.003257f
C7813 VDPWR.n1617 VSS 0.003115f
C7814 VDPWR.n1618 VSS 0.002164f
C7815 VDPWR.n1619 VSS 0.013477f
C7816 VDPWR.n1620 VSS 0.013477f
C7817 VDPWR.n1621 VSS 0.013038f
C7818 VDPWR.n1622 VSS 0.00622f
C7819 VDPWR.n1623 VSS 0.00509f
C7820 VDPWR.n1624 VSS 0.004977f
C7821 VDPWR.n1625 VSS 0.005646f
C7822 VDPWR.n1626 VSS 0.00622f
C7823 VDPWR.n1627 VSS 0.013038f
C7824 VDPWR.n1628 VSS 0.013477f
C7825 VDPWR.n1629 VSS 0.010328f
C7826 VDPWR.n1630 VSS 0.00622f
C7827 VDPWR.n1631 VSS 0.00622f
C7828 VDPWR.n1632 VSS 0.009888f
C7829 VDPWR.n1633 VSS 0.013477f
C7830 VDPWR.n1634 VSS 0.013477f
C7831 VDPWR.n1635 VSS 0.00622f
C7832 VDPWR.n1636 VSS 0.00622f
C7833 VDPWR.n1637 VSS 0.002366f
C7834 VDPWR.n1638 VSS 0.002085f
C7835 VDPWR.n1639 VSS 0.003595f
C7836 VDPWR.n1640 VSS 0.003257f
C7837 VDPWR.n1641 VSS 0.002912f
C7838 VDPWR.n1642 VSS 0.003854f
C7839 VDPWR.n1643 VSS 0.013477f
C7840 VDPWR.n1644 VSS 0.013477f
C7841 VDPWR.t872 VSS 0.005792f
C7842 VDPWR.n1645 VSS 0.004785f
C7843 VDPWR.t1028 VSS 0.005792f
C7844 VDPWR.n1646 VSS 0.007899f
C7845 VDPWR.n1647 VSS 0.013038f
C7846 VDPWR.n1648 VSS 0.002164f
C7847 VDPWR.n1649 VSS 0.00311f
C7848 VDPWR.n1650 VSS 0.002085f
C7849 VDPWR.n1651 VSS 0.001668f
C7850 VDPWR.n1652 VSS 0.003719f
C7851 VDPWR.n1653 VSS 0.003595f
C7852 VDPWR.n1654 VSS 0.003257f
C7853 VDPWR.n1655 VSS 5.79e-19
C7854 VDPWR.n1656 VSS 0.003347f
C7855 VDPWR.n1657 VSS 0.002366f
C7856 VDPWR.n1658 VSS 0.001735f
C7857 VDPWR.n1659 VSS 0.003194f
C7858 VDPWR.n1660 VSS 0.0024f
C7859 VDPWR.n1661 VSS 0.004665f
C7860 VDPWR.n1662 VSS 0.009163f
C7861 VDPWR.t1090 VSS 0.005265f
C7862 VDPWR.n1663 VSS 0.012091f
C7863 VDPWR.n1664 VSS 0.015997f
C7864 VDPWR.n1665 VSS 0.055357f
C7865 VDPWR.t1222 VSS 0.076721f
C7866 VDPWR.n1666 VSS 0.042898f
C7867 VDPWR.n1667 VSS 0.011102f
C7868 VDPWR.n1668 VSS 0.00622f
C7869 VDPWR.n1669 VSS 0.00622f
C7870 VDPWR.n1670 VSS 0.00622f
C7871 VDPWR.n1671 VSS 0.021966f
C7872 VDPWR.n1672 VSS 0.021966f
C7873 VDPWR.t1091 VSS 0.005265f
C7874 VDPWR.n1673 VSS 0.012091f
C7875 VDPWR.n1674 VSS 0.021249f
C7876 VDPWR.n1675 VSS 0.00622f
C7877 VDPWR.n1676 VSS 0.003685f
C7878 VDPWR.n1677 VSS 0.002085f
C7879 VDPWR.n1678 VSS 0.003595f
C7880 VDPWR.n1679 VSS 0.003257f
C7881 VDPWR.n1680 VSS 0.00156f
C7882 VDPWR.n1681 VSS 0.001859f
C7883 VDPWR.n1682 VSS 0.007471f
C7884 VDPWR.n1683 VSS 0.014368f
C7885 VDPWR.n1684 VSS 0.002164f
C7886 VDPWR.n1685 VSS 0.002231f
C7887 VDPWR.n1686 VSS 0.002085f
C7888 VDPWR.n1687 VSS 0.001668f
C7889 VDPWR.n1688 VSS 0.003719f
C7890 VDPWR.n1689 VSS 0.003595f
C7891 VDPWR.n1690 VSS 0.003257f
C7892 VDPWR.n1691 VSS 9.85e-19
C7893 VDPWR.n1692 VSS 0.001589f
C7894 VDPWR.n1693 VSS 0.0031f
C7895 VDPWR.n1694 VSS 0.005006f
C7896 VDPWR.n1695 VSS 0.004665f
C7897 VDPWR.n1696 VSS 0.00622f
C7898 VDPWR.n1697 VSS 0.013038f
C7899 VDPWR.n1698 VSS 0.013477f
C7900 VDPWR.n1699 VSS 0.010328f
C7901 VDPWR.n1700 VSS 0.00622f
C7902 VDPWR.n1701 VSS 0.00622f
C7903 VDPWR.n1702 VSS 0.009888f
C7904 VDPWR.n1703 VSS 0.013477f
C7905 VDPWR.n1704 VSS 0.013477f
C7906 VDPWR.n1705 VSS 0.00622f
C7907 VDPWR.n1706 VSS 0.00622f
C7908 VDPWR.n1707 VSS 0.00622f
C7909 VDPWR.n1708 VSS 0.013477f
C7910 VDPWR.n1709 VSS 0.013477f
C7911 VDPWR.t866 VSS 0.005792f
C7912 VDPWR.t1014 VSS 0.005792f
C7913 VDPWR.n1710 VSS 0.007899f
C7914 VDPWR.n1711 VSS 0.013038f
C7915 VDPWR.n1712 VSS 0.006018f
C7916 VDPWR.n1713 VSS 7.78e-19
C7917 VDPWR.n1714 VSS 0.003115f
C7918 VDPWR.n1715 VSS 0.003257f
C7919 VDPWR.n1716 VSS 0.001668f
C7920 VDPWR.n1717 VSS 0.002085f
C7921 VDPWR.n1718 VSS 0.002535f
C7922 VDPWR.n1719 VSS 0.00311f
C7923 VDPWR.n1720 VSS 0.002164f
C7924 VDPWR.t1053 VSS 0.005308f
C7925 VDPWR.t1226 VSS 0.011265f
C7926 VDPWR.n1722 VSS 0.028883f
C7927 VDPWR.t1054 VSS 0.005308f
C7928 VDPWR.n1723 VSS 0.015733f
C7929 VDPWR.n1724 VSS 0.013263f
C7930 VDPWR.n1725 VSS 0.001454f
C7931 VDPWR.n1726 VSS 0.003047f
C7932 VDPWR.n1727 VSS 0.002231f
C7933 VDPWR.n1728 VSS 0.002085f
C7934 VDPWR.n1729 VSS 0.001668f
C7935 VDPWR.n1730 VSS 0.003719f
C7936 VDPWR.n1731 VSS 0.003595f
C7937 VDPWR.n1732 VSS 0.259227f
C7938 VDPWR.n1733 VSS 0.248273f
C7939 VDPWR.n1734 VSS 0.003719f
C7940 VDPWR.n1735 VSS 0.007285f
C7941 VDPWR.n1736 VSS 0.003595f
C7942 VDPWR.n1737 VSS 0.003257f
C7943 VDPWR.n1738 VSS 0.001555f
C7944 VDPWR.n1739 VSS 0.002085f
C7945 VDPWR.n1740 VSS 0.001668f
C7946 VDPWR.n1741 VSS 0.00311f
C7947 VDPWR.n1742 VSS 0.002085f
C7948 VDPWR.n1743 VSS 0.001668f
C7949 VDPWR.n1744 VSS 0.003719f
C7950 VDPWR.n1745 VSS 0.003595f
C7951 VDPWR.n1746 VSS 0.003257f
C7952 VDPWR.n1747 VSS 0.003047f
C7953 VDPWR.n1748 VSS 0.001454f
C7954 VDPWR.n1749 VSS 0.012953f
C7955 VDPWR.n1750 VSS 0.019039f
C7956 VDPWR.n1751 VSS 0.001856f
C7957 VDPWR.n1752 VSS 0.002366f
C7958 VDPWR.n1753 VSS 0.003685f
C7959 VDPWR.n1754 VSS 0.00622f
C7960 VDPWR.n1755 VSS 0.001197f
C7961 VDPWR.n1756 VSS 0.005459f
C7962 VDPWR.n1757 VSS 0.004755f
C7963 VDPWR.n1758 VSS 9.94e-19
C7964 VDPWR.n1759 VSS 0.007321f
C7965 VDPWR.n1760 VSS 0.00622f
C7966 VDPWR.n1761 VSS 0.00622f
C7967 VDPWR.n1762 VSS 0.001317f
C7968 VDPWR.n1763 VSS 0.002203f
C7969 VDPWR.n1764 VSS 0.002084f
C7970 VDPWR.n1765 VSS 0.005071f
C7971 VDPWR.n1766 VSS 0.00254f
C7972 VDPWR.n1767 VSS 0.003257f
C7973 VDPWR.n1768 VSS 0.003595f
C7974 VDPWR.n1769 VSS 0.245208f
C7975 VDPWR.n1770 VSS 0.003595f
C7976 VDPWR.n1771 VSS 0.003257f
C7977 VDPWR.n1772 VSS 0.003115f
C7978 VDPWR.n1773 VSS 0.004936f
C7979 VDPWR.n1774 VSS 0.00784f
C7980 VDPWR.n1775 VSS 0.00784f
C7981 VDPWR.n1776 VSS 0.004218f
C7982 VDPWR.n1777 VSS 0.00622f
C7983 VDPWR.n1778 VSS 0.00622f
C7984 VDPWR.n1779 VSS 0.005646f
C7985 VDPWR.n1780 VSS 0.004005f
C7986 VDPWR.n1781 VSS 0.006407f
C7987 VDPWR.n1782 VSS 0.03575f
C7988 VDPWR.n1783 VSS 0.004772f
C7989 VDPWR.n1784 VSS 0.00213f
C7990 VDPWR.n1785 VSS 0.006452f
C7991 VDPWR.n1786 VSS 0.00213f
C7992 VDPWR.n1787 VSS 0.002431f
C7993 VDPWR.n1788 VSS 0.006613f
C7994 VDPWR.n1789 VSS 0.016847f
C7995 VDPWR.n1790 VSS 0.003347f
C7996 VDPWR.n1791 VSS 5.79e-19
C7997 VDPWR.n1792 VSS 0.003257f
C7998 VDPWR.n1793 VSS 0.003595f
C7999 VDPWR.n1794 VSS 0.245208f
C8000 VDPWR.n1795 VSS 0.003595f
C8001 VDPWR.n1796 VSS 0.003257f
C8002 VDPWR.n1797 VSS 0.002912f
C8003 VDPWR.n1798 VSS 0.003854f
C8004 VDPWR.n1799 VSS 0.013477f
C8005 VDPWR.n1800 VSS 0.013477f
C8006 VDPWR.n1801 VSS 0.009888f
C8007 VDPWR.n1802 VSS 0.00622f
C8008 VDPWR.n1803 VSS 0.00622f
C8009 VDPWR.n1804 VSS 0.010328f
C8010 VDPWR.n1805 VSS 0.009888f
C8011 VDPWR.n1806 VSS 0.038654f
C8012 VDPWR.n1807 VSS 0.009888f
C8013 VDPWR.n1808 VSS 0.00622f
C8014 VDPWR.n1809 VSS 0.005646f
C8015 VDPWR.n1810 VSS 0.004907f
C8016 VDPWR.n1811 VSS 0.011783f
C8017 VDPWR.n1812 VSS 0.004565f
C8018 VDPWR.n1813 VSS 0.00449f
C8019 VDPWR.n1814 VSS 0.003685f
C8020 VDPWR.n1815 VSS 0.005003f
C8021 VDPWR.t1159 VSS 0.005792f
C8022 VDPWR.n1816 VSS 0.007319f
C8023 VDPWR.n1817 VSS 0.013038f
C8024 VDPWR.n1818 VSS 0.013477f
C8025 VDPWR.n1819 VSS 0.004124f
C8026 VDPWR.n1820 VSS 0.003115f
C8027 VDPWR.n1821 VSS 0.003257f
C8028 VDPWR.n1822 VSS 0.003595f
C8029 VDPWR.n1823 VSS 0.245208f
C8030 VDPWR.n1824 VSS 0.003595f
C8031 VDPWR.n1825 VSS 0.003257f
C8032 VDPWR.n1826 VSS 0.003115f
C8033 VDPWR.n1827 VSS 0.005882f
C8034 VDPWR.n1828 VSS 0.010328f
C8035 VDPWR.n1829 VSS 0.009888f
C8036 VDPWR.n1830 VSS 0.038654f
C8037 VDPWR.n1831 VSS 0.009888f
C8038 VDPWR.n1832 VSS 0.00622f
C8039 VDPWR.n1833 VSS 0.004665f
C8040 VDPWR.n1834 VSS 0.004907f
C8041 VDPWR.n1835 VSS 0.011783f
C8042 VDPWR.n1836 VSS 0.007446f
C8043 VDPWR.t1131 VSS 0.005344f
C8044 VDPWR.n1837 VSS 0.015593f
C8045 VDPWR.n1838 VSS 0.016558f
C8046 VDPWR.t1189 VSS 0.022315f
C8047 VDPWR.n1839 VSS 0.022091f
C8048 VDPWR.t1130 VSS 0.005265f
C8049 VDPWR.n1840 VSS 0.006338f
C8050 VDPWR.t957 VSS 0.00581f
C8051 VDPWR.n1841 VSS 0.011909f
C8052 VDPWR.n1842 VSS 0.006339f
C8053 VDPWR.n1843 VSS 0.003323f
C8054 VDPWR.n1844 VSS 0.002366f
C8055 VDPWR.n1845 VSS 0.003347f
C8056 VDPWR.n1846 VSS 0.018083f
C8057 VDPWR.n1847 VSS 0.006356f
C8058 VDPWR.n1848 VSS 0.002671f
C8059 VDPWR.n1849 VSS 0.003115f
C8060 VDPWR.n1850 VSS 0.003257f
C8061 VDPWR.n1851 VSS 0.003595f
C8062 VDPWR.n1852 VSS 0.003719f
C8063 VDPWR.n1853 VSS 0.003719f
C8064 VDPWR.n1854 VSS 0.003595f
C8065 VDPWR.n1855 VSS 0.003257f
C8066 VDPWR.n1856 VSS 0.003115f
C8067 VDPWR.n1857 VSS 0.0048f
C8068 VDPWR.n1858 VSS 0.00622f
C8069 VDPWR.n1859 VSS 0.013477f
C8070 VDPWR.n1860 VSS 0.013038f
C8071 VDPWR.t956 VSS 0.005792f
C8072 VDPWR.n1861 VSS 0.007319f
C8073 VDPWR.n1862 VSS 0.003026f
C8074 VDPWR.n1863 VSS 0.005646f
C8075 VDPWR.n1864 VSS 0.003685f
C8076 VDPWR.n1865 VSS 0.00339f
C8077 VDPWR.t987 VSS 0.005792f
C8078 VDPWR.n1866 VSS 0.007319f
C8079 VDPWR.n1867 VSS 0.013038f
C8080 VDPWR.n1868 VSS 0.013038f
C8081 VDPWR.n1869 VSS 0.00622f
C8082 VDPWR.n1870 VSS 0.004665f
C8083 VDPWR.n1871 VSS 0.005928f
C8084 VDPWR.n1872 VSS 0.009235f
C8085 VDPWR.n1873 VSS 0.003685f
C8086 VDPWR.n1874 VSS 0.00622f
C8087 VDPWR.n1875 VSS 0.021249f
C8088 VDPWR.n1876 VSS 0.021966f
C8089 VDPWR.n1877 VSS 0.016116f
C8090 VDPWR.n1878 VSS 0.003178f
C8091 VDPWR.n1879 VSS 0.002236f
C8092 VDPWR.n1880 VSS 0.002085f
C8093 VDPWR.n1881 VSS 0.003719f
C8094 VDPWR.n1882 VSS 0.001668f
C8095 VDPWR.n1883 VSS 0.003257f
C8096 VDPWR.n1884 VSS 0.002085f
C8097 VDPWR.n1885 VSS 0.003043f
C8098 VDPWR.n1886 VSS 0.002164f
C8099 VDPWR.n1887 VSS 0.016832f
C8100 VDPWR.n1888 VSS 0.016116f
C8101 VDPWR.n1889 VSS 0.002164f
C8102 VDPWR.n1890 VSS 0.002502f
C8103 VDPWR.n1891 VSS 0.002085f
C8104 VDPWR.n1892 VSS 0.003257f
C8105 VDPWR.n1893 VSS 0.003595f
C8106 VDPWR.n1894 VSS 0.245208f
C8107 VDPWR.n1895 VSS 0.003719f
C8108 VDPWR.n1896 VSS 0.002777f
C8109 VDPWR.n1897 VSS 0.001668f
C8110 VDPWR.n1898 VSS 0.001668f
C8111 VDPWR.n1899 VSS 0.002085f
C8112 VDPWR.n1900 VSS 0.00311f
C8113 VDPWR.n1901 VSS 0.016116f
C8114 VDPWR.t983 VSS 0.005792f
C8115 VDPWR.t883 VSS 0.005265f
C8116 VDPWR.n1902 VSS 0.012671f
C8117 VDPWR.n1903 VSS 0.004059f
C8118 VDPWR.t1022 VSS 0.005308f
C8119 VDPWR.t1186 VSS 0.011265f
C8120 VDPWR.n1905 VSS 0.028883f
C8121 VDPWR.t1023 VSS 0.005308f
C8122 VDPWR.n1906 VSS 0.015733f
C8123 VDPWR.n1907 VSS 0.003719f
C8124 VDPWR.n1908 VSS 0.004665f
C8125 VDPWR.n1909 VSS 0.005237f
C8126 VDPWR.t1099 VSS 0.005308f
C8127 VDPWR.t1169 VSS 0.011265f
C8128 VDPWR.n1911 VSS 0.028883f
C8129 VDPWR.t1100 VSS 0.005308f
C8130 VDPWR.n1912 VSS 0.015733f
C8131 VDPWR.t847 VSS 0.005308f
C8132 VDPWR.t1251 VSS 0.011265f
C8133 VDPWR.n1914 VSS 0.028883f
C8134 VDPWR.t848 VSS 0.005308f
C8135 VDPWR.n1915 VSS 0.015733f
C8136 VDPWR.n1916 VSS 0.004061f
C8137 VDPWR.t939 VSS 0.005308f
C8138 VDPWR.t1229 VSS 0.011265f
C8139 VDPWR.n1918 VSS 0.028883f
C8140 VDPWR.t940 VSS 0.005308f
C8141 VDPWR.n1919 VSS 0.015733f
C8142 VDPWR.n1920 VSS 0.012962f
C8143 VDPWR.n1921 VSS 0.014221f
C8144 VDPWR.n1922 VSS 0.003497f
C8145 VDPWR.t1241 VSS 0.038277f
C8146 VDPWR.n1923 VSS 0.028878f
C8147 VDPWR.n1924 VSS 0.027133f
C8148 VDPWR.n1925 VSS 0.002164f
C8149 VDPWR.n1926 VSS 0.016832f
C8150 VDPWR.n1927 VSS 0.016116f
C8151 VDPWR.n1928 VSS 0.002164f
C8152 VDPWR.n1929 VSS 0.002502f
C8153 VDPWR.n1930 VSS 0.002085f
C8154 VDPWR.n1931 VSS 0.003257f
C8155 VDPWR.n1932 VSS 0.003595f
C8156 VDPWR.n1933 VSS 0.245208f
C8157 VDPWR.n1934 VSS 0.003595f
C8158 VDPWR.n1935 VSS 0.003257f
C8159 VDPWR.n1936 VSS 0.002236f
C8160 VDPWR.n1937 VSS 0.003178f
C8161 VDPWR.n1938 VSS 0.016116f
C8162 VDPWR.n1939 VSS 0.021966f
C8163 VDPWR.t884 VSS 0.005265f
C8164 VDPWR.n1940 VSS 0.012091f
C8165 VDPWR.n1941 VSS 0.021249f
C8166 VDPWR.n1942 VSS 0.00622f
C8167 VDPWR.n1943 VSS 0.003685f
C8168 VDPWR.n1944 VSS 0.004665f
C8169 VDPWR.n1945 VSS 0.005928f
C8170 VDPWR.t965 VSS 0.005792f
C8171 VDPWR.n1946 VSS 0.007319f
C8172 VDPWR.n1947 VSS 0.013038f
C8173 VDPWR.n1948 VSS 0.013038f
C8174 VDPWR.n1949 VSS 0.00622f
C8175 VDPWR.n1950 VSS 0.003685f
C8176 VDPWR.n1951 VSS 0.00339f
C8177 VDPWR.t1208 VSS 0.078173f
C8178 VDPWR.n1952 VSS 0.036257f
C8179 VDPWR.n1953 VSS 0.003026f
C8180 VDPWR.t951 VSS 0.005792f
C8181 VDPWR.n1954 VSS 0.007319f
C8182 VDPWR.n1955 VSS 0.013038f
C8183 VDPWR.n1956 VSS 0.00622f
C8184 VDPWR.n1957 VSS 0.00622f
C8185 VDPWR.n1958 VSS 0.0048f
C8186 VDPWR.n1959 VSS 0.010328f
C8187 VDPWR.n1960 VSS 0.038654f
C8188 VDPWR.n1961 VSS 0.009888f
C8189 VDPWR.n1962 VSS 0.013477f
C8190 VDPWR.n1963 VSS 0.016847f
C8191 VDPWR.t952 VSS 0.005809f
C8192 VDPWR.n1964 VSS 0.017223f
C8193 VDPWR.n1965 VSS 0.010226f
C8194 VDPWR.n1966 VSS 0.00622f
C8195 VDPWR.n1967 VSS 0.01126f
C8196 VDPWR.n1968 VSS 0.016832f
C8197 VDPWR.t1271 VSS 0.076721f
C8198 VDPWR.n1969 VSS 0.042181f
C8199 VDPWR.t854 VSS 0.005265f
C8200 VDPWR.n1970 VSS 0.006241f
C8201 VDPWR.t1070 VSS 0.005792f
C8202 VDPWR.n1971 VSS 0.007319f
C8203 VDPWR.n1972 VSS 0.002164f
C8204 VDPWR.n1973 VSS 0.002085f
C8205 VDPWR.n1974 VSS 0.001668f
C8206 VDPWR.n1975 VSS 0.001668f
C8207 VDPWR.n1976 VSS 0.002085f
C8208 VDPWR.n1977 VSS 0.002164f
C8209 VDPWR.n1978 VSS 0.00622f
C8210 VDPWR.t1172 VSS 0.076721f
C8211 VDPWR.n1979 VSS 0.013038f
C8212 VDPWR.n1980 VSS 0.00311f
C8213 VDPWR.n1981 VSS 0.002231f
C8214 VDPWR.n1982 VSS 0.002085f
C8215 VDPWR.n1983 VSS 0.003043f
C8216 VDPWR.n1984 VSS 0.002164f
C8217 VDPWR.n1985 VSS 0.013477f
C8218 VDPWR.n1986 VSS 0.010328f
C8219 VDPWR.n1987 VSS 0.038654f
C8220 VDPWR.n1988 VSS 0.006081f
C8221 VDPWR.n1989 VSS 0.00622f
C8222 VDPWR.t1049 VSS 0.005792f
C8223 VDPWR.n1990 VSS 0.007319f
C8224 VDPWR.t1184 VSS 0.076721f
C8225 VDPWR.n1991 VSS 0.038215f
C8226 VDPWR.t1071 VSS 0.005792f
C8227 VDPWR.n1992 VSS 0.00373f
C8228 VDPWR.t1064 VSS 0.005792f
C8229 VDPWR.n1993 VSS 0.007319f
C8230 VDPWR.n1994 VSS 0.00622f
C8231 VDPWR.t1174 VSS 0.076721f
C8232 VDPWR.n1995 VSS 0.038654f
C8233 VDPWR.n1996 VSS 0.002366f
C8234 VDPWR.n1997 VSS 0.002085f
C8235 VDPWR.n1998 VSS 0.001668f
C8236 VDPWR.n1999 VSS 0.001668f
C8237 VDPWR.n2000 VSS 0.002085f
C8238 VDPWR.n2001 VSS 0.002164f
C8239 VDPWR.t846 VSS 0.06996f
C8240 VDPWR.t1021 VSS 0.076737f
C8241 VDPWR.t882 VSS 0.115803f
C8242 VDPWR.t982 VSS 0.067568f
C8243 VDPWR.t964 VSS 0.115803f
C8244 VDPWR.t950 VSS 0.104242f
C8245 VDPWR.n2002 VSS 0.076594f
C8246 VDPWR.t852 VSS 0.091685f
C8247 VDPWR.t1154 VSS 0.115803f
C8248 VDPWR.t1069 VSS 0.104242f
C8249 VDPWR.t1048 VSS 0.115803f
C8250 VDPWR.t1063 VSS 0.104242f
C8251 VDPWR.t918 VSS 0.055011f
C8252 VDPWR.t210 VSS 0.048833f
C8253 VDPWR.t436 VSS 0.03488f
C8254 VDPWR.t479 VSS 0.018337f
C8255 VDPWR.t1010 VSS 0.006976f
C8256 VDPWR.t183 VSS 0.050028f
C8257 VDPWR.t181 VSS 0.040461f
C8258 VDPWR.t185 VSS 0.012955f
C8259 VDPWR.t438 VSS 0.022722f
C8260 VDPWR.t735 VSS 0.016743f
C8261 VDPWR.t454 VSS 0.016743f
C8262 VDPWR.t284 VSS 0.018536f
C8263 VDPWR.t207 VSS 0.018935f
C8264 VDPWR.t367 VSS 0.018935f
C8265 VDPWR.t73 VSS 0.02631f
C8266 VDPWR.t653 VSS 0.024516f
C8267 VDPWR.t687 VSS 0.013753f
C8268 VDPWR.t283 VSS 0.018935f
C8269 VDPWR.t11 VSS 0.018935f
C8270 VDPWR.t736 VSS 0.016743f
C8271 VDPWR.t13 VSS 0.016942f
C8272 VDPWR.t675 VSS 0.024715f
C8273 VDPWR.t760 VSS 0.013554f
C8274 VDPWR.t285 VSS 0.014351f
C8275 VDPWR.t505 VSS 0.016743f
C8276 VDPWR.t86 VSS 0.009368f
C8277 VDPWR.t1144 VSS 0.076737f
C8278 VDPWR.n2003 VSS 0.064037f
C8279 VDPWR.n2004 VSS 0.009888f
C8280 VDPWR.n2005 VSS 0.002164f
C8281 VDPWR.n2006 VSS 0.002085f
C8282 VDPWR.n2007 VSS 0.00311f
C8283 VDPWR.n2008 VSS 0.00311f
C8284 VDPWR.n2009 VSS 0.002164f
C8285 VDPWR.n2010 VSS 0.013038f
C8286 VDPWR.t1050 VSS 0.005792f
C8287 VDPWR.n2011 VSS 0.007319f
C8288 VDPWR.n2012 VSS 0.006356f
C8289 VDPWR.t1145 VSS 0.005265f
C8290 VDPWR.n2013 VSS 0.006599f
C8291 VDPWR.n2014 VSS 0.00622f
C8292 VDPWR.t1275 VSS 0.021971f
C8293 VDPWR.n2015 VSS 0.022507f
C8294 VDPWR.t1146 VSS 0.005265f
C8295 VDPWR.t506 VSS 0.007592f
C8296 VDPWR.n2016 VSS 0.012849f
C8297 VDPWR.n2017 VSS 0.003651f
C8298 VDPWR.t676 VSS 0.002909f
C8299 VDPWR.t14 VSS 0.00665f
C8300 VDPWR.n2018 VSS 0.005788f
C8301 VDPWR.n2019 VSS 0.004936f
C8302 VDPWR.n2020 VSS 0.001688f
C8303 VDPWR.n2021 VSS 0.003115f
C8304 VDPWR.n2022 VSS 0.003257f
C8305 VDPWR.n2023 VSS 0.002085f
C8306 VDPWR.n2024 VSS 0.001668f
C8307 VDPWR.n2025 VSS 0.002085f
C8308 VDPWR.n2026 VSS 0.001555f
C8309 VDPWR.n2027 VSS 0.002164f
C8310 VDPWR.n2028 VSS 0.00311f
C8311 VDPWR.n2029 VSS 0.002164f
C8312 VDPWR.n2030 VSS 0.005137f
C8313 VDPWR.t208 VSS 0.001183f
C8314 VDPWR.t74 VSS -0.001244f
C8315 VDPWR.n2031 VSS 0.007877f
C8316 VDPWR.t654 VSS 0.002942f
C8317 VDPWR.t368 VSS 0.001426f
C8318 VDPWR.n2032 VSS 0.00599f
C8319 VDPWR.n2033 VSS 0.004582f
C8320 VDPWR.n2034 VSS 0.004627f
C8321 VDPWR.n2035 VSS 0.001173f
C8322 VDPWR.t182 VSS 0.001902f
C8323 VDPWR.t184 VSS 0.001902f
C8324 VDPWR.n2036 VSS 0.004272f
C8325 VDPWR.n2037 VSS 0.018084f
C8326 VDPWR.t186 VSS 0.002994f
C8327 VDPWR.n2038 VSS 0.00622f
C8328 VDPWR.n2039 VSS 0.013554f
C8329 VDPWR.t1196 VSS 0.039499f
C8330 VDPWR.t1011 VSS 0.005265f
C8331 VDPWR.n2040 VSS 0.06614f
C8332 VDPWR.n2041 VSS 0.017376f
C8333 VDPWR.t437 VSS 0.001972f
C8334 VDPWR.t211 VSS 0.002183f
C8335 VDPWR.n2042 VSS 0.004205f
C8336 VDPWR.t1012 VSS 0.005265f
C8337 VDPWR.n2043 VSS 0.009272f
C8338 VDPWR.n2044 VSS 7.78e-19
C8339 VDPWR.n2045 VSS 0.002085f
C8340 VDPWR.n2046 VSS 0.003719f
C8341 VDPWR.n2047 VSS 0.001668f
C8342 VDPWR.n2048 VSS 0.001555f
C8343 VDPWR.n2049 VSS 0.002164f
C8344 VDPWR.n2050 VSS 0.002231f
C8345 VDPWR.n2051 VSS 0.005779f
C8346 VDPWR.t919 VSS 0.005308f
C8347 VDPWR.t1232 VSS 0.011265f
C8348 VDPWR.n2053 VSS 0.028883f
C8349 VDPWR.t920 VSS 0.005308f
C8350 VDPWR.n2054 VSS 0.015733f
C8351 VDPWR.t997 VSS 0.005308f
C8352 VDPWR.t1203 VSS 0.011265f
C8353 VDPWR.n2056 VSS 0.028883f
C8354 VDPWR.t998 VSS 0.005308f
C8355 VDPWR.n2057 VSS 0.015733f
C8356 VDPWR.n2058 VSS 0.002085f
C8357 VDPWR.n2059 VSS 0.003595f
C8358 VDPWR.n2060 VSS 0.003257f
C8359 VDPWR.n2061 VSS 0.003047f
C8360 VDPWR.n2062 VSS 0.001454f
C8361 VDPWR.n2063 VSS 0.013261f
C8362 VDPWR.n2064 VSS 0.002164f
C8363 VDPWR.n2065 VSS 0.00311f
C8364 VDPWR.n2066 VSS 0.002085f
C8365 VDPWR.n2067 VSS 0.001668f
C8366 VDPWR.n2068 VSS 0.003719f
C8367 VDPWR.n2069 VSS 0.003595f
C8368 VDPWR.n2070 VSS 0.003257f
C8369 VDPWR.n2071 VSS 0.00156f
C8370 VDPWR.n2072 VSS 0.004665f
C8371 VDPWR.n2073 VSS 0.015796f
C8372 VDPWR.n2074 VSS 0.008342f
C8373 VDPWR.n2075 VSS 0.010531f
C8374 VDPWR.n2076 VSS 0.013222f
C8375 VDPWR.n2077 VSS 0.005646f
C8376 VDPWR.n2078 VSS 0.00213f
C8377 VDPWR.n2079 VSS 0.006585f
C8378 VDPWR.n2080 VSS 0.002366f
C8379 VDPWR.n2081 VSS 0.006842f
C8380 VDPWR.t455 VSS 7.99e-19
C8381 VDPWR.t439 VSS 7.99e-19
C8382 VDPWR.n2082 VSS 0.001849f
C8383 VDPWR.n2083 VSS 0.017477f
C8384 VDPWR.n2084 VSS 0.002203f
C8385 VDPWR.n2085 VSS 0.007147f
C8386 VDPWR.n2086 VSS 0.003115f
C8387 VDPWR.n2087 VSS 0.003257f
C8388 VDPWR.n2088 VSS 0.003595f
C8389 VDPWR.n2089 VSS 0.003719f
C8390 VDPWR.n2090 VSS 0.003595f
C8391 VDPWR.n2091 VSS 0.003719f
C8392 VDPWR.n2092 VSS 0.001668f
C8393 VDPWR.n2093 VSS 0.002085f
C8394 VDPWR.n2094 VSS 9.8e-19
C8395 VDPWR.n2095 VSS 0.001808f
C8396 VDPWR.t12 VSS 0.002606f
C8397 VDPWR.t688 VSS 0.001972f
C8398 VDPWR.n2096 VSS 0.004954f
C8399 VDPWR.n2097 VSS 0.009868f
C8400 VDPWR.n2098 VSS 0.001736f
C8401 VDPWR.n2099 VSS 0.00622f
C8402 VDPWR.n2100 VSS 0.004665f
C8403 VDPWR.n2101 VSS 1.56e-19
C8404 VDPWR.n2102 VSS 0.004702f
C8405 VDPWR.n2103 VSS 0.001748f
C8406 VDPWR.t87 VSS 0.001217f
C8407 VDPWR.t286 VSS 0.001217f
C8408 VDPWR.n2104 VSS 0.002534f
C8409 VDPWR.n2105 VSS 0.007075f
C8410 VDPWR.n2106 VSS 0.005646f
C8411 VDPWR.n2107 VSS 0.00213f
C8412 VDPWR.n2108 VSS 0.003685f
C8413 VDPWR.n2109 VSS 0.00778f
C8414 VDPWR.t1065 VSS 0.005792f
C8415 VDPWR.n2110 VSS 0.012671f
C8416 VDPWR.n2111 VSS 0.021249f
C8417 VDPWR.n2112 VSS 0.016474f
C8418 VDPWR.n2113 VSS 0.00622f
C8419 VDPWR.n2114 VSS 0.004665f
C8420 VDPWR.n2115 VSS 0.009456f
C8421 VDPWR.n2116 VSS 0.017714f
C8422 VDPWR.n2117 VSS 0.003347f
C8423 VDPWR.n2118 VSS 5.79e-19
C8424 VDPWR.n2119 VSS 0.003257f
C8425 VDPWR.n2120 VSS 0.003595f
C8426 VDPWR.n2121 VSS 0.003719f
C8427 VDPWR.n2122 VSS 0.003719f
C8428 VDPWR.n2123 VSS 0.003595f
C8429 VDPWR.n2124 VSS 0.003257f
C8430 VDPWR.n2125 VSS 0.002912f
C8431 VDPWR.n2126 VSS 0.003854f
C8432 VDPWR.n2127 VSS 0.010328f
C8433 VDPWR.n2128 VSS 0.013477f
C8434 VDPWR.n2129 VSS 0.013038f
C8435 VDPWR.n2130 VSS 0.00622f
C8436 VDPWR.n2131 VSS 0.005646f
C8437 VDPWR.n2132 VSS 0.006081f
C8438 VDPWR.n2133 VSS 0.00613f
C8439 VDPWR.n2134 VSS 0.003685f
C8440 VDPWR.n2135 VSS 0.00622f
C8441 VDPWR.n2136 VSS 0.010328f
C8442 VDPWR.n2137 VSS 0.013477f
C8443 VDPWR.n2138 VSS 0.013038f
C8444 VDPWR.n2139 VSS 0.00622f
C8445 VDPWR.n2140 VSS 0.005646f
C8446 VDPWR.n2141 VSS 0.003685f
C8447 VDPWR.n2142 VSS 0.00613f
C8448 VDPWR.t1156 VSS 0.005792f
C8449 VDPWR.n2143 VSS 0.007319f
C8450 VDPWR.n2144 VSS 0.013038f
C8451 VDPWR.n2145 VSS 0.009888f
C8452 VDPWR.n2146 VSS 0.004124f
C8453 VDPWR.n2147 VSS 0.003115f
C8454 VDPWR.n2148 VSS 0.003257f
C8455 VDPWR.n2149 VSS 0.003595f
C8456 VDPWR.n2150 VSS 0.003719f
C8457 VDPWR.n2151 VSS 0.003719f
C8458 VDPWR.n2152 VSS 0.003595f
C8459 VDPWR.n2153 VSS 0.003257f
C8460 VDPWR.n2154 VSS 0.003115f
C8461 VDPWR.n2155 VSS 0.004327f
C8462 VDPWR.n2156 VSS 0.005928f
C8463 VDPWR.n2157 VSS 0.009235f
C8464 VDPWR.n2158 VSS 0.003685f
C8465 VDPWR.n2159 VSS 0.00622f
C8466 VDPWR.n2160 VSS 0.00622f
C8467 VDPWR.n2161 VSS 0.021966f
C8468 VDPWR.n2162 VSS 0.021249f
C8469 VDPWR.t1155 VSS 0.005792f
C8470 VDPWR.n2163 VSS 0.011204f
C8471 VDPWR.n2164 VSS 0.0143f
C8472 VDPWR.t853 VSS 0.005265f
C8473 VDPWR.n2165 VSS 0.031587f
C8474 VDPWR.t1249 VSS 0.018514f
C8475 VDPWR.n2166 VSS 0.035885f
C8476 VDPWR.n2167 VSS 0.008189f
C8477 VDPWR.n2168 VSS 0.001833f
C8478 VDPWR.n2169 VSS 0.010417f
C8479 VDPWR.n2170 VSS 0.005646f
C8480 VDPWR.n2171 VSS 0.005232f
C8481 VDPWR.n2172 VSS 0.003347f
C8482 VDPWR.n2173 VSS 0.002671f
C8483 VDPWR.n2174 VSS 0.006356f
C8484 VDPWR.t966 VSS 0.005792f
C8485 VDPWR.n2175 VSS 0.007319f
C8486 VDPWR.n2176 VSS 0.013038f
C8487 VDPWR.n2177 VSS 0.002164f
C8488 VDPWR.n2178 VSS 0.00311f
C8489 VDPWR.n2179 VSS 0.002085f
C8490 VDPWR.n2180 VSS 0.003719f
C8491 VDPWR.n2181 VSS 0.001668f
C8492 VDPWR.n2182 VSS 0.002085f
C8493 VDPWR.n2183 VSS 0.002366f
C8494 VDPWR.n2184 VSS 0.002907f
C8495 VDPWR.n2185 VSS 0.002085f
C8496 VDPWR.n2186 VSS 0.003257f
C8497 VDPWR.n2187 VSS 0.003595f
C8498 VDPWR.n2188 VSS 0.245208f
C8499 VDPWR.n2189 VSS 0.003719f
C8500 VDPWR.n2190 VSS 0.003115f
C8501 VDPWR.n2191 VSS 0.001668f
C8502 VDPWR.t1279 VSS 0.076721f
C8503 VDPWR.n2192 VSS 0.038654f
C8504 VDPWR.n2193 VSS 0.00622f
C8505 VDPWR.t1209 VSS 0.076721f
C8506 VDPWR.n2194 VSS 0.038215f
C8507 VDPWR.t899 VSS 0.005792f
C8508 VDPWR.n2195 VSS 0.007319f
C8509 VDPWR.n2196 VSS 0.004665f
C8510 VDPWR.t963 VSS 0.005265f
C8511 VDPWR.n2197 VSS 0.012091f
C8512 VDPWR.n2198 VSS 0.00622f
C8513 VDPWR.n2199 VSS 0.016116f
C8514 VDPWR.n2200 VSS 0.003043f
C8515 VDPWR.n2201 VSS 0.002085f
C8516 VDPWR.n2202 VSS 0.003719f
C8517 VDPWR.n2203 VSS 0.001668f
C8518 VDPWR.n2204 VSS 0.002502f
C8519 VDPWR.t1243 VSS 0.038955f
C8520 VDPWR.t962 VSS 0.005265f
C8521 VDPWR.n2205 VSS 0.012091f
C8522 VDPWR.t1085 VSS 0.005389f
C8523 VDPWR.n2206 VSS 0.002259f
C8524 VDPWR.n2207 VSS 0.012313f
C8525 VDPWR.t1188 VSS 0.011303f
C8526 VDPWR.n2208 VSS 0.021734f
C8527 VDPWR.t1084 VSS 0.005308f
C8528 VDPWR.n2209 VSS 0.007681f
C8529 VDPWR.n2210 VSS 0.007573f
C8530 VDPWR.t931 VSS 0.005308f
C8531 VDPWR.t1254 VSS 0.011265f
C8532 VDPWR.n2212 VSS 0.028883f
C8533 VDPWR.t932 VSS 0.005308f
C8534 VDPWR.n2213 VSS 0.015733f
C8535 VDPWR.t1040 VSS 0.005308f
C8536 VDPWR.t1183 VSS 0.011265f
C8537 VDPWR.n2215 VSS 0.028883f
C8538 VDPWR.t1041 VSS 0.005308f
C8539 VDPWR.n2216 VSS 0.015733f
C8540 VDPWR.n2217 VSS 0.012962f
C8541 VDPWR.n2218 VSS 0.004061f
C8542 VDPWR.n2219 VSS 0.003721f
C8543 VDPWR.n2220 VSS 0.00213f
C8544 VDPWR.n2221 VSS 0.002918f
C8545 VDPWR.t898 VSS 0.005813f
C8546 VDPWR.n2222 VSS 0.006446f
C8547 VDPWR.n2223 VSS 0.007942f
C8548 VDPWR.n2224 VSS 0.004665f
C8549 VDPWR.n2225 VSS 0.002085f
C8550 VDPWR.n2226 VSS 0.003595f
C8551 VDPWR.n2227 VSS 0.003257f
C8552 VDPWR.n2228 VSS 0.002777f
C8553 VDPWR.n2229 VSS 0.003719f
C8554 VDPWR.n2230 VSS 0.015997f
C8555 VDPWR.n2231 VSS 0.055357f
C8556 VDPWR.t1238 VSS 0.076721f
C8557 VDPWR.n2232 VSS 0.042898f
C8558 VDPWR.n2233 VSS 0.011102f
C8559 VDPWR.n2234 VSS 0.002164f
C8560 VDPWR.n2235 VSS 0.002164f
C8561 VDPWR.n2236 VSS 0.00311f
C8562 VDPWR.n2237 VSS 0.002085f
C8563 VDPWR.n2238 VSS 0.001668f
C8564 VDPWR.n2239 VSS 0.003719f
C8565 VDPWR.n2240 VSS 0.003595f
C8566 VDPWR.n2241 VSS 0.003257f
C8567 VDPWR.n2242 VSS 0.002236f
C8568 VDPWR.n2243 VSS 0.003178f
C8569 VDPWR.n2244 VSS 0.021966f
C8570 VDPWR.n2245 VSS 0.021966f
C8571 VDPWR.n2246 VSS 0.021249f
C8572 VDPWR.n2247 VSS 0.00622f
C8573 VDPWR.n2248 VSS 0.003685f
C8574 VDPWR.n2249 VSS 0.009235f
C8575 VDPWR.n2250 VSS 0.005928f
C8576 VDPWR.t1046 VSS 0.005792f
C8577 VDPWR.n2251 VSS 0.007319f
C8578 VDPWR.n2252 VSS 0.012598f
C8579 VDPWR.n2253 VSS 0.00622f
C8580 VDPWR.n2254 VSS 0.003685f
C8581 VDPWR.n2255 VSS 0.00613f
C8582 VDPWR.t1110 VSS 0.005792f
C8583 VDPWR.n2256 VSS 0.004169f
C8584 VDPWR.n2257 VSS 0.006081f
C8585 VDPWR.n2258 VSS 0.005646f
C8586 VDPWR.n2259 VSS 0.00622f
C8587 VDPWR.n2260 VSS 0.009888f
C8588 VDPWR.n2261 VSS 0.013477f
C8589 VDPWR.n2262 VSS 0.010328f
C8590 VDPWR.n2263 VSS 0.00622f
C8591 VDPWR.n2264 VSS 0.0048f
C8592 VDPWR.n2265 VSS 0.009888f
C8593 VDPWR.n2266 VSS 0.013477f
C8594 VDPWR.n2267 VSS 0.002164f
C8595 VDPWR.n2268 VSS 0.002085f
C8596 VDPWR.n2269 VSS 0.002366f
C8597 VDPWR.n2270 VSS 0.002907f
C8598 VDPWR.n2271 VSS 0.002085f
C8599 VDPWR.n2272 VSS 0.003257f
C8600 VDPWR.n2273 VSS 0.003595f
C8601 VDPWR.n2274 VSS 0.245208f
C8602 VDPWR.n2275 VSS 0.003595f
C8603 VDPWR.n2276 VSS 0.003257f
C8604 VDPWR.n2277 VSS 0.002085f
C8605 VDPWR.n2278 VSS 0.00311f
C8606 VDPWR.n2279 VSS 0.002164f
C8607 VDPWR.n2280 VSS 0.013038f
C8608 VDPWR.t1047 VSS 0.005792f
C8609 VDPWR.n2281 VSS 0.007319f
C8610 VDPWR.n2282 VSS 0.006356f
C8611 VDPWR.n2283 VSS 0.002671f
C8612 VDPWR.n2284 VSS 0.003347f
C8613 VDPWR.n2285 VSS 0.002366f
C8614 VDPWR.n2286 VSS 0.006604f
C8615 VDPWR.t1111 VSS 0.005813f
C8616 VDPWR.n2287 VSS 0.006593f
C8617 VDPWR.n2288 VSS 0.002451f
C8618 VDPWR.n2289 VSS 0.00213f
C8619 VDPWR.n2290 VSS 0.00311f
C8620 VDPWR.n2291 VSS 0.001775f
C8621 VDPWR.n2292 VSS 0.015074f
C8622 VDPWR.t63 VSS 0.001972f
C8623 VDPWR.t476 VSS 0.001972f
C8624 VDPWR.n2293 VSS 0.004238f
C8625 VDPWR.t969 VSS 0.005265f
C8626 VDPWR.n2294 VSS 0.014912f
C8627 VDPWR.n2295 VSS 0.01553f
C8628 VDPWR.n2296 VSS 0.005646f
C8629 VDPWR.n2297 VSS 0.003685f
C8630 VDPWR.n2298 VSS 0.004665f
C8631 VDPWR.n2299 VSS 0.00304f
C8632 VDPWR.t838 VSS 0.005792f
C8633 VDPWR.n2300 VSS 0.003731f
C8634 VDPWR.n2301 VSS 0.009231f
C8635 VDPWR.n2302 VSS 0.004726f
C8636 VDPWR.n2303 VSS 0.006616f
C8637 VDPWR.n2304 VSS 0.00622f
C8638 VDPWR.n2305 VSS 0.005882f
C8639 VDPWR.n2306 VSS 0.003394f
C8640 VDPWR.n2307 VSS 0.035868f
C8641 VDPWR.n2308 VSS 0.003995f
C8642 VDPWR.n2309 VSS 0.009136f
C8643 VDPWR.t794 VSS 0.001972f
C8644 VDPWR.t816 VSS 0.001972f
C8645 VDPWR.n2310 VSS 0.004071f
C8646 VDPWR.n2311 VSS 0.009136f
C8647 VDPWR.n2312 VSS 0.005585f
C8648 VDPWR.n2313 VSS 0.005757f
C8649 VDPWR.n2314 VSS 0.002164f
C8650 VDPWR.n2315 VSS 0.00311f
C8651 VDPWR.n2316 VSS 0.002085f
C8652 VDPWR.n2317 VSS 0.003257f
C8653 VDPWR.n2318 VSS 0.003595f
C8654 VDPWR.n2319 VSS 0.245208f
C8655 VDPWR.n2320 VSS 0.003595f
C8656 VDPWR.n2321 VSS 0.003257f
C8657 VDPWR.n2322 VSS 0.003115f
C8658 VDPWR.n2323 VSS 0.004124f
C8659 VDPWR.n2324 VSS 0.00622f
C8660 VDPWR.n2325 VSS 0.005027f
C8661 VDPWR.n2326 VSS 0.00883f
C8662 VDPWR.n2327 VSS 0.006831f
C8663 VDPWR.t796 VSS 0.001972f
C8664 VDPWR.t806 VSS 0.001972f
C8665 VDPWR.n2328 VSS 0.004071f
C8666 VDPWR.n2329 VSS 0.008572f
C8667 VDPWR.n2330 VSS 0.004511f
C8668 VDPWR.n2331 VSS 0.00622f
C8669 VDPWR.n2332 VSS 0.003685f
C8670 VDPWR.n2333 VSS 0.003165f
C8671 VDPWR.n2334 VSS 0.002896f
C8672 VDPWR.n2335 VSS 0.005135f
C8673 VDPWR.t1142 VSS 0.005792f
C8674 VDPWR.n2336 VSS 0.00449f
C8675 VDPWR.n2337 VSS 0.007218f
C8676 VDPWR.n2338 VSS 0.00622f
C8677 VDPWR.n2339 VSS 0.00622f
C8678 VDPWR.n2340 VSS 0.004364f
C8679 VDPWR.n2341 VSS 0.006004f
C8680 VDPWR.n2342 VSS 0.035153f
C8681 VDPWR.n2343 VSS 0.008035f
C8682 VDPWR.n2344 VSS 0.004602f
C8683 VDPWR.n2345 VSS 0.004665f
C8684 VDPWR.n2346 VSS 0.002366f
C8685 VDPWR.n2347 VSS 0.002299f
C8686 VDPWR.n2348 VSS 0.009456f
C8687 VDPWR.t1133 VSS 0.005265f
C8688 VDPWR.n2349 VSS 0.006599f
C8689 VDPWR.n2350 VSS 0.022507f
C8690 VDPWR.n2351 VSS 0.002164f
C8691 VDPWR.n2352 VSS 0.021249f
C8692 VDPWR.n2353 VSS 0.016474f
C8693 VDPWR.n2354 VSS 0.002164f
C8694 VDPWR.n2355 VSS 0.002366f
C8695 VDPWR.n2356 VSS 0.002085f
C8696 VDPWR.n2357 VSS 0.003257f
C8697 VDPWR.n2358 VSS 0.003595f
C8698 VDPWR.n2359 VSS 0.245208f
C8699 VDPWR.n2360 VSS 0.003595f
C8700 VDPWR.n2361 VSS 0.003257f
C8701 VDPWR.n2362 VSS 5.79e-19
C8702 VDPWR.n2363 VSS 0.002164f
C8703 VDPWR.n2364 VSS 0.009456f
C8704 VDPWR.n2365 VSS 0.017679f
C8705 VDPWR.n2366 VSS 0.002366f
C8706 VDPWR.n2367 VSS 0.00213f
C8707 VDPWR.n2368 VSS 0.00313f
C8708 VDPWR.t494 VSS 0.007287f
C8709 VDPWR.n2369 VSS 0.007165f
C8710 VDPWR.n2370 VSS 0.002948f
C8711 VDPWR.n2371 VSS 0.00213f
C8712 VDPWR.n2372 VSS 0.005646f
C8713 VDPWR.n2373 VSS 0.007329f
C8714 VDPWR.n2374 VSS 0.00956f
C8715 VDPWR.n2375 VSS 0.004176f
C8716 VDPWR.t492 VSS 0.001972f
C8717 VDPWR.t294 VSS 0.001972f
C8718 VDPWR.n2376 VSS 0.004228f
C8719 VDPWR.n2377 VSS 0.008964f
C8720 VDPWR.t1216 VSS 0.077619f
C8721 VDPWR.n2378 VSS 0.03183f
C8722 VDPWR.n2379 VSS 0.00678f
C8723 VDPWR.n2380 VSS 0.00622f
C8724 VDPWR.n2381 VSS 0.00622f
C8725 VDPWR.n2382 VSS 0.00622f
C8726 VDPWR.n2383 VSS 0.006616f
C8727 VDPWR.n2384 VSS 0.009136f
C8728 VDPWR.n2385 VSS 0.005241f
C8729 VDPWR.n2386 VSS 0.006101f
C8730 VDPWR.n2387 VSS 0.00622f
C8731 VDPWR.n2388 VSS 0.004936f
C8732 VDPWR.n2389 VSS 0.005757f
C8733 VDPWR.t302 VSS 0.001972f
C8734 VDPWR.t306 VSS 0.001972f
C8735 VDPWR.n2390 VSS 0.004071f
C8736 VDPWR.n2391 VSS 0.006015f
C8737 VDPWR.n2392 VSS 0.009136f
C8738 VDPWR.n2393 VSS 0.005585f
C8739 VDPWR.n2394 VSS 0.002164f
C8740 VDPWR.n2395 VSS 0.002085f
C8741 VDPWR.n2396 VSS 0.002231f
C8742 VDPWR.n2397 VSS 0.003043f
C8743 VDPWR.n2398 VSS 0.002085f
C8744 VDPWR.n2399 VSS 0.003227f
C8745 VDPWR.n2400 VSS 0.003626f
C8746 VDPWR.n2401 VSS 0.245208f
C8747 VDPWR.n2402 VSS 0.003626f
C8748 VDPWR.n2403 VSS 0.003227f
C8749 VDPWR.n2404 VSS 0.002085f
C8750 VDPWR.n2405 VSS 0.00311f
C8751 VDPWR.n2406 VSS 0.001589f
C8752 VDPWR.n2407 VSS 0.001396f
C8753 VDPWR.n2408 VSS 0.007166f
C8754 VDPWR.n2409 VSS 0.002578f
C8755 VDPWR.n2410 VSS 0.005071f
C8756 VDPWR.n2411 VSS 0.00622f
C8757 VDPWR.n2412 VSS 0.004253f
C8758 VDPWR.n2413 VSS 0.00883f
C8759 VDPWR.n2414 VSS 0.007347f
C8760 VDPWR.t292 VSS 0.001972f
C8761 VDPWR.t316 VSS 0.001972f
C8762 VDPWR.n2415 VSS 0.004071f
C8763 VDPWR.n2416 VSS 0.006982f
C8764 VDPWR.n2417 VSS 0.003995f
C8765 VDPWR.n2418 VSS 0.00622f
C8766 VDPWR.n2419 VSS 0.00622f
C8767 VDPWR.n2420 VSS 0.00537f
C8768 VDPWR.n2421 VSS 0.009034f
C8769 VDPWR.n2422 VSS 0.004364f
C8770 VDPWR.t314 VSS 0.006928f
C8771 VDPWR.n2423 VSS 0.010124f
C8772 VDPWR.n2424 VSS 0.007155f
C8773 VDPWR.n2425 VSS 0.00622f
C8774 VDPWR.n2426 VSS 0.004665f
C8775 VDPWR.n2427 VSS 0.004665f
C8776 VDPWR.n2428 VSS 0.009456f
C8777 VDPWR.t1102 VSS 0.005265f
C8778 VDPWR.n2429 VSS 0.006599f
C8779 VDPWR.n2430 VSS 0.022507f
C8780 VDPWR.n2431 VSS 0.016474f
C8781 VDPWR.t1103 VSS 0.005265f
C8782 VDPWR.t996 VSS 0.005792f
C8783 VDPWR.n2432 VSS 0.012671f
C8784 VDPWR.n2433 VSS 0.021249f
C8785 VDPWR.n2434 VSS 0.006018f
C8786 VDPWR.n2435 VSS 7.78e-19
C8787 VDPWR.n2436 VSS 0.003115f
C8788 VDPWR.n2437 VSS 0.003257f
C8789 VDPWR.n2438 VSS 0.001668f
C8790 VDPWR.n2439 VSS 0.002085f
C8791 VDPWR.n2440 VSS 0.001555f
C8792 VDPWR.n2441 VSS 0.00311f
C8793 VDPWR.n2442 VSS 0.002164f
C8794 VDPWR.t1097 VSS 0.005308f
C8795 VDPWR.t1167 VSS 0.011265f
C8796 VDPWR.n2444 VSS 0.028883f
C8797 VDPWR.t1098 VSS 0.005308f
C8798 VDPWR.n2445 VSS 0.015733f
C8799 VDPWR.n2446 VSS 0.013258f
C8800 VDPWR.n2447 VSS 0.001454f
C8801 VDPWR.n2448 VSS 0.003047f
C8802 VDPWR.n2449 VSS 0.002231f
C8803 VDPWR.n2450 VSS 0.002085f
C8804 VDPWR.n2451 VSS 0.001668f
C8805 VDPWR.n2452 VSS 0.003719f
C8806 VDPWR.n2453 VSS 0.003595f
C8807 VDPWR.n2454 VSS 0.248273f
C8808 VDPWR.n2455 VSS 0.248273f
C8809 VDPWR.n2456 VSS 0.003719f
C8810 VDPWR.n2457 VSS 0.001668f
C8811 VDPWR.n2458 VSS 0.001555f
C8812 VDPWR.n2459 VSS 0.002164f
C8813 VDPWR.n2460 VSS 0.002231f
C8814 VDPWR.t869 VSS 0.005265f
C8815 VDPWR.t1094 VSS 0.005792f
C8816 VDPWR.n2461 VSS 0.012671f
C8817 VDPWR.n2462 VSS 0.007742f
C8818 VDPWR.t1081 VSS 0.005308f
C8819 VDPWR.t1190 VSS 0.011265f
C8820 VDPWR.n2464 VSS 0.028883f
C8821 VDPWR.t1082 VSS 0.005308f
C8822 VDPWR.n2465 VSS 0.015733f
C8823 VDPWR.t850 VSS 0.005308f
C8824 VDPWR.t1253 VSS 0.011265f
C8825 VDPWR.n2467 VSS 0.028883f
C8826 VDPWR.t851 VSS 0.005308f
C8827 VDPWR.n2468 VSS 0.015733f
C8828 VDPWR.n2469 VSS 0.002085f
C8829 VDPWR.n2470 VSS 0.003595f
C8830 VDPWR.n2471 VSS 0.003257f
C8831 VDPWR.n2472 VSS 0.003047f
C8832 VDPWR.n2473 VSS 0.001454f
C8833 VDPWR.n2474 VSS 0.013258f
C8834 VDPWR.n2475 VSS 0.002164f
C8835 VDPWR.n2476 VSS 0.00311f
C8836 VDPWR.n2477 VSS 0.002085f
C8837 VDPWR.n2478 VSS 0.001668f
C8838 VDPWR.n2479 VSS 0.003719f
C8839 VDPWR.n2480 VSS 0.003595f
C8840 VDPWR.n2481 VSS 0.003257f
C8841 VDPWR.n2482 VSS 0.003115f
C8842 VDPWR.n2483 VSS 0.006018f
C8843 VDPWR.n2484 VSS 0.00622f
C8844 VDPWR.n2485 VSS 0.021966f
C8845 VDPWR.n2486 VSS 0.021966f
C8846 VDPWR.n2487 VSS 0.047471f
C8847 VDPWR.n2488 VSS 0.00622f
C8848 VDPWR.n2489 VSS 0.004665f
C8849 VDPWR.n2490 VSS 0.009456f
C8850 VDPWR.n2491 VSS 0.007471f
C8851 VDPWR.n2492 VSS 0.005752f
C8852 VDPWR.n2493 VSS 0.00622f
C8853 VDPWR.n2494 VSS 0.004665f
C8854 VDPWR.n2495 VSS 0.003685f
C8855 VDPWR.n2496 VSS 0.007755f
C8856 VDPWR.n2497 VSS 0.008496f
C8857 VDPWR.n2498 VSS 0.00375f
C8858 VDPWR.t1093 VSS 0.005792f
C8859 VDPWR.n2499 VSS 0.0045f
C8860 VDPWR.n2500 VSS 0.002941f
C8861 VDPWR.n2501 VSS 0.005071f
C8862 VDPWR.n2502 VSS 0.00254f
C8863 VDPWR.n2503 VSS 0.003257f
C8864 VDPWR.n2504 VSS 0.003595f
C8865 VDPWR.n2505 VSS 0.003719f
C8866 VDPWR.n2506 VSS 0.003595f
C8867 VDPWR.n2507 VSS 0.003719f
C8868 VDPWR.n2508 VSS 0.001668f
C8869 VDPWR.n2509 VSS 0.002085f
C8870 VDPWR.n2510 VSS 0.003043f
C8871 VDPWR.n2511 VSS 0.002164f
C8872 VDPWR.n2512 VSS 0.00784f
C8873 VDPWR.n2513 VSS 0.00784f
C8874 VDPWR.n2514 VSS 0.006008f
C8875 VDPWR.n2515 VSS 0.00622f
C8876 VDPWR.n2516 VSS 0.00622f
C8877 VDPWR.n2517 VSS 0.005752f
C8878 VDPWR.n2518 VSS 0.00784f
C8879 VDPWR.n2519 VSS 0.005752f
C8880 VDPWR.n2520 VSS 0.00622f
C8881 VDPWR.n2521 VSS 0.00622f
C8882 VDPWR.n2522 VSS 0.005112f
C8883 VDPWR.n2523 VSS 0.008523f
C8884 VDPWR.n2524 VSS 0.004815f
C8885 VDPWR.n2525 VSS 0.007499f
C8886 VDPWR.n2526 VSS 0.00622f
C8887 VDPWR.n2527 VSS 0.004665f
C8888 VDPWR.n2528 VSS 0.0024f
C8889 VDPWR.n2529 VSS 0.001735f
C8890 VDPWR.n2530 VSS 0.013131f
C8891 VDPWR.t849 VSS 0.055011f
C8892 VDPWR.t867 VSS 0.104242f
C8893 VDPWR.t1092 VSS 0.060991f
C8894 VDPWR.t490 VSS 0.027107f
C8895 VDPWR.t637 VSS 0.042056f
C8896 VDPWR.t58 VSS 0.02631f
C8897 VDPWR.t561 VSS 0.042056f
C8898 VDPWR.t578 VSS 0.0291f
C8899 VDPWR.t514 VSS 0.035877f
C8900 VDPWR.t563 VSS 0.039465f
C8901 VDPWR.t71 VSS 0.046839f
C8902 VDPWR.t69 VSS 0.035678f
C8903 VDPWR.t1119 VSS 0.018935f
C8904 VDPWR.t564 VSS 0.02631f
C8905 VDPWR.t513 VSS 0.039465f
C8906 VDPWR.t92 VSS 0.064578f
C8907 VDPWR.t565 VSS 0.058599f
C8908 VDPWR.t90 VSS 0.024715f
C8909 VDPWR.n2531 VSS 0.040309f
C8910 VDPWR.t819 VSS 0.030894f
C8911 VDPWR.t906 VSS 0.019533f
C8912 VDPWR.t95 VSS 0.019134f
C8913 VDPWR.t693 VSS 0.041258f
C8914 VDPWR.t199 VSS 0.039066f
C8915 VDPWR.t77 VSS 0.039465f
C8916 VDPWR.t222 VSS 0.014351f
C8917 VDPWR.t821 VSS 0.016743f
C8918 VDPWR.t603 VSS 0.019134f
C8919 VDPWR.t569 VSS 0.041856f
C8920 VDPWR.t224 VSS 0.045045f
C8921 VDPWR.t731 VSS 0.022722f
C8922 VDPWR.t606 VSS 0.022523f
C8923 VDPWR.t410 VSS 0.013753f
C8924 VDPWR.t237 VSS 0.021925f
C8925 VDPWR.t779 VSS 0.028303f
C8926 VDPWR.t733 VSS 0.023719f
C8927 VDPWR.t165 VSS 0.016942f
C8928 VDPWR.t446 VSS 0.018736f
C8929 VDPWR.t364 VSS 0.02053f
C8930 VDPWR.t234 VSS 0.02332f
C8931 VDPWR.t605 VSS 0.030495f
C8932 VDPWR.t592 VSS 0.016942f
C8933 VDPWR.t770 VSS 0.021925f
C8934 VDPWR.t719 VSS 0.035877f
C8935 VDPWR.t600 VSS 0.020928f
C8936 VDPWR.t235 VSS 0.005979f
C8937 VDPWR.t537 VSS 0.018536f
C8938 VDPWR.t741 VSS 0.026908f
C8939 VDPWR.t743 VSS 0.018138f
C8940 VDPWR.t268 VSS 0.017141f
C8941 VDPWR.t739 VSS 0.01754f
C8942 VDPWR.t201 VSS 0.007574f
C8943 VDPWR.t495 VSS 0.018138f
C8944 VDPWR.t386 VSS 0.025712f
C8945 VDPWR.t384 VSS 0.031691f
C8946 VDPWR.n2532 VSS 0.020387f
C8947 VDPWR.n2533 VSS 0.011966f
C8948 VDPWR.n2534 VSS 0.001195f
C8949 VDPWR.n2535 VSS 0.002671f
C8950 VDPWR.n2536 VSS 0.003115f
C8951 VDPWR.n2537 VSS 0.003257f
C8952 VDPWR.n2538 VSS 0.003595f
C8953 VDPWR.n2539 VSS 0.003719f
C8954 VDPWR.n2540 VSS 0.003595f
C8955 VDPWR.n2541 VSS 0.003719f
C8956 VDPWR.n2542 VSS 0.001668f
C8957 VDPWR.n2543 VSS 0.002085f
C8958 VDPWR.n2544 VSS 0.002907f
C8959 VDPWR.n2545 VSS 0.002164f
C8960 VDPWR.n2546 VSS 0.001799f
C8961 VDPWR.n2547 VSS 0.00143f
C8962 VDPWR.n2548 VSS 0.005839f
C8963 VDPWR.n2549 VSS 0.007983f
C8964 VDPWR.n2550 VSS 0.001158f
C8965 VDPWR.n2551 VSS 0.00622f
C8966 VDPWR.n2552 VSS 0.004682f
C8967 VDPWR.n2553 VSS 0.003685f
C8968 VDPWR.n2554 VSS 0.00138f
C8969 VDPWR.n2555 VSS 0.007116f
C8970 VDPWR.n2556 VSS 0.001442f
C8971 VDPWR.n2557 VSS 0.006361f
C8972 VDPWR.t7 VSS 0.004499f
C8973 VDPWR.n2558 VSS 0.004141f
C8974 VDPWR.t678 VSS 0.001094f
C8975 VDPWR.n2559 VSS 0.003115f
C8976 VDPWR.n2560 VSS 0.006107f
C8977 VDPWR.n2561 VSS 0.00622f
C8978 VDPWR.n2562 VSS 0.00622f
C8979 VDPWR.n2563 VSS 0.002588f
C8980 VDPWR.n2564 VSS 0.00885f
C8981 VDPWR.n2565 VSS 0.006078f
C8982 VDPWR.n2566 VSS 0.003685f
C8983 VDPWR.n2567 VSS 0.005646f
C8984 VDPWR.n2568 VSS 0.02258f
C8985 VDPWR.n2569 VSS 0.013755f
C8986 VDPWR.n2570 VSS 6.42e-19
C8987 VDPWR.n2571 VSS 0.00156f
C8988 VDPWR.n2572 VSS 0.003257f
C8989 VDPWR.n2573 VSS 0.002085f
C8990 VDPWR.n2574 VSS 9.8e-19
C8991 VDPWR.n2575 VSS 0.001859f
C8992 VDPWR.n2576 VSS 0.022802f
C8993 VDPWR.n2577 VSS 0.002164f
C8994 VDPWR.n2578 VSS 0.002502f
C8995 VDPWR.n2579 VSS 0.002085f
C8996 VDPWR.n2580 VSS 0.003257f
C8997 VDPWR.n2581 VSS 0.003595f
C8998 VDPWR.n2582 VSS 0.245208f
C8999 VDPWR.n2584 VSS 0.003719f
C9000 VDPWR.n2585 VSS 0.002777f
C9001 VDPWR.n2586 VSS 0.002085f
C9002 VDPWR.n2587 VSS 0.001668f
C9003 VDPWR.t1125 VSS 0.005265f
C9004 VDPWR.t1176 VSS 0.022165f
C9005 VDPWR.n2589 VSS 0.038508f
C9006 VDPWR.t1126 VSS 0.005265f
C9007 VDPWR.n2590 VSS 0.022096f
C9008 VDPWR.t904 VSS 0.005265f
C9009 VDPWR.t1276 VSS 0.022165f
C9010 VDPWR.n2592 VSS 0.038508f
C9011 VDPWR.t905 VSS 0.005265f
C9012 VDPWR.n2593 VSS 0.022096f
C9013 VDPWR.n2594 VSS 0.019039f
C9014 VDPWR.t1112 VSS 0.005308f
C9015 VDPWR.t1179 VSS 0.011265f
C9016 VDPWR.n2596 VSS 0.028883f
C9017 VDPWR.t1113 VSS 0.005308f
C9018 VDPWR.n2597 VSS 0.015733f
C9019 VDPWR.t895 VSS 0.005308f
C9020 VDPWR.t1278 VSS 0.011265f
C9021 VDPWR.n2599 VSS 0.028883f
C9022 VDPWR.t896 VSS 0.005308f
C9023 VDPWR.n2600 VSS 0.015733f
C9024 VDPWR.n2601 VSS 0.012962f
C9025 VDPWR.n2602 VSS 0.004061f
C9026 VDPWR.n2603 VSS 0.007291f
C9027 VDPWR.n2604 VSS 0.002164f
C9028 VDPWR.n2605 VSS 0.001856f
C9029 VDPWR.n2606 VSS 0.001197f
C9030 VDPWR.n2607 VSS 0.002164f
C9031 VDPWR.n2608 VSS 0.002502f
C9032 VDPWR.n2609 VSS 0.002085f
C9033 VDPWR.n2610 VSS 0.003227f
C9034 VDPWR.n2611 VSS 0.003626f
C9035 VDPWR.n2612 VSS 0.132183f
C9036 VDPWR.n2613 VSS 0.310241f
C9037 VDPWR.n2614 VSS 0.130999f
C9038 VDPWR.n2615 VSS 0.001668f
C9039 VDPWR.n2616 VSS 0.001668f
C9040 VDPWR.n2617 VSS 0.003227f
C9041 VDPWR.n2618 VSS 0.451964f
C9042 VDPWR.n2619 VSS 0.002085f
C9043 VDPWR.n2620 VSS 0.003043f
C9044 VDPWR.n2621 VSS 0.004665f
C9045 VDPWR.t1269 VSS 0.021971f
C9046 VDPWR.t826 VSS 0.006676f
C9047 VDPWR.n2622 VSS 0.006469f
C9048 VDPWR.n2623 VSS 0.002085f
C9049 VDPWR.n2624 VSS 0.002502f
C9050 VDPWR.t377 VSS 0.001902f
C9051 VDPWR.t374 VSS 0.001902f
C9052 VDPWR.n2625 VSS 0.004166f
C9053 VDPWR.n2626 VSS 0.002777f
C9054 VDPWR.n2627 VSS 0.003719f
C9055 VDPWR.t169 VSS 0.001614f
C9056 VDPWR.t376 VSS 0.001614f
C9057 VDPWR.n2628 VSS 0.003585f
C9058 VDPWR.n2629 VSS 0.001808f
C9059 VDPWR.t129 VSS 0.001614f
C9060 VDPWR.t353 VSS 0.001614f
C9061 VDPWR.n2630 VSS 0.003585f
C9062 VDPWR.t880 VSS 0.005308f
C9063 VDPWR.t1274 VSS 0.011265f
C9064 VDPWR.n2632 VSS 0.028883f
C9065 VDPWR.t881 VSS 0.005308f
C9066 VDPWR.n2633 VSS 0.015733f
C9067 VDPWR.t999 VSS 0.005308f
C9068 VDPWR.t1211 VSS 0.011265f
C9069 VDPWR.n2635 VSS 0.028883f
C9070 VDPWR.t1000 VSS 0.005308f
C9071 VDPWR.n2636 VSS 0.015733f
C9072 VDPWR.n2637 VSS 0.013309f
C9073 VDPWR.n2638 VSS 0.004061f
C9074 VDPWR.n2639 VSS 0.00213f
C9075 VDPWR.n2640 VSS 0.001461f
C9076 VDPWR.n2641 VSS 0.009701f
C9077 VDPWR.n2642 VSS 0.003381f
C9078 VDPWR.n2643 VSS 0.00213f
C9079 VDPWR.n2644 VSS 0.004665f
C9080 VDPWR.n2645 VSS 0.001808f
C9081 VDPWR.n2646 VSS 0.013409f
C9082 VDPWR.n2647 VSS 0.001509f
C9083 VDPWR.n2648 VSS 9.13e-19
C9084 VDPWR.n2649 VSS 0.002085f
C9085 VDPWR.n2650 VSS 0.001555f
C9086 VDPWR.n2651 VSS 0.002164f
C9087 VDPWR.n2652 VSS 0.003008f
C9088 VDPWR.t844 VSS 0.005265f
C9089 VDPWR.n2653 VSS 0.00519f
C9090 VDPWR.n2654 VSS 0.019873f
C9091 VDPWR.t453 VSS 0.002395f
C9092 VDPWR.t595 VSS 0.002465f
C9093 VDPWR.n2655 VSS 0.005792f
C9094 VDPWR.n2656 VSS 0.009409f
C9095 VDPWR.n2657 VSS 0.004665f
C9096 VDPWR.n2658 VSS 0.006239f
C9097 VDPWR.t1194 VSS 0.030953f
C9098 VDPWR.t1043 VSS 0.005265f
C9099 VDPWR.n2659 VSS 0.009272f
C9100 VDPWR.t127 VSS 0.002895f
C9101 VDPWR.n2660 VSS 0.011931f
C9102 VDPWR.n2661 VSS 0.0048f
C9103 VDPWR.t487 VSS 0.001094f
C9104 VDPWR.t30 VSS 0.001094f
C9105 VDPWR.n2662 VSS 0.002291f
C9106 VDPWR.n2663 VSS 0.001883f
C9107 VDPWR.n2664 VSS 0.003115f
C9108 VDPWR.n2665 VSS 0.003227f
C9109 VDPWR.n2666 VSS 0.002085f
C9110 VDPWR.n2667 VSS 0.003227f
C9111 VDPWR.n2668 VSS 0.001555f
C9112 VDPWR.n2669 VSS 7.78e-19
C9113 VDPWR.n2670 VSS 0.003115f
C9114 VDPWR.t84 VSS 0.001614f
C9115 VDPWR.t761 VSS 0.001614f
C9116 VDPWR.n2671 VSS 0.003509f
C9117 VDPWR.t597 VSS 0.004145f
C9118 VDPWR.t622 VSS 0.003028f
C9119 VDPWR.n2672 VSS 0.010723f
C9120 VDPWR.n2673 VSS 0.008247f
C9121 VDPWR.t879 VSS 0.055011f
C9122 VDPWR.t128 VSS 0.018536f
C9123 VDPWR.t352 VSS 0.018138f
C9124 VDPWR.t824 VSS 0.024516f
C9125 VDPWR.t168 VSS 0.033485f
C9126 VDPWR.t373 VSS 0.01754f
C9127 VDPWR.t375 VSS 0.013753f
C9128 VDPWR.t825 VSS 0.040461f
C9129 VDPWR.t431 VSS 0.039465f
C9130 VDPWR.t843 VSS 0.032887f
C9131 VDPWR.t452 VSS 0.018138f
C9132 VDPWR.t161 VSS 0.007773f
C9133 VDPWR.t594 VSS 0.01754f
C9134 VDPWR.t166 VSS 0.018736f
C9135 VDPWR.t25 VSS 0.021925f
C9136 VDPWR.t153 VSS 0.028104f
C9137 VDPWR.t130 VSS 0.05541f
C9138 VDPWR.t1042 VSS 0.006179f
C9139 VDPWR.t126 VSS 0.02033f
C9140 VDPWR.t486 VSS 0.040661f
C9141 VDPWR.t29 VSS 0.028901f
C9142 VDPWR.t596 VSS 0.018337f
C9143 VDPWR.t83 VSS 0.023719f
C9144 VDPWR.t621 VSS 0.045444f
C9145 VDPWR.t21 VSS 0.020131f
C9146 VDPWR.t635 VSS 0.01754f
C9147 VDPWR.t745 VSS 0.016543f
C9148 VDPWR.t747 VSS 0.018337f
C9149 VDPWR.t762 VSS 0.030894f
C9150 VDPWR.t1138 VSS 0.033286f
C9151 VDPWR.t258 VSS 0.048434f
C9152 VDPWR.t249 VSS 0.023719f
C9153 VDPWR.t915 VSS 0.018337f
C9154 VDPWR.t1075 VSS 0.109823f
C9155 VDPWR.t220 VSS 0.048434f
C9156 VDPWR.t666 VSS 0.018337f
C9157 VDPWR.t672 VSS 0.006179f
C9158 VDPWR.t163 VSS 0.026509f
C9159 VDPWR.t81 VSS 0.03787f
C9160 VDPWR.t670 VSS 0.022722f
C9161 VDPWR.t885 VSS 0.019932f
C9162 VDPWR.t576 VSS 0.024117f
C9163 VDPWR.n2674 VSS 0.056102f
C9164 VDPWR.n2675 VSS 0.023403f
C9165 VDPWR.t1255 VSS 0.030953f
C9166 VDPWR.t577 VSS 0.002895f
C9167 VDPWR.n2676 VSS 0.011931f
C9168 VDPWR.n2677 VSS 0.00622f
C9169 VDPWR.t671 VSS 0.001094f
C9170 VDPWR.t82 VSS 0.001094f
C9171 VDPWR.n2678 VSS 0.002291f
C9172 VDPWR.t887 VSS 0.005265f
C9173 VDPWR.n2679 VSS 0.009272f
C9174 VDPWR.t164 VSS 0.004145f
C9175 VDPWR.t673 VSS 0.003028f
C9176 VDPWR.n2680 VSS 0.010803f
C9177 VDPWR.n2681 VSS 0.00213f
C9178 VDPWR.n2682 VSS 0.004091f
C9179 VDPWR.t667 VSS 0.001614f
C9180 VDPWR.t221 VSS 0.001614f
C9181 VDPWR.n2683 VSS 0.003585f
C9182 VDPWR.n2684 VSS 0.002647f
C9183 VDPWR.n2685 VSS 0.001149f
C9184 VDPWR.n2686 VSS 0.002085f
C9185 VDPWR.n2687 VSS 0.001668f
C9186 VDPWR.n2688 VSS 0.003227f
C9187 VDPWR.n2689 VSS 0.001555f
C9188 VDPWR.n2690 VSS 0.002164f
C9189 VDPWR.n2691 VSS 0.003115f
C9190 VDPWR.t1076 VSS 0.005265f
C9191 VDPWR.t916 VSS 0.005792f
C9192 VDPWR.n2692 VSS 0.012671f
C9193 VDPWR.n2693 VSS 0.004059f
C9194 VDPWR.n2694 VSS 0.003481f
C9195 VDPWR.t1182 VSS 0.030748f
C9196 VDPWR.n2695 VSS 0.01614f
C9197 VDPWR.n2696 VSS 0.016832f
C9198 VDPWR.n2697 VSS 0.003685f
C9199 VDPWR.t1264 VSS 0.076721f
C9200 VDPWR.n2698 VSS 0.042898f
C9201 VDPWR.t250 VSS 0.001614f
C9202 VDPWR.t259 VSS 0.001614f
C9203 VDPWR.n2699 VSS 0.003509f
C9204 VDPWR.n2700 VSS 0.014624f
C9205 VDPWR.t917 VSS 0.005811f
C9206 VDPWR.n2701 VSS 0.011961f
C9207 VDPWR.n2702 VSS 0.00449f
C9208 VDPWR.t748 VSS 0.001598f
C9209 VDPWR.t763 VSS 5.96e-19
C9210 VDPWR.n2703 VSS 0.007345f
C9211 VDPWR.t746 VSS 0.001614f
C9212 VDPWR.t22 VSS 0.001614f
C9213 VDPWR.n2704 VSS 0.003509f
C9214 VDPWR.n2705 VSS 0.00852f
C9215 VDPWR.n2706 VSS 9.85e-19
C9216 VDPWR.n2707 VSS 0.002085f
C9217 VDPWR.n2708 VSS 0.001555f
C9218 VDPWR.n2709 VSS 0.002535f
C9219 VDPWR.n2710 VSS 7.78e-19
C9220 VDPWR.n2711 VSS 0.001305f
C9221 VDPWR.n2712 VSS 0.016368f
C9222 VDPWR.t1140 VSS 0.005343f
C9223 VDPWR.n2713 VSS 0.006246f
C9224 VDPWR.n2714 VSS 0.024304f
C9225 VDPWR.t1280 VSS 0.022315f
C9226 VDPWR.n2715 VSS 0.022091f
C9227 VDPWR.t1139 VSS 0.005265f
C9228 VDPWR.n2716 VSS 0.006338f
C9229 VDPWR.n2717 VSS 0.006286f
C9230 VDPWR.n2718 VSS 0.003323f
C9231 VDPWR.n2719 VSS 0.002366f
C9232 VDPWR.n2720 VSS 0.006604f
C9233 VDPWR.n2721 VSS 0.00784f
C9234 VDPWR.n2722 VSS 0.004665f
C9235 VDPWR.n2723 VSS 0.005646f
C9236 VDPWR.n2724 VSS 0.00213f
C9237 VDPWR.n2725 VSS 0.007471f
C9238 VDPWR.n2726 VSS 0.009456f
C9239 VDPWR.t1077 VSS 0.005265f
C9240 VDPWR.n2727 VSS 0.012091f
C9241 VDPWR.n2728 VSS 0.0154f
C9242 VDPWR.n2729 VSS 0.00622f
C9243 VDPWR.n2730 VSS 0.00622f
C9244 VDPWR.n2731 VSS 0.004124f
C9245 VDPWR.n2732 VSS 0.021846f
C9246 VDPWR.n2733 VSS 0.021271f
C9247 VDPWR.n2734 VSS 0.010386f
C9248 VDPWR.n2735 VSS 0.002164f
C9249 VDPWR.n2736 VSS 0.002085f
C9250 VDPWR.n2737 VSS 0.002231f
C9251 VDPWR.n2738 VSS 0.003043f
C9252 VDPWR.n2739 VSS 0.002085f
C9253 VDPWR.n2740 VSS 0.001668f
C9254 VDPWR.n2741 VSS 0.083366f
C9255 VDPWR.n2742 VSS 0.003227f
C9256 VDPWR.n2743 VSS 0.00156f
C9257 VDPWR.n2744 VSS 0.00311f
C9258 VDPWR.n2745 VSS 0.001808f
C9259 VDPWR.n2746 VSS 0.009474f
C9260 VDPWR.n2747 VSS 0.00986f
C9261 VDPWR.n2748 VSS 0.005328f
C9262 VDPWR.n2749 VSS 0.003685f
C9263 VDPWR.n2750 VSS 0.00622f
C9264 VDPWR.n2751 VSS 0.014376f
C9265 VDPWR.n2752 VSS 0.014756f
C9266 VDPWR.n2753 VSS 0.009584f
C9267 VDPWR.n2754 VSS 0.015796f
C9268 VDPWR.n2755 VSS 0.005646f
C9269 VDPWR.n2756 VSS 0.00213f
C9270 VDPWR.n2757 VSS 0.034386f
C9271 VDPWR.t886 VSS 0.005265f
C9272 VDPWR.n2758 VSS 0.009272f
C9273 VDPWR.n2759 VSS 0.005779f
C9274 VDPWR.n2760 VSS 0.002366f
C9275 VDPWR.n2761 VSS 0.002366f
C9276 VDPWR.n2762 VSS 0.003651f
C9277 VDPWR.n2763 VSS 0.001856f
C9278 VDPWR.n2764 VSS 0.008053f
C9279 VDPWR.n2765 VSS 0.002164f
C9280 VDPWR.n2766 VSS 0.002535f
C9281 VDPWR.n2767 VSS 0.002085f
C9282 VDPWR.n2768 VSS 0.001668f
C9283 VDPWR.n2769 VSS 0.085924f
C9284 VDPWR.n2770 VSS 0.001668f
C9285 VDPWR.n2771 VSS 0.002085f
C9286 VDPWR.n2772 VSS 9.8e-19
C9287 VDPWR.n2773 VSS 0.001995f
C9288 VDPWR.n2774 VSS 0.006239f
C9289 VDPWR.t1044 VSS 0.005265f
C9290 VDPWR.n2775 VSS 0.007852f
C9291 VDPWR.n2776 VSS 0.014223f
C9292 VDPWR.n2777 VSS 0.009584f
C9293 VDPWR.n2778 VSS 0.015796f
C9294 VDPWR.n2779 VSS 0.005646f
C9295 VDPWR.n2780 VSS 0.00213f
C9296 VDPWR.n2781 VSS 0.008697f
C9297 VDPWR.n2782 VSS 0.042017f
C9298 VDPWR.n2783 VSS 0.004665f
C9299 VDPWR.n2784 VSS 0.004665f
C9300 VDPWR.n2785 VSS 0.002366f
C9301 VDPWR.n2786 VSS 0.001488f
C9302 VDPWR.t26 VSS 0.002324f
C9303 VDPWR.t154 VSS 0.002324f
C9304 VDPWR.n2787 VSS 0.004738f
C9305 VDPWR.n2788 VSS 0.006878f
C9306 VDPWR.t162 VSS 0.001614f
C9307 VDPWR.t167 VSS 0.001614f
C9308 VDPWR.n2789 VSS 0.003585f
C9309 VDPWR.n2790 VSS 0.009102f
C9310 VDPWR.n2791 VSS 0.005646f
C9311 VDPWR.n2792 VSS 0.00213f
C9312 VDPWR.n2793 VSS 0.00213f
C9313 VDPWR.n2794 VSS 0.005953f
C9314 VDPWR.t845 VSS 0.005265f
C9315 VDPWR.n2795 VSS 0.009272f
C9316 VDPWR.n2796 VSS 0.015796f
C9317 VDPWR.n2797 VSS 0.012246f
C9318 VDPWR.n2798 VSS 0.003178f
C9319 VDPWR.n2799 VSS 0.002236f
C9320 VDPWR.n2800 VSS 0.003227f
C9321 VDPWR.n2801 VSS 0.259182f
C9322 VDPWR.n2802 VSS 0.12621f
C9323 VDPWR.n2803 VSS 0.245208f
C9324 VDPWR.n2804 VSS 0.003626f
C9325 VDPWR.n2805 VSS 0.003227f
C9326 VDPWR.n2806 VSS 0.002085f
C9327 VDPWR.n2807 VSS 0.003043f
C9328 VDPWR.n2808 VSS 0.002164f
C9329 VDPWR.n2809 VSS 0.001976f
C9330 VDPWR.t123 VSS 0.002994f
C9331 VDPWR.t828 VSS 0.002994f
C9332 VDPWR.n2810 VSS 0.012115f
C9333 VDPWR.n2811 VSS 0.00158f
C9334 VDPWR.n2812 VSS 0.00622f
C9335 VDPWR.n2813 VSS 0.00622f
C9336 VDPWR.n2814 VSS 0.00622f
C9337 VDPWR.n2815 VSS 0.002203f
C9338 VDPWR.n2816 VSS 0.001616f
C9339 VDPWR.n2817 VSS 0.008207f
C9340 VDPWR.n2818 VSS 0.001688f
C9341 VDPWR.n2819 VSS 0.00622f
C9342 VDPWR.n2820 VSS 0.00622f
C9343 VDPWR.n2821 VSS 0.00622f
C9344 VDPWR.n2822 VSS 0.002203f
C9345 VDPWR.n2823 VSS 0.001976f
C9346 VDPWR.t152 VSS 0.002933f
C9347 VDPWR.t257 VSS 0.002933f
C9348 VDPWR.n2824 VSS 0.009993f
C9349 VDPWR.n2825 VSS 0.00622f
C9350 VDPWR.n2826 VSS 0.00622f
C9351 VDPWR.n2827 VSS 0.0048f
C9352 VDPWR.t241 VSS 0.001217f
C9353 VDPWR.t540 VSS 0.001217f
C9354 VDPWR.n2828 VSS 0.002534f
C9355 VDPWR.n2829 VSS 0.01209f
C9356 VDPWR.n2830 VSS 0.001437f
C9357 VDPWR.n2831 VSS 0.001995f
C9358 VDPWR.n2832 VSS 0.00311f
C9359 VDPWR.n2833 VSS 0.002164f
C9360 VDPWR.n2834 VSS 0.001668f
C9361 VDPWR.n2835 VSS 0.002085f
C9362 VDPWR.n2836 VSS 0.001555f
C9363 VDPWR.n2837 VSS 9.8e-19
C9364 VDPWR.n2838 VSS 0.002085f
C9365 VDPWR.n2839 VSS 0.003257f
C9366 VDPWR.n2840 VSS 0.003595f
C9367 VDPWR.n2841 VSS 0.245208f
C9368 VDPWR.n2842 VSS 0.003595f
C9369 VDPWR.n2843 VSS 0.003257f
C9370 VDPWR.n2844 VSS 0.003115f
C9371 VDPWR.n2845 VSS 0.002671f
C9372 VDPWR.n2846 VSS 0.002366f
C9373 VDPWR.t894 VSS 0.079129f
C9374 VDPWR.t903 VSS 0.095074f
C9375 VDPWR.t124 VSS 0.043252f
C9376 VDPWR.t332 VSS 0.058599f
C9377 VDPWR.t122 VSS 0.064578f
C9378 VDPWR.t159 VSS 0.039465f
C9379 VDPWR.t243 VSS 0.035678f
C9380 VDPWR.t270 VSS 0.045245f
C9381 VDPWR.t191 VSS 0.046839f
C9382 VDPWR.t242 VSS 0.039465f
C9383 VDPWR.t160 VSS 0.035877f
C9384 VDPWR.t151 VSS 0.054413f
C9385 VDPWR.t240 VSS 0.054214f
C9386 VDPWR.t539 VSS 0.02631f
C9387 VDPWR.t336 VSS 0.033286f
C9388 VDPWR.t900 VSS 0.016743f
C9389 VDPWR.t141 VSS 0.021726f
C9390 VDPWR.t831 VSS 0.055011f
C9391 VDPWR.t641 VSS 0.030495f
C9392 VDPWR.t692 VSS 0.02033f
C9393 VDPWR.t958 VSS 0.018536f
C9394 VDPWR.t60 VSS 0.02631f
C9395 VDPWR.t1163 VSS 0.042056f
C9396 VDPWR.t586 VSS 0.009567f
C9397 VDPWR.t88 VSS 0.016942f
C9398 VDPWR.t121 VSS 0.016743f
C9399 VDPWR.t508 VSS 0.018935f
C9400 VDPWR.t1162 VSS 0.037471f
C9401 VDPWR.t681 VSS 0.02053f
C9402 VDPWR.t545 VSS 0.016942f
C9403 VDPWR.t512 VSS 0.02631f
C9404 VDPWR.t275 VSS 0.018935f
C9405 VDPWR.t507 VSS 0.018935f
C9406 VDPWR.t1165 VSS 0.02053f
C9407 VDPWR.t99 VSS 0.016743f
C9408 VDPWR.t120 VSS 0.02631f
C9409 VDPWR.t97 VSS 0.022722f
C9410 VDPWR.t193 VSS 0.018935f
C9411 VDPWR.t510 VSS 0.032289f
C9412 VDPWR.t511 VSS 0.02631f
C9413 VDPWR.t277 VSS 0.022722f
C9414 VDPWR.t114 VSS 0.016743f
C9415 VDPWR.t195 VSS 0.041856f
C9416 VDPWR.t319 VSS 0.041059f
C9417 VDPWR.t674 VSS 0.016743f
C9418 VDPWR.t112 VSS 0.037471f
C9419 VDPWR.t721 VSS 0.026509f
C9420 VDPWR.t729 VSS 0.021726f
C9421 VDPWR.t1135 VSS 0.016743f
C9422 VDPWR.t448 VSS 0.025512f
C9423 VDPWR.t85 VSS 0.024516f
C9424 VDPWR.n2847 VSS 0.021773f
C9425 VDPWR.t155 VSS 0.030894f
C9426 VDPWR.t888 VSS 0.016743f
C9427 VDPWR.t27 VSS 0.027506f
C9428 VDPWR.t255 VSS 0.036674f
C9429 VDPWR.t695 VSS 0.018138f
C9430 VDPWR.t503 VSS 0.01455f
C9431 VDPWR.t31 VSS 0.016743f
C9432 VDPWR.t23 VSS 0.018736f
C9433 VDPWR.t501 VSS 0.018536f
C9434 VDPWR.t149 VSS 0.019134f
C9435 VDPWR.t727 VSS 0.018935f
C9436 VDPWR.t157 VSS 0.019134f
C9437 VDPWR.t663 VSS 0.037471f
C9438 VDPWR.t65 VSS 0.038468f
C9439 VDPWR.t541 VSS 0.010165f
C9440 VDPWR.t79 VSS 0.016743f
C9441 VDPWR.t413 VSS 0.018536f
C9442 VDPWR.t664 VSS 0.019134f
C9443 VDPWR.t574 VSS 0.022921f
C9444 VDPWR.t580 VSS 0.018337f
C9445 VDPWR.t829 VSS 0.009567f
C9446 VDPWR.t643 VSS 0.018935f
C9447 VDPWR.t412 VSS 0.037272f
C9448 VDPWR.t232 VSS 0.037471f
C9449 VDPWR.t543 VSS 0.02631f
C9450 VDPWR.t572 VSS 0.016942f
C9451 VDPWR.t139 VSS 0.018935f
C9452 VDPWR.t415 VSS 0.018935f
C9453 VDPWR.t559 VSS 0.016743f
C9454 VDPWR.t830 VSS 0.02053f
C9455 VDPWR.t338 VSS 0.022722f
C9456 VDPWR.t187 VSS 0.02631f
C9457 VDPWR.t348 VSS 0.033884f
C9458 VDPWR.t558 VSS 0.026908f
C9459 VDPWR.t785 VSS 0.016743f
C9460 VDPWR.t140 VSS 0.016743f
C9461 VDPWR.t189 VSS 0.022722f
C9462 VDPWR.t334 VSS 0.029897f
C9463 VDPWR.n2848 VSS 0.033342f
C9464 VDPWR.n2849 VSS 0.011469f
C9465 VDPWR.n2850 VSS 0.005706f
C9466 VDPWR.n2851 VSS 0.001952f
C9467 VDPWR.t190 VSS 0.001902f
C9468 VDPWR.t786 VSS 0.001902f
C9469 VDPWR.n2852 VSS 0.004259f
C9470 VDPWR.n2853 VSS 0.005483f
C9471 VDPWR.n2854 VSS 0.001197f
C9472 VDPWR.n2855 VSS 0.00622f
C9473 VDPWR.n2856 VSS 0.00622f
C9474 VDPWR.n2857 VSS 0.00622f
C9475 VDPWR.n2858 VSS 0.001353f
C9476 VDPWR.n2859 VSS 0.005119f
C9477 VDPWR.n2860 VSS 0.004403f
C9478 VDPWR.n2861 VSS 0.001688f
C9479 VDPWR.n2862 VSS 0.002203f
C9480 VDPWR.n2863 VSS 0.00622f
C9481 VDPWR.n2864 VSS 0.00622f
C9482 VDPWR.n2865 VSS 0.00622f
C9483 VDPWR.n2866 VSS 0.001616f
C9484 VDPWR.n2867 VSS 0.004427f
C9485 VDPWR.n2868 VSS 0.0059f
C9486 VDPWR.n2869 VSS 0.001425f
C9487 VDPWR.n2870 VSS 0.002164f
C9488 VDPWR.n2871 VSS 0.001668f
C9489 VDPWR.n2872 VSS 0.002085f
C9490 VDPWR.n2873 VSS 0.003043f
C9491 VDPWR.n2874 VSS 0.002164f
C9492 VDPWR.n2875 VSS 0.00311f
C9493 VDPWR.n2876 VSS 0.002085f
C9494 VDPWR.n2877 VSS 0.003257f
C9495 VDPWR.n2878 VSS 0.003595f
C9496 VDPWR.n2879 VSS 0.245208f
C9497 VDPWR.n2880 VSS 0.003595f
C9498 VDPWR.n2881 VSS 0.003257f
C9499 VDPWR.n2882 VSS 0.00156f
C9500 VDPWR.n2883 VSS 6.42e-19
C9501 VDPWR.n2884 VSS 0.001437f
C9502 VDPWR.n2885 VSS 0.021317f
C9503 VDPWR.n2886 VSS 0.007314f
C9504 VDPWR.n2887 VSS 0.006481f
C9505 VDPWR.n2888 VSS 0.003685f
C9506 VDPWR.n2889 VSS 0.00311f
C9507 VDPWR.n2890 VSS 0.004665f
C9508 VDPWR.n2891 VSS 0.00182f
C9509 VDPWR.n2892 VSS 0.006337f
C9510 VDPWR.n2893 VSS 0.007045f
C9511 VDPWR.t24 VSS 7.99e-19
C9512 VDPWR.t504 VSS 7.99e-19
C9513 VDPWR.n2894 VSS 0.001849f
C9514 VDPWR.n2895 VSS 0.025049f
C9515 VDPWR.n2896 VSS 0.005137f
C9516 VDPWR.n2897 VSS 0.002096f
C9517 VDPWR.n2898 VSS 0.002299f
C9518 VDPWR.n2899 VSS 0.006239f
C9519 VDPWR.t889 VSS 0.005265f
C9520 VDPWR.n2900 VSS 0.004835f
C9521 VDPWR.n2901 VSS 0.010139f
C9522 VDPWR.n2902 VSS 0.016678f
C9523 VDPWR.t156 VSS 0.003189f
C9524 VDPWR.n2903 VSS 0.005779f
C9525 VDPWR.t890 VSS 0.005265f
C9526 VDPWR.n2904 VSS 0.004569f
C9527 VDPWR.n2905 VSS 0.013041f
C9528 VDPWR.n2906 VSS 0.00311f
C9529 VDPWR.n2907 VSS 0.002164f
C9530 VDPWR.n2908 VSS 0.012868f
C9531 VDPWR.n2909 VSS 0.012246f
C9532 VDPWR.n2910 VSS 0.002164f
C9533 VDPWR.n2911 VSS 0.002366f
C9534 VDPWR.n2912 VSS 0.002085f
C9535 VDPWR.n2913 VSS 0.003257f
C9536 VDPWR.n2914 VSS 0.003595f
C9537 VDPWR.n2915 VSS 0.245208f
C9538 VDPWR.n2916 VSS 0.003595f
C9539 VDPWR.n2917 VSS 0.003257f
C9540 VDPWR.n2918 VSS 5.79e-19
C9541 VDPWR.n2919 VSS 0.00213f
C9542 VDPWR.n2920 VSS 0.005237f
C9543 VDPWR.t1136 VSS 0.005308f
C9544 VDPWR.t1180 VSS 0.011265f
C9545 VDPWR.n2922 VSS 0.028883f
C9546 VDPWR.t1137 VSS 0.005308f
C9547 VDPWR.n2923 VSS 0.015733f
C9548 VDPWR.n2924 VSS 0.014055f
C9549 VDPWR.n2925 VSS 0.003845f
C9550 VDPWR.n2926 VSS 0.001317f
C9551 VDPWR.n2927 VSS 0.001197f
C9552 VDPWR.n2928 VSS 0.00622f
C9553 VDPWR.n2929 VSS 0.004665f
C9554 VDPWR.n2930 VSS 0.001976f
C9555 VDPWR.t115 VSS 0.002994f
C9556 VDPWR.n2931 VSS 0.007536f
C9557 VDPWR.t196 VSS 0.001902f
C9558 VDPWR.t278 VSS 0.001902f
C9559 VDPWR.n2932 VSS 0.004259f
C9560 VDPWR.n2933 VSS 0.005483f
C9561 VDPWR.n2934 VSS 5.75e-19
C9562 VDPWR.n2935 VSS 0.00622f
C9563 VDPWR.n2936 VSS 0.00622f
C9564 VDPWR.n2937 VSS 0.004936f
C9565 VDPWR.n2938 VSS 0.007536f
C9566 VDPWR.n2939 VSS 9.94e-19
C9567 VDPWR.n2940 VSS 0.004654f
C9568 VDPWR.n2941 VSS 0.001688f
C9569 VDPWR.t276 VSS 0.001426f
C9570 VDPWR.t546 VSS 0.002942f
C9571 VDPWR.n2942 VSS 0.00599f
C9572 VDPWR.n2943 VSS 0.004654f
C9573 VDPWR.n2944 VSS 0.00622f
C9574 VDPWR.t682 VSS 0.002933f
C9575 VDPWR.t509 VSS 0.001217f
C9576 VDPWR.t89 VSS 0.001217f
C9577 VDPWR.n2945 VSS 0.002534f
C9578 VDPWR.n2946 VSS 0.007314f
C9579 VDPWR.t587 VSS 0.002933f
C9580 VDPWR.t959 VSS 0.005265f
C9581 VDPWR.n2947 VSS 0.009272f
C9582 VDPWR.n2948 VSS 0.003685f
C9583 VDPWR.t1250 VSS 0.030953f
C9584 VDPWR.t1164 VSS 0.001217f
C9585 VDPWR.t61 VSS 0.001217f
C9586 VDPWR.n2949 VSS 0.002507f
C9587 VDPWR.n2950 VSS 0.015796f
C9588 VDPWR.n2951 VSS 7.78e-19
C9589 VDPWR.n2952 VSS 0.002085f
C9590 VDPWR.n2953 VSS 0.001668f
C9591 VDPWR.n2954 VSS 0.001668f
C9592 VDPWR.n2955 VSS 0.002085f
C9593 VDPWR.n2956 VSS 0.002231f
C9594 VDPWR.t642 VSS 0.007445f
C9595 VDPWR.t960 VSS 0.005265f
C9596 VDPWR.n2957 VSS 0.019751f
C9597 VDPWR.n2958 VSS 0.005779f
C9598 VDPWR.t832 VSS 0.005308f
C9599 VDPWR.t1285 VSS 0.011265f
C9600 VDPWR.n2960 VSS 0.028883f
C9601 VDPWR.t833 VSS 0.005308f
C9602 VDPWR.n2961 VSS 0.015733f
C9603 VDPWR.n2962 VSS 0.001555f
C9604 VDPWR.n2963 VSS 0.002164f
C9605 VDPWR.n2964 VSS 0.002085f
C9606 VDPWR.n2965 VSS 0.00311f
C9607 VDPWR.n2966 VSS 0.002164f
C9608 VDPWR.t953 VSS 0.005308f
C9609 VDPWR.t1256 VSS 0.011265f
C9610 VDPWR.n2968 VSS 0.028883f
C9611 VDPWR.t954 VSS 0.005308f
C9612 VDPWR.n2969 VSS 0.015733f
C9613 VDPWR.n2970 VSS 0.013261f
C9614 VDPWR.n2971 VSS 0.001454f
C9615 VDPWR.n2972 VSS 0.003047f
C9616 VDPWR.n2973 VSS 0.003257f
C9617 VDPWR.n2974 VSS 0.003595f
C9618 VDPWR.n2975 VSS 0.003719f
C9619 VDPWR.n2976 VSS 0.003719f
C9620 VDPWR.n2977 VSS 0.003595f
C9621 VDPWR.n2978 VSS 0.003257f
C9622 VDPWR.n2979 VSS 0.003115f
C9623 VDPWR.n2980 VSS 0.005409f
C9624 VDPWR.n2981 VSS 0.002164f
C9625 VDPWR.n2982 VSS 0.016328f
C9626 VDPWR.n2983 VSS 0.016151f
C9627 VDPWR.n2984 VSS 0.01274f
C9628 VDPWR.n2985 VSS 0.034031f
C9629 VDPWR.n2986 VSS 0.00622f
C9630 VDPWR.n2987 VSS 0.004665f
C9631 VDPWR.n2988 VSS 0.005679f
C9632 VDPWR.n2989 VSS 0.005996f
C9633 VDPWR.n2990 VSS 0.003685f
C9634 VDPWR.n2991 VSS 0.00622f
C9635 VDPWR.n2992 VSS 0.00622f
C9636 VDPWR.n2993 VSS 0.001425f
C9637 VDPWR.n2994 VSS 0.006415f
C9638 VDPWR.n2995 VSS 0.001461f
C9639 VDPWR.n2996 VSS 0.00622f
C9640 VDPWR.n2997 VSS 0.005071f
C9641 VDPWR.n2998 VSS 0.001616f
C9642 VDPWR.n2999 VSS 0.002203f
C9643 VDPWR.n3000 VSS 0.002164f
C9644 VDPWR.n3001 VSS 0.00311f
C9645 VDPWR.n3002 VSS 0.002085f
C9646 VDPWR.n3003 VSS 0.003719f
C9647 VDPWR.n3004 VSS 0.001668f
C9648 VDPWR.n3005 VSS 0.002085f
C9649 VDPWR.n3006 VSS 0.002231f
C9650 VDPWR.n3007 VSS 0.003043f
C9651 VDPWR.n3008 VSS 0.002085f
C9652 VDPWR.n3009 VSS 0.003257f
C9653 VDPWR.n3010 VSS 0.003595f
C9654 VDPWR.n3011 VSS 0.245208f
C9655 VDPWR.n3012 VSS 0.13021f
C9656 VDPWR.n3013 VSS 0.12621f
C9657 VDPWR.n3014 VSS 0.083273f
C9658 VDPWR.n3015 VSS 0.003227f
C9659 VDPWR.n3016 VSS 0.003115f
C9660 VDPWR.n3017 VSS 0.004361f
C9661 VDPWR.n3018 VSS 0.00213f
C9662 VDPWR.n3019 VSS 0.00205f
C9663 VDPWR.n3020 VSS 0.006239f
C9664 VDPWR.n3021 VSS 0.003685f
C9665 VDPWR.n3022 VSS 0.004665f
C9666 VDPWR.n3023 VSS 0.012335f
C9667 VDPWR.n3024 VSS 0.016328f
C9668 VDPWR.n3025 VSS 0.011891f
C9669 VDPWR.n3026 VSS 0.00622f
C9670 VDPWR.n3027 VSS 0.00622f
C9671 VDPWR.n3028 VSS 0.005646f
C9672 VDPWR.n3029 VSS 0.012069f
C9673 VDPWR.n3030 VSS 0.049078f
C9674 VDPWR.n3031 VSS 0.009669f
C9675 VDPWR.n3032 VSS 0.011093f
C9676 VDPWR.n3033 VSS 0.00213f
C9677 VDPWR.n3034 VSS 0.0024f
C9678 VDPWR.n3035 VSS 0.005779f
C9679 VDPWR.n3036 VSS 0.013131f
C9680 VDPWR.n3037 VSS 0.001221f
C9681 VDPWR.n3038 VSS 0.002164f
C9682 VDPWR.n3039 VSS 0.00311f
C9683 VDPWR.n3040 VSS 0.002085f
C9684 VDPWR.n3041 VSS 0.001668f
C9685 VDPWR.n3042 VSS 0.082828f
C9686 VDPWR.n3043 VSS 0.287656f
C9687 VDPWR.n3044 VSS 0.147111f
C9688 VDPWR.n3045 VSS 0.147111f
C9689 VDPWR.n3046 VSS 0.221779f
C9690 VDPWR.n3047 VSS 0.309233f
C9691 VDPWR.n3048 VSS 0.190419f
C9692 VDPWR.n3049 VSS 0.070292f
C9693 VDPWR.n3050 VSS 0.188943f
C9694 VDPWR.n3051 VSS 0.026863f
C9695 VDPWR.n3052 VSS 0.071815f
C9696 VDPWR.n3053 VSS 1.66323f
C9697 VDPWR.n3054 VSS 5.0056f
C9698 VDPWR.n3055 VSS 1.54201f
C9699 VDPWR.n3056 VSS 0.41281f
C9700 VDPWR.n3057 VSS 0.037257f
C9701 VDPWR.n3058 VSS 0.120941f
C9702 VDPWR.n3059 VSS 0.058602f
C9703 VDPWR.n3060 VSS 0.058602f
C9704 VDPWR.n3061 VSS 0.058411f
C9705 VDPWR.n3062 VSS 0.080977f
C9706 VDPWR.n3063 VSS 0.261065f
C9707 VDPWR.t363 VSS 0.376779f
C9708 VDPWR.n3064 VSS 0.363781f
C9709 VDPWR.t463 VSS 0.376779f
C9710 VDPWR.n3065 VSS 0.261065f
C9711 VDPWR.n3066 VSS 2.51e-19
C9712 VDPWR.n3067 VSS 0.006628f
C9713 VDPWR.n3068 VSS 0.064054f
C9714 VDPWR.n3069 VSS 0.019206f
C9715 VDPWR.n3070 VSS 0.032407f
C9716 VDPWR.n3071 VSS 0.164857f
C9717 VDPWR.n3072 VSS 0.178603f
C9718 VDPWR.n3073 VSS 0.037221f
C9719 VDPWR.n3074 VSS 0.120941f
C9720 VDPWR.n3075 VSS 0.004701f
C9721 VDPWR.n3076 VSS 0.058602f
C9722 VDPWR.n3077 VSS 0.058602f
C9723 VDPWR.n3078 VSS 0.058411f
C9724 VDPWR.n3079 VSS 0.080977f
C9725 VDPWR.n3080 VSS 0.261065f
C9726 VDPWR.t556 VSS 0.376779f
C9727 VDPWR.n3081 VSS 0.363781f
C9728 VDPWR.t557 VSS 0.376779f
C9729 VDPWR.n3082 VSS 0.261065f
C9730 VDPWR.n3083 VSS 0.002139f
C9731 VDPWR.n3084 VSS 0.064116f
C9732 VDPWR.n3085 VSS 0.019206f
C9733 VDPWR.n3086 VSS 0.030813f
C9734 VDPWR.n3087 VSS 0.169973f
C9735 VDPWR.n3088 VSS 0.193894f
C9736 VDPWR.n3089 VSS 0.037101f
C9737 VDPWR.n3090 VSS 0.120941f
C9738 VDPWR.n3091 VSS 0.004709f
C9739 VDPWR.n3092 VSS 0.058602f
C9740 VDPWR.n3093 VSS 0.058602f
C9741 VDPWR.n3094 VSS 0.058411f
C9742 VDPWR.n3095 VSS 0.080977f
C9743 VDPWR.n3096 VSS 0.261065f
C9744 VDPWR.t470 VSS 0.376779f
C9745 VDPWR.n3097 VSS 0.363781f
C9746 VDPWR.t64 VSS 0.376779f
C9747 VDPWR.n3098 VSS 0.261065f
C9748 VDPWR.n3099 VSS 0.002259f
C9749 VDPWR.n3100 VSS 0.064116f
C9750 VDPWR.n3101 VSS 0.019206f
C9751 VDPWR.n3102 VSS 0.030813f
C9752 VDPWR.n3103 VSS 0.171881f
C9753 VDPWR.n3104 VSS 0.176051f
C9754 VDPWR.n3105 VSS 0.006609f
C9755 VDPWR.n3106 VSS 0.064079f
C9756 VDPWR.n3107 VSS 0.019206f
C9757 VDPWR.n3108 VSS 0.031091f
C9758 VDPWR.n3109 VSS 0.063632f
C9759 VDPWR.n3110 VSS 0.712985f
C9760 VDPWR.t702 VSS 0.002958f
C9761 VDPWR.t1212 VSS 0.001743f
C9762 VDPWR.t705 VSS 0.002958f
C9763 VDPWR.t1206 VSS 0.001743f
C9764 VDPWR.n3111 VSS 0.004963f
C9765 VDPWR.n3112 VSS 0.007338f
C9766 VDPWR.n3113 VSS 0.007288f
C9767 VDPWR.n3114 VSS 0.031849f
C9768 VDPWR.n3115 VSS 0.097815f
C9769 VDPWR.n3116 VSS 0.039528f
C9770 ringtest_0.x4.net2.t7 VSS 0.015381f
C9771 ringtest_0.x4.net2.t8 VSS 0.026101f
C9772 ringtest_0.x4.net2.n0 VSS 0.037026f
C9773 ringtest_0.x4.net2.t4 VSS 0.015381f
C9774 ringtest_0.x4.net2.t3 VSS 0.026101f
C9775 ringtest_0.x4.net2.n1 VSS 0.033335f
C9776 ringtest_0.x4.net2.n2 VSS 0.017289f
C9777 ringtest_0.x4.net2.n3 VSS 0.0837f
C9778 ringtest_0.x4.net2.t5 VSS 0.026101f
C9779 ringtest_0.x4.net2.t2 VSS 0.016278f
C9780 ringtest_0.x4.net2.n4 VSS 0.052479f
C9781 ringtest_0.x4.net2.n5 VSS 0.259642f
C9782 ringtest_0.x4.net2.t9 VSS 0.013842f
C9783 ringtest_0.x4.net2.t11 VSS 0.011454f
C9784 ringtest_0.x4.net2.n6 VSS 0.060494f
C9785 ringtest_0.x4.net2.n7 VSS 0.03533f
C9786 ringtest_0.x4.net2.n8 VSS 0.650991f
C9787 ringtest_0.x4.net2.t6 VSS 0.017756f
C9788 ringtest_0.x4.net2.t10 VSS 0.028277f
C9789 ringtest_0.x4.net2.n9 VSS 0.038818f
C9790 ringtest_0.x4.net2.n10 VSS 0.03575f
C9791 ringtest_0.x4.net2.n11 VSS 0.11929f
C9792 ringtest_0.x4.net2.n12 VSS 0.278364f
C9793 ringtest_0.x4.net2.n13 VSS 0.037886f
C9794 ringtest_0.x4.net2.t1 VSS 0.08709f
C9795 ringtest_0.x4.net2.n14 VSS 0.10636f
C9796 ringtest_0.x4.net2.t0 VSS 0.032833f
.ends

