magic
tech sky130A
magscale 1 2
timestamp 1728162076
<< metal1 >>
rect 4142 774 4194 776
rect 4138 770 4198 774
rect 4138 718 4142 770
rect 4194 718 4198 770
rect 3898 643 3950 648
rect 3895 642 3953 643
rect 3895 586 3898 642
rect 3950 586 3953 642
rect 3088 502 3140 506
rect 3084 500 3144 502
rect 3084 444 3088 500
rect 3140 444 3144 500
rect 2858 367 2910 372
rect 2856 366 2913 367
rect 2856 310 2858 366
rect 2910 310 2913 366
rect 2040 238 2092 242
rect 2038 236 2094 238
rect 2038 184 2040 236
rect 2092 184 2094 236
rect 1804 116 1856 120
rect 1801 114 1860 116
rect 1801 58 1804 114
rect 1856 58 1860 114
rect 998 14 1050 20
rect 1050 -42 1051 13
rect 754 -88 806 -84
rect 752 -90 808 -88
rect 752 -142 754 -90
rect 806 -142 808 -90
rect 752 -384 808 -142
rect 998 -344 1051 -42
rect 1801 -387 1860 58
rect 2038 -358 2094 184
rect 2856 -382 2913 310
rect 3084 -380 3144 444
rect 3895 -369 3953 586
rect 4138 -324 4198 718
<< via1 >>
rect 4142 718 4194 770
rect 3898 586 3950 642
rect 3088 444 3140 500
rect 2858 310 2910 366
rect 2040 184 2092 236
rect 1804 58 1856 114
rect 998 -42 1050 14
rect 754 -142 806 -90
<< metal2 >>
rect -3614 770 -3558 772
rect -3614 718 4142 770
rect 4194 718 4200 770
rect -3614 -372 -3558 718
rect -3062 586 3898 642
rect 3950 586 3956 642
rect -3062 584 -2826 586
rect -3062 -396 -3006 584
rect -2510 444 3088 500
rect 3140 444 3146 500
rect -2510 -424 -2454 444
rect -1958 310 2858 366
rect 2910 310 2916 366
rect -1958 -382 -1902 310
rect -1406 236 2096 238
rect -1406 184 2040 236
rect 2092 184 2098 236
rect -1406 182 2096 184
rect -1406 -396 -1350 182
rect -854 58 1804 114
rect 1856 58 1862 114
rect -854 -404 -798 58
rect -302 -42 998 14
rect 1050 -42 1056 14
rect -302 -366 -246 -42
rect 250 -90 806 -89
rect 250 -142 754 -90
rect 806 -142 812 -90
rect 250 -146 806 -142
rect 250 -356 306 -146
rect -3494 -4912 -3322 -4754
rect -2106 -4920 -1934 -4762
rect -554 -4894 -368 -4892
rect -554 -4902 848 -4894
rect -368 -5056 848 -4902
rect -554 -5066 848 -5056
rect -546 -5094 848 -5066
<< via2 >>
rect -554 -5056 -368 -4902
<< metal3 >>
rect -1145 -208 1434 -10
rect -1145 -930 -947 -208
rect 1236 -422 1434 -208
rect -2562 -968 -916 -930
rect -2562 -1070 -2540 -968
rect -2240 -1070 -1236 -968
rect -936 -1070 -916 -968
rect -2562 -1106 -916 -1070
rect -2562 -1268 -2248 -1106
rect -1246 -1274 -928 -1106
rect -1902 -4110 -1592 -3904
rect -588 -4110 -278 -3890
rect -3230 -4114 -244 -4110
rect -3230 -4244 -3218 -4114
rect -2928 -4124 -244 -4114
rect -2928 -4132 -584 -4124
rect -2928 -4244 -1888 -4132
rect -3230 -4256 -1888 -4244
rect -1902 -4262 -1888 -4256
rect -1598 -4254 -584 -4132
rect -294 -4254 -244 -4124
rect -1598 -4256 -244 -4254
rect -1598 -4262 -1588 -4256
rect -1902 -4266 -1592 -4262
rect -566 -4902 -328 -4256
rect -566 -5056 -554 -4902
rect -368 -5056 -328 -4902
rect -566 -5084 -328 -5056
<< via3 >>
rect -2540 -1070 -2240 -968
rect -1236 -1070 -936 -968
rect -3218 -4244 -2928 -4114
rect -1888 -4262 -1598 -4132
rect -584 -4254 -294 -4124
<< metal4 >>
rect -2556 -968 -2238 -950
rect -2556 -1070 -2540 -968
rect -2240 -1070 -2238 -968
rect -2556 -1264 -2238 -1070
rect -1246 -968 -928 -960
rect -1246 -1070 -1236 -968
rect -936 -1070 -928 -968
rect -1246 -1274 -928 -1070
rect -3226 -4114 -2918 -3850
rect -3226 -4244 -3218 -4114
rect -2928 -4244 -2918 -4114
rect -585 -4124 -293 -4123
rect -3226 -4252 -2918 -4244
rect -1889 -4132 -1597 -4131
rect -1889 -4262 -1888 -4132
rect -1598 -4262 -1597 -4132
rect -585 -4254 -584 -4124
rect -294 -4254 -293 -4124
rect -585 -4255 -293 -4254
rect -1889 -4263 -1597 -4262
use passgatesCtrl  passgatesCtrl_0
timestamp 1728160187
transform -1 0 878 0 -1 950
box 566 1232 4494 5870
use passgatex4  passgatex4_0
timestamp 1725644236
transform 1 0 -10990 0 1 -4896
box 11366 -356 15589 4682
<< labels >>
flabel metal2 -2106 -4920 -1934 -4762 0 FreeSans 1600 0 0 0 select0
port 1 nsew
flabel metal2 -3494 -4912 -3322 -4754 0 FreeSans 1600 0 0 0 select1
port 2 nsew
flabel metal1 452 -422 652 -222 0 FreeSans 1600 0 0 0 A1
port 3 nsew
flabel metal1 1508 -424 1708 -224 0 FreeSans 1600 0 0 0 A2
port 4 nsew
flabel metal1 2552 -428 2752 -228 0 FreeSans 1600 0 0 0 A3
port 5 nsew
flabel metal1 3582 -414 3782 -214 0 FreeSans 1600 0 0 0 A4
port 6 nsew
flabel metal1 424 -5158 624 -4794 0 FreeSans 1600 0 0 0 Z1
port 7 nsew
flabel metal1 1492 -5154 1692 -4954 0 FreeSans 1600 0 0 0 Z2
port 8 nsew
flabel metal1 2562 -5190 2762 -4990 0 FreeSans 1600 0 0 0 Z3
port 9 nsew
flabel metal1 3620 -5192 3820 -4790 0 FreeSans 1600 0 0 0 Z4
port 10 nsew
flabel metal1 -568 -5090 -330 -4814 0 FreeSans 1600 0 0 0 VDD
port 11 nsew
flabel metal1 -1148 -214 -956 -22 0 FreeSans 1600 0 0 0 VSS
port 12 nsew
<< end >>
