* NGSPICE file created from mux4onehot_b_parax.ext - technology: sky130A

.subckt mux4onehot_b_parax select1 select2 A1 A3 Z1 A2 A4 select0 Z4 Z3 VDD Z2 VSS
+ nselect2
X0 A2.t1 x2.GP2.t4 Z2.t0 VDD.t19 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1 VDD.t5 a_5275_n4059# a_5275_n4235# VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 A1.t2 x2.GP1.t4 Z1.t2 VDD.t53 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X3 VSS.t56 select0.t0 a_5275_n3507# VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 a_5275_n3683# a_5275_n3507# a_5301_n3555# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X5 A4.t3 x2.GP4.t4 Z4.t2 VDD.t3 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X6 VSS.t17 select1.t0 x1.nSEL1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VSS.t32 x2.GN2 x2.GP2.t3 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 x1.nSEL0 select0.t1 VSS.t54 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VSS.t27 a_5275_n4651# x2.GN1.t1 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VDD.t52 select0.t2 x1.nSEL0 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 x2.GP1.t0 x2.GN1.t2 VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VSS.t43 x2.GN1.t3 x2.GP1.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 x2.GP4.t0 x2.GN4.t2 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 VDD.t63 x2.GN4.t3 x2.GP4.t3 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 a_5275_n4059# select1.t1 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X16 VSS.t11 VDD.t71 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X17 a_5301_n4107# select0.t3 VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X18 VSS.t61 a_5275_n4235# x2.GN2 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_5275_n4651# x1.nSEL1 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X20 VSS.t8 VDD.t72 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X21 a_5275_n3507# select0.t4 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X22 a_5275_n4235# select0.t5 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X23 VDD.t42 x1.nSEL0 a_5275_n4651# VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VDD.t50 a_5275_n3507# a_5275_n3683# VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X25 VDD.t48 a_5275_n3683# x2.GN3 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X26 VSS.t39 a_5275_n2995# x2.GN4.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X27 nselect2.t1 select2.t0 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 A3.t3 x2.GP3 Z3.t2 VDD.t70 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X29 VSS.t50 select0.t6 x1.nSEL0 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 Z3.t0 x2.GN3 A3.t1 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X31 Z3.t1 x2.GN3 A3.t0 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X32 VDD.t65 select2.t1 nselect2.t0 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 x2.GP4.t1 x2.GN4.t4 VSS.t45 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X34 x2.GP3 x2.GN3 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 x1.nSEL1 select1.t2 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 x2.GP2.t0 x2.GN2 VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X37 VDD.t12 VSS.t68 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X38 VSS.t65 x2.GN4.t5 x2.GP4.t2 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 VSS.t5 VDD.t73 VSS.t4 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X40 a_5329_n4513# x1.nSEL1 VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X41 VDD.t2 VSS.t69 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X42 a_5275_n4651# x1.nSEL0 a_5329_n4513# VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 A4.t2 x2.GP4.t5 Z4.t3 VDD.t3 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X44 a_5275_n2995# select0.t7 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X45 VDD.t28 x2.GN3 x2.GP3 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X46 VDD.t32 a_5275_n4651# x2.GN1.t0 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X47 Z4.t1 x2.GN4.t6 A4.t1 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X48 VSS.t2 VDD.t74 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X49 Z4.t0 x2.GN4.t7 A4.t0 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X50 VDD.t7 select1.t3 a_5275_n2995# VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X51 a_5275_n3683# select1.t4 VDD.t56 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X52 nselect2.t3 select2.t2 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 a_5275_n4235# a_5275_n4059# a_5301_n4107# VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X54 VSS.t35 select2.t3 nselect2.t2 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 x2.GP3 x2.GN3 VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X56 VDD.t59 VSS.t70 VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X57 A2.t0 x2.GP2.t5 Z2.t1 VDD.t19 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X58 VDD.t61 select1.t5 x1.nSEL1 VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X59 x1.nSEL1 select1.t6 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 x2.GP2.t2 x2.GN2 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X61 VDD.t55 a_5275_n4235# x2.GN2 VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X62 Z2.t2 x2.GN2 A2.t3 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X63 a_5329_n2857# select0.t8 VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X64 A1.t1 x2.GP1.t5 Z1.t1 VDD.t53 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X65 Z2.t3 x2.GN2 A2.t2 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X66 VDD.t38 a_5275_n2995# x2.GN4.t0 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X67 VDD.t24 VSS.t71 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X68 VSS.t22 x2.GN3 x2.GP3 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X69 VDD.t34 x2.GN2 x2.GP2.t1 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X70 x1.nSEL0 select0.t9 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X71 Z1.t3 x2.GN1.t4 A1.t3 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X72 x2.GP1.t2 x2.GN1.t5 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 Z1.t0 x2.GN1.t6 A1.t0 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X74 a_5275_n2995# select1.t7 a_5329_n2857# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 a_5301_n3555# select1.t8 VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X76 VSS.t58 a_5275_n3683# x2.GN3 VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X77 VSS.t63 select1.t9 a_5275_n4059# VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X78 VDD.t69 x2.GN1.t7 x2.GP1.t3 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X79 A3.t2 x2.GP3 Z3.t3 VDD.t70 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
R0 x2.GP2.n4 x2.GP2.t4 450.938
R1 x2.GP2.n4 x2.GP2.t5 445.666
R2 x2.GP2.n5 x2.GP2.n3 195.958
R3 x2.GP2.n1 x2.GP2.n0 101.49
R4 x2.GP2.n3 x2.GP2.t1 26.5955
R5 x2.GP2.n3 x2.GP2.t0 26.5955
R6 x2.GP2.n0 x2.GP2.t3 24.9236
R7 x2.GP2.n0 x2.GP2.t2 24.9236
R8 x1.gpo1 x2.x2.GP 13.129
R9 x2.GP2.n5 x1.gpo1 11.995
R10 x2.GP2.n2 x1.x12.Y 10.7525
R11 x1.x12.Y x2.GP2.n5 7.96524
R12 x2.GP2.n2 x1.x12.Y 6.6565
R13 x1.x12.Y x2.GP2.n2 5.04292
R14 x2.x2.GP x2.GP2.n4 2.94361
R15 x1.x12.Y x2.GP2.n1 2.5605
R16 x2.GP2.n1 x1.x12.Y 1.93989
R17 Z2.n1 Z2.t1 23.6581
R18 Z2.n3 Z2.t0 23.3739
R19 Z2.n1 Z2.t2 10.7528
R20 Z2.n0 Z2.t3 10.6417
R21 Z2.n2 Z2.n1 1.30064
R22 Z2.n5 Z2.n4 0.936641
R23 Z2.n3 Z2.n2 0.726502
R24 Z2.n2 Z2.n0 0.512491
R25 Z2.n4 Z2.n0 0.359663
R26 Z2.n4 Z2.n3 0.216071
R27 Z2.n5 Z2 0.0776605
R28 Z2 Z2.n5 0.0561931
R29 A2.n1 A2.t1 26.3998
R30 A2.n1 A2.t0 23.5483
R31 A2.n0 A2.t2 12.7127
R32 A2.n0 A2.t3 10.8578
R33 A2.n2 A2.n1 3.12177
R34 A2.n2 A2.n0 1.81453
R35 A2.n3 A2.n2 1.1255
R36 A2.n3 A2 0.219402
R37 A2 A2.n3 0.0655
R38 VDD.n57 VDD.n55 8629.41
R39 VDD.n60 VDD.n54 8629.41
R40 VDD.n40 VDD.n39 8629.41
R41 VDD.n42 VDD.n37 8629.41
R42 VDD.n23 VDD.n22 8629.41
R43 VDD.n25 VDD.n20 8629.41
R44 VDD.n6 VDD.n4 8629.41
R45 VDD.n9 VDD.n3 8629.41
R46 VDD.n56 VDD.n53 920.471
R47 VDD.n43 VDD.n36 920.471
R48 VDD.n26 VDD.n19 920.471
R49 VDD.n5 VDD.n2 920.471
R50 VDD.n62 VDD.n53 914.447
R51 VDD.n45 VDD.n43 914.447
R52 VDD.n28 VDD.n26 914.447
R53 VDD.n11 VDD.n2 914.447
R54 VDD.t58 VDD.n127 804.731
R55 VDD.n129 VDD.t58 751.692
R56 VDD.n101 VDD.t7 671.408
R57 VDD.n90 VDD.t42 671.408
R58 VDD VDD.t57 630.375
R59 VDD.n160 VDD.n159 602.456
R60 VDD.n182 VDD.n70 602.456
R61 VDD.n74 VDD.n73 585
R62 VDD.n76 VDD.n75 585
R63 VDD.n56 VDD.n51 480.764
R64 VDD.n36 VDD.n34 480.764
R65 VDD.n19 VDD.n17 480.764
R66 VDD.n5 VDD.n1 480.764
R67 VDD VDD.t22 458.724
R68 VDD.t57 VDD 458.724
R69 VDD.n122 VDD.t64 420.25
R70 VDD.n118 VDD.t23 388.656
R71 VDD.n153 VDD.t24 388.656
R72 VDD.n131 VDD.t59 388.656
R73 VDD.n104 VDD.t1 388.656
R74 VDD.n113 VDD.t2 388.656
R75 VDD.n78 VDD.t11 388.656
R76 VDD.n83 VDD.t12 388.656
R77 VDD.n64 VDD.n51 379.2
R78 VDD.n47 VDD.n34 379.2
R79 VDD.n30 VDD.n17 379.2
R80 VDD.n13 VDD.n1 379.2
R81 VDD VDD.t60 369.938
R82 VDD VDD.t51 369.938
R83 VDD.n107 VDD.n100 322.329
R84 VDD.n85 VDD.n81 322.329
R85 VDD.n164 VDD.n162 259.697
R86 VDD.n140 VDD.t52 255.905
R87 VDD.n145 VDD.t61 255.905
R88 VDD.n121 VDD.t65 255.905
R89 VDD.n161 VDD.t28 255.905
R90 VDD.n111 VDD.t63 254.475
R91 VDD.n136 VDD.t26 252.95
R92 VDD.n141 VDD.t67 252.95
R93 VDD.n146 VDD.t40 252.95
R94 VDD.n181 VDD.t36 252.95
R95 VDD.n160 VDD.t9 251.516
R96 VDD.n71 VDD.t69 250.724
R97 VDD.n69 VDD.t34 250.724
R98 VDD.t64 VDD.t39 248.599
R99 VDD.t60 VDD.t66 248.599
R100 VDD.t51 VDD.t25 248.599
R101 VDD.n176 VDD.t46 248.219
R102 VDD.n163 VDD.t30 248.219
R103 VDD.n122 VDD 221.964
R104 VDD.n129 VDD.t73 215.827
R105 VDD.n111 VDD.n110 213.119
R106 VDD.n151 VDD.n122 213.119
R107 VDD.n119 VDD.t74 210.964
R108 VDD.n105 VDD.t72 210.964
R109 VDD.n80 VDD.t71 210.964
R110 VDD.n171 VDD.n170 209.368
R111 VDD.t39 VDD 198.287
R112 VDD.t66 VDD 198.287
R113 VDD.t25 VDD 198.287
R114 VDD.n173 VDD.n172 183.673
R115 VDD VDD.t37 182.952
R116 VDD VDD.n171 182.952
R117 VDD.t31 VDD 182.952
R118 VDD.n75 VDD.n74 159.476
R119 VDD.n162 VDD.t56 157.014
R120 VDD.t68 VDD.t43 154.417
R121 VDD.t49 VDD.t27 147.703
R122 VDD.t20 VDD.t6 140.989
R123 VDD.t27 VDD.t29 140.989
R124 VDD.t35 VDD.t33 140.989
R125 VDD.t45 VDD.t68 140.989
R126 VDD.t41 VDD.t13 140.989
R127 VDD.n162 VDD.t48 137.079
R128 VDD.n110 VDD 125.883
R129 VDD.n172 VDD 125.883
R130 VDD.n100 VDD.t21 116.341
R131 VDD.n81 VDD.t14 116.341
R132 VDD.t6 VDD 112.457
R133 VDD.t29 VDD 112.457
R134 VDD VDD.t41 112.457
R135 VDD VDD.t54 109.1
R136 VDD.t0 VDD.t20 104.064
R137 VDD.t13 VDD.t10 104.064
R138 VDD.t15 VDD 102.385
R139 VDD.t62 VDD 99.0288
R140 VDD.n159 VDD.t50 96.1553
R141 VDD.n70 VDD.t5 96.1553
R142 VDD VDD.t4 92.315
R143 VDD.n74 VDD.t44 86.7743
R144 VDD.n110 VDD.t62 83.9228
R145 VDD.n171 VDD.t47 80.5659
R146 VDD.t37 VDD.t0 77.209
R147 VDD.t10 VDD.t31 77.209
R148 VDD.n75 VDD.t55 66.8398
R149 VDD.n63 VDD.n62 66.6358
R150 VDD.n46 VDD.n45 66.6358
R151 VDD.n29 VDD.n28 66.6358
R152 VDD.n12 VDD.n11 66.6358
R153 VDD.n159 VDD.t16 63.3219
R154 VDD.n70 VDD.t18 63.3219
R155 VDD VDD.t49 62.103
R156 VDD.n57 VDD.n56 61.6672
R157 VDD.n61 VDD.n60 61.6672
R158 VDD.n40 VDD.n36 61.6672
R159 VDD.n37 VDD.n35 61.6672
R160 VDD.n23 VDD.n19 61.6672
R161 VDD.n20 VDD.n18 61.6672
R162 VDD.n6 VDD.n5 61.6672
R163 VDD.n10 VDD.n9 61.6672
R164 VDD.n58 VDD.n57 60.9564
R165 VDD.n60 VDD.n59 60.9564
R166 VDD.n41 VDD.n40 60.9564
R167 VDD.n38 VDD.n37 60.9564
R168 VDD.n24 VDD.n23 60.9564
R169 VDD.n21 VDD.n20 60.9564
R170 VDD.n7 VDD.n6 60.9564
R171 VDD.n9 VDD.n8 60.9564
R172 VDD.n46 VDD.n35 60.6123
R173 VDD.n29 VDD.n18 60.6123
R174 VDD.n63 VDD.n52 59.4829
R175 VDD.n12 VDD.n0 58.7299
R176 VDD.t43 VDD 55.3892
R177 VDD.t17 VDD 52.0323
R178 VDD VDD.t47 45.3185
R179 VDD VDD.t8 41.9616
R180 VDD.n58 VDD.n54 38.5759
R181 VDD.n59 VDD.n55 38.5759
R182 VDD.n42 VDD.n41 38.5759
R183 VDD.n39 VDD.n38 38.5759
R184 VDD.n25 VDD.n24 38.5759
R185 VDD.n22 VDD.n21 38.5759
R186 VDD.n7 VDD.n3 38.5759
R187 VDD.n8 VDD.n4 38.5759
R188 VDD.n170 VDD.n92 34.6358
R189 VDD.n170 VDD.n93 34.6358
R190 VDD.n175 VDD.n174 34.6358
R191 VDD.n172 VDD 28.5341
R192 VDD.n100 VDD.t38 28.4453
R193 VDD.n81 VDD.t32 28.4453
R194 VDD.n177 VDD.n176 28.3534
R195 VDD.n174 VDD.n173 25.6953
R196 VDD.n140 VDD.n125 25.224
R197 VDD.n136 VDD.n125 25.224
R198 VDD.n145 VDD.n124 25.224
R199 VDD.n141 VDD.n124 25.224
R200 VDD.n147 VDD.n121 25.224
R201 VDD.n147 VDD.n146 25.224
R202 VDD.n165 VDD.n161 25.224
R203 VDD.n111 VDD.n95 23.7181
R204 VDD VDD.n101 23.252
R205 VDD.n160 VDD.n95 21.4593
R206 VDD.n141 VDD.n140 20.3299
R207 VDD.n146 VDD.n145 20.3299
R208 VDD.t4 VDD.t35 20.1418
R209 VDD.n182 VDD.n69 19.9534
R210 VDD.n181 VDD.n180 19.8181
R211 VDD.n151 VDD.n121 17.3181
R212 VDD.n164 VDD.n163 17.3181
R213 VDD.n161 VDD.n160 16.5652
R214 VDD.n165 VDD.n164 16.5652
R215 VDD.n136 VDD.n135 15.8123
R216 VDD.n152 VDD.n151 14.2735
R217 VDD.n112 VDD.n111 14.2735
R218 VDD.n174 VDD.n90 13.9299
R219 VDD.n67 VDD.n66 13.6791
R220 VDD.n182 VDD.n181 13.5534
R221 VDD.n117 VDD.n116 11.4366
R222 VDD.n65 VDD.n64 11.3235
R223 VDD.n48 VDD.n47 11.3235
R224 VDD.n31 VDD.n30 11.3235
R225 VDD.n14 VDD.n13 11.3235
R226 VDD.n173 VDD.n91 11.2937
R227 VDD.n157 VDD.n156 11.2737
R228 VDD.t8 VDD.t15 10.0712
R229 VDD.n131 VDD.n128 9.60526
R230 VDD.n118 VDD.n117 9.60526
R231 VDD.n83 VDD.n82 9.60526
R232 VDD.n120 VDD.n96 9.3005
R233 VDD.n155 VDD.n154 9.3005
R234 VDD.n152 VDD.n97 9.3005
R235 VDD.n151 VDD.n150 9.3005
R236 VDD.n146 VDD.n123 9.3005
R237 VDD.n142 VDD.n141 9.3005
R238 VDD.n137 VDD.n136 9.3005
R239 VDD.n133 VDD.n132 9.3005
R240 VDD.n138 VDD.n125 9.3005
R241 VDD.n140 VDD.n139 9.3005
R242 VDD.n143 VDD.n124 9.3005
R243 VDD.n145 VDD.n144 9.3005
R244 VDD.n148 VDD.n147 9.3005
R245 VDD.n149 VDD.n121 9.3005
R246 VDD.n178 VDD.n177 9.3005
R247 VDD.n183 VDD.n182 9.3005
R248 VDD.n167 VDD.n92 9.3005
R249 VDD.n160 VDD.n158 9.3005
R250 VDD.n111 VDD.n109 9.3005
R251 VDD.n103 VDD.n102 9.3005
R252 VDD.n106 VDD.n98 9.3005
R253 VDD.n115 VDD.n114 9.3005
R254 VDD.n112 VDD.n99 9.3005
R255 VDD.n108 VDD.n95 9.3005
R256 VDD.n161 VDD.n94 9.3005
R257 VDD.n166 VDD.n165 9.3005
R258 VDD.n170 VDD.n169 9.3005
R259 VDD.n168 VDD.n93 9.3005
R260 VDD.n181 VDD.n68 9.3005
R261 VDD.n180 VDD.n179 9.3005
R262 VDD.n175 VDD.n72 9.3005
R263 VDD.n174 VDD.n77 9.3005
R264 VDD.n89 VDD.n88 9.3005
R265 VDD.n87 VDD.n86 9.3005
R266 VDD.n84 VDD.n79 9.3005
R267 VDD.n15 VDD.n0 8.23557
R268 VDD.n76 VDD.n73 6.8005
R269 VDD.n135 VDD.n127 6.48583
R270 VDD.n62 VDD.n61 6.02403
R271 VDD.n11 VDD.n10 6.02403
R272 VDD.n130 VDD.n129 5.8885
R273 VDD.n44 VDD.n35 4.89462
R274 VDD.n28 VDD.n27 4.89462
R275 VDD.n154 VDD.n120 4.67352
R276 VDD.n135 VDD.n134 4.62124
R277 VDD.n132 VDD.n131 4.36875
R278 VDD.n154 VDD.n153 4.36875
R279 VDD.n114 VDD.n113 4.36875
R280 VDD.n84 VDD.n83 4.36875
R281 VDD.t33 VDD.t17 3.35739
R282 VDD.t54 VDD.t45 3.35739
R283 VDD.n44 VDD.n33 3.23917
R284 VDD.n27 VDD.n16 3.23136
R285 VDD.n52 VDD.n50 3.22655
R286 VDD.n132 VDD.n130 3.2005
R287 VDD.n54 VDD.n53 2.84665
R288 VDD.n55 VDD.n51 2.84665
R289 VDD.n43 VDD.n42 2.84665
R290 VDD.n39 VDD.n34 2.84665
R291 VDD.n26 VDD.n25 2.84665
R292 VDD.n22 VDD.n17 2.84665
R293 VDD.n3 VDD.n2 2.84665
R294 VDD.n4 VDD.n1 2.84665
R295 VDD.n130 VDD.n127 2.8165
R296 VDD.n107 VDD.n106 2.54018
R297 VDD.n86 VDD.n85 2.54018
R298 VDD.n120 VDD.n119 2.33701
R299 VDD.n106 VDD.n105 2.33701
R300 VDD.n86 VDD.n80 2.33701
R301 VDD.n64 VDD.n63 2.28169
R302 VDD.n47 VDD.n46 2.28169
R303 VDD.n30 VDD.n29 2.28169
R304 VDD.n13 VDD.n12 2.28169
R305 VDD.n114 VDD.n107 2.13383
R306 VDD.n85 VDD.n84 2.13383
R307 VDD.n119 VDD.n118 2.03225
R308 VDD.n105 VDD.n104 2.03225
R309 VDD.n80 VDD.n78 2.03225
R310 VDD.n10 VDD.n0 1.88285
R311 VDD.n185 VDD.n184 1.753
R312 VDD.n93 VDD.n69 1.50638
R313 VDD.n177 VDD.n76 1.4005
R314 VDD.n103 VDD.n101 1.37193
R315 VDD.n90 VDD.n89 1.37193
R316 VDD.n49 VDD.n48 1.143
R317 VDD.n32 VDD.n31 1.143
R318 VDD.n66 VDD.n65 1.13925
R319 VDD.n15 VDD.n14 1.13675
R320 VDD.n61 VDD.n52 1.12991
R321 VDD.n45 VDD.n44 1.12991
R322 VDD.n27 VDD.n18 1.12991
R323 VDD.n126 VDD 1.06099
R324 VDD.n33 VDD.n32 0.862816
R325 VDD.n16 VDD.n15 0.770881
R326 VDD.n163 VDD.n92 0.753441
R327 VDD.n176 VDD.n175 0.753441
R328 VDD.n50 VDD.n49 0.729231
R329 VDD.n73 VDD.n71 0.6005
R330 VDD.n185 VDD.n67 0.511794
R331 VDD VDD.n185 0.460219
R332 VDD.n66 VDD.n50 0.405788
R333 VDD.n180 VDD.n71 0.4005
R334 VDD.n32 VDD.n16 0.392323
R335 VDD.n49 VDD.n33 0.360318
R336 VDD.n153 VDD.n152 0.305262
R337 VDD.n104 VDD.n103 0.305262
R338 VDD.n113 VDD.n112 0.305262
R339 VDD.n89 VDD.n78 0.305262
R340 VDD.t53 VDD.n58 0.27666
R341 VDD.n59 VDD.t53 0.27666
R342 VDD.n41 VDD.t19 0.27666
R343 VDD.n38 VDD.t19 0.27666
R344 VDD.n24 VDD.t70 0.27666
R345 VDD.n21 VDD.t70 0.27666
R346 VDD.t3 VDD.n7 0.27666
R347 VDD.n8 VDD.t3 0.27666
R348 VDD.n134 VDD.n133 0.180304
R349 VDD.n134 VDD 0.120408
R350 VDD.n117 VDD.n96 0.120292
R351 VDD.n155 VDD.n97 0.120292
R352 VDD.n149 VDD.n148 0.120292
R353 VDD.n148 VDD.n123 0.120292
R354 VDD.n144 VDD.n143 0.120292
R355 VDD.n143 VDD.n142 0.120292
R356 VDD.n139 VDD.n138 0.120292
R357 VDD.n138 VDD.n137 0.120292
R358 VDD.n133 VDD.n128 0.120292
R359 VDD.n102 VDD.n98 0.120292
R360 VDD.n115 VDD.n99 0.120292
R361 VDD.n166 VDD.n94 0.120292
R362 VDD.n167 VDD.n166 0.120292
R363 VDD.n183 VDD.n68 0.120292
R364 VDD.n179 VDD.n178 0.120292
R365 VDD.n178 VDD.n72 0.120292
R366 VDD.n88 VDD.n87 0.120292
R367 VDD.n87 VDD.n79 0.120292
R368 VDD.n82 VDD.n79 0.120292
R369 VDD.n156 VDD.n96 0.11899
R370 VDD.n102 VDD 0.0981562
R371 VDD.n157 VDD 0.0955521
R372 VDD.n116 VDD.n98 0.0916458
R373 VDD.n65 VDD 0.06425
R374 VDD.n48 VDD 0.06425
R375 VDD.n31 VDD 0.06425
R376 VDD.n14 VDD 0.06425
R377 VDD.n150 VDD 0.0603958
R378 VDD VDD.n149 0.0603958
R379 VDD.n144 VDD 0.0603958
R380 VDD.n139 VDD 0.0603958
R381 VDD.n109 VDD 0.0603958
R382 VDD VDD.n108 0.0603958
R383 VDD VDD.n94 0.0603958
R384 VDD.n169 VDD 0.0603958
R385 VDD VDD.n168 0.0603958
R386 VDD.n179 VDD 0.0603958
R387 VDD.n88 VDD 0.0603958
R388 VDD.n91 VDD 0.0590938
R389 VDD.n184 VDD 0.0525833
R390 VDD.n184 VDD.n183 0.0460729
R391 VDD.n109 VDD 0.0382604
R392 VDD VDD.n126 0.0369583
R393 VDD.n150 VDD 0.03175
R394 VDD.n169 VDD 0.03175
R395 VDD.n116 VDD.n115 0.0291458
R396 VDD.n67 VDD 0.0236148
R397 VDD VDD.n97 0.0226354
R398 VDD VDD.n123 0.0226354
R399 VDD.n142 VDD 0.0226354
R400 VDD.n137 VDD 0.0226354
R401 VDD.n128 VDD 0.0226354
R402 VDD VDD.n99 0.0226354
R403 VDD.n108 VDD 0.0226354
R404 VDD.n158 VDD 0.0226354
R405 VDD VDD.n167 0.0226354
R406 VDD.n168 VDD 0.0226354
R407 VDD VDD.n68 0.0226354
R408 VDD VDD.n72 0.0226354
R409 VDD VDD.n77 0.0226354
R410 VDD.n82 VDD 0.0226354
R411 VDD.n158 VDD.n157 0.00310417
R412 VDD.n156 VDD.n155 0.00180208
R413 VDD.n126 VDD 0.00180208
R414 VDD.n91 VDD.n77 0.00180208
R415 x2.GP1.n4 x2.GP1.t4 450.938
R416 x2.GP1.n4 x2.GP1.t5 445.666
R417 x2.GP1.n5 x2.GP1.n3 195.832
R418 x2.GP1.n1 x2.GP1.n0 101.49
R419 x2.GP1.n3 x2.GP1.t3 26.5955
R420 x2.GP1.n3 x2.GP1.t2 26.5955
R421 x2.GP1.n0 x2.GP1.t1 24.9236
R422 x2.GP1.n0 x2.GP1.t0 24.9236
R423 x2.GP1.n5 x1.gpo0 11.8923
R424 x1.gpo0 x2.x1.GP 11.5413
R425 x2.GP1.n2 x1.x11.Y 10.7525
R426 x1.x11.Y x2.GP1.n5 8.09215
R427 x2.GP1.n2 x1.x11.Y 6.6565
R428 x1.x11.Y x2.GP1.n2 5.04292
R429 x2.x1.GP x2.GP1.n4 2.90754
R430 x1.x11.Y x2.GP1.n1 2.5605
R431 x2.GP1.n1 x1.x11.Y 1.93989
R432 Z1.n1 Z1.t1 23.6581
R433 Z1.n3 Z1.t2 23.3739
R434 Z1.n1 Z1.t3 10.7528
R435 Z1.n0 Z1.t0 10.6417
R436 Z1.n2 Z1.n1 1.30064
R437 Z1 Z1.n4 0.983856
R438 Z1.n3 Z1.n2 0.726502
R439 Z1.n2 Z1.n0 0.512491
R440 Z1.n4 Z1.n0 0.359663
R441 Z1.n4 Z1.n3 0.216071
R442 A1.n1 A1.t2 26.3998
R443 A1.n1 A1.t1 23.5483
R444 A1.n0 A1.t0 12.7127
R445 A1.n0 A1.t3 10.8578
R446 A1.n2 A1.n1 3.12177
R447 A1.n2 A1.n0 1.81453
R448 A1.n3 A1.n2 1.1255
R449 A1.n3 A1 0.21174
R450 A1 A1.n3 0.0655
R451 select0.n5 select0.t4 327.99
R452 select0.n9 select0.t3 293.969
R453 select0.n3 select0.t7 261.887
R454 select0.n1 select0.t9 212.081
R455 select0.n0 select0.t2 212.081
R456 select0.n5 select0.t0 199.457
R457 select0.n2 select0.n1 183.185
R458 select0.n3 select0.t8 155.847
R459 select0 select0.n9 154.065
R460 select0.n6 select0.n5 152
R461 select0.n4 select0.n3 152
R462 select0.n1 select0.t1 139.78
R463 select0.n0 select0.t6 139.78
R464 select0.n9 select0.t5 138.338
R465 select0.n1 select0.n0 61.346
R466 select0.n10 select0 13.4199
R467 select0.n8 select0.n4 11.9062
R468 select0.n11 select0.n8 11.7395
R469 select0.n12 select0.n11 11.5949
R470 select0.n12 select0.n2 9.68118
R471 select0.n7 select0 9.17383
R472 select0.n2 select0 5.8885
R473 select0.n10 select0 5.57469
R474 select0.n8 select0.n7 4.6505
R475 select0.n11 select0.n10 4.6505
R476 select0.n7 select0.n6 2.98717
R477 select0.n6 select0 2.34717
R478 select0.n4 select0 2.07109
R479 select0 select0.n12 0.559212
R480 VSS.n182 VSS.n181 545142
R481 VSS.n42 VSS.n41 20148.7
R482 VSS.n55 VSS.n10 19433.3
R483 VSS.n49 VSS.n48 19054.3
R484 VSS VSS.n180 11981.2
R485 VSS.n50 VSS.n11 11744.7
R486 VSS.n54 VSS.n11 11744.7
R487 VSS.n50 VSS.n12 11744.7
R488 VSS.n54 VSS.n12 11744.7
R489 VSS.n36 VSS.n22 11744.7
R490 VSS.n40 VSS.n22 11744.7
R491 VSS.n36 VSS.n23 11744.7
R492 VSS.n40 VSS.n23 11744.7
R493 VSS.n43 VSS.n16 11744.7
R494 VSS.n47 VSS.n16 11744.7
R495 VSS.n43 VSS.n17 11744.7
R496 VSS.n47 VSS.n17 11744.7
R497 VSS.n184 VSS.n4 11744.7
R498 VSS.n184 VSS.n5 11744.7
R499 VSS.n9 VSS.n5 11744.7
R500 VSS.n9 VSS.n4 11744.7
R501 VSS.n56 VSS.n7 5416.06
R502 VSS.n21 VSS.n7 5357.62
R503 VSS.n180 VSS.n56 3878.48
R504 VSS.n183 VSS.n182 2174.55
R505 VSS VSS.t55 1289.66
R506 VSS.n179 VSS.n178 1198.25
R507 VSS.n137 VSS.n135 1198.25
R508 VSS.n146 VSS.n6 1194.5
R509 VSS.n165 VSS.n164 1171.32
R510 VSS VSS.n6 918.774
R511 VSS.t26 VSS 918.774
R512 VSS.t40 VSS.t57 826.054
R513 VSS.t51 VSS.t60 826.054
R514 VSS.t62 VSS.t16 792.337
R515 VSS.n45 VSS.n44 767.294
R516 VSS.n8 VSS.n3 767.294
R517 VSS.n52 VSS.n51 763.106
R518 VSS.n38 VSS.n37 763.106
R519 VSS.n51 VSS.n15 732.236
R520 VSS.n37 VSS.n34 732.236
R521 VSS.n44 VSS.n20 732.236
R522 VSS.n8 VSS.n1 732.236
R523 VSS.n181 VSS.n6 708.047
R524 VSS.t34 VSS.t19 708.047
R525 VSS.t16 VSS.t66 708.047
R526 VSS.t49 VSS.t53 708.047
R527 VSS.t46 VSS.t14 708.047
R528 VSS.n164 VSS.t9 681.482
R529 VSS.t19 VSS 564.751
R530 VSS.t53 VSS 564.751
R531 VSS VSS.t46 564.751
R532 VSS.n182 VSS 564.751
R533 VSS.t38 VSS.t47 554.492
R534 VSS.t14 VSS.t3 522.606
R535 VSS.n181 VSS.t38 513.419
R536 VSS.t13 VSS 480.461
R537 VSS.t6 VSS 459.26
R538 VSS.t9 VSS 459.26
R539 VSS.t47 VSS.t33 431.272
R540 VSS.t3 VSS.t26 387.74
R541 VSS VSS.t64 370.37
R542 VSS VSS.t21 370.37
R543 VSS.t42 VSS 370.37
R544 VSS.t33 VSS 343.991
R545 VSS.n135 VSS.t59 337.166
R546 VSS.n179 VSS.n57 334.815
R547 VSS.n46 VSS.n45 325.502
R548 VSS.n185 VSS.n3 325.502
R549 VSS.n135 VSS.t40 320.307
R550 VSS.n53 VSS.n52 304.204
R551 VSS.n39 VSS.n38 304.204
R552 VSS.t59 VSS 295.019
R553 VSS.n180 VSS.t6 278.519
R554 VSS VSS.t62 261.303
R555 VSS.t64 VSS.t44 248.889
R556 VSS.t21 VSS.t23 248.889
R557 VSS.t29 VSS.t31 248.889
R558 VSS.t36 VSS.t42 248.889
R559 VSS.t0 VSS 244.445
R560 VSS.n53 VSS.n13 242.448
R561 VSS.n39 VSS.n24 242.448
R562 VSS.n46 VSS.n18 242.448
R563 VSS.n186 VSS.n185 242.448
R564 VSS.n10 VSS.t18 241.579
R565 VSS.n153 VSS.t63 240.575
R566 VSS.n133 VSS.t56 237.327
R567 VSS VSS.n179 222.222
R568 VSS.n164 VSS 222.222
R569 VSS.n112 VSS.t68 218.308
R570 VSS.n88 VSS.t69 218.308
R571 VSS.n70 VSS.t70 218.308
R572 VSS.n140 VSS.t71 218.308
R573 VSS.n109 VSS.t10 214.456
R574 VSS.n111 VSS.t11 214.456
R575 VSS.n122 VSS.t7 214.456
R576 VSS.n89 VSS.t8 214.456
R577 VSS.n65 VSS.t4 214.456
R578 VSS.n69 VSS.t5 214.456
R579 VSS.n145 VSS.t1 214.456
R580 VSS.n139 VSS.t2 214.456
R581 VSS.n127 VSS.n126 204.457
R582 VSS.n78 VSS.n77 200.231
R583 VSS.n83 VSS.n82 200.231
R584 VSS.n72 VSS.n67 200.105
R585 VSS.t44 VSS 198.519
R586 VSS.t23 VSS 198.519
R587 VSS VSS.t29 198.519
R588 VSS VSS.t36 198.519
R589 VSS.n45 VSS.n17 195
R590 VSS.t25 VSS.n17 195
R591 VSS.n19 VSS.n16 195
R592 VSS.t25 VSS.n16 195
R593 VSS.n38 VSS.n23 195
R594 VSS.t12 VSS.n23 195
R595 VSS.n33 VSS.n22 195
R596 VSS.t12 VSS.n22 195
R597 VSS.n52 VSS.n12 195
R598 VSS.n12 VSS.t28 195
R599 VSS.n14 VSS.n11 195
R600 VSS.n11 VSS.t28 195
R601 VSS.n4 VSS.n2 195
R602 VSS.n57 VSS.n4 195
R603 VSS.n5 VSS.n3 195
R604 VSS.t18 VSS.n5 195
R605 VSS VSS.t51 177.012
R606 VSS.n36 VSS.n35 174.921
R607 VSS.n42 VSS.t25 163.988
R608 VSS.n49 VSS.t28 163.85
R609 VSS.n100 VSS.t65 162.471
R610 VSS.n95 VSS.t22 162.471
R611 VSS.n177 VSS.t32 162.471
R612 VSS.n172 VSS.t43 162.471
R613 VSS.n154 VSS.t17 162.471
R614 VSS.n78 VSS.t50 160.046
R615 VSS.n83 VSS.t35 160.046
R616 VSS.n91 VSS.t45 160.017
R617 VSS.n58 VSS.t24 160.017
R618 VSS.n61 VSS.t30 160.017
R619 VSS.n170 VSS.t37 160.017
R620 VSS.n161 VSS.t54 160.017
R621 VSS.n156 VSS.t67 160.017
R622 VSS.n153 VSS.t20 158.534
R623 VSS.n184 VSS.n183 152.552
R624 VSS VSS.t18 121.481
R625 VSS.n41 VSS.n21 105.025
R626 VSS.n48 VSS.n7 98.5767
R627 VSS.n56 VSS.n55 98.4942
R628 VSS.t31 VSS.n57 85.9264
R629 VSS.t66 VSS.t13 84.2917
R630 VSS.n67 VSS.t15 72.8576
R631 VSS.n126 VSS.t48 72.8576
R632 VSS.t25 VSS.n7 65.4109
R633 VSS.n56 VSS.t28 65.3562
R634 VSS.n35 VSS.n21 58.925
R635 VSS.n77 VSS.t52 58.5719
R636 VSS.n82 VSS.t41 58.5719
R637 VSS.t57 VSS.t34 50.5752
R638 VSS.t60 VSS.t49 50.5752
R639 VSS.n125 VSS 43.9579
R640 VSS.n128 VSS.n125 34.6358
R641 VSS.n132 VSS.n85 34.6358
R642 VSS.n15 VSS.n14 30.8711
R643 VSS.n34 VSS.n33 30.8711
R644 VSS.n20 VSS.n19 30.8711
R645 VSS.n2 VSS.n1 30.8711
R646 VSS.n165 VSS.n63 26.9246
R647 VSS.n146 VSS.n132 25.6926
R648 VSS.n77 VSS.t61 25.4291
R649 VSS.n82 VSS.t58 25.4291
R650 VSS.n100 VSS.n99 25.224
R651 VSS.n99 VSS.n91 25.224
R652 VSS.n95 VSS.n94 25.224
R653 VSS.n94 VSS.n58 25.224
R654 VSS.n177 VSS.n176 25.224
R655 VSS.n176 VSS.n61 25.224
R656 VSS.n172 VSS.n171 25.224
R657 VSS.n171 VSS.n170 25.224
R658 VSS.n161 VSS.n160 25.224
R659 VSS.n155 VSS.n154 25.224
R660 VSS.n156 VSS.n155 25.224
R661 VSS.n183 VSS.t18 24.1956
R662 VSS.n153 VSS.n152 24.0946
R663 VSS.n67 VSS.t27 22.3257
R664 VSS.n126 VSS.t39 22.3257
R665 VSS.n160 VSS.n78 21.4593
R666 VSS.n152 VSS.n83 21.4593
R667 VSS.n95 VSS.n91 20.3299
R668 VSS.n172 VSS.n61 20.3299
R669 VSS.n101 VSS.n100 19.2926
R670 VSS.n161 VSS.n76 17.7867
R671 VSS.n178 VSS.n177 17.3181
R672 VSS.t55 VSS.t0 16.8587
R673 VSS.n178 VSS.n58 15.8123
R674 VSS.n170 VSS.n63 15.8123
R675 VSS.n108 VSS.n63 14.775
R676 VSS.n138 VSS.n137 14.775
R677 VSS.n154 VSS.n153 13.5534
R678 VSS.n124 VSS.n123 11.2844
R679 VSS.n47 VSS.n46 11.0382
R680 VSS.n48 VSS.n47 11.0382
R681 VSS.n44 VSS.n43 11.0382
R682 VSS.n43 VSS.n42 11.0382
R683 VSS.n40 VSS.n39 11.0382
R684 VSS.n41 VSS.n40 11.0382
R685 VSS.n37 VSS.n36 11.0382
R686 VSS.n54 VSS.n53 11.0382
R687 VSS.n55 VSS.n54 11.0382
R688 VSS.n51 VSS.n50 11.0382
R689 VSS.n50 VSS.n49 11.0382
R690 VSS.n9 VSS.n8 11.0382
R691 VSS.n10 VSS.n9 11.0382
R692 VSS.n185 VSS.n184 11.0382
R693 VSS.n14 VSS.n13 10.9181
R694 VSS.n33 VSS.n24 10.9181
R695 VSS.n19 VSS.n18 10.9181
R696 VSS.n186 VSS.n2 10.9181
R697 VSS.n27 VSS.n15 10.4476
R698 VSS.n34 VSS.n32 10.4476
R699 VSS.n25 VSS.n20 10.4476
R700 VSS.n187 VSS.n1 10.4476
R701 VSS.n156 VSS.n78 10.1652
R702 VSS.n111 VSS.n106 9.70901
R703 VSS.n123 VSS.n122 9.70901
R704 VSS.n69 VSS.n68 9.70901
R705 VSS.n127 VSS.n85 9.41227
R706 VSS.n166 VSS.n165 9.3005
R707 VSS.n170 VSS.n169 9.3005
R708 VSS.n174 VSS.n61 9.3005
R709 VSS.n178 VSS.n59 9.3005
R710 VSS.n92 VSS.n58 9.3005
R711 VSS.n97 VSS.n91 9.3005
R712 VSS.n102 VSS.n101 9.3005
R713 VSS.n120 VSS.n119 9.3005
R714 VSS.n121 VSS.n87 9.3005
R715 VSS.n100 VSS.n90 9.3005
R716 VSS.n99 VSS.n98 9.3005
R717 VSS.n96 VSS.n95 9.3005
R718 VSS.n94 VSS.n93 9.3005
R719 VSS.n177 VSS.n60 9.3005
R720 VSS.n176 VSS.n175 9.3005
R721 VSS.n173 VSS.n172 9.3005
R722 VSS.n171 VSS.n62 9.3005
R723 VSS.n114 VSS.n113 9.3005
R724 VSS.n110 VSS.n105 9.3005
R725 VSS.n108 VSS.n107 9.3005
R726 VSS.n168 VSS.n63 9.3005
R727 VSS.n147 VSS.n146 9.3005
R728 VSS.n144 VSS.n143 9.3005
R729 VSS.n84 VSS.n83 9.3005
R730 VSS.n153 VSS.n81 9.3005
R731 VSS.n158 VSS.n78 9.3005
R732 VSS.n71 VSS.n66 9.3005
R733 VSS.n74 VSS.n73 9.3005
R734 VSS.n76 VSS.n75 9.3005
R735 VSS.n162 VSS.n161 9.3005
R736 VSS.n160 VSS.n159 9.3005
R737 VSS.n157 VSS.n156 9.3005
R738 VSS.n155 VSS.n79 9.3005
R739 VSS.n154 VSS.n80 9.3005
R740 VSS.n152 VSS.n151 9.3005
R741 VSS.n138 VSS.n134 9.3005
R742 VSS.n142 VSS.n141 9.3005
R743 VSS.n132 VSS.n131 9.3005
R744 VSS.n130 VSS.n85 9.3005
R745 VSS.n129 VSS.n128 9.3005
R746 VSS.n125 VSS.n86 9.3005
R747 VSS.n137 VSS.n136 9.3005
R748 VSS.n31 VSS.n30 8.45078
R749 VSS.n188 VSS.n0 8.30267
R750 VSS.n29 VSS.n28 7.97888
R751 VSS.n30 VSS.n26 7.97601
R752 VSS.n28 VSS.n27 7.16724
R753 VSS.n32 VSS.n31 7.16724
R754 VSS.n26 VSS.n25 7.16724
R755 VSS.n188 VSS.n187 7.16724
R756 VSS.n137 VSS.n83 7.15344
R757 VSS.n167 VSS.n163 6.50373
R758 VSS.n128 VSS.n127 6.4005
R759 VSS.n113 VSS.n110 6.26433
R760 VSS.n121 VSS.n120 6.26433
R761 VSS.n110 VSS.n109 5.85582
R762 VSS.n122 VSS.n121 5.85582
R763 VSS.n73 VSS.n65 5.85582
R764 VSS.n145 VSS.n144 5.85582
R765 VSS.n141 VSS.n133 5.85582
R766 VSS.n168 VSS.n167 4.788
R767 VSS.n27 VSS.n13 4.73093
R768 VSS.n32 VSS.n24 4.73093
R769 VSS.n25 VSS.n18 4.73093
R770 VSS.n187 VSS.n186 4.73093
R771 VSS.n167 VSS.n166 4.50726
R772 VSS.n103 VSS 4.01425
R773 VSS.n72 VSS.n71 3.40476
R774 VSS.n113 VSS.n112 3.13241
R775 VSS.n120 VSS.n88 3.13241
R776 VSS.n71 VSS.n70 3.13241
R777 VSS.n141 VSS.n140 3.13241
R778 VSS.n149 VSS.n148 2.88636
R779 VSS.n73 VSS.n72 2.86007
R780 VSS.n112 VSS.n111 2.7239
R781 VSS.n89 VSS.n88 2.7239
R782 VSS.n70 VSS.n69 2.7239
R783 VSS.n140 VSS.n139 2.7239
R784 VSS.n118 VSS.n117 1.753
R785 VSS.n116 VSS.n115 1.753
R786 VSS.n150 VSS.n149 1.21169
R787 VSS.n117 VSS.n116 0.761313
R788 VSS.n117 VSS.n104 0.591917
R789 VSS.n149 VSS 0.531208
R790 VSS.n104 VSS.n103 0.506165
R791 VSS.n30 VSS.n29 0.467019
R792 VSS.n109 VSS.n108 0.409011
R793 VSS.n101 VSS.n89 0.409011
R794 VSS.n76 VSS.n65 0.409011
R795 VSS.n146 VSS.n145 0.409011
R796 VSS.n144 VSS.n133 0.409011
R797 VSS.n139 VSS.n138 0.409011
R798 VSS.n103 VSS.n0 0.198729
R799 VSS.n166 VSS.n64 0.1255
R800 VSS.n123 VSS.n87 0.120292
R801 VSS.n119 VSS.n87 0.120292
R802 VSS.n98 VSS.n90 0.120292
R803 VSS.n98 VSS.n97 0.120292
R804 VSS.n96 VSS.n93 0.120292
R805 VSS.n93 VSS.n92 0.120292
R806 VSS.n175 VSS.n60 0.120292
R807 VSS.n175 VSS.n174 0.120292
R808 VSS.n173 VSS.n62 0.120292
R809 VSS.n169 VSS.n62 0.120292
R810 VSS.n107 VSS.n105 0.120292
R811 VSS.n114 VSS.n106 0.120292
R812 VSS.n129 VSS.n86 0.120292
R813 VSS.n130 VSS.n129 0.120292
R814 VSS.n131 VSS.n130 0.120292
R815 VSS.n142 VSS.n134 0.120292
R816 VSS.n80 VSS.n79 0.120292
R817 VSS.n157 VSS.n79 0.120292
R818 VSS.n159 VSS.n158 0.120292
R819 VSS.n75 VSS.n74 0.120292
R820 VSS.n74 VSS.n66 0.120292
R821 VSS.n68 VSS.n66 0.120292
R822 VSS VSS.n142 0.0981562
R823 VSS VSS.n124 0.09425
R824 VSS.n116 VSS 0.0881354
R825 VSS.n29 VSS.n0 0.0766574
R826 VSS.n115 VSS.n114 0.0721146
R827 VSS.n151 VSS.n150 0.0708125
R828 VSS.n28 VSS 0.064875
R829 VSS.n26 VSS 0.064875
R830 VSS VSS.n188 0.064875
R831 VSS.n31 VSS 0.063625
R832 VSS.n119 VSS.n118 0.0616979
R833 VSS.n90 VSS 0.0603958
R834 VSS VSS.n96 0.0603958
R835 VSS VSS.n59 0.0603958
R836 VSS.n60 VSS 0.0603958
R837 VSS VSS.n173 0.0603958
R838 VSS VSS.n168 0.0603958
R839 VSS.n107 VSS 0.0603958
R840 VSS.n131 VSS 0.0603958
R841 VSS.n143 VSS 0.0603958
R842 VSS.n136 VSS 0.0603958
R843 VSS VSS.n84 0.0603958
R844 VSS.n151 VSS 0.0603958
R845 VSS VSS.n81 0.0603958
R846 VSS VSS.n80 0.0603958
R847 VSS.n158 VSS 0.0603958
R848 VSS.n159 VSS 0.0603958
R849 VSS.n75 VSS 0.0603958
R850 VSS.n118 VSS.n102 0.0590938
R851 VSS.n163 VSS 0.0590938
R852 VSS.n150 VSS.n84 0.0499792
R853 VSS.n115 VSS.n105 0.0486771
R854 VSS.n148 VSS 0.0460729
R855 VSS.n147 VSS 0.0343542
R856 VSS VSS.n59 0.0330521
R857 VSS.n136 VSS 0.0330521
R858 VSS VSS.n64 0.03175
R859 VSS.n104 VSS 0.0292529
R860 VSS.n35 VSS.t12 0.028591
R861 VSS.n102 VSS 0.0226354
R862 VSS.n97 VSS 0.0226354
R863 VSS.n92 VSS 0.0226354
R864 VSS.n174 VSS 0.0226354
R865 VSS.n169 VSS 0.0226354
R866 VSS.n106 VSS 0.0226354
R867 VSS.n143 VSS 0.0226354
R868 VSS VSS.n134 0.0226354
R869 VSS.n81 VSS 0.0226354
R870 VSS VSS.n157 0.0226354
R871 VSS.n162 VSS 0.0226354
R872 VSS.n68 VSS 0.0226354
R873 VSS.n148 VSS.n147 0.0148229
R874 VSS.n124 VSS.n86 0.00440625
R875 VSS.n168 VSS.n64 0.00180208
R876 VSS.n163 VSS.n162 0.00180208
R877 x2.GP4.n2 x2.GP4.t4 450.938
R878 x2.GP4.n2 x2.GP4.t5 445.666
R879 x1.x14.Y x2.GP4.n4 203.923
R880 x2.GP4.n0 x2.GP4.n1 101.49
R881 x2.GP4.n4 x2.GP4.t3 26.5955
R882 x2.GP4.n4 x2.GP4.t0 26.5955
R883 x2.GP4.n1 x2.GP4.t2 24.9236
R884 x2.GP4.n1 x2.GP4.t1 24.9236
R885 x1.gpo3 x2.x4.GP 16.5752
R886 x2.GP4.n3 x1.x14.Y 10.7525
R887 x2.GP4.n0 x1.gpo3 7.7042
R888 x2.GP4.n3 x1.x14.Y 6.6565
R889 x1.x14.Y x2.GP4.n3 5.04292
R890 x2.x4.GP x2.GP4.n2 2.95993
R891 x1.x14.Y x2.GP4.n0 2.5605
R892 x2.GP4.n0 x1.x14.Y 1.93989
R893 Z4.n1 Z4.t3 23.6581
R894 Z4.n3 Z4.t2 23.3739
R895 Z4.n1 Z4.t0 10.7528
R896 Z4.n0 Z4.t1 10.6417
R897 Z4.n2 Z4.n1 1.30064
R898 Z4 Z4.n4 0.983856
R899 Z4.n3 Z4.n2 0.726502
R900 Z4.n2 Z4.n0 0.512491
R901 Z4.n4 Z4.n0 0.359663
R902 Z4.n4 Z4.n3 0.216071
R903 A4.n1 A4.t3 26.3998
R904 A4.n1 A4.t2 23.5483
R905 A4.n0 A4.t1 12.7127
R906 A4.n0 A4.t0 10.8578
R907 A4.n2 A4.n1 3.12177
R908 A4.n2 A4.n0 1.81453
R909 A4.n3 A4.n2 1.1255
R910 A4 A4.n3 0.203263
R911 A4.n3 A4 0.0655
R912 select1.n10 select1.t1 327.99
R913 select1.n3 select1.t8 293.969
R914 select1.n6 select1.t3 256.07
R915 select1.n1 select1.t2 212.081
R916 select1.n0 select1.t5 212.081
R917 select1.n10 select1.t9 199.457
R918 select1.n2 select1.n1 182.929
R919 select1 select1.n3 154.065
R920 select1.n11 select1.n10 152
R921 select1.n7 select1.n6 152
R922 select1.n6 select1.t7 150.03
R923 select1.n1 select1.t6 139.78
R924 select1.n0 select1.t0 139.78
R925 select1.n3 select1.t4 138.338
R926 select1.n1 select1.n0 61.346
R927 select1.n5 select1 22.1096
R928 select1.n14 select1.n13 14.6836
R929 select1.n13 select1.n12 14.6704
R930 select1.n12 select1 13.8672
R931 select1.n4 select1 13.8328
R932 select1.n11 select1 12.1605
R933 select1.n14 select1.n2 10.6811
R934 select1.n7 select1.n5 10.4374
R935 select1.n9 select1.n8 8.15359
R936 select1.n2 select1 6.1445
R937 select1.n4 select1 5.16179
R938 select1.n9 select1.n4 4.65206
R939 select1.n8 select1 3.93896
R940 select1 select1.n11 2.34717
R941 select1.n5 select1 2.16665
R942 select1.n8 select1.n7 1.57588
R943 select1.n13 select1.n9 0.79438
R944 select1.n12 select1 0.6405
R945 select1 select1.n14 0.248606
R946 x2.GN1.n1 x2.GN1.t6 377.486
R947 x2.GN1.n1 x2.GN1.t4 374.202
R948 x2.GN1.n7 x2.GN1.t0 339.418
R949 x2.GN1.n0 x2.GN1.t1 274.06
R950 x2.GN1.n4 x2.GN1.t5 212.081
R951 x2.GN1.n3 x2.GN1.t7 212.081
R952 x2.GN1.n5 x2.GN1.n4 182.673
R953 x2.GN1.n4 x2.GN1.t2 139.78
R954 x2.GN1.n3 x2.GN1.t3 139.78
R955 x2.GN1.n4 x2.GN1.n3 61.346
R956 x2.GN1 x2.GN1.n5 15.8606
R957 x2.GN1 x2.GN1.n6 13.8044
R958 x2.GN1.n2 x2.GN1 11.5859
R959 x2.GN1 x2.GN1.n0 11.0989
R960 x2.GN1 x2.GN1.n2 10.8756
R961 x2.GN1.n6 x2.GN1 8.1246
R962 x2.GN1.n8 x2.GN1 6.6565
R963 x2.GN1.n5 x2.GN1 6.4005
R964 x2.GN1.n0 x2.GN1 6.1445
R965 x2.GN1.n2 x2.GN1 4.55738
R966 x2.GN1.n8 x2.GN1.n7 4.0914
R967 x2.GN1 x2.GN1.n8 3.61789
R968 x2.GN1.n6 x2.GN1 3.26325
R969 x2.GN1.n0 x2.GN1 2.86947
R970 x2.GN1 x2.GN1.n1 2.04102
R971 x2.GN1.n7 x2.GN1 1.74382
R972 x2.GN4.n1 x2.GN4.t6 377.486
R973 x2.GN4.n1 x2.GN4.t7 374.202
R974 x2.GN4.n7 x2.GN4.t0 339.418
R975 x2.GN4.n0 x2.GN4.t1 274.06
R976 x2.GN4.n4 x2.GN4.t2 212.081
R977 x2.GN4.n3 x2.GN4.t3 212.081
R978 x2.GN4.n5 x2.GN4.n4 184.977
R979 x2.GN4.n4 x2.GN4.t4 139.78
R980 x2.GN4.n3 x2.GN4.t5 139.78
R981 x2.GN4.n4 x2.GN4.n3 61.346
R982 x2.GN4.n6 x2.GN4 18.2601
R983 x2.GN4 x2.GN4.n2 17.2682
R984 x2.GN4 x2.GN4.n5 15.0136
R985 x2.GN4 x2.GN4.n0 11.2645
R986 x2.GN4 x2.GN4.n6 8.9605
R987 x2.GN4.n6 x2.GN4 8.4485
R988 x2.GN4.n2 x2.GN4 8.16743
R989 x2.GN4.n8 x2.GN4 6.6565
R990 x2.GN4.n0 x2.GN4 6.1445
R991 x2.GN4.n2 x2.GN4 4.58237
R992 x2.GN4.n5 x2.GN4 4.0965
R993 x2.GN4.n8 x2.GN4.n7 4.0914
R994 x2.GN4 x2.GN4.n8 3.61789
R995 x2.GN4.n0 x2.GN4 2.86947
R996 x2.GN4 x2.GN4.n1 2.04102
R997 x2.GN4.n7 x2.GN4 1.74382
R998 select2.n1 select2.t0 212.081
R999 select2.n0 select2.t1 212.081
R1000 select2.n2 select2.n1 183.441
R1001 select2.n1 select2.t2 139.78
R1002 select2.n0 select2.t3 139.78
R1003 select2.n1 select2.n0 61.346
R1004 select2 select2.n2 11.4331
R1005 select2.n2 select2 5.6325
R1006 nselect2.n5 nselect2.n4 196.339
R1007 nselect2.n1 nselect2.n0 101.49
R1008 nselect2.n4 nselect2.t0 26.5955
R1009 nselect2.n4 nselect2.t1 26.5955
R1010 nselect2.n0 nselect2.t2 24.9236
R1011 nselect2.n0 nselect2.t3 24.9236
R1012 nselect2.n2 nselect2 13.5685
R1013 nselect2.n3 nselect2 10.7525
R1014 nselect2.n6 nselect2.n2 9.50196
R1015 nselect2.n6 nselect2.n5 7.64514
R1016 nselect2.n5 nselect2 7.58449
R1017 nselect2.n3 nselect2 6.6565
R1018 nselect2 nselect2.n3 5.04292
R1019 nselect2 nselect2.n2 3.8405
R1020 nselect2 nselect2.n1 2.5605
R1021 nselect2.n1 nselect2 1.93989
R1022 nselect2 nselect2.n6 1.81877
R1023 Z3.n1 Z3.t2 23.6581
R1024 Z3.n3 Z3.t3 23.3739
R1025 Z3.n1 Z3.t0 10.7528
R1026 Z3.n0 Z3.t1 10.6417
R1027 Z3.n2 Z3.n1 1.30064
R1028 Z3.n5 Z3.n4 0.924585
R1029 Z3.n3 Z3.n2 0.726502
R1030 Z3.n2 Z3.n0 0.512491
R1031 Z3.n4 Z3.n0 0.359663
R1032 Z3.n4 Z3.n3 0.216071
R1033 Z3.n5 Z3 0.0656042
R1034 Z3 Z3.n5 0.0376287
R1035 A3.n1 A3.t2 26.3998
R1036 A3.n1 A3.t3 23.5483
R1037 A3.n0 A3.t0 12.7127
R1038 A3.n0 A3.t1 10.8578
R1039 A3.n2 A3.n1 3.12177
R1040 A3.n2 A3.n0 1.81453
R1041 A3.n3 A3.n2 1.1255
R1042 A3.n3 A3 0.210543
R1043 A3 A3.n3 0.0655
C0 x2.GN1 x2.GN3 0.00286f
C1 x2.GN3 a_5275_n2995# 1.07e-20
C2 a_5275_n3507# A1 5.02e-20
C3 x2.GN2 x1.nSEL0 0.154394f
C4 x2.GN1 x1.nSEL1 0.034891f
C5 a_5275_n4059# x1.nSEL0 0.001174f
C6 select0 select2 0.368835f
C7 x2.GN2 a_5275_n4235# 0.106186f
C8 select1 x2.GN2 0.108649f
C9 A4 x2.GN4 3.83736f
C10 a_5275_n4059# a_5275_n4235# 0.185422f
C11 a_5275_n4059# select1 0.254026f
C12 x1.nSEL0 x2.GN4 2.26e-20
C13 A4 VDD 1.54289f
C14 x1.nSEL0 VDD 0.391764f
C15 m3_8196_n3226# x2.GN3 0.001446f
C16 x2.GN3 a_5301_n4107# 5.17e-20
C17 A2 A1 1.81909f
C18 select1 x2.GN4 0.059813f
C19 select1 VDD 2.64545f
C20 a_5275_n4235# VDD 0.161854f
C21 A4 A3 2.08862f
C22 x2.GN3 select2 0.001055f
C23 m3_8196_n3226# m3_9240_n3230# 0.003764f
C24 m2_5406_n4650# select0 0.130999f
C25 x1.nSEL1 a_5301_n4107# 9.57e-19
C26 x1.nSEL1 select2 0.164723f
C27 x2.GN3 Z2 0.00126f
C28 a_5329_n4513# a_5275_n4651# 0.006584f
C29 nselect2 a_5275_n3507# 6.01e-20
C30 x2.GP3 a_5275_n3507# 5.21e-19
C31 Z3 x2.GN3 0.427085f
C32 x2.GN2 select0 0.114345f
C33 a_5275_n4059# select0 0.143958f
C34 x2.GP3 A1 0.001277f
C35 x1.nSEL1 m2_5406_n4650# 0.00815f
C36 x2.GN4 select0 0.218396f
C37 select0 VDD 1.09594f
C38 a_5275_n3683# a_5275_n3507# 0.185422f
C39 a_5275_n3683# A1 1.55e-21
C40 a_5301_n3555# x2.GP3 4.39e-19
C41 A2 x2.GP3 0.001826f
C42 x2.GN2 x2.GN3 0.067572f
C43 a_5275_n4059# x2.GN3 0.048646f
C44 x2.GN3 x2.GN4 0.07149f
C45 x2.GN3 VDD 0.649708f
C46 x1.nSEL1 x2.GN2 0.209956f
C47 a_5301_n3555# a_5275_n3683# 0.004764f
C48 x1.nSEL1 a_5275_n4059# 0.041068f
C49 x2.GN1 a_5275_n3507# 3.78e-20
C50 m3_9240_n3230# x2.GN2 0.016745f
C51 x2.GN1 A1 4.61808f
C52 x2.GN4 m3_10270_n3216# 0.084813f
C53 x2.GN3 A3 3.80482f
C54 Z1 select0 4.1e-22
C55 x1.nSEL1 VDD 0.481997f
C56 m3_9240_n3230# x2.GN4 7.07e-19
C57 select1 x1.nSEL0 0.137403f
C58 x1.nSEL0 a_5275_n4235# 0.03096f
C59 x2.GN1 a_5275_n4651# 0.12869f
C60 x2.GN1 A2 1.78e-19
C61 m3_9240_n3230# A3 0.097296f
C62 Z4 x2.GP3 0.071646f
C63 select1 a_5275_n4235# 0.03417f
C64 x2.GN3 Z1 4.42e-20
C65 x2.GN1 a_5329_n4513# 0.001144f
C66 nselect2 a_5275_n3683# 1.29e-19
C67 x2.GP3 a_5275_n3683# 0.00144f
C68 m3_8196_n3226# A2 0.1002f
C69 Z2 A1 0.004942f
C70 x2.GN1 x2.GP3 0.002439f
C71 x1.nSEL0 select0 0.324538f
C72 nselect2 a_5275_n2995# 9.77e-20
C73 Z3 A1 4.74e-21
C74 select1 select0 1.66811f
C75 a_5275_n4235# select0 0.246189f
C76 Z2 A2 4.51569f
C77 x2.GN1 a_5275_n3683# 6.43e-20
C78 a_5329_n2857# a_5275_n2995# 0.006584f
C79 A4 x2.GN3 0.004656f
C80 m2_5406_n4650# a_5275_n4651# 0.01297f
C81 x2.GN3 x1.nSEL0 4.01e-20
C82 m3_8196_n3226# x2.GP3 9.67e-19
C83 Z3 A2 0.004565f
C84 x2.GN2 a_5275_n3507# 5.62e-20
C85 nselect2 select2 0.150826f
C86 A4 m3_10270_n3216# 0.091998f
C87 select1 x2.GN3 0.272312f
C88 x2.GN2 A1 0.157008f
C89 x2.GN3 a_5275_n4235# 6.68e-19
C90 x1.nSEL1 x1.nSEL0 0.352716f
C91 A4 m3_9240_n3230# 6.07e-21
C92 x2.GN4 a_5275_n3507# 0.003699f
C93 a_5275_n3507# VDD 0.262185f
C94 x2.GN4 A1 0.001437f
C95 VDD A1 1.98654f
C96 x1.nSEL1 a_5275_n4235# 0.073392f
C97 x1.nSEL1 select1 0.272823f
C98 x2.GN2 a_5275_n4651# 0.039612f
C99 x2.GN2 A2 3.81441f
C100 x2.GN2 a_5301_n3555# 3.11e-20
C101 a_5275_n3683# select2 0.009143f
C102 Z2 x2.GP3 1.03e-20
C103 x2.GN2 a_5329_n4513# 8.86e-19
C104 x2.GN4 A2 3.42e-19
C105 a_5301_n3555# x2.GN4 3.22e-19
C106 a_5275_n4651# VDD 0.210313f
C107 A2 VDD 1.61513f
C108 a_5301_n3555# VDD 0.001496f
C109 x2.GN1 m3_8196_n3226# 6.03e-20
C110 Z3 x2.GP3 0.278332f
C111 x2.GN1 a_5301_n4107# 1.22e-20
C112 Z3 Z4 0.002229f
C113 x2.GN1 select2 0.009187f
C114 A2 A3 1.81997f
C115 a_5329_n4513# VDD 9.09e-19
C116 Z1 A1 4.51491f
C117 x2.GN3 select0 0.254198f
C118 x2.GN2 x2.GP3 0.004319f
C119 x2.GN1 Z2 4.77e-21
C120 x1.nSEL1 select0 0.168464f
C121 x2.GN2 a_5329_n2857# 8.14e-21
C122 nselect2 x2.GN4 1.53e-20
C123 nselect2 VDD 1.06761f
C124 x2.GN4 x2.GP3 3.44338f
C125 x2.GN1 m2_5406_n4650# 0.06935f
C126 x2.GP3 VDD 1.78272f
C127 Z4 x2.GN4 0.443708f
C128 Z4 VDD 2.81281f
C129 x2.GN2 a_5275_n3683# 1.63e-19
C130 a_5275_n4059# a_5275_n3683# 3.02e-19
C131 x2.GN4 a_5329_n2857# 0.001562f
C132 a_5329_n2857# VDD 8.97e-19
C133 x2.GN3 m3_10270_n3216# 0.016026f
C134 x2.GP3 A3 4.01143f
C135 Z4 A3 0.005563f
C136 x1.nSEL1 x2.GN3 0.012418f
C137 x2.GN4 a_5275_n3683# 6.84e-19
C138 m3_9240_n3230# x2.GN3 0.087318f
C139 a_5275_n3683# VDD 0.171441f
C140 m3_9240_n3230# m3_10270_n3216# 0.003741f
C141 x2.GN1 x2.GN2 0.065209f
C142 x2.GN1 a_5275_n4059# 1.46e-19
C143 x1.nSEL0 a_5275_n3507# 1.21e-20
C144 Z1 x2.GP3 7.56e-20
C145 x1.nSEL0 A1 1.93e-21
C146 m2_5406_n4650# select2 4.4e-19
C147 x2.GN1 x2.GN4 0.001075f
C148 select1 a_5275_n3507# 0.127717f
C149 x2.GN2 a_5275_n2995# 7.58e-21
C150 x2.GN1 VDD 1.36505f
C151 select1 A1 1.45e-21
C152 x1.nSEL0 a_5275_n4651# 0.081627f
C153 A4 A2 2.39e-19
C154 x2.GN4 a_5275_n2995# 0.134079f
C155 a_5275_n2995# VDD 0.217381f
C156 m3_8196_n3226# x2.GN2 0.099332f
C157 x2.GN2 a_5301_n4107# 0.002418f
C158 a_5275_n4235# a_5275_n4651# 0.002207f
C159 select1 a_5275_n4651# 0.02803f
C160 Z3 Z2 7.65e-19
C161 x2.GN2 select2 0.001308f
C162 a_5275_n4059# select2 1.67e-19
C163 m3_8196_n3226# x2.GN4 7.17e-19
C164 a_5301_n4107# VDD 4.32e-19
C165 x2.GN1 Z1 0.428262f
C166 VDD select2 0.231538f
C167 x2.GN2 Z2 0.427019f
C168 select0 a_5275_n3507# 0.279858f
C169 A4 x2.GP3 0.161499f
C170 A4 Z4 4.51497f
C171 select0 A1 3.49e-20
C172 Z2 VDD 2.85288f
C173 select1 nselect2 0.001177f
C174 Z3 x2.GN2 2.12e-20
C175 select1 x2.GP3 0.003386f
C176 m2_5406_n4650# VDD 0.139545f
C177 Z2 A3 1.49e-20
C178 x1.nSEL0 a_5275_n3683# 1.91e-20
C179 a_5275_n4651# select0 0.048888f
C180 select1 a_5329_n2857# 8.84e-19
C181 Z3 x2.GN4 0.00128f
C182 a_5301_n3555# select0 0.001558f
C183 x2.GN3 a_5275_n3507# 0.004288f
C184 Z3 VDD 2.85668f
C185 x2.GN3 A1 0.002069f
C186 select1 a_5275_n3683# 0.261734f
C187 a_5329_n4513# select0 9.55e-19
C188 Z3 A3 4.51555f
C189 a_5275_n4059# x2.GN2 0.017018f
C190 x1.nSEL1 a_5275_n3507# 1.59e-19
C191 x2.GN1 x1.nSEL0 0.004383f
C192 x2.GN3 a_5301_n3555# 0.001073f
C193 x2.GN3 A2 0.164396f
C194 x2.GN2 x2.GN4 8.84e-19
C195 x2.GN2 VDD 0.600374f
C196 a_5275_n4059# VDD 0.19314f
C197 x2.GN1 a_5275_n4235# 0.012466f
C198 x2.GN1 select1 0.312198f
C199 x2.GN2 A3 0.004147f
C200 x1.nSEL1 a_5275_n4651# 0.193944f
C201 x2.GN4 VDD 1.23434f
C202 x1.nSEL1 a_5301_n3555# 4.08e-19
C203 nselect2 select0 1.88e-19
C204 select0 x2.GP3 2.82e-19
C205 select1 a_5275_n2995# 0.125445f
C206 x1.nSEL1 a_5329_n4513# 0.00175f
C207 x2.GN4 A3 0.187073f
C208 A3 VDD 1.61205f
C209 a_5329_n2857# select0 1.4e-19
C210 x1.nSEL0 a_5301_n4107# 2.51e-19
C211 x2.GN2 Z1 7.73e-19
C212 select0 a_5275_n3683# 0.086353f
C213 x1.nSEL0 select2 0.131218f
C214 nselect2 x2.GN3 7.39e-21
C215 x2.GN3 x2.GP3 2.868f
C216 a_5301_n4107# a_5275_n4235# 0.004764f
C217 Z4 x2.GN3 1.95e-20
C218 a_5275_n4235# select2 8.66e-20
C219 select1 select2 0.139336f
C220 x2.GN3 a_5329_n2857# 1.07e-20
C221 Z1 VDD 2.90992f
C222 m3_10270_n3216# x2.GP3 0.006132f
C223 x1.nSEL1 nselect2 0.047548f
C224 x2.GN3 a_5275_n3683# 0.104343f
C225 m3_9240_n3230# x2.GP3 0.002824f
C226 x2.GN1 select0 0.020307f
C227 x1.nSEL0 m2_5406_n4650# 3.43e-19
C228 a_5275_n2995# select0 0.220366f
C229 x1.nSEL1 a_5275_n3683# 7.84e-19
C230 select1 m2_5406_n4650# 0.183786f
C231 Z4 VSS 2.703709f
C232 A4 VSS 3.673923f
C233 Z3 VSS 2.48903f
C234 A3 VSS 3.139328f
C235 Z2 VSS 2.454758f
C236 A2 VSS 3.238628f
C237 Z1 VSS 2.838278f
C238 A1 VSS 3.972252f
C239 nselect2 VSS 0.47102f
C240 select2 VSS 1.16504f
C241 select0 VSS 1.41757f
C242 select1 VSS 1.610708f
C243 VDD VSS 56.37729f
C244 m3_10270_n3216# VSS 0.090191f $ **FLOATING
C245 m3_9240_n3230# VSS 0.086003f $ **FLOATING
C246 m3_8196_n3226# VSS 0.168273f $ **FLOATING
C247 m2_5406_n4650# VSS 0.065655f $ **FLOATING
C248 a_5329_n4513# VSS 0.006505f
C249 a_5275_n4651# VSS 0.266782f
C250 x1.nSEL0 VSS 0.649982f
C251 x2.GN1 VSS 6.355386f
C252 a_5301_n4107# VSS 0.004461f
C253 a_5275_n4235# VSS 0.220868f
C254 x1.nSEL1 VSS 0.69132f
C255 x2.GN2 VSS 3.93258f
C256 a_5275_n4059# VSS 0.23458f
C257 x2.GP3 VSS 1.67788f
C258 a_5301_n3555# VSS 0.006801f
C259 x2.GN3 VSS 3.65509f
C260 a_5275_n3683# VSS 0.232764f
C261 a_5275_n3507# VSS 0.249604f
C262 x2.GN4 VSS 7.590769f
C263 a_5329_n2857# VSS 0.006439f
C264 a_5275_n2995# VSS 0.306675f
C265 A3.t0 VSS 0.893857f
C266 A3.t1 VSS 0.513146f
C267 A3.n0 VSS 4.9699f
C268 A3.t2 VSS 0.925152f
C269 A3.t3 VSS 0.654459f
C270 A3.n1 VSS 5.08132f
C271 A3.n2 VSS 0.803733f
C272 A3.n3 VSS 0.264783f
C273 Z3.t1 VSS 0.362117f
C274 Z3.n0 VSS 0.540706f
C275 Z3.t0 VSS 0.369386f
C276 Z3.t2 VSS 0.490183f
C277 Z3.n1 VSS 2.47361f
C278 Z3.n2 VSS 0.836966f
C279 Z3.t3 VSS 0.477048f
C280 Z3.n3 VSS 0.593305f
C281 Z3.n4 VSS 0.728891f
C282 Z3.n5 VSS 0.331987f
C283 x2.GN4.t1 VSS 0.06076f
C284 x2.GN4.n0 VSS 0.070042f
C285 x2.GN4.t6 VSS 0.686652f
C286 x2.GN4.t7 VSS 0.670085f
C287 x2.GN4.n1 VSS 3.00641f
C288 x2.GN4.n2 VSS 1.54718f
C289 x2.GN4.t2 VSS 0.038143f
C290 x2.GN4.t4 VSS 0.022477f
C291 x2.GN4.t3 VSS 0.038143f
C292 x2.GN4.t5 VSS 0.022477f
C293 x2.GN4.n3 VSS 0.063998f
C294 x2.GN4.n4 VSS 0.094806f
C295 x2.GN4.n5 VSS 0.042443f
C296 x2.GN4.n6 VSS 0.343794f
C297 x2.GN4.t0 VSS 0.155177f
C298 x2.GN4.n7 VSS 0.027911f
C299 x2.GN4.n8 VSS 0.031268f
C300 x2.GN1.t1 VSS 0.029997f
C301 x2.GN1.n0 VSS 0.034614f
C302 x2.GN1.t6 VSS 0.338995f
C303 x2.GN1.t4 VSS 0.330816f
C304 x2.GN1.n1 VSS 1.48424f
C305 x2.GN1.n2 VSS 0.51776f
C306 x2.GN1.t5 VSS 0.018831f
C307 x2.GN1.t2 VSS 0.011097f
C308 x2.GN1.t7 VSS 0.018831f
C309 x2.GN1.t3 VSS 0.011097f
C310 x2.GN1.n3 VSS 0.031595f
C311 x2.GN1.n4 VSS 0.046667f
C312 x2.GN1.n5 VSS 0.045389f
C313 x2.GN1.n6 VSS 0.098587f
C314 x2.GN1.t0 VSS 0.076609f
C315 x2.GN1.n7 VSS 0.013779f
C316 x2.GN1.n8 VSS 0.015437f
C317 select1.t2 VSS 0.032343f
C318 select1.t6 VSS 0.019059f
C319 select1.t5 VSS 0.032343f
C320 select1.t0 VSS 0.019059f
C321 select1.n0 VSS 0.054267f
C322 select1.n1 VSS 0.080179f
C323 select1.n2 VSS 0.048819f
C324 select1.t4 VSS 0.014966f
C325 select1.t8 VSS 0.031563f
C326 select1.n3 VSS 0.113336f
C327 select1.n4 VSS 0.021975f
C328 select1.n5 VSS 0.018928f
C329 select1.t3 VSS 0.022802f
C330 select1.t7 VSS 0.015669f
C331 select1.n6 VSS 0.06626f
C332 select1.n7 VSS 0.015263f
C333 select1.n8 VSS 0.109332f
C334 select1.n9 VSS 0.396f
C335 select1.t1 VSS 0.02778f
C336 select1.t9 VSS 0.018863f
C337 select1.n10 VSS 0.065634f
C338 select1.n11 VSS 0.01571f
C339 select1.n12 VSS 0.101902f
C340 select1.n13 VSS 0.457083f
C341 select1.n14 VSS 0.597136f
C342 A4.t1 VSS 0.893325f
C343 A4.t0 VSS 0.512841f
C344 A4.n0 VSS 4.96695f
C345 A4.t3 VSS 0.924602f
C346 A4.t2 VSS 0.65407f
C347 A4.n1 VSS 5.0783f
C348 A4.n2 VSS 0.803255f
C349 A4.n3 VSS 0.258761f
C350 Z4.t1 VSS 0.356817f
C351 Z4.n0 VSS 0.532792f
C352 Z4.t0 VSS 0.363979f
C353 Z4.t3 VSS 0.483009f
C354 Z4.n1 VSS 2.43741f
C355 Z4.n2 VSS 0.824716f
C356 Z4.t2 VSS 0.470066f
C357 Z4.n3 VSS 0.584621f
C358 Z4.n4 VSS 0.742893f
C359 x2.GP4.n0 VSS 0.095571f
C360 x2.x4.GP VSS 2.50543f
C361 x1.gpo3 VSS 1.18077f
C362 x2.GP4.t2 VSS 0.012052f
C363 x2.GP4.t1 VSS 0.012052f
C364 x2.GP4.n1 VSS 0.028739f
C365 x1.x14.Y VSS 0.104168f
C366 x2.GP4.t5 VSS 0.609957f
C367 x2.GP4.t4 VSS 0.626965f
C368 x2.GP4.n2 VSS 2.22891f
C369 x2.GP4.n3 VSS 0.017567f
C370 x2.GP4.t3 VSS 0.018542f
C371 x2.GP4.t0 VSS 0.018542f
C372 x2.GP4.n4 VSS 0.040723f
C373 A1.t0 VSS 0.813767f
C374 A1.t3 VSS 0.467169f
C375 A1.n0 VSS 4.5246f
C376 A1.t2 VSS 0.842259f
C377 A1.t1 VSS 0.59582f
C378 A1.n1 VSS 4.62603f
C379 A1.n2 VSS 0.731718f
C380 A1.n3 VSS 0.224671f
C381 Z1.t0 VSS 0.363377f
C382 Z1.n0 VSS 0.542586f
C383 Z1.t3 VSS 0.370671f
C384 Z1.t1 VSS 0.491889f
C385 Z1.n1 VSS 2.48222f
C386 Z1.n2 VSS 0.839878f
C387 Z1.t2 VSS 0.478707f
C388 Z1.n3 VSS 0.595368f
C389 Z1.n4 VSS 0.756551f
C390 x2.x1.GP VSS 1.98566f
C391 x2.GP1.t1 VSS 0.012716f
C392 x2.GP1.t0 VSS 0.012716f
C393 x2.GP1.n0 VSS 0.03032f
C394 x1.x11.Y VSS 0.046385f
C395 x2.GP1.n1 VSS 0.059566f
C396 x2.GP1.n2 VSS 0.018534f
C397 x2.GP1.t3 VSS 0.019563f
C398 x2.GP1.t2 VSS 0.019563f
C399 x2.GP1.n3 VSS 0.040309f
C400 x2.GP1.t5 VSS 0.643518f
C401 x2.GP1.t4 VSS 0.661463f
C402 x2.GP1.n4 VSS 2.33672f
C403 x1.gpo0 VSS 0.626909f
C404 x2.GP1.n5 VSS 0.086057f
C405 VDD.n0 VSS 0.03081f
C406 VDD.n1 VSS 0.137121f
C407 VDD.n2 VSS 0.066225f
C408 VDD.n3 VSS 0.557756f
C409 VDD.n4 VSS 0.557756f
C410 VDD.n5 VSS 0.091797f
C411 VDD.n6 VSS 0.067234f
C412 VDD.t3 VSS 0.741619f
C413 VDD.n9 VSS 0.067234f
C414 VDD.n10 VSS 2.85e-19
C415 VDD.n11 VSS 0.040828f
C416 VDD.n12 VSS 0.007424f
C417 VDD.n13 VSS 0.080708f
C418 VDD.n14 VSS 0.043153f
C419 VDD.n15 VSS 0.08763f
C420 VDD.n16 VSS 0.101662f
C421 VDD.n17 VSS 0.137121f
C422 VDD.n18 VSS 0.002226f
C423 VDD.n19 VSS 0.091797f
C424 VDD.n20 VSS 0.067234f
C425 VDD.t70 VSS 0.741619f
C426 VDD.n22 VSS 0.557756f
C427 VDD.n23 VSS 0.067234f
C428 VDD.n25 VSS 0.557756f
C429 VDD.n26 VSS 0.066225f
C430 VDD.n27 VSS 0.00533f
C431 VDD.n28 VSS 0.040787f
C432 VDD.n29 VSS 0.007491f
C433 VDD.n30 VSS 0.080708f
C434 VDD.n31 VSS 0.042812f
C435 VDD.n32 VSS 0.069384f
C436 VDD.n33 VSS 0.099666f
C437 VDD.n34 VSS 0.137121f
C438 VDD.n35 VSS 0.002362f
C439 VDD.n36 VSS 0.091797f
C440 VDD.n37 VSS 0.067234f
C441 VDD.t19 VSS 0.741619f
C442 VDD.n39 VSS 0.557756f
C443 VDD.n40 VSS 0.067234f
C444 VDD.n42 VSS 0.557756f
C445 VDD.n43 VSS 0.066225f
C446 VDD.n44 VSS 0.005339f
C447 VDD.n45 VSS 0.040651f
C448 VDD.n46 VSS 0.007491f
C449 VDD.n47 VSS 0.080708f
C450 VDD.n48 VSS 0.042812f
C451 VDD.n49 VSS 0.067641f
C452 VDD.n50 VSS 0.103727f
C453 VDD.n51 VSS 0.137121f
C454 VDD.n52 VSS 0.007292f
C455 VDD.n53 VSS 0.066225f
C456 VDD.n54 VSS 0.557756f
C457 VDD.n55 VSS 0.557756f
C458 VDD.n56 VSS 0.091797f
C459 VDD.n57 VSS 0.067234f
C460 VDD.t53 VSS 0.741619f
C461 VDD.n60 VSS 0.067234f
C462 VDD.n61 VSS 2.58e-19
C463 VDD.n62 VSS 0.040828f
C464 VDD.n63 VSS 0.007451f
C465 VDD.n64 VSS 0.080708f
C466 VDD.n65 VSS 0.043126f
C467 VDD.n66 VSS 0.246672f
C468 VDD.n67 VSS 0.187384f
C469 VDD.n68 VSS 0.004178f
C470 VDD.t34 VSS 0.008431f
C471 VDD.n69 VSS 0.008293f
C472 VDD.t18 VSS 9.05e-19
C473 VDD.t5 VSS 0.001375f
C474 VDD.n70 VSS 0.002375f
C475 VDD.t36 VSS 0.008593f
C476 VDD.t69 VSS 0.008431f
C477 VDD.n71 VSS 0.008031f
C478 VDD.n72 VSS 0.004178f
C479 VDD.n73 VSS 0.003782f
C480 VDD.t44 VSS 0.001241f
C481 VDD.n74 VSS 0.003521f
C482 VDD.t55 VSS 0.005101f
C483 VDD.n75 VSS 0.004695f
C484 VDD.n76 VSS 0.00419f
C485 VDD.t46 VSS 0.008433f
C486 VDD.n77 VSS 6.9e-19
C487 VDD.t42 VSS 0.003616f
C488 VDD.t11 VSS 0.005969f
C489 VDD.n78 VSS 0.005884f
C490 VDD.n79 VSS 0.007052f
C491 VDD.t71 VSS 0.024909f
C492 VDD.n80 VSS 0.02253f
C493 VDD.t32 VSS 6.76e-19
C494 VDD.t14 VSS 0.001812f
C495 VDD.n81 VSS 0.008269f
C496 VDD.t12 VSS 0.005969f
C497 VDD.n82 VSS 0.004367f
C498 VDD.n83 VSS 0.0163f
C499 VDD.n84 VSS 0.012878f
C500 VDD.n85 VSS 0.016727f
C501 VDD.n86 VSS 0.009658f
C502 VDD.n87 VSS 0.007052f
C503 VDD.n88 VSS 0.005289f
C504 VDD.n89 VSS 0.00332f
C505 VDD.n90 VSS 0.010459f
C506 VDD.n91 VSS 0.016397f
C507 VDD.t47 VSS 0.016948f
C508 VDD.n92 VSS 0.001276f
C509 VDD.n93 VSS 0.001303f
C510 VDD.n94 VSS 0.005289f
C511 VDD.n95 VSS 0.001629f
C512 VDD.t9 VSS 0.008547f
C513 VDD.n96 VSS 0.007014f
C514 VDD.n97 VSS 0.004178f
C515 VDD.t74 VSS 0.024909f
C516 VDD.n98 VSS 0.006209f
C517 VDD.n99 VSS 0.004178f
C518 VDD.t38 VSS 6.76e-19
C519 VDD.t21 VSS 0.001812f
C520 VDD.n100 VSS 0.008269f
C521 VDD.t72 VSS 0.024909f
C522 VDD.t7 VSS 0.003616f
C523 VDD.n101 VSS 0.011165f
C524 VDD.n102 VSS 0.006401f
C525 VDD.n103 VSS 0.00332f
C526 VDD.t1 VSS 0.005969f
C527 VDD.n104 VSS 0.005884f
C528 VDD.n105 VSS 0.02253f
C529 VDD.n106 VSS 0.009658f
C530 VDD.n107 VSS 0.016727f
C531 VDD.t2 VSS 0.005969f
C532 VDD.t63 VSS 0.008548f
C533 VDD.n108 VSS 0.002415f
C534 VDD.n109 VSS 0.002875f
C535 VDD.t6 VSS 0.034122f
C536 VDD.t20 VSS 0.032992f
C537 VDD.t0 VSS 0.024405f
C538 VDD.t37 VSS 0.035026f
C539 VDD.t29 VSS 0.034122f
C540 VDD.t27 VSS 0.038867f
C541 VDD.t49 VSS 0.028246f
C542 VDD.t15 VSS 0.01514f
C543 VDD.t8 VSS 0.007005f
C544 VDD.t62 VSS 0.024631f
C545 VDD.n110 VSS 0.032141f
C546 VDD.n111 VSS 0.02229f
C547 VDD.n112 VSS 0.006552f
C548 VDD.n113 VSS 0.010512f
C549 VDD.n114 VSS 0.012878f
C550 VDD.n115 VSS 0.004369f
C551 VDD.n116 VSS 0.034804f
C552 VDD.n117 VSS 0.047342f
C553 VDD.t23 VSS 0.005969f
C554 VDD.n118 VSS 0.011672f
C555 VDD.n119 VSS 0.02253f
C556 VDD.n120 VSS 0.013884f
C557 VDD.t24 VSS 0.005969f
C558 VDD.t65 VSS 0.008589f
C559 VDD.n121 VSS 0.010036f
C560 VDD.t22 VSS 0.076766f
C561 VDD.t57 VSS 0.047161f
C562 VDD.t25 VSS 0.019351f
C563 VDD.t51 VSS 0.026784f
C564 VDD.t66 VSS 0.019351f
C565 VDD.t60 VSS 0.026784f
C566 VDD.t39 VSS 0.019351f
C567 VDD.t64 VSS 0.028963f
C568 VDD.n122 VSS 0.031705f
C569 VDD.n123 VSS 0.004178f
C570 VDD.n124 VSS 0.001819f
C571 VDD.t61 VSS 0.008589f
C572 VDD.n125 VSS 0.001819f
C573 VDD.t52 VSS 0.008589f
C574 VDD.n126 VSS 0.122759f
C575 VDD.n127 VSS 0.007185f
C576 VDD.n128 VSS 0.004367f
C577 VDD.t73 VSS 0.025299f
C578 VDD.t58 VSS 0.005969f
C579 VDD.n129 VSS 0.025046f
C580 VDD.n130 VSS 0.012447f
C581 VDD.t59 VSS 0.005969f
C582 VDD.n131 VSS 0.0163f
C583 VDD.n132 VSS 0.014991f
C584 VDD.n133 VSS 0.009406f
C585 VDD.n134 VSS 0.00734f
C586 VDD.n135 VSS 0.007158f
C587 VDD.t26 VSS 0.008593f
C588 VDD.n136 VSS 0.010814f
C589 VDD.n137 VSS 0.004178f
C590 VDD.n138 VSS 0.007052f
C591 VDD.n139 VSS 0.005289f
C592 VDD.n140 VSS 0.010144f
C593 VDD.t67 VSS 0.008593f
C594 VDD.n141 VSS 0.010977f
C595 VDD.n142 VSS 0.004178f
C596 VDD.n143 VSS 0.007052f
C597 VDD.n144 VSS 0.005289f
C598 VDD.n145 VSS 0.010144f
C599 VDD.t40 VSS 0.008593f
C600 VDD.n146 VSS 0.010977f
C601 VDD.n147 VSS 0.001819f
C602 VDD.n148 VSS 0.007052f
C603 VDD.n149 VSS 0.005289f
C604 VDD.n150 VSS 0.002683f
C605 VDD.n151 VSS 0.014656f
C606 VDD.n152 VSS 0.006552f
C607 VDD.n153 VSS 0.010512f
C608 VDD.n154 VSS 0.017908f
C609 VDD.n155 VSS 0.003564f
C610 VDD.n156 VSS 0.032389f
C611 VDD.n157 VSS 0.031406f
C612 VDD.n158 VSS 7.28e-19
C613 VDD.t16 VSS 9.05e-19
C614 VDD.t50 VSS 0.001375f
C615 VDD.n159 VSS 0.002375f
C616 VDD.n160 VSS 0.015943f
C617 VDD.t28 VSS 0.008589f
C618 VDD.n161 VSS 0.010009f
C619 VDD.t56 VSS 0.00283f
C620 VDD.t48 VSS 0.007522f
C621 VDD.n162 VSS 0.004267f
C622 VDD.t30 VSS 0.008433f
C623 VDD.n163 VSS 0.008897f
C624 VDD.n164 VSS 0.011444f
C625 VDD.n165 VSS 0.001507f
C626 VDD.n166 VSS 0.007052f
C627 VDD.n167 VSS 0.004178f
C628 VDD.n168 VSS 0.002415f
C629 VDD.n169 VSS 0.002683f
C630 VDD.n170 VSS 0.01436f
C631 VDD.n171 VSS 0.039157f
C632 VDD.t17 VSS 0.007457f
C633 VDD.t33 VSS 0.019434f
C634 VDD.t35 VSS 0.021693f
C635 VDD.t4 VSS 0.01514f
C636 VDD.t43 VSS 0.028246f
C637 VDD.t68 VSS 0.039771f
C638 VDD.t45 VSS 0.019434f
C639 VDD.t54 VSS 0.01514f
C640 VDD.t31 VSS 0.035026f
C641 VDD.t10 VSS 0.024405f
C642 VDD.t13 VSS 0.032992f
C643 VDD.t41 VSS 0.034122f
C644 VDD.n172 VSS 0.023237f
C645 VDD.n173 VSS 0.006751f
C646 VDD.n174 VSS 0.004805f
C647 VDD.n175 VSS 0.001276f
C648 VDD.n176 VSS 0.009362f
C649 VDD.n177 VSS 0.003571f
C650 VDD.n178 VSS 0.007052f
C651 VDD.n179 VSS 0.005289f
C652 VDD.n180 VSS 0.003144f
C653 VDD.n181 VSS 0.010688f
C654 VDD.n182 VSS 0.007648f
C655 VDD.n183 VSS 0.004868f
C656 VDD.n184 VSS 0.013764f
C657 VDD.n185 VSS 0.087548f
C658 A2.t2 VSS 0.763965f
C659 A2.t3 VSS 0.438578f
C660 A2.n0 VSS 4.2477f
C661 A2.t1 VSS 0.790712f
C662 A2.t0 VSS 0.559356f
C663 A2.n1 VSS 4.34292f
C664 A2.n2 VSS 0.686937f
C665 A2.n3 VSS 0.222065f
C666 Z2.t3 VSS 0.363425f
C667 Z2.n0 VSS 0.542659f
C668 Z2.t2 VSS 0.37072f
C669 Z2.t1 VSS 0.491954f
C670 Z2.n1 VSS 2.48255f
C671 Z2.n2 VSS 0.83999f
C672 Z2.t0 VSS 0.478771f
C673 Z2.n3 VSS 0.595448f
C674 Z2.n4 VSS 0.733795f
C675 Z2.n5 VSS 0.3243f
C676 x2.x2.GP VSS 2.76866f
C677 x1.gpo1 VSS 0.998586f
C678 x2.GP2.t3 VSS 0.016016f
C679 x2.GP2.t2 VSS 0.016016f
C680 x2.GP2.n0 VSS 0.03819f
C681 x1.x12.Y VSS 0.058128f
C682 x2.GP2.n1 VSS 0.075027f
C683 x2.GP2.n2 VSS 0.023344f
C684 x2.GP2.t1 VSS 0.02464f
C685 x2.GP2.t0 VSS 0.02464f
C686 x2.GP2.n3 VSS 0.050813f
C687 x2.GP2.t5 VSS 0.810542f
C688 x2.GP2.t4 VSS 0.833144f
C689 x2.GP2.n4 VSS 2.95587f
C690 x2.GP2.n5 VSS 0.106388f
.ends

