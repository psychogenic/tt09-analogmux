* NGSPICE file created from simplecounter_parax.ext - technology: sky130A

.subckt simplecounter_parax clk enable counter[1] counter[3] counter[5] counter[6]
+ counter[7] counter[8] counter[0] counter[2] counter[4] counter[9] VPWR VGND
X0 a_2431_7497# a_2302_7241# a_2011_7351# VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1 VGND.t700 a_2502_7396# a_2431_7497# VGND.t699 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X2 VPWR.t386 a_4329_5461# clknet_0_clk.t15 VPWR.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VGND.t440 VPWR.t829 VGND.t439 VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X4 clknet_0_clk.t31 a_4329_5461# VGND.t693 VGND.t692 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR.t687 VGND.t817 VPWR.t686 VPWR.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6 VGND.t538 a_5814_4399# clknet_1_1__leaf_clk.t31 VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR.t332 _05_ a_5333_5321# VPWR.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X8 VGND.t443 VPWR.t830 VGND.t442 VGND.t441 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X9 _17_ a_6375_5309# VGND.t595 VGND.t594 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X10 VGND.t445 VPWR.t831 VGND.t444 VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X11 VPWR.t118 a_6425_2388# counter[6].t0 VPWR.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X12 VGND.t328 VPWR.t832 VGND.t327 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X13 VPWR.t684 VGND.t818 VPWR.t683 VPWR.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X14 VGND.t477 clknet_0_clk.t32 a_5814_4399# VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 VGND.t331 VPWR.t833 VGND.t330 VGND.t329 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X16 a_2673_4233# a_1683_3861# a_2547_3855# VGND.t599 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X17 VPWR.t749 net1 a_1499_7119# VPWR.t748 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X18 a_4454_4649# _17_ a_4382_4649# VPWR.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X19 a_3225_4399# a_2235_4399# a_3099_4765# VGND.t263 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 _04_ a_3215_3829# VGND.t765 VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X21 a_2471_2741# a_2614_2883# VPWR.t320 VPWR.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X22 net10 a_7683_3829# VPWR.t240 VPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND.t334 VPWR.t834 VGND.t333 VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X24 VPWR.t681 VGND.t819 VPWR.t680 VPWR.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X25 VGND.t691 a_4329_5461# clknet_0_clk.t30 VGND.t690 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 VPWR.t342 _23_ a_7019_4943# VPWR.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_4413_3311# _15_ a_4341_3311# VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_5599_2741# net7 VPWR.t352 VPWR.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X29 VGND.t695 a_3849_2388# counter[3].t1 VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X30 VGND.t337 VPWR.t835 VGND.t336 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X31 VPWR.t678 VGND.t820 VPWR.t677 VPWR.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X32 clknet_1_0__leaf_clk.t31 a_1845_5461# VGND.t584 VGND.t583 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 a_2840_3087# net5 VGND.t548 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 a_4349_3855# _15_ VPWR.t305 VPWR.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X35 a_7199_4943# a_7019_4943# VPWR.t316 VPWR.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X36 a_6427_2741# _11_.t4 VPWR.t120 VPWR.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X37 VPWR.t307 _17_ a_3799_4943# VPWR.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X38 VPWR.t303 _15_ a_6427_2741# VPWR.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 VGND.t340 VPWR.t836 VGND.t339 VGND.t338 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X40 VPWR.t29 a_2745_2388# counter[2].t0 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X41 VPWR.t384 a_4329_5461# clknet_0_clk.t14 VPWR.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X42 VPWR.t675 VGND.t821 VPWR.t674 VPWR.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X43 VPWR.t94 clknet_1_1__leaf_clk.t32 a_6651_3861# VPWR.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X44 a_1845_5461# clknet_0_clk.t33 VPWR.t769 VPWR.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X45 VPWR.t672 VGND.t822 VPWR.t671 VPWR.t670 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X46 a_3979_4943# a_3799_4943# VPWR.t56 VPWR.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X47 VGND.t281 a_3267_4667# a_3225_4399# VGND.t280 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X48 VPWR.t138 a_1457_2388# counter[0].t0 VPWR.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X49 VGND.t427 a_5675_3855# a_5843_3829# VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X50 net11 a_7683_3579# VGND.t230 VGND.t229 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X51 clknet_1_1__leaf_clk.t15 a_5814_4399# VPWR.t228 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X52 a_2125_8527# net2.t2 VGND.t414 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X53 VPWR.t723 a_2502_7637# a_2431_7663# VPWR.t722 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X54 a_1825_2388# net3.t2 VPWR.t96 VPWR.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X55 a_7363_3087# _15_ a_7267_3087# VGND.t612 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X56 VPWR.t719 a_7258_3829# a_7185_3855# VPWR.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X57 VGND.t723 _21_ a_4995_4399# VGND.t722 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X58 VPWR.t272 a_1845_5461# clknet_1_0__leaf_clk.t15 VPWR.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X59 a_7753_2767# _23_ VPWR.t340 VPWR.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 VPWR.t669 VGND.t823 VPWR.t668 VPWR.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X61 a_6043_3677# a_5345_3311# a_5786_3423# VGND.t746 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X62 a_2823_3677# a_1959_3311# a_2566_3423# VPWR.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X63 clknet_1_1__leaf_clk.t30 a_5814_4399# VGND.t536 VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X64 VPWR.t667 VGND.t824 VPWR.t666 VPWR.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X65 a_7185_3855# a_6651_3861# a_7090_3855# VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X66 a_4329_5461# clk.t0 VPWR.t751 VPWR.t750 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X67 a_1915_7351# a_2011_7351# VPWR.t392 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X68 VPWR.t665 VGND.t825 VPWR.t664 VPWR.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X69 VGND.t362 _16_.t2 a_5436_4399# VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.06615 ps=0.735 w=0.42 l=0.15
X70 VGND.t343 VPWR.t837 VGND.t342 VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X71 VGND.t689 a_4329_5461# clknet_0_clk.t29 VGND.t688 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X72 VGND.t31 _14_ _02_ VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X73 a_2823_3677# a_2125_3311# a_2566_3423# VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X74 VPWR.t662 VGND.t826 VPWR.t661 VPWR.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X75 VGND.t346 VPWR.t838 VGND.t345 VGND.t344 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X76 VGND.t297 a_6425_2388# counter[6].t1 VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X77 VGND.t349 VPWR.t839 VGND.t348 VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X78 VPWR.t791 a_2991_3579# a_2907_3677# VPWR.t790 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X79 VGND.t239 _22_ a_7363_3087# VGND.t238 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X80 VPWR.t132 clknet_1_0__leaf_clk.t32 a_1683_3861# VPWR.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X81 VPWR.t689 a_2502_7396# a_2431_7497# VPWR.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X82 VPWR.t382 a_4329_5461# clknet_0_clk.t13 VPWR.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X83 VGND.t352 VPWR.t840 VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X84 VGND.t304 VPWR.t841 VGND.t303 VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X85 clknet_0_clk.t28 a_4329_5461# VGND.t687 VGND.t686 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X86 a_6375_5309# net6.t2 VPWR.t136 VPWR.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X87 VPWR.t660 VGND.t827 VPWR.t659 VPWR.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X88 _24_ a_7077_2767# VGND.t789 VGND.t788 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X89 a_5801_4233# a_4811_3861# a_5675_3855# VGND.t643 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X90 VGND.t582 a_1845_5461# clknet_1_0__leaf_clk.t30 VGND.t581 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X91 a_7171_2767# net10 a_7077_2767# VPWR.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X92 VPWR.t658 VGND.t828 VPWR.t657 VPWR.t656 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X93 _00_ a_1875_8207# a_2125_8207# VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X94 VPWR.t270 a_1845_5461# clknet_1_0__leaf_clk.t14 VPWR.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X95 VPWR.t35 a_8265_2388# counter[8].t0 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X96 VPWR.t655 VGND.t829 VPWR.t654 VPWR.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X97 VPWR.t653 VGND.t830 VPWR.t652 VPWR.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X98 a_7619_5162# _25_ VPWR.t805 VPWR.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X99 a_2217_3855# a_1683_3861# a_2122_3855# VPWR.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X100 VGND.t307 VPWR.t842 VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X101 clknet_0_clk.t3 a_4329_5461# VPWR.t380 VPWR.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X102 a_5077_4721# _21_ VPWR.t718 VPWR.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X103 VPWR.t80 net6.t3 a_5599_2741# VPWR.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X104 VGND.t52 a_2745_2388# counter[2].t1 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X105 VGND.t310 VPWR.t843 VGND.t309 VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X106 a_2125_3311# a_1959_3311# VGND.t814 VGND.t813 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X107 a_7515_3677# a_6651_3311# a_7258_3423# VPWR.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X108 a_7345_2388# net9 VPWR.t728 VPWR.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X109 a_4779_5161# clknet_1_1__leaf_clk.t33 VGND.t275 VGND.t274 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X110 VPWR.t650 VGND.t831 VPWR.t649 VPWR.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X111 VPWR.t647 VGND.t832 VPWR.t646 VPWR.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X112 VGND.t410 a_1457_2388# counter[0].t1 VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X113 clknet_1_0__leaf_clk.t13 a_1845_5461# VPWR.t268 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X114 a_1825_2388# net3.t3 VGND.t506 VGND.t505 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X115 a_7005_3855# _08_ VGND.t418 VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X116 VPWR.t644 VGND.t833 VPWR.t643 VPWR.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X117 a_2295_7337# clknet_1_0__leaf_clk.t33 VPWR.t176 VPWR.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X118 VGND.t312 VPWR.t844 VGND.t311 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X119 VGND.t314 VPWR.t845 VGND.t313 VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X120 VPWR.t106 net11 a_7939_2223# VPWR.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X121 a_7515_3677# a_6817_3311# a_7258_3423# VGND.t416 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X122 VPWR.t301 _15_ a_3831_3339# VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 _12_ net3.t4 a_1499_7119# VPWR.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X124 VPWR.t641 VGND.t834 VPWR.t640 VPWR.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X125 VGND.t534 a_5814_4399# clknet_1_1__leaf_clk.t29 VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X126 VPWR.t110 a_1915_7351# net3.t0 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X127 net4 a_2715_3829# VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X128 VPWR.t700 a_4585_2388# counter[4].t0 VPWR.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X129 VPWR.t60 a_7683_3579# a_7599_3677# VPWR.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X130 a_4737_4943# a_4399_5175# VPWR.t116 VPWR.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X131 a_7258_3423# a_7090_3677# VPWR.t752 VPWR.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X132 net10 a_7683_3829# VGND.t552 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X133 a_3917_3105# net4 a_3831_3105# VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X134 VGND.t316 VPWR.t846 VGND.t315 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X135 VGND.t705 _20_ a_4413_3311# VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X136 VPWR.t638 VGND.t835 VPWR.t637 VPWR.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X137 a_7005_3311# _09_ VGND.t729 VGND.t728 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X138 VGND.t56 _24_ a_7289_5309# VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X139 VPWR.t716 _21_ a_4520_4373# VPWR.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.1176 ps=1.4 w=0.42 l=0.15
X140 VPWR.t314 a_2561_9514# net1 VPWR.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X141 clknet_0_clk.t2 a_4329_5461# VPWR.t378 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X142 a_4915_5321# a_4779_5161# a_4495_5175# VPWR.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X143 a_5345_3311# a_5179_3311# VPWR.t46 VPWR.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X144 VGND.t319 VPWR.t847 VGND.t318 VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X145 VGND.t322 VPWR.t848 VGND.t321 VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X146 VGND.t277 clknet_1_1__leaf_clk.t34 a_5179_3311# VGND.t276 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X147 VGND.t727 a_6427_2741# _23_ VGND.t726 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X148 VGND.t29 _14_ a_2840_3087# VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X149 a_5250_3855# a_4977_3861# a_5165_3855# VPWR.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X150 a_7619_5162# _25_ VGND.t796 VGND.t795 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X151 a_1915_7351# a_2011_7351# VGND.t696 VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X152 a_4399_5175# a_4495_5175# VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X153 VPWR.t86 clknet_1_1__leaf_clk.t35 a_4811_3861# VPWR.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X154 VGND.t58 a_8265_2388# counter[8].t1 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X155 VGND.t325 VPWR.t849 VGND.t324 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X156 VPWR.t636 VGND.t836 VPWR.t635 VPWR.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X157 VPWR.t376 a_4329_5461# clknet_0_clk.t1 VPWR.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X158 VPWR.t633 VGND.t837 VPWR.t632 VPWR.t534 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X159 VGND.t532 a_5814_4399# clknet_1_1__leaf_clk.t28 VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X160 a_7345_2388# net9 VGND.t738 VGND.t737 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X161 VPWR.t178 clknet_1_0__leaf_clk.t34 a_1959_3311# VPWR.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X162 VGND.t63 VPWR.t850 VGND.t62 VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X163 VGND.t580 a_1845_5461# clknet_1_0__leaf_clk.t29 VGND.t579 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X164 VGND.t810 net8 a_4287_4399# VGND.t809 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X165 a_5599_2741# net9 VPWR.t726 VPWR.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X166 VPWR.t266 a_1845_5461# clknet_1_0__leaf_clk.t12 VPWR.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X167 a_2317_6575# net2.t3 a_2235_6575# VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X168 VPWR.t631 VGND.t838 VPWR.t630 VPWR.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X169 VGND.t287 net11 a_7939_2223# VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X170 a_3215_3829# _16_.t3 a_3601_3855# VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X171 a_6427_2741# _22_ VPWR.t70 VPWR.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X172 VGND.t639 _05_ a_5333_5321# VGND.t638 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X173 _25_ a_7199_4943# VPWR.t698 VPWR.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X174 a_5786_3423# a_5618_3677# VPWR.t40 VPWR.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X175 a_5786_3423# a_5618_3677# VGND.t208 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X176 _16_.t0 a_3831_3339# VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X177 a_4329_5461# clk.t1 VPWR.t322 VPWR.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X178 VGND.t270 clknet_1_1__leaf_clk.t36 a_6651_3861# VGND.t269 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X179 clknet_1_1__leaf_clk.t27 a_5814_4399# VGND.t530 VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X180 VPWR.t629 VGND.t839 VPWR.t628 VPWR.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X181 VPWR.t626 VGND.t840 VPWR.t625 VPWR.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X182 _19_ a_3979_4943# VGND.t787 VGND.t786 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X183 _06_ a_4454_4649# VGND.t603 VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X184 VGND.t709 a_4585_2388# counter[4].t1 VGND.t708 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X185 VPWR.t696 _20_ a_4259_3311# VPWR.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X186 VPWR.t624 VGND.t841 VPWR.t623 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X187 VPWR.t622 VGND.t842 VPWR.t621 VPWR.t620 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X188 VPWR.t619 VGND.t843 VPWR.t618 VPWR.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X189 VGND.t780 a_2295_7637# a_2302_7937# VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X190 a_2041_4649# _11_.t5 _13_ VPWR.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X191 VPWR.t812 a_5871_5162# _05_ VPWR.t811 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X192 a_2547_3855# a_1683_3861# a_2290_3829# VPWR.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X193 a_7019_4943# _23_ VGND.t650 VGND.t649 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X194 a_2401_4399# a_2235_4399# VGND.t262 VGND.t261 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X195 VGND.t792 a_2290_3829# a_2248_4233# VGND.t791 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X196 VGND.t66 VPWR.t851 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X197 _21_ a_4259_3311# VPWR.t42 VPWR.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X198 VGND.t731 clknet_0_clk.t34 a_5814_4399# VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X199 VGND.t43 clknet_0_clk.t35 a_1845_5461# VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X200 net8 a_5843_3829# VPWR.t50 VPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X201 a_5135_5309# a_4915_5321# VGND.t601 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X202 a_3831_3105# net4 VPWR.t710 VPWR.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X203 VPWR.t616 VGND.t844 VPWR.t615 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X204 a_3849_2388# net5 VPWR.t238 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X205 VPWR.t614 VGND.t845 VPWR.t613 VPWR.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X206 VGND.t622 a_2561_9514# net1 VGND.t621 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X207 a_3799_4943# _17_ VGND.t617 VGND.t616 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X208 a_6719_3133# _15_ a_6623_3133# VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X209 a_2253_8029# a_1915_7815# VPWR.t21 VPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X210 VGND.t289 a_1915_7351# net3.t1 VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X211 a_5149_4721# net9 a_5077_4721# VPWR.t724 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0441 ps=0.63 w=0.42 l=0.15
X212 clknet_0_clk.t0 a_4329_5461# VPWR.t374 VPWR.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X213 VGND.t299 clknet_1_1__leaf_clk.t37 a_6651_3311# VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X214 VPWR.t11 a_2715_3829# a_2631_3855# VPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X215 VGND.t69 VPWR.t852 VGND.t68 VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X216 clknet_1_0__leaf_clk.t28 a_1845_5461# VGND.t578 VGND.t577 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X217 a_2037_3855# _02_ VGND.t740 VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X218 VGND.t72 VPWR.t853 VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X219 VPWR.t264 a_1845_5461# clknet_1_0__leaf_clk.t11 VPWR.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X220 a_5505_2388# net7 VPWR.t350 VPWR.t349 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X221 VPWR.t226 a_5814_4399# clknet_1_1__leaf_clk.t14 VPWR.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X222 VPWR.t611 VGND.t846 VPWR.t610 VPWR.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X223 clknet_1_0__leaf_clk.t27 a_1845_5461# VGND.t576 VGND.t575 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X224 VGND.t659 net7 a_4220_3829# VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X225 VGND.t540 clknet_1_0__leaf_clk.t35 a_1683_3861# VGND.t539 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X226 clknet_0_clk.t8 a_4329_5461# VPWR.t372 VPWR.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X227 a_2614_2883# _16_.t4 VGND.t60 VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X228 net11 a_7683_3579# VPWR.t58 VPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X229 VPWR.t166 a_4220_3829# _18_ VPWR.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X230 VPWR.t609 VGND.t847 VPWR.t608 VPWR.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X231 VGND.t37 a_2842_4511# a_2800_4399# VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X232 clknet_1_1__leaf_clk.t26 a_5814_4399# VGND.t528 VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X233 VGND.t75 VPWR.t854 VGND.t74 VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X234 a_7267_3087# _11_.t6 a_7077_2767# VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X235 a_2431_7663# a_2295_7637# a_2011_7637# VPWR.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X236 a_6169_3311# a_5179_3311# a_6043_3677# VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X237 a_1505_3855# _13_ VPWR.t123 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X238 VGND.t78 VPWR.t855 VGND.t77 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X239 VGND.t81 VPWR.t856 VGND.t80 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X240 VPWR.t606 VGND.t848 VPWR.t605 VPWR.t604 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X241 VPWR.t820 net8 a_5599_2741# VPWR.t819 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X242 a_2253_7119# a_1915_7351# VPWR.t108 VPWR.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X243 clknet_1_0__leaf_clk.t10 a_1845_5461# VPWR.t262 VPWR.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X244 a_7090_3855# a_6817_3861# a_7005_3855# VPWR.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X245 clknet_1_1__leaf_clk.t13 a_5814_4399# VPWR.t224 VPWR.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X246 VPWR.t603 VGND.t849 VPWR.t602 VPWR.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X247 VPWR.t600 VGND.t850 VPWR.t599 VPWR.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X248 a_2235_6575# net3.t5 VPWR.t196 VPWR.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 VGND.t285 net11 a_7941_3087# VGND.t284 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X250 VPWR.t82 net6.t4 a_3245_3855# VPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 a_5618_3677# a_5345_3311# a_5533_3311# VPWR.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X252 VGND.t526 a_5814_4399# clknet_1_1__leaf_clk.t25 VGND.t525 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X253 a_5814_4399# clknet_0_clk.t36 VPWR.t767 VPWR.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X254 a_7005_3311# _09_ VPWR.t721 VPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X255 a_2949_3311# a_1959_3311# a_2823_3677# VGND.t812 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X256 VPWR.t72 clk.t2 a_4329_5461# VPWR.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X257 a_7289_5309# a_7019_4943# a_7199_4943# VGND.t623 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X258 a_2589_4399# _04_ VGND.t625 VGND.t624 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X259 a_6427_2741# net10 a_6825_3133# VGND.t589 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X260 VGND.t84 VPWR.t857 VGND.t83 VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X261 VPWR.t597 VGND.t851 VPWR.t596 VPWR.t595 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X262 VGND.t803 a_5871_5162# _05_ VGND.t802 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X263 VGND.t2 VPWR.t858 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X264 VGND.t775 a_2695_6575# _11_.t3 VGND.t774 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X265 a_8109_2767# net11 VPWR.t104 VPWR.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X266 a_2431_7497# a_2295_7337# a_2011_7351# VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X267 a_6457_5309# net6.t5 a_6375_5309# VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X268 a_3099_4765# a_2235_4399# a_2842_4511# VPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X269 VPWR.t594 VGND.t852 VPWR.t593 VPWR.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X270 VGND.t5 VPWR.t859 VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X271 VGND.t779 a_6211_3579# a_6169_3311# VGND.t778 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X272 VPWR.t7 a_5786_3423# a_5713_3677# VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X273 VPWR.t148 _11_.t7 a_4349_3855# VPWR.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X274 a_4454_4649# a_4520_4373# a_4287_4399# VGND.t219 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X275 a_1499_7119# net2.t4 VPWR.t158 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X276 _07_ a_5149_4721# VPWR.t170 VPWR.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14575 ps=1.335 w=1 l=0.15
X277 VGND.t8 VPWR.t860 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X278 _15_ a_3831_3105# VGND.t620 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X279 a_3849_2388# net5 VGND.t546 VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X280 net5 a_2991_3579# VGND.t785 VGND.t784 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X281 a_5713_3677# a_5179_3311# a_5618_3677# VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X282 VPWR.t591 VGND.t853 VPWR.t590 VPWR.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X283 VPWR.t589 VGND.t854 VPWR.t588 VPWR.t587 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X284 a_5675_3855# a_4811_3861# a_5418_3829# VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X285 VPWR.t586 VGND.t855 VPWR.t585 VPWR.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X286 VGND.t801 a_5418_3829# a_5376_4233# VGND.t800 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X287 a_2122_3855# a_1849_3861# a_2037_3855# VPWR.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X288 VPWR.t370 a_4329_5461# clknet_0_clk.t7 VPWR.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X289 _10_ a_2235_6575# VPWR.t25 VPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X290 VPWR.t100 a_3267_4667# a_3183_4765# VPWR.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X291 clknet_1_0__leaf_clk.t9 a_1845_5461# VPWR.t260 VPWR.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X292 VGND.t574 a_1845_5461# clknet_1_0__leaf_clk.t26 VGND.t573 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X293 VGND.t716 net4 _13_ VGND.t715 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X294 a_2614_2883# _16_.t5 VPWR.t38 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X295 a_3215_2999# net4 a_3389_3105# VGND.t714 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X296 a_4399_5175# a_4495_5175# VGND.t54 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X297 a_5505_2388# net7 VGND.t657 VGND.t656 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X298 VPWR.t584 VGND.t856 VPWR.t583 VPWR.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X299 VGND.t572 a_1845_5461# clknet_1_0__leaf_clk.t25 VGND.t571 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X300 VGND.t11 VPWR.t861 VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X301 VPWR.t150 _11_.t8 a_4259_3311# VPWR.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X302 _17_ a_6375_5309# VPWR.t283 VPWR.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X303 VGND.t524 a_5814_4399# clknet_1_1__leaf_clk.t24 VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X304 a_2389_6575# net3.t6 a_2317_6575# VGND.t471 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X305 VPWR.t48 a_5843_3829# a_5759_3855# VPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X306 a_3433_4175# _16_.t6 _04_ VGND.t271 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X307 VGND.t14 VPWR.t862 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X308 _09_ a_7723_2741# VGND.t798 VGND.t797 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X309 VPWR.t801 a_2290_3829# a_2217_3855# VPWR.t800 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X310 VPWR.t738 a_4779_5161# a_4786_5065# VPWR.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X311 a_4767_3463# net8 VPWR.t818 VPWR.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X312 a_2230_7485# a_1915_7351# VGND.t288 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X313 VGND.t17 VPWR.t863 VGND.t16 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X314 a_5165_3855# _06_ VGND.t483 VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X315 a_6651_5309# _11_.t9 a_6545_5309# VGND.t633 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X316 VGND.t19 VPWR.t864 VGND.t18 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X317 VGND.t550 a_7683_3829# a_7641_4233# VGND.t549 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X318 VGND.t301 clknet_1_1__leaf_clk.t38 a_4811_3861# VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X319 VPWR.t230 clknet_1_0__leaf_clk.t36 a_2235_4399# VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X320 VPWR.t222 a_5814_4399# clknet_1_1__leaf_clk.t12 VPWR.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X321 VGND.t242 VPWR.t865 VGND.t241 VGND.t240 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X322 a_5001_3311# net7 a_4929_3311# VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X323 VPWR.t582 VGND.t857 VPWR.t581 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X324 a_6127_3677# a_5345_3311# a_6043_3677# VPWR.t734 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X325 clknet_1_1__leaf_clk.t23 a_5814_4399# VGND.t522 VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X326 VPWR.t579 VGND.t858 VPWR.t578 VPWR.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X327 VGND.t245 VPWR.t866 VGND.t244 VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X328 VPWR.t576 VGND.t859 VPWR.t575 VPWR.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X329 VGND.t248 VPWR.t867 VGND.t247 VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X330 VPWR.t573 VGND.t860 VPWR.t572 VPWR.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X331 net8 a_5843_3829# VGND.t218 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X332 a_3245_3855# a_3215_3829# _04_ VPWR.t753 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X333 _00_ net1 a_2125_8527# VGND.t761 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X334 VPWR.t368 a_4329_5461# clknet_0_clk.t6 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X335 VGND.t711 a_6043_3677# a_6211_3579# VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X336 VPWR.t88 _16_.t7 a_5213_4664# VPWR.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.129 ps=1.18 w=0.42 l=0.15
X337 a_2398_3677# a_1959_3311# a_2313_3311# VGND.t811 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X338 a_2907_3677# a_2125_3311# a_2823_3677# VPWR.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X339 VPWR.t571 VGND.t861 VPWR.t570 VPWR.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X340 VGND.t423 clknet_0_clk.t37 a_1845_5461# VGND.t422 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X341 a_5814_4399# clknet_0_clk.t38 VPWR.t765 VPWR.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X342 VGND.t251 VPWR.t868 VGND.t250 VGND.t249 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X343 VGND.t228 a_7683_3579# a_7641_3311# VGND.t227 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X344 a_2524_3311# a_2125_3311# a_2398_3677# VGND.t541 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X345 VGND.t254 VPWR.t869 VGND.t253 VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X346 VGND.t256 VPWR.t870 VGND.t255 VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X347 VPWR.t15 clk.t3 a_4329_5461# VPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X348 a_2678_8029# a_2431_7663# VPWR.t714 VPWR.t713 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X349 a_7171_2767# _15_ VPWR.t299 VPWR.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X350 VPWR.t742 _10_ a_2695_6575# VPWR.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X351 VGND.t259 VPWR.t871 VGND.t258 VGND.t257 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X352 VGND.t35 a_2715_3829# a_2673_4233# VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X353 VGND.t149 VPWR.t872 VGND.t148 VGND.t147 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X354 VGND.t492 a_2566_3423# a_2524_3311# VGND.t491 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X355 VPWR.t568 VGND.t862 VPWR.t567 VPWR.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X356 VPWR.t565 VGND.t863 VPWR.t564 VPWR.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X357 VGND.t152 VPWR.t873 VGND.t151 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X358 VGND.t155 VPWR.t874 VGND.t154 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X359 clknet_0_clk.t5 a_4329_5461# VPWR.t366 VPWR.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X360 a_7258_3829# a_7090_3855# VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X361 a_1849_3861# a_1683_3861# VPWR.t285 VPWR.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X362 VGND.t619 a_5599_2741# _22_ VGND.t618 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X363 a_1845_5461# clknet_0_clk.t39 VGND.t225 VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X364 VPWR.t562 VGND.t864 VPWR.t561 VPWR.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X365 net6.t0 a_3267_4667# VPWR.t98 VPWR.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X366 _02_ _14_ a_1505_3855# VPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X367 clknet_1_1__leaf_clk.t22 a_5814_4399# VGND.t520 VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X368 a_2849_7663# a_2302_7937# a_2502_7637# VPWR.t180 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X369 VPWR.t559 VGND.t865 VPWR.t558 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X370 VPWR.t556 VGND.t866 VPWR.t555 VPWR.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X371 VPWR.t553 VGND.t867 VPWR.t552 VPWR.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X372 a_4495_5175# a_4779_5161# a_4714_5309# VGND.t750 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X373 VGND.t732 a_2502_7637# a_2431_7663# VGND.t699 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X374 a_2678_7119# a_2431_7497# VPWR.t394 VPWR.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X375 a_3145_6825# _12_ _01_ VPWR.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X376 VPWR.t708 net4 a_3215_2999# VPWR.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X377 VPWR.t68 _22_ a_7171_2767# VPWR.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X378 a_7515_3855# a_6651_3861# a_7258_3829# VPWR.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X379 VPWR.t550 VGND.t868 VPWR.t549 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X380 VGND.t158 VPWR.t875 VGND.t157 VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X381 a_2313_3311# _03_ VGND.t45 VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X382 VGND.t725 a_7258_3829# a_7216_4233# VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X383 _11_.t1 a_2695_6575# VPWR.t777 VPWR.t776 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X384 clknet_1_0__leaf_clk.t8 a_1845_5461# VPWR.t258 VPWR.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X385 net6.t1 a_3267_4667# VGND.t279 VGND.t278 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X386 clknet_1_1__leaf_clk.t11 a_5814_4399# VPWR.t220 VPWR.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X387 VPWR.t164 a_5505_2388# counter[5].t0 VPWR.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X388 a_7090_3677# a_6651_3311# a_7005_3311# VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X389 _24_ a_7077_2767# VPWR.t795 VPWR.t794 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X390 a_2125_8207# net2.t5 VPWR.t160 VPWR.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X391 a_7599_3677# a_6817_3311# a_7515_3677# VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X392 VPWR.t548 VGND.t869 VPWR.t547 VPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X393 a_2290_3829# a_2122_3855# VPWR.t826 VPWR.t825 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X394 VGND.t161 VPWR.t876 VGND.t160 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X395 VGND.t164 VPWR.t877 VGND.t163 VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X396 a_7216_3311# a_6817_3311# a_7090_3677# VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X397 a_2290_3829# a_2122_3855# VGND.t816 VGND.t815 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X398 VPWR.t239 a_7683_3829# a_7599_3855# VPWR.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X399 a_2849_7497# a_2302_7241# a_2502_7396# VPWR.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X400 clknet_0_clk.t4 a_4329_5461# VPWR.t364 VPWR.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X401 VGND.t386 net2.t6 a_1875_8207# VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X402 VPWR.t218 a_5814_4399# clknet_1_1__leaf_clk.t10 VPWR.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X403 VPWR.t763 clknet_0_clk.t40 a_5814_4399# VPWR.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X404 VPWR.t337 a_2547_3855# a_2715_3829# VPWR.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X405 VPWR.t546 VGND.t870 VPWR.t545 VPWR.t544 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X406 VPWR.t543 VGND.t871 VPWR.t542 VPWR.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X407 VGND.t718 a_7258_3423# a_7216_3311# VGND.t717 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X408 a_7515_3855# a_6817_3861# a_7258_3829# VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X409 VPWR.t541 VGND.t872 VPWR.t540 VPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X410 VPWR.t182 a_1825_2388# counter[1].t0 VPWR.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X411 VGND.t167 VPWR.t878 VGND.t166 VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X412 a_2295_7637# clknet_1_0__leaf_clk.t37 VPWR.t156 VPWR.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X413 VPWR.t362 a_4329_5461# clknet_0_clk.t12 VPWR.t361 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X414 a_4220_3829# net6.t6 a_4443_4175# VGND.t431 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X415 clknet_0_clk.t27 a_4329_5461# VGND.t685 VGND.t684 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X416 a_2589_4399# _04_ VPWR.t318 VPWR.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X417 VGND.t188 VPWR.t879 VGND.t187 VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X418 clknet_1_0__leaf_clk.t7 a_1845_5461# VPWR.t256 VPWR.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X419 VPWR.t538 VGND.t873 VPWR.t537 VPWR.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X420 a_2295_7337# clknet_1_0__leaf_clk.t38 VGND.t429 VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X421 a_5891_3133# net8 a_5795_3133# VGND.t808 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X422 a_6817_3311# a_6651_3311# VPWR.t2 VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X423 VGND.t799 _01_ a_2849_7497# VGND.t741 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X424 a_2674_4765# a_2235_4399# a_2589_4399# VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X425 VGND.t216 a_5843_3829# a_5801_4233# VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X426 VGND.t518 a_5814_4399# clknet_1_1__leaf_clk.t21 VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X427 VGND.t190 VPWR.t880 VGND.t189 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X428 clknet_1_0__leaf_clk.t24 a_1845_5461# VGND.t570 VGND.t569 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X429 VPWR.t536 VGND.t874 VPWR.t535 VPWR.t534 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X430 a_5345_3311# a_5179_3311# VGND.t213 VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X431 _16_.t1 a_3831_3339# VGND.t25 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X432 a_4977_3861# a_4811_3861# VPWR.t334 VPWR.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X433 a_2800_4399# a_2401_4399# a_2674_4765# VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X434 VGND.t683 a_4329_5461# clknet_0_clk.t26 VGND.t682 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X435 VPWR.t533 VGND.t875 VPWR.t532 VPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X436 VGND.t192 VPWR.t881 VGND.t191 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X437 a_2547_3855# a_1849_3861# a_2290_3829# VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X438 VGND.t767 _18_ a_4069_5309# VGND.t766 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X439 a_3099_4765# a_2401_4399# a_2842_4511# VGND.t424 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X440 VGND.t435 a_5505_2388# counter[5].t1 VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X441 VGND.t195 VPWR.t882 VGND.t194 VGND.t193 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X442 VGND.t197 VPWR.t883 VGND.t196 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X443 VPWR.t720 a_6427_2741# _23_ VPWR.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X444 VPWR.t530 VGND.t876 VPWR.t529 VPWR.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X445 VGND.t200 VPWR.t884 VGND.t199 VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X446 _21_ a_4259_3311# VGND.t210 VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X447 a_3215_3829# net6.t7 VGND.t433 VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X448 clknet_1_1__leaf_clk.t9 a_5814_4399# VPWR.t216 VPWR.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X449 a_2936_2767# _14_ a_2471_2741# VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X450 VGND.t468 clknet_1_0__leaf_clk.t39 a_1959_3311# VGND.t467 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X451 a_5436_4399# _22_ a_5213_4664# VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.1092 ps=1.36 w=0.42 l=0.15
X452 a_2651_7485# a_2431_7497# VGND.t698 VGND.t697 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X453 VPWR.t527 VGND.t877 VPWR.t526 VPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X454 a_1875_8207# net1 VGND.t760 VGND.t759 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X455 a_4287_4399# _17_ VGND.t615 VGND.t614 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X456 VPWR.t63 a_2295_7337# a_2302_7241# VPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X457 VGND.t749 a_4779_5161# a_4786_5065# VGND.t748 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X458 VPWR.t125 a_7619_5162# _08_ VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X459 VPWR.t524 VGND.t878 VPWR.t523 VPWR.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X460 net4 a_2715_3829# VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X461 VGND.t202 VPWR.t885 VGND.t201 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X462 VPWR.t360 a_4329_5461# clknet_0_clk.t11 VPWR.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X463 VGND.t128 VPWR.t886 VGND.t127 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X464 VPWR.t92 a_4986_5220# a_4915_5321# VPWR.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X465 VPWR.t787 a_5213_4664# a_5149_4721# VPWR.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.0672 ps=0.74 w=0.42 l=0.15
X466 net5 a_2991_3579# VPWR.t789 VPWR.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X467 VGND.t131 VPWR.t887 VGND.t130 VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X468 VGND.t134 VPWR.t888 VGND.t133 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X469 VGND.t137 VPWR.t889 VGND.t136 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X470 a_3831_3339# _11_.t10 VPWR.t326 VPWR.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X471 VGND.t635 _11_.t11 _01_ VGND.t634 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X472 VGND.t648 _23_ a_7723_2741# VGND.t647 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X473 a_5418_3829# a_5250_3855# VPWR.t78 VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X474 VPWR.t354 a_7345_2388# counter[7].t0 VPWR.t353 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X475 a_5418_3829# a_5250_3855# VGND.t265 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X476 VGND.t490 a_1825_2388# counter[1].t1 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X477 VGND.t610 _15_ a_3917_3339# VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X478 VPWR.t521 VGND.t879 VPWR.t520 VPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X479 clknet_0_clk.t10 a_4329_5461# VPWR.t358 VPWR.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X480 VPWR.t193 a_4767_3463# _20_ VPWR.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X481 VGND.t721 _21_ a_4520_4373# VGND.t720 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X482 a_1915_7815# a_2011_7637# VPWR.t189 VPWR.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X483 VGND.t140 VPWR.t890 VGND.t139 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X484 a_6425_2388# net8 VPWR.t816 VPWR.t815 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X485 VGND.t681 a_4329_5461# clknet_0_clk.t25 VGND.t680 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X486 VPWR.t254 a_1845_5461# clknet_1_0__leaf_clk.t6 VPWR.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X487 a_1845_5461# clknet_0_clk.t41 VGND.t628 VGND.t627 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X488 a_2313_3311# _03_ VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X489 _19_ a_3979_4943# VPWR.t793 VPWR.t792 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X490 VPWR.t518 VGND.t880 VPWR.t517 VPWR.t516 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X491 VGND.t498 a_3215_2999# _14_ VGND.t497 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X492 a_2566_3423# a_2398_3677# VGND.t502 VGND.t501 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X493 VPWR.t747 net1 a_2235_6575# VPWR.t746 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X494 a_4767_3463# net6.t8 VPWR.t162 VPWR.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X495 clknet_1_1__leaf_clk.t20 a_5814_4399# VGND.t516 VGND.t515 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X496 a_2122_3855# a_1683_3861# a_2037_3855# VGND.t598 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X497 VGND.t143 VPWR.t891 VGND.t142 VGND.t141 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X498 VGND.t146 VPWR.t892 VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X499 VGND.t568 a_1845_5461# clknet_1_0__leaf_clk.t23 VGND.t567 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X500 VGND.t390 VPWR.t893 VGND.t389 VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X501 VPWR.t33 _24_ a_7199_4943# VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X502 a_2248_4233# a_1849_3861# a_2122_3855# VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X503 VPWR.t515 VGND.t881 VPWR.t514 VPWR.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X504 a_4329_5461# clk.t4 VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X505 VPWR.t114 a_4399_5175# net7 VPWR.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X506 a_1849_3861# a_1683_3861# VGND.t597 VGND.t596 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X507 a_2769_4765# a_2235_4399# a_2674_4765# VPWR.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X508 VPWR.t512 VGND.t882 VPWR.t511 VPWR.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X509 a_2745_2388# net4 VPWR.t706 VPWR.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X510 a_1582_7439# net1 VGND.t758 VGND.t757 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X511 VPWR.t702 a_6043_3677# a_6211_3579# VPWR.t701 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X512 a_1915_7815# a_2011_7637# VGND.t500 VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X513 VGND.t645 a_2547_3855# a_2715_3829# VGND.t644 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X514 VPWR.t214 a_5814_4399# clknet_1_1__leaf_clk.t8 VPWR.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X515 VPWR.t509 VGND.t883 VPWR.t508 VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X516 a_1457_2388# net2.t7 VPWR.t134 VPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X517 a_7005_3855# _08_ VPWR.t144 VPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X518 VGND.t356 a_7619_5162# _08_ VGND.t355 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X519 a_4220_3829# net7 a_4349_3855# VPWR.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X520 a_2849_7663# a_2295_7637# a_2502_7637# VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X521 VGND.t393 VPWR.t894 VGND.t392 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X522 a_7641_3311# a_6651_3311# a_7515_3677# VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X523 VGND.t679 a_4329_5461# clknet_0_clk.t24 VGND.t678 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X524 a_4341_3311# _11_.t12 a_4259_3311# VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X525 a_5675_3855# a_4977_3861# a_5418_3829# VGND.t630 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X526 VPWR.t704 net4 a_2041_4649# VPWR.t703 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X527 VPWR.t84 _11_.t13 a_7171_2767# VPWR.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X528 a_6817_3861# a_6651_3861# VPWR.t185 VPWR.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X529 VPWR.t506 VGND.t884 VPWR.t505 VPWR.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X530 VGND.t396 VPWR.t895 VGND.t395 VGND.t394 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X531 a_5599_2741# net6.t9 a_5997_3133# VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X532 VGND.t661 a_7345_2388# counter[7].t1 VGND.t660 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X533 VPWR.t504 VGND.t885 VPWR.t503 VPWR.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X534 VGND.t399 VPWR.t896 VGND.t398 VGND.t397 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X535 VPWR.t19 a_1915_7815# net2.t0 VPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X536 VGND.t566 a_1845_5461# clknet_1_0__leaf_clk.t22 VGND.t565 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X537 a_7258_3423# a_7090_3677# VGND.t763 VGND.t762 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X538 VPWR.t102 net11 a_7753_2767# VPWR.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X539 clknet_0_clk.t23 a_4329_5461# VGND.t677 VGND.t676 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X540 VGND.t402 VPWR.t897 VGND.t401 VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X541 VGND.t470 clknet_1_0__leaf_clk.t40 a_2235_4399# VGND.t469 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X542 a_4995_4399# net9 VGND.t736 VGND.t735 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X543 VPWR.t501 VGND.t886 VPWR.t500 VPWR.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X544 a_6425_2388# net8 VGND.t807 VGND.t806 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X545 VPWR.t347 net7 a_4767_3463# VPWR.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X546 a_2398_3677# a_2125_3311# a_2313_3311# VPWR.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X547 a_2502_7637# a_2295_7637# a_2678_8029# VPWR.t784 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X548 VPWR.t498 VGND.t887 VPWR.t497 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X549 clknet_1_0__leaf_clk.t21 a_1845_5461# VGND.t564 VGND.t563 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X550 a_4069_5309# a_3799_4943# a_3979_4943# VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X551 VPWR.t495 VGND.t888 VPWR.t494 VPWR.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X552 VGND.t405 VPWR.t898 VGND.t404 VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X553 a_2840_3087# a_2614_2883# a_2471_2741# VGND.t626 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X554 a_7258_3829# a_7090_3855# VPWR.t54 VPWR.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X555 a_5759_3855# a_4977_3861# a_5675_3855# VPWR.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X556 VPWR.t212 a_5814_4399# clknet_1_1__leaf_clk.t7 VPWR.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X557 VPWR.t492 VGND.t889 VPWR.t491 VPWR.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X558 VPWR.t297 _15_ a_6375_5309# VPWR.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X559 VGND.t408 VPWR.t899 VGND.t407 VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X560 VGND.t447 VPWR.t900 VGND.t446 VGND.t394 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X561 a_2849_7497# a_2295_7337# a_2502_7396# VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X562 VPWR.t252 a_1845_5461# clknet_1_0__leaf_clk.t5 VPWR.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X563 _15_ a_3831_3105# VPWR.t312 VPWR.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X564 VGND.t783 a_2991_3579# a_2949_3311# VGND.t782 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X565 VPWR.t184 a_2566_3423# a_2493_3677# VPWR.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X566 a_4349_4175# _15_ VGND.t609 VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X567 a_8265_2388# net10 VPWR.t276 VPWR.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X568 a_2230_7663# a_1915_7815# VGND.t41 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X569 VPWR.t740 a_7515_3855# a_7683_3829# VPWR.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X570 VGND.t39 a_1915_7815# net2.t1 VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X571 a_5250_3855# a_4811_3861# a_5165_3855# VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X572 VGND.t450 VPWR.t901 VGND.t449 VGND.t448 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X573 VGND.t453 VPWR.t902 VGND.t452 VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X574 a_2745_2388# net4 VGND.t713 VGND.t712 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X575 a_2842_4511# a_2674_4765# VGND.t420 VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X576 a_2493_3677# a_1959_3311# a_2398_3677# VPWR.t823 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X577 a_2502_7396# a_2295_7337# a_2678_7119# VPWR.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X578 a_2011_7637# a_2302_7937# a_2253_8029# VPWR.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X579 a_1457_2388# net2.t8 VGND.t388 VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X580 a_5376_4233# a_4977_3861# a_5250_3855# VGND.t629 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X581 clknet_1_1__leaf_clk.t6 a_5814_4399# VPWR.t210 VPWR.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X582 a_4977_3861# a_4811_3861# VGND.t641 VGND.t640 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X583 VPWR.t489 VGND.t890 VPWR.t488 VPWR.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X584 VPWR.t486 VGND.t891 VPWR.t485 VPWR.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X585 VPWR.t797 net2.t9 a_2235_6575# VPWR.t796 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X586 clknet_0_clk.t22 a_4329_5461# VGND.t675 VGND.t674 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X587 a_7941_3087# _23_ _09_ VGND.t646 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X588 a_2011_7637# a_2295_7637# a_2230_7663# VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X589 a_3245_3855# _16_.t8 VPWR.t90 VPWR.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X590 VPWR.t483 VGND.t892 VPWR.t482 VPWR.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X591 VPWR.t761 clknet_0_clk.t42 a_5814_4399# VPWR.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X592 VPWR.t759 clknet_0_clk.t43 a_1845_5461# VPWR.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X593 a_4585_2388# net6.t10 VPWR.t27 VPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X594 VGND.t291 a_7515_3677# a_7683_3579# VGND.t290 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X595 net9 a_6211_3579# VGND.t777 VGND.t776 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X596 VGND.t456 VPWR.t903 VGND.t455 VGND.t454 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X597 VPWR.t480 VGND.t893 VPWR.t479 VPWR.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X598 VGND.t673 a_4329_5461# clknet_0_clk.t21 VGND.t672 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X599 a_5795_3133# net9 VGND.t734 VGND.t733 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X600 VGND.t458 VPWR.t904 VGND.t457 VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X601 a_2011_7351# a_2302_7241# a_2253_7119# VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X602 a_5997_3133# net7 a_5891_3133# VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X603 VGND.t461 VPWR.t905 VGND.t460 VGND.t459 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X604 VGND.t652 a_1875_8207# _00_ VGND.t651 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X605 a_6623_3133# _22_ VGND.t236 VGND.t235 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X606 clknet_1_0__leaf_clk.t4 a_1845_5461# VPWR.t250 VPWR.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X607 a_7753_2767# a_7723_2741# _09_ VPWR.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X608 a_6825_3133# _11_.t14 a_6719_3133# VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X609 VGND.t464 VPWR.t906 VGND.t463 VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X610 VGND.t108 VPWR.t907 VGND.t107 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X611 VPWR.t712 a_7258_3423# a_7185_3677# VPWR.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X612 a_2561_9514# enable.t0 VPWR.t168 VPWR.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X613 clknet_1_0__leaf_clk.t3 a_1845_5461# VPWR.t248 VPWR.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X614 VGND.t562 a_1845_5461# clknet_1_0__leaf_clk.t20 VGND.t561 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X615 VGND.t473 net3.t7 _12_ VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X616 VGND.t544 net5 a_3917_3105# VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X617 VGND.t605 a_2823_3677# a_2991_3579# VGND.t604 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X618 _02_ _13_ VGND.t354 VGND.t353 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X619 clknet_1_1__leaf_clk.t5 a_5814_4399# VPWR.t208 VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X620 VPWR.t477 VGND.t894 VPWR.t476 VPWR.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X621 VPWR.t474 VGND.t895 VPWR.t473 VPWR.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X622 VGND.t591 a_2471_2741# _03_ VGND.t590 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X623 a_7185_3677# a_6651_3311# a_7090_3677# VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X624 a_2037_3855# _02_ VPWR.t730 VPWR.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X625 a_4329_5461# clk.t5 VGND.t364 VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X626 a_3389_3105# _11_.t15 VGND.t358 VGND.t357 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X627 VPWR.t471 VGND.t896 VPWR.t470 VPWR.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X628 a_7077_2767# net10 VGND.t588 VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X629 a_8265_2388# net10 VGND.t586 VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X630 VGND.t756 net1 a_2389_6575# VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X631 VPWR.t468 VGND.t897 VPWR.t467 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X632 _13_ _11_.t16 VGND.t360 VGND.t359 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X633 VGND.t295 a_4399_5175# net7 VGND.t294 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X634 a_2011_7351# a_2295_7337# a_2230_7485# VGND.t233 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X635 VPWR.t206 a_5814_4399# clknet_1_1__leaf_clk.t4 VPWR.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X636 VPWR.t732 _00_ a_2849_7663# VPWR.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X637 VGND.t111 VPWR.t908 VGND.t110 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X638 VPWR.t310 a_5599_2741# _22_ VPWR.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X639 a_7599_3855# a_6817_3861# a_7515_3855# VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X640 VPWR.t466 VGND.t898 VPWR.t465 VPWR.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X641 VPWR.t775 a_2695_6575# _11_.t0 VPWR.t774 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X642 VGND.t113 VPWR.t909 VGND.t112 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X643 a_5618_3677# a_5179_3311# a_5533_3311# VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X644 VPWR.t463 VGND.t899 VPWR.t462 VPWR.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X645 a_2125_3311# a_1959_3311# VPWR.t822 VPWR.t821 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X646 VPWR.t745 net1 a_2125_8207# VPWR.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X647 counter[9].t0 a_7939_2223# VPWR.t694 VPWR.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X648 VPWR.t460 VGND.t900 VPWR.t459 VPWR.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X649 clknet_0_clk.t20 a_4329_5461# VGND.t671 VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X650 VPWR.t274 net10 a_6427_2741# VPWR.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X651 VGND.t116 VPWR.t910 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X652 VPWR.t52 a_4520_4373# a_4454_4649# VPWR.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X653 VPWR.t457 VGND.t901 VPWR.t456 VPWR.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X654 a_7090_3855# a_6651_3861# a_7005_3855# VGND.t496 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X655 a_6043_3677# a_5179_3311# a_5786_3423# VPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X656 VGND.t119 VPWR.t911 VGND.t118 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X657 a_4585_2388# net6.t11 VGND.t50 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X658 a_5744_3311# a_5345_3311# a_5618_3677# VGND.t745 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X659 VGND.t560 a_1845_5461# clknet_1_0__leaf_clk.t19 VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X660 VGND.t122 VPWR.t912 VGND.t121 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X661 VPWR.t454 VGND.t902 VPWR.t453 VPWR.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X662 VGND.t514 a_5814_4399# clknet_1_1__leaf_clk.t19 VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X663 VPWR.t808 _01_ a_2849_7497# VPWR.t807 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X664 a_5871_5162# _19_ VPWR.t803 VPWR.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X665 a_7216_4233# a_6817_3861# a_7090_3855# VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X666 clknet_0_clk.t19 a_4329_5461# VGND.t669 VGND.t668 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X667 VPWR.t451 VGND.t903 VPWR.t450 VPWR.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X668 VPWR.t448 VGND.t904 VPWR.t447 VPWR.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X669 VPWR.t445 VGND.t905 VPWR.t444 VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X670 VPWR.t442 VGND.t906 VPWR.t441 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X671 VGND.t27 a_5786_3423# a_5744_3311# VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X672 a_6817_3861# a_6651_3861# VGND.t495 VGND.t494 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X673 VPWR.t439 VGND.t907 VPWR.t438 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X674 VGND.t125 VPWR.t913 VGND.t124 VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X675 VGND.t169 VPWR.t914 VGND.t168 VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X676 VPWR.t246 a_1845_5461# clknet_1_0__leaf_clk.t2 VPWR.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X677 VPWR.t436 VGND.t908 VPWR.t435 VPWR.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X678 VPWR.t433 VGND.t909 VPWR.t432 VPWR.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X679 VPWR.t781 a_6211_3579# a_6127_3677# VPWR.t780 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X680 VGND.t752 a_7515_3855# a_7683_3829# VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X681 clknet_1_0__leaf_clk.t18 a_1845_5461# VGND.t558 VGND.t557 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X682 clknet_1_1__leaf_clk.t18 a_5814_4399# VGND.t512 VGND.t511 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X683 a_2561_9514# enable.t1 VGND.t475 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X684 VGND.t172 VPWR.t915 VGND.t171 VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X685 VPWR.t244 a_1845_5461# clknet_1_0__leaf_clk.t1 VPWR.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X686 a_2295_7637# clknet_1_0__leaf_clk.t41 VGND.t636 VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X687 VPWR.t204 a_5814_4399# clknet_1_1__leaf_clk.t3 VPWR.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X688 a_2631_3855# a_1849_3861# a_2547_3855# VPWR.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X689 a_5814_4399# clknet_0_clk.t44 VGND.t485 VGND.t484 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X690 VGND.t742 _00_ a_2849_7663# VGND.t741 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X691 VPWR.t430 VGND.t910 VPWR.t429 VPWR.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X692 a_2674_4765# a_2401_4399# a_2589_4399# VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X693 VPWR.t427 VGND.t911 VPWR.t426 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X694 VGND.t174 VPWR.t916 VGND.t173 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X695 a_2566_3423# a_2398_3677# VPWR.t191 VPWR.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X696 VGND.t176 VPWR.t917 VGND.t175 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X697 VGND.t366 clk.t6 a_4329_5461# VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X698 VPWR.t127 _11_.t17 a_3145_6825# VPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X699 a_5533_3311# _07_ VGND.t771 VGND.t770 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X700 VPWR.t424 VGND.t912 VPWR.t423 VPWR.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X701 VGND.t179 VPWR.t918 VGND.t178 VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X702 VPWR.t281 a_3099_4765# a_3267_4667# VPWR.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X703 VPWR.t236 net5 a_3831_3105# VPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X704 a_6817_3311# a_6651_3311# VGND.t21 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X705 a_4349_3855# net6.t12 VPWR.t328 VPWR.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X706 a_4495_5175# a_4786_5065# a_4737_4943# VPWR.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X707 VPWR.t421 VGND.t913 VPWR.t420 VPWR.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X708 VPWR.t129 clknet_1_1__leaf_clk.t39 a_5179_3311# VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X709 clknet_1_1__leaf_clk.t2 a_5814_4399# VPWR.t202 VPWR.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X710 a_5165_3855# _06_ VPWR.t174 VPWR.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X711 a_6375_5309# _11_.t18 VPWR.t691 VPWR.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X712 a_3215_2999# _11_.t19 VPWR.t693 VPWR.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X713 VGND.t182 VPWR.t919 VGND.t181 VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X714 VGND.t185 VPWR.t920 VGND.t184 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X715 VPWR.t17 a_2842_4511# a_2769_4765# VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X716 a_4767_3463# net6.t13 a_5001_3311# VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X717 VGND.t87 VPWR.t921 VGND.t86 VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X718 a_2651_7663# a_2431_7663# VGND.t719 VGND.t697 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X719 VGND.t273 a_4986_5220# a_4915_5321# VGND.t272 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X720 VPWR.t345 net7 a_6375_5309# VPWR.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X721 VGND.t593 a_3099_4765# a_3267_4667# VGND.t592 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X722 VGND.t504 a_4767_3463# _20_ VGND.t503 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X723 _07_ a_5149_4721# VGND.t479 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.098625 ps=0.98 w=0.65 l=0.15
X724 _06_ a_4454_4649# VPWR.t291 VPWR.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.18575 ps=1.415 w=1 l=0.15
X725 counter[9].t1 a_7939_2223# VGND.t703 VGND.t702 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X726 VGND.t466 _16_.t9 a_3215_3829# VGND.t465 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X727 VPWR.t757 clknet_0_clk.t45 a_1845_5461# VPWR.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X728 VGND.t90 VPWR.t922 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X729 a_2502_7637# a_2302_7937# a_2651_7663# VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X730 VGND.t667 a_4329_5461# clknet_0_clk.t18 VGND.t666 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X731 _25_ a_7199_4943# VGND.t707 VGND.t706 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X732 a_4382_4649# net8 VPWR.t814 VPWR.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X733 _10_ a_2235_6575# VGND.t47 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X734 VGND.t93 VPWR.t923 VGND.t92 VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X735 VPWR.t799 net2.t10 a_1957_8207# VPWR.t798 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X736 VGND.t96 VPWR.t924 VGND.t95 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X737 a_5871_5162# _19_ VGND.t794 VGND.t793 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X738 clknet_1_0__leaf_clk.t17 a_1845_5461# VGND.t556 VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X739 VGND.t99 VPWR.t925 VGND.t98 VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X740 a_3601_3855# net6.t14 VPWR.t330 VPWR.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X741 a_6545_5309# net7 a_6457_5309# VGND.t653 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X742 VGND.t607 _15_ a_6651_5309# VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X743 a_4986_5220# a_4779_5161# a_5162_4943# VPWR.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X744 a_1845_5461# clknet_0_clk.t46 VPWR.t755 VPWR.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X745 VPWR.t783 a_2295_7637# a_2302_7937# VPWR.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X746 VPWR.t418 VGND.t914 VPWR.t417 VPWR.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X747 a_5162_4943# a_4915_5321# VPWR.t289 VPWR.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X748 VGND.t510 a_5814_4399# clknet_1_1__leaf_clk.t17 VGND.t509 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X749 clknet_1_1__leaf_clk.t1 a_5814_4399# VPWR.t200 VPWR.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X750 a_7723_2741# _23_ a_8109_2767# VPWR.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X751 VGND.t102 VPWR.t926 VGND.t101 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X752 VGND.t105 VPWR.t927 VGND.t104 VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X753 VGND.t369 VPWR.t928 VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X754 a_3183_4765# a_2401_4399# a_3099_4765# VPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X755 VPWR.t415 VGND.t915 VPWR.t414 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X756 VGND.t232 a_2295_7337# a_2302_7241# VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X757 VPWR.t412 VGND.t916 VPWR.t411 VPWR.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X758 a_4915_5321# a_4786_5065# a_4495_5175# VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X759 VPWR.t154 a_5675_3855# a_5843_3829# VPWR.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X760 VPWR.t409 VGND.t917 VPWR.t408 VPWR.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X761 VGND.t665 a_4329_5461# clknet_0_clk.t17 VGND.t664 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X762 VGND.t372 VPWR.t929 VGND.t371 VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X763 _12_ net2.t11 a_1582_7439# VGND.t790 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X764 a_2502_7396# a_2302_7241# a_2651_7485# VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X765 VPWR.t406 VGND.t918 VPWR.t405 VPWR.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X766 VGND.t437 a_4220_3829# _18_ VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X767 a_5333_5321# a_4786_5065# a_4986_5220# VPWR.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X768 VPWR.t130 clknet_1_1__leaf_clk.t40 a_6651_3311# VPWR.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X769 a_5814_4399# clknet_0_clk.t47 VGND.t204 VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X770 VPWR.t187 a_3215_2999# _14_ VPWR.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X771 VPWR.t234 net5 a_2936_2767# VPWR.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X772 VGND.t375 VPWR.t930 VGND.t374 VGND.t373 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X773 VPWR.t403 VGND.t919 VPWR.t402 VPWR.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X774 a_4986_5220# a_4786_5065# a_5135_5309# VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X775 VPWR.t400 VGND.t920 VPWR.t399 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X776 VGND.t632 clk.t7 a_4329_5461# VGND.t631 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X777 a_5213_4664# _22_ VPWR.t66 VPWR.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.20925 ps=1.345 w=0.42 l=0.15
X778 VPWR.t279 a_2471_2741# _03_ VPWR.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
X779 a_4259_3311# _15_ VPWR.t295 VPWR.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X780 a_2431_7663# a_2302_7937# a_2011_7637# VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X781 VGND.t754 _10_ a_2695_6575# VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X782 a_1957_8207# net1 a_1875_8207# VPWR.t743 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X783 VPWR.t112 a_7515_3677# a_7683_3579# VPWR.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X784 a_5333_5321# a_4779_5161# a_4986_5220# VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X785 VPWR.t388 a_3849_2388# counter[3].t0 VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X786 VPWR.t397 VGND.t921 VPWR.t396 VPWR.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X787 net9 a_6211_3579# VPWR.t779 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X788 VGND.t223 net6.t15 a_3433_4175# VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X789 a_4779_5161# clknet_1_1__leaf_clk.t41 VPWR.t828 VPWR.t827 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X790 clknet_0_clk.t16 a_4329_5461# VGND.t663 VGND.t662 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X791 a_2842_4511# a_2674_4765# VPWR.t146 VPWR.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X792 VPWR.t810 a_5418_3829# a_5345_3855# VPWR.t809 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X793 VPWR.t771 _18_ a_3979_4943# VPWR.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X794 a_2401_4399# a_2235_4399# VPWR.t74 VPWR.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X795 a_7641_4233# a_6651_3861# a_7515_3855# VGND.t493 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X796 a_5345_3855# a_4811_3861# a_5250_3855# VPWR.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X797 clknet_0_clk.t9 a_4329_5461# VPWR.t356 VPWR.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X798 a_7723_2741# net11 VGND.t283 VGND.t282 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X799 a_5533_3311# _07_ VPWR.t773 VPWR.t772 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X800 VPWR.t293 a_2823_3677# a_2991_3579# VPWR.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X801 a_4443_4175# _11_.t20 a_4349_4175# VGND.t701 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X802 VGND.t378 VPWR.t931 VGND.t377 VGND.t376 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X803 VGND.t381 VPWR.t932 VGND.t380 VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X804 a_4929_3311# net8 VGND.t805 VGND.t804 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X805 _01_ _12_ VGND.t744 VGND.t743 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X806 a_7090_3677# a_6817_3311# a_7005_3311# VPWR.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X807 VGND.t384 VPWR.t933 VGND.t383 VGND.t382 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X808 a_3917_3339# _11_.t21 a_3831_3339# VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X809 _11_.t2 a_2695_6575# VGND.t773 VGND.t772 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X810 clknet_1_0__leaf_clk.t16 a_1845_5461# VGND.t554 VGND.t553 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X811 clknet_1_0__leaf_clk.t0 a_1845_5461# VPWR.t242 VPWR.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X812 clknet_1_1__leaf_clk.t16 a_5814_4399# VGND.t508 VGND.t507 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X813 a_5149_4721# a_5213_4664# a_4995_4399# VGND.t781 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X814 VPWR.t198 a_5814_4399# clknet_1_1__leaf_clk.t0 VPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X815 a_4714_5309# a_4399_5175# VGND.t293 VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 VGND.n1259 VGND 8722.05
R1 VGND.n1025 VGND 8664.24
R2 VGND VGND.n1097 8611.64
R3 VGND.n1090 VGND 8561.42
R4 VGND.n1263 VGND.n1025 7881.01
R5 VGND.n1093 VGND.n1091 7881.01
R6 VGND.n1091 VGND.n1090 7881.01
R7 VGND.n1262 VGND.n1261 7881.01
R8 VGND.n1263 VGND.n1262 7881.01
R9 VGND.n1096 VGND.n1094 7881.01
R10 VGND.n1094 VGND.n1093 7881.01
R11 VGND.n1260 VGND.n1259 7881.01
R12 VGND.n1261 VGND.n1260 7881.01
R13 VGND.n1097 VGND.n1096 7881.01
R14 VGND.t394 VGND 4888.89
R15 VGND VGND.t394 4408.43
R16 VGND.t441 VGND.t335 3877.39
R17 VGND.t12 VGND.t243 3877.39
R18 VGND VGND.t3 3346.36
R19 VGND VGND.t462 3346.36
R20 VGND VGND.t350 3346.36
R21 VGND VGND.t82 3346.36
R22 VGND VGND.t144 3346.36
R23 VGND VGND.t0 3346.36
R24 VGND VGND.t403 3346.36
R25 VGND.t150 VGND.t454 3101.92
R26 VGND.t252 VGND.t326 3101.92
R27 VGND.t448 VGND.t79 3101.92
R28 VGND.t367 VGND 2857.47
R29 VGND.t329 VGND 2857.47
R30 VGND VGND.t61 2857.47
R31 VGND VGND.t400 2857.47
R32 VGND.t317 VGND 2857.47
R33 VGND.t73 VGND 2857.47
R34 VGND.t370 VGND.t575 2495.02
R35 VGND VGND.n196 2469.73
R36 VGND.t6 VGND 2452.87
R37 VGND VGND.t180 2452.87
R38 VGND.t153 VGND.t70 2326.44
R39 VGND.t156 VGND.t126 2326.44
R40 VGND.t451 VGND.t117 2326.44
R41 VGND.n1025 VGND 2183.14
R42 VGND VGND.n1263 2183.14
R43 VGND.n1262 VGND 2183.14
R44 VGND.n1261 VGND 2183.14
R45 VGND.n1260 VGND 2183.14
R46 VGND.n1259 VGND 2183.14
R47 VGND.t621 VGND.t332 2097.71
R48 VGND VGND.t257 2081.99
R49 VGND.t162 VGND 2081.99
R50 VGND.t249 VGND.n1095 1938.7
R51 VGND.n1090 VGND 1896.55
R52 VGND.n1091 VGND 1896.55
R53 VGND.n1093 VGND 1896.55
R54 VGND.n1094 VGND 1896.55
R55 VGND.n1096 VGND 1896.55
R56 VGND.n1097 VGND 1896.55
R57 VGND VGND.t376 1886.64
R58 VGND.t132 VGND 1886.64
R59 VGND.t103 VGND 1886.64
R60 VGND VGND.t162 1812.26
R61 VGND.t240 VGND 1795.4
R62 VGND VGND.t150 1795.4
R63 VGND VGND.t252 1795.4
R64 VGND VGND.t448 1795.4
R65 VGND VGND.t114 1786.97
R66 VGND.t159 VGND 1786.97
R67 VGND.t459 VGND 1786.97
R68 VGND.t94 VGND 1702.68
R69 VGND.t376 VGND 1698.3
R70 VGND VGND.t132 1698.3
R71 VGND VGND.t103 1698.3
R72 VGND.t332 VGND 1698.3
R73 VGND VGND.n434 1677.39
R74 VGND.t782 VGND.t604 1593.1
R75 VGND.t549 VGND.t751 1593.1
R76 VGND.t499 VGND.t40 1593.1
R77 VGND.t355 VGND.t706 1584.67
R78 VGND.t741 VGND.t231 1584.67
R79 VGND.t141 VGND.t209 1567.82
R80 VGND.t3 VGND.t391 1550.96
R81 VGND.t462 VGND.t367 1550.96
R82 VGND.t350 VGND.t329 1550.96
R83 VGND.t61 VGND.t159 1550.96
R84 VGND.t82 VGND.t100 1550.96
R85 VGND.t144 VGND.t323 1550.96
R86 VGND.t0 VGND.t317 1550.96
R87 VGND.t403 VGND.t73 1550.96
R88 VGND.t761 VGND.t651 1550.96
R89 VGND.t290 VGND.t797 1416.09
R90 VGND VGND.t24 1407.66
R91 VGND.t106 VGND 1407.66
R92 VGND.t67 VGND 1407.66
R93 VGND.t76 VGND 1407.66
R94 VGND.t138 VGND 1407.66
R95 VGND.t302 VGND 1407.66
R96 VGND.t594 VGND.t606 1399.23
R97 VGND.t85 VGND 1399.23
R98 VGND VGND.t38 1390.8
R99 VGND VGND.t147 1306.51
R100 VGND.t114 VGND 1306.51
R101 VGND VGND.t370 1306.51
R102 VGND.t391 VGND 1306.51
R103 VGND.t454 VGND 1306.51
R104 VGND.t135 VGND 1306.51
R105 VGND VGND.t305 1306.51
R106 VGND.t100 VGND 1306.51
R107 VGND.t326 VGND 1306.51
R108 VGND VGND.t249 1306.51
R109 VGND VGND.t165 1306.51
R110 VGND.t323 VGND 1306.51
R111 VGND.t79 VGND 1306.51
R112 VGND.t170 VGND 1306.51
R113 VGND VGND.t459 1306.51
R114 VGND VGND.t129 1295.65
R115 VGND.n2474 VGND.n64 1294.86
R116 VGND VGND.t91 1289.15
R117 VGND.t770 VGND 1272.8
R118 VGND.t9 VGND.n821 1251.96
R119 VGND.n1110 VGND.n1098 1198.25
R120 VGND.n1092 VGND.n485 1198.25
R121 VGND.n1611 VGND.n697 1198.25
R122 VGND.n1513 VGND.n821 1198.25
R123 VGND.n1441 VGND.n847 1198.25
R124 VGND.n1258 VGND.n1257 1198.25
R125 VGND.n1095 VGND.n161 1196.22
R126 VGND.n2201 VGND.n196 1196.22
R127 VGND.n2439 VGND.n78 1194.5
R128 VGND.n2375 VGND.n117 1194.5
R129 VGND.n1973 VGND.n337 1194.5
R130 VGND.n2038 VGND.n300 1194.5
R131 VGND.n1875 VGND.n434 1194.5
R132 VGND.n1713 VGND.n617 1194.5
R133 VGND.n1294 VGND.n1264 1194.5
R134 VGND.n1024 VGND.n1023 1194.5
R135 VGND.t720 VGND.t658 1188.51
R136 VGND.t710 VGND.n1024 1146.36
R137 VGND.t651 VGND 1137.93
R138 VGND.t551 VGND 1104.21
R139 VGND.t91 VGND 1100.81
R140 VGND.t129 VGND 1100.81
R141 VGND.t804 VGND.t503 1078.93
R142 VGND.t209 VGND.t704 1078.93
R143 VGND.t596 VGND 1078.93
R144 VGND.t634 VGND 1070.5
R145 VGND VGND.t594 1036.78
R146 VGND.t46 VGND 1036.78
R147 VGND VGND.t9 1025.15
R148 VGND.t305 VGND 1019.92
R149 VGND.t400 VGND 1019.92
R150 VGND.t335 VGND 1019.92
R151 VGND.t243 VGND 1019.92
R152 VGND.t491 VGND.t501 1003.07
R153 VGND VGND.t649 1003.07
R154 VGND.t699 VGND.t697 1003.07
R155 VGND.n2330 VGND.n2329 999.607
R156 VGND.n2156 VGND.n2155 999.607
R157 VGND.n1928 VGND.n1927 999.607
R158 VGND.n847 VGND.t406 973.746
R159 VGND.t786 VGND.t670 960.92
R160 VGND.t280 VGND.t271 952.49
R161 VGND.t23 VGND.t728 944.062
R162 VGND.t44 VGND.t811 944.062
R163 VGND.t234 VGND.t741 944.062
R164 VGND.n337 VGND 927.203
R165 VGND.n117 VGND 927.203
R166 VGND VGND.t382 919.313
R167 VGND VGND.t308 919.313
R168 VGND.t120 VGND 919.313
R169 VGND VGND.t177 918.774
R170 VGND VGND.t106 918.774
R171 VGND VGND.t67 918.774
R172 VGND VGND.t76 918.774
R173 VGND.t70 VGND 918.774
R174 VGND VGND.n300 918.774
R175 VGND VGND.t138 918.774
R176 VGND.t126 VGND 918.774
R177 VGND VGND.t85 918.774
R178 VGND.t117 VGND 918.774
R179 VGND VGND.n78 918.774
R180 VGND VGND.t302 918.774
R181 VGND.t24 VGND.t543 910.346
R182 VGND VGND.n697 901.917
R183 VGND VGND.n1092 901.917
R184 VGND.t379 VGND.t341 896.236
R185 VGND.t424 VGND.t263 893.487
R186 VGND.t233 VGND.t487 893.487
R187 VGND.n1807 VGND.n1806 870.4
R188 VGND.t486 VGND 851.341
R189 VGND.t815 VGND.t412 851.341
R190 VGND.t487 VGND.t699 851.341
R191 VGND.t722 VGND.t640 842.913
R192 VGND.t745 VGND.t211 834.484
R193 VGND.t629 VGND.t642 834.484
R194 VGND.t608 VGND.t436 834.484
R195 VGND.t425 VGND.t36 834.484
R196 VGND.t598 VGND.t411 834.484
R197 VGND.t488 VGND.t234 834.484
R198 VGND.t697 VGND.t488 834.484
R199 VGND.t501 VGND.t626 826.054
R200 VGND.t706 VGND.t55 826.054
R201 VGND.t123 VGND.t226 826.054
R202 VGND.t618 VGND.t770 809.196
R203 VGND.t606 VGND.t633 809.196
R204 VGND.t227 VGND.t22 800.766
R205 VGND.t493 VGND.t549 800.766
R206 VGND.t753 VGND.t772 800.766
R207 VGND.t40 VGND.t233 800.766
R208 VGND.t64 VGND.t653 792.337
R209 VGND.t774 VGND.t15 792.337
R210 VGND.t542 VGND.t28 783.909
R211 VGND.t257 VGND.t240 775.48
R212 VGND.t541 VGND.t59 758.621
R213 VGND.t616 VGND.t123 758.621
R214 VGND.t757 VGND.t790 750.192
R215 VGND.t382 VGND 746.942
R216 VGND.t406 VGND 746.942
R217 VGND.t308 VGND 746.942
R218 VGND VGND.t120 746.942
R219 VGND.t589 VGND.t268 741.763
R220 VGND.t513 VGND.t769 741.763
R221 VGND.t795 VGND.t355 741.763
R222 VGND.t653 VGND.t266 741.763
R223 VGND.t235 VGND.t776 724.904
R224 VGND.t515 VGND.t537 724.904
R225 VGND.t519 VGND.t517 724.904
R226 VGND.t521 VGND.t531 724.904
R227 VGND.t730 VGND.t484 724.904
R228 VGND.t484 VGND.t476 724.904
R229 VGND.t363 VGND.t365 724.904
R230 VGND.t678 VGND.t674 724.904
R231 VGND.t684 VGND.t680 724.904
R232 VGND.t690 VGND.t686 724.904
R233 VGND.t662 VGND.t690 724.904
R234 VGND.t627 VGND.t422 724.904
R235 VGND.t42 VGND.t627 724.904
R236 VGND.t224 VGND.t42 724.904
R237 VGND.t573 VGND.t224 724.904
R238 VGND.t577 VGND.t573 724.904
R239 VGND.t583 VGND.t581 724.904
R240 VGND.t579 VGND.t583 724.904
R241 VGND.t555 VGND.t579 724.904
R242 VGND.t559 VGND.t555 724.904
R243 VGND.t553 VGND.t559 724.904
R244 VGND.t557 VGND.t565 724.904
R245 VGND.t561 VGND.t557 724.904
R246 VGND.t563 VGND.t561 724.904
R247 VGND.t567 VGND.t563 724.904
R248 VGND.t569 VGND.t567 724.904
R249 VGND.t571 VGND.t569 724.904
R250 VGND.t790 VGND.t472 724.904
R251 VGND.t525 VGND.t183 716.476
R252 VGND.t658 VGND.t219 716.476
R253 VGND.t431 VGND.t614 716.476
R254 VGND.t631 VGND.t802 716.476
R255 VGND.t282 VGND.t284 708.047
R256 VGND.t20 VGND.t298 708.047
R257 VGND.t212 VGND.t276 708.047
R258 VGND.t543 VGND.t486 708.047
R259 VGND.t467 VGND.t813 708.047
R260 VGND.t735 VGND.t722 708.047
R261 VGND.t432 VGND.t465 708.047
R262 VGND.t624 VGND.t599 708.047
R263 VGND.t359 VGND.t715 708.047
R264 VGND.t539 VGND.t596 708.047
R265 VGND.t353 VGND.t30 708.047
R266 VGND.t743 VGND.t634 708.047
R267 VGND.t772 VGND.t774 708.047
R268 VGND.t231 VGND.t428 708.047
R269 VGND.t38 VGND.t499 708.047
R270 VGND.t413 VGND.t761 708.047
R271 VGND.t385 VGND.t413 708.047
R272 VGND.t759 VGND.t385 708.047
R273 VGND.t186 VGND.t409 701.582
R274 VGND.t600 VGND.t676 699.617
R275 VGND.t338 VGND.t551 691.188
R276 VGND.t215 VGND.t203 691.188
R277 VGND.t670 VGND.t294 691.188
R278 VGND VGND.t590 682.76
R279 VGND.t776 VGND.t726 674.331
R280 VGND.t531 VGND 674.331
R281 VGND.t781 VGND.t482 674.331
R282 VGND.t666 VGND.t53 674.331
R283 VGND.t416 VGND.t238 657.471
R284 VGND.t32 VGND.t424 657.471
R285 VGND.t55 VGND.t623 657.471
R286 VGND.t226 VGND.t766 657.471
R287 VGND VGND.t193 650.173
R288 VGND.t88 VGND 649.043
R289 VGND.n1098 VGND 646.199
R290 VGND VGND.t438 641.101
R291 VGND.t222 VGND.t278 640.614
R292 VGND.t271 VGND.t592 640.614
R293 VGND VGND.t6 632.184
R294 VGND VGND.n697 632.184
R295 VGND.t180 VGND 632.184
R296 VGND.t533 VGND.t217 632.184
R297 VGND VGND.n617 632.184
R298 VGND VGND.t94 632.184
R299 VGND VGND.n434 632.184
R300 VGND.t292 VGND.t664 632.184
R301 VGND.n1092 VGND 632.184
R302 VGND VGND.t153 632.184
R303 VGND VGND.n337 632.184
R304 VGND VGND.n300 632.184
R305 VGND VGND.t156 632.184
R306 VGND VGND.n196 632.184
R307 VGND.n1095 VGND 632.184
R308 VGND VGND.t451 632.184
R309 VGND VGND.n117 632.184
R310 VGND VGND.n78 632.184
R311 VGND.t517 VGND.t417 623.755
R312 VGND.t507 VGND.t220 615.327
R313 VGND.n1264 VGND.t533 615.327
R314 VGND.t535 VGND.t426 615.327
R315 VGND.t701 VGND.t809 615.327
R316 VGND.t347 VGND 613.884
R317 VGND.t637 VGND.t655 606.898
R318 VGND.t655 VGND.t804 606.898
R319 VGND.t704 VGND.t613 606.898
R320 VGND.t613 VGND.t267 606.898
R321 VGND.t784 VGND.t357 606.898
R322 VGND.t496 VGND.t511 606.898
R323 VGND.t575 VGND.t320 606.898
R324 VGND.t471 VGND.t755 606.898
R325 VGND.t430 VGND.t471 606.898
R326 VGND.t762 VGND.t612 598.467
R327 VGND.t207 VGND.t808 598.467
R328 VGND.t812 VGND.t547 598.467
R329 VGND.t764 VGND.t280 598.467
R330 VGND.t674 VGND.t748 598.467
R331 VGND.n1258 VGND.t198 597.491
R332 VGND.t480 VGND.t672 590.038
R333 VGND VGND.t353 581.61
R334 VGND.t623 VGND 581.61
R335 VGND.t682 VGND.t274 581.61
R336 VGND.t229 VGND.t646 573.181
R337 VGND.t57 VGND.t702 568.523
R338 VGND.t714 VGND 564.751
R339 VGND.t260 VGND.t34 564.751
R340 VGND.t755 VGND 564.751
R341 VGND.t746 VGND.t654 556.322
R342 VGND.t750 VGND.t692 556.322
R343 VGND VGND.t753 556.322
R344 VGND.t267 VGND 547.894
R345 VGND.t264 VGND.t361 547.894
R346 VGND.t436 VGND 547.894
R347 VGND.t261 VGND.t815 547.894
R348 VGND.t649 VGND 547.894
R349 VGND.t266 VGND 547.894
R350 VGND VGND.t616 547.894
R351 VGND VGND.t430 547.894
R352 VGND VGND.t246 542.288
R353 VGND VGND.t397 539.465
R354 VGND VGND.t743 539.465
R355 VGND.t373 VGND 531.034
R356 VGND VGND.t441 531.034
R357 VGND VGND.t12 531.034
R358 VGND VGND.t109 531.034
R359 VGND.t529 VGND 522.606
R360 VGND VGND.t786 522.606
R361 VGND.t728 VGND 514.177
R362 VGND.t644 VGND.t419 514.177
R363 VGND VGND.t46 514.177
R364 VGND.t237 VGND.t629 505.748
R365 VGND VGND.t739 505.748
R366 VGND.t357 VGND 497.318
R367 VGND.t768 VGND.t509 497.318
R368 VGND.t581 VGND.t344 497.318
R369 VGND.t36 VGND.t644 488.889
R370 VGND.t778 VGND 480.461
R371 VGND.t523 VGND.t494 480.461
R372 VGND.t640 VGND 480.461
R373 VGND.t747 VGND.t668 480.461
R374 VGND.t660 VGND 477.801
R375 VGND.t434 VGND 477.801
R376 VGND.t708 VGND 477.801
R377 VGND VGND.t51 477.801
R378 VGND VGND.t489 477.801
R379 VGND.t193 VGND 468.729
R380 VGND.t438 VGND 468.729
R381 VGND VGND.t631 463.603
R382 VGND.t668 VGND.t638 463.603
R383 VGND.t688 VGND.t272 463.603
R384 VGND.t22 VGND 455.173
R385 VGND.t587 VGND.t23 455.173
R386 VGND.t361 VGND.t800 455.173
R387 VGND.t791 VGND.t261 455.173
R388 VGND.t647 VGND 446.743
R389 VGND.n1024 VGND.t778 446.743
R390 VGND.t214 VGND 446.743
R391 VGND VGND.t493 446.743
R392 VGND.t769 VGND 446.743
R393 VGND VGND.t630 446.743
R394 VGND VGND.t720 438.315
R395 VGND.t421 VGND.t415 429.885
R396 VGND.t733 VGND.t745 429.885
R397 VGND.t565 VGND 429.885
R398 VGND.t296 VGND.n847 423.368
R399 VGND.t694 VGND.n821 423.368
R400 VGND.t612 VGND.t717 404.599
R401 VGND.t717 VGND.t421 404.599
R402 VGND.t808 VGND.t26 404.599
R403 VGND.t26 VGND.t733 404.599
R404 VGND.t276 VGND 404.599
R405 VGND.t604 VGND.t497 404.599
R406 VGND VGND.t467 404.599
R407 VGND VGND.t269 404.599
R408 VGND VGND.t469 404.599
R409 VGND VGND.t539 404.599
R410 VGND.t724 VGND.t507 387.74
R411 VGND.t481 VGND.t688 387.74
R412 VGND.t415 VGND.t587 379.31
R413 VGND VGND.t235 379.31
R414 VGND.t177 VGND.t44 370.882
R415 VGND.t341 VGND 353.949
R416 VGND VGND.t198 353.949
R417 VGND.t246 VGND 353.949
R418 VGND.n736 VGND.n727 352
R419 VGND.t509 VGND.t724 337.166
R420 VGND.t630 VGND 337.166
R421 VGND.t692 VGND.t481 337.166
R422 VGND VGND.t186 329.623
R423 VGND VGND.t647 328.736
R424 VGND.t800 VGND.t237 328.736
R425 VGND.t465 VGND 328.736
R426 VGND VGND.t214 320.307
R427 VGND VGND.t212 311.877
R428 VGND.t497 VGND.t784 303.449
R429 VGND.t643 VGND 303.449
R430 VGND.t766 VGND 303.449
R431 VGND.t654 VGND.t207 295.019
R432 VGND.t813 VGND 295.019
R433 VGND.t611 VGND 286.591
R434 VGND VGND.t553 286.591
R435 VGND.t472 VGND 286.591
R436 VGND.t474 VGND.t621 285.757
R437 VGND.n240 VGND.t473 281.25
R438 VGND.n133 VGND.t833 276.531
R439 VGND.n2127 VGND.t902 276.531
R440 VGND.n1937 VGND.t907 276.531
R441 VGND.n2512 VGND.t760 275.293
R442 VGND.n616 VGND.t466 275.293
R443 VGND.n896 VGND.t648 275.293
R444 VGND.t642 VGND.t781 269.733
R445 VGND.t34 VGND.t425 269.733
R446 VGND.t422 VGND 269.733
R447 VGND.n195 VGND.t914 269.488
R448 VGND.n2280 VGND.t857 269.445
R449 VGND.t585 VGND.t57 266.118
R450 VGND.t702 VGND.t286 266.118
R451 VGND.t737 VGND.t660 266.118
R452 VGND.t806 VGND.t296 266.118
R453 VGND.t656 VGND.t434 266.118
R454 VGND.t49 VGND.t708 266.118
R455 VGND.t545 VGND.t694 266.118
R456 VGND.t51 VGND.t712 266.118
R457 VGND.t489 VGND.t505 266.118
R458 VGND.t409 VGND.t387 266.118
R459 VGND.n2488 VGND.t892 265.317
R460 VGND.n575 VGND.t834 265.317
R461 VGND.n118 VGND.t843 265.298
R462 VGND.n338 VGND.t916 265.298
R463 VGND.n137 VGND.t889 262.784
R464 VGND.n138 VGND.t891 262.784
R465 VGND.n140 VGND.t898 262.784
R466 VGND.n2328 VGND.t906 262.784
R467 VGND.n2491 VGND.t826 262.784
R468 VGND.n2492 VGND.t829 262.784
R469 VGND.n245 VGND.t895 262.784
R470 VGND.n247 VGND.t911 262.784
R471 VGND.n2131 VGND.t855 262.784
R472 VGND.n2132 VGND.t863 262.784
R473 VGND.n2134 VGND.t868 262.784
R474 VGND.n2154 VGND.t875 262.784
R475 VGND.n2088 VGND.t897 262.784
R476 VGND.n2090 VGND.t913 262.784
R477 VGND.n354 VGND.t856 262.784
R478 VGND.n355 VGND.t866 262.784
R479 VGND.n357 VGND.t869 262.784
R480 VGND.n1926 VGND.t877 262.784
R481 VGND.n387 VGND.t824 262.784
R482 VGND.n388 VGND.t827 262.784
R483 VGND.n562 VGND.t871 262.784
R484 VGND.n563 VGND.t874 262.784
R485 VGND.n936 VGND.t899 262.784
R486 VGND.n955 VGND.t908 262.784
R487 VGND.n1767 VGND.t837 262.784
R488 VGND.n1768 VGND.t841 262.784
R489 VGND.n881 VGND.t873 262.784
R490 VGND.n894 VGND.t876 262.784
R491 VGND.n750 VGND.t915 262.784
R492 VGND.n751 VGND.t921 262.784
R493 VGND.n36 VGND.t846 262.719
R494 VGND.n1087 VGND.t835 262.719
R495 VGND.n1144 VGND.t904 262.719
R496 VGND.n2364 VGND.t890 262.719
R497 VGND.n98 VGND.t844 262.719
R498 VGND.n2404 VGND.t836 262.719
R499 VGND.n81 VGND.t882 262.719
R500 VGND.n2434 VGND.t849 262.719
R501 VGND.n67 VGND.t886 262.719
R502 VGND.n67 VGND.t883 262.719
R503 VGND.n2190 VGND.t862 262.719
R504 VGND.n180 VGND.t917 262.719
R505 VGND.n177 VGND.t819 262.719
R506 VGND.n164 VGND.t847 262.719
R507 VGND.n2086 VGND.t870 262.719
R508 VGND.n2063 VGND.t859 262.719
R509 VGND.n1962 VGND.t865 262.719
R510 VGND.n319 VGND.t919 262.719
R511 VGND.n2002 VGND.t918 262.719
R512 VGND.n303 VGND.t848 262.719
R513 VGND.n2032 VGND.t820 262.719
R514 VGND.n534 VGND.t822 262.719
R515 VGND.n419 VGND.t825 262.719
R516 VGND.n1877 VGND.t867 262.719
R517 VGND.n684 VGND.t901 262.719
R518 VGND.n1030 VGND.t839 262.719
R519 VGND VGND.t373 261.303
R520 VGND VGND.t282 261.303
R521 VGND VGND.t788 261.303
R522 VGND VGND.t589 261.303
R523 VGND VGND.t48 261.303
R524 VGND VGND.t637 261.303
R525 VGND.t147 VGND 261.303
R526 VGND.t478 VGND.t264 261.303
R527 VGND.t793 VGND 261.303
R528 VGND.t638 VGND.t678 261.303
R529 VGND.t428 VGND 261.303
R530 VGND.n25 VGND.t885 259.082
R531 VGND.n1053 VGND.t900 259.082
R532 VGND.n1297 VGND.t909 259.082
R533 VGND.n1606 VGND.t817 259.082
R534 VGND.n774 VGND.t821 259.082
R535 VGND.n1376 VGND.t838 259.082
R536 VGND.n1578 VGND.t884 259.082
R537 VGND.n1221 VGND.t853 259.082
R538 VGND.n1167 VGND.t840 259.082
R539 VGND VGND.t478 252.875
R540 VGND.t469 VGND.t791 252.875
R541 VGND.t30 VGND 252.875
R542 VGND.t272 VGND.t684 252.875
R543 VGND.t15 VGND 252.875
R544 VGND.n237 VGND.t41 251
R545 VGND.n237 VGND.t288 251
R546 VGND.n1720 VGND.t281 251
R547 VGND.n1743 VGND.t35 251
R548 VGND.n1350 VGND.t228 251
R549 VGND.n792 VGND.t783 251
R550 VGND.n1835 VGND.t293 245.82
R551 VGND.n972 VGND.t550 245.82
R552 VGND.n1272 VGND.t216 245.82
R553 VGND.n997 VGND.t779 245.82
R554 VGND.t397 VGND 244.445
R555 VGND VGND.t97 244.445
R556 VGND.t672 VGND.t747 244.445
R557 VGND VGND.t135 244.445
R558 VGND VGND.t170 244.445
R559 VGND VGND.t379 243.542
R560 VGND VGND.n1258 243.542
R561 VGND.n1098 VGND 243.542
R562 VGND.n224 VGND.t742 243.028
R563 VGND.n224 VGND.t799 243.028
R564 VGND.n1682 VGND.t483 243.028
R565 VGND.n1748 VGND.t625 243.028
R566 VGND.n1005 VGND.t729 243.028
R567 VGND.n1651 VGND.t771 243.028
R568 VGND.n1822 VGND.t671 242.067
R569 VGND.n926 VGND.t514 242.067
R570 VGND.n1870 VGND.t366 240.948
R571 VGND.n642 VGND.t204 240.948
R572 VGND.n458 VGND.t639 238.675
R573 VGND.n1311 VGND.t418 238.675
R574 VGND.n1785 VGND.t740 238.675
R575 VGND.n775 VGND.t45 238.675
R576 VGND.n558 VGND.t576 238.44
R577 VGND.n1813 VGND.t617 237.327
R578 VGND.n1890 VGND.t650 237.327
R579 VGND.t494 VGND.t519 236.016
R580 VGND.t602 VGND 236.016
R581 VGND.t599 VGND.t260 236.016
R582 VGND.n2062 VGND.t775 235.607
R583 VGND.n672 VGND.n669 234.667
R584 VGND.n1692 VGND.t659 230.977
R585 VGND.n910 VGND.t588 230.977
R586 VGND.n253 VGND.t758 229.833
R587 VGND.n636 VGND.n635 228.294
R588 VGND.n783 VGND.n724 228.294
R589 VGND.t511 VGND.t768 227.587
R590 VGND.t269 VGND.t523 227.587
R591 VGND VGND.t300 227.587
R592 VGND.t344 VGND.t577 227.587
R593 VGND.n2213 VGND.t336 227.256
R594 VGND VGND.t347 226.804
R595 VGND.n1806 VGND.t423 226.708
R596 VGND.n959 VGND.t858 224.196
R597 VGND.n103 VGND.t912 224.102
R598 VGND.n324 VGND.t879 224.102
R599 VGND.n2039 VGND.t331 223.282
R600 VGND.n1824 VGND.n479 222.691
R601 VGND.n297 VGND.t851 221.972
R602 VGND.n1719 VGND.n1717 221.804
R603 VGND.n619 VGND.t893 220.952
R604 VGND.n1711 VGND.t896 220.952
R605 VGND.n299 VGND.t306 219.972
R606 VGND.n239 VGND.n213 218.506
R607 VGND.n239 VGND.n214 218.506
R608 VGND.n967 VGND.n932 218.506
R609 VGND.n1289 VGND.n1268 218.506
R610 VGND.n606 VGND.n605 218.506
R611 VGND.n902 VGND.n901 218.506
R612 VGND.n1014 VGND.n1013 218.506
R613 VGND.n718 VGND.n706 218.506
R614 VGND.n2489 VGND.t894 218.308
R615 VGND.n243 VGND.t860 218.308
R616 VGND.n2287 VGND.t850 218.308
R617 VGND.n569 VGND.t830 218.308
R618 VGND.n1815 VGND.t818 218.308
R619 VGND.n897 VGND.t823 218.308
R620 VGND.n1404 VGND.t888 218.308
R621 VGND.n1502 VGND.t831 218.308
R622 VGND.n1673 VGND.n641 218.13
R623 VGND.n2411 VGND.t404 217.977
R624 VGND.n2390 VGND.t1 217.977
R625 VGND.n2009 VGND.t351 217.977
R626 VGND.n1988 VGND.t463 217.977
R627 VGND.n116 VGND.t81 217.953
R628 VGND.n336 VGND.t456 217.953
R629 VGND.n2409 VGND.t319 217.892
R630 VGND.n2007 VGND.t369 217.892
R631 VGND.n406 VGND.t163 216.933
R632 VGND.n104 VGND.t171 216.589
R633 VGND.n325 VGND.t136 216.589
R634 VGND.n2044 VGND.t16 216.579
R635 VGND.n933 VGND.t339 215.992
R636 VGND.n103 VGND.t172 214.487
R637 VGND.n324 VGND.t137 214.487
R638 VGND.n1099 VGND.t130 214.456
R639 VGND.n2536 VGND.t131 214.456
R640 VGND.n21 VGND.t334 214.456
R641 VGND.n2559 VGND.t333 214.456
R642 VGND.n24 VGND.t248 214.456
R643 VGND.n22 VGND.t247 214.456
R644 VGND.n1163 VGND.t381 214.456
R645 VGND.n1168 VGND.t380 214.456
R646 VGND.n1220 VGND.t343 214.456
R647 VGND.n1223 VGND.t342 214.456
R648 VGND.n1182 VGND.t92 214.456
R649 VGND.n1205 VGND.t93 214.456
R650 VGND.n1028 VGND.t378 214.456
R651 VGND.n1191 VGND.t377 214.456
R652 VGND.n1052 VGND.t200 214.456
R653 VGND.n1051 VGND.t199 214.456
R654 VGND.n1138 VGND.t134 214.456
R655 VGND.n1066 VGND.t133 214.456
R656 VGND.n1088 VGND.t105 214.456
R657 VGND.n1071 VGND.t104 214.456
R658 VGND.n2490 VGND.t111 214.456
R659 VGND.n2490 VGND.t461 214.456
R660 VGND.n2500 VGND.t460 214.456
R661 VGND.n2477 VGND.t110 214.456
R662 VGND.n65 VGND.t447 214.456
R663 VGND.n2443 VGND.t446 214.456
R664 VGND.n65 VGND.t396 214.456
R665 VGND.n2443 VGND.t395 214.456
R666 VGND.n77 VGND.t75 214.456
R667 VGND.n79 VGND.t405 214.456
R668 VGND.n2414 VGND.t74 214.456
R669 VGND.n96 VGND.t2 214.456
R670 VGND.n2392 VGND.t318 214.456
R671 VGND.n122 VGND.t80 214.456
R672 VGND.n2371 VGND.t450 214.456
R673 VGND.n123 VGND.t325 214.456
R674 VGND.n2342 VGND.t449 214.456
R675 VGND.n2335 VGND.t146 214.456
R676 VGND.n136 VGND.t324 214.456
R677 VGND.n136 VGND.t145 214.456
R678 VGND.n137 VGND.t458 214.456
R679 VGND.n137 VGND.t457 214.456
R680 VGND.n138 VGND.t453 214.456
R681 VGND.n138 VGND.t452 214.456
R682 VGND.n140 VGND.t176 214.456
R683 VGND.n140 VGND.t175 214.456
R684 VGND.n2328 VGND.t119 214.456
R685 VGND.n2328 VGND.t118 214.456
R686 VGND.n2491 VGND.t314 214.456
R687 VGND.n2491 VGND.t313 214.456
R688 VGND.n2492 VGND.t304 214.456
R689 VGND.n2492 VGND.t303 214.456
R690 VGND.n162 VGND.t245 214.456
R691 VGND.n2267 VGND.t13 214.456
R692 VGND.n2288 VGND.t251 214.456
R693 VGND.n2281 VGND.t250 214.456
R694 VGND.n2288 VGND.t14 214.456
R695 VGND.n244 VGND.t167 214.456
R696 VGND.n255 VGND.t166 214.456
R697 VGND.n245 VGND.t87 214.456
R698 VGND.n245 VGND.t86 214.456
R699 VGND.n247 VGND.t169 214.456
R700 VGND.n247 VGND.t168 214.456
R701 VGND.n2246 VGND.t244 214.456
R702 VGND.n2251 VGND.t443 214.456
R703 VGND.n178 VGND.t337 214.456
R704 VGND.n2235 VGND.t442 214.456
R705 VGND.n185 VGND.t402 214.456
R706 VGND.n2207 VGND.t328 214.456
R707 VGND.n194 VGND.t401 214.456
R708 VGND.n200 VGND.t327 214.456
R709 VGND.n2197 VGND.t254 214.456
R710 VGND.n201 VGND.t102 214.456
R711 VGND.n2168 VGND.t253 214.456
R712 VGND.n2161 VGND.t84 214.456
R713 VGND.n2130 VGND.t101 214.456
R714 VGND.n2130 VGND.t83 214.456
R715 VGND.n2131 VGND.t158 214.456
R716 VGND.n2131 VGND.t157 214.456
R717 VGND.n2132 VGND.t256 214.456
R718 VGND.n2132 VGND.t255 214.456
R719 VGND.n2134 VGND.t128 214.456
R720 VGND.n2134 VGND.t127 214.456
R721 VGND.n2154 VGND.t190 214.456
R722 VGND.n2154 VGND.t189 214.456
R723 VGND.n2033 VGND.t352 214.456
R724 VGND.n2012 VGND.t330 214.456
R725 VGND.n297 VGND.t307 214.456
R726 VGND.n283 VGND.t17 214.456
R727 VGND.n2075 VGND.t160 214.456
R728 VGND.n2087 VGND.t63 214.456
R729 VGND.n2082 VGND.t62 214.456
R730 VGND.n2087 VGND.t161 214.456
R731 VGND.n2088 VGND.t140 214.456
R732 VGND.n2088 VGND.t139 214.456
R733 VGND.n2090 VGND.t174 214.456
R734 VGND.n2090 VGND.t173 214.456
R735 VGND.n317 VGND.t464 214.456
R736 VGND.n1990 VGND.t368 214.456
R737 VGND.n342 VGND.t455 214.456
R738 VGND.n1969 VGND.t152 214.456
R739 VGND.n343 VGND.t393 214.456
R740 VGND.n349 VGND.t151 214.456
R741 VGND.n350 VGND.t5 214.456
R742 VGND.n353 VGND.t392 214.456
R743 VGND.n353 VGND.t4 214.456
R744 VGND.n354 VGND.t316 214.456
R745 VGND.n354 VGND.t315 214.456
R746 VGND.n355 VGND.t155 214.456
R747 VGND.n355 VGND.t154 214.456
R748 VGND.n357 VGND.t72 214.456
R749 VGND.n357 VGND.t71 214.456
R750 VGND.n1926 VGND.t192 214.456
R751 VGND.n1926 VGND.t191 214.456
R752 VGND.n387 VGND.t96 214.456
R753 VGND.n387 VGND.t95 214.456
R754 VGND.n388 VGND.t312 214.456
R755 VGND.n388 VGND.t311 214.456
R756 VGND.n1814 VGND.t125 214.456
R757 VGND.n484 VGND.t124 214.456
R758 VGND.n506 VGND.t346 214.456
R759 VGND.n1804 VGND.t345 214.456
R760 VGND.n548 VGND.t321 214.456
R761 VGND.n568 VGND.t372 214.456
R762 VGND.n560 VGND.t371 214.456
R763 VGND.n568 VGND.t322 214.456
R764 VGND.n562 VGND.t78 214.456
R765 VGND.n562 VGND.t77 214.456
R766 VGND.n563 VGND.t202 214.456
R767 VGND.n563 VGND.t201 214.456
R768 VGND.n436 VGND.t66 214.456
R769 VGND.n1891 VGND.t65 214.456
R770 VGND.n427 VGND.t99 214.456
R771 VGND.n380 VGND.t98 214.456
R772 VGND.n412 VGND.t164 214.456
R773 VGND.n1763 VGND.t399 214.456
R774 VGND.n1759 VGND.t398 214.456
R775 VGND.n1296 VGND.t185 214.456
R776 VGND.n993 VGND.t184 214.456
R777 VGND.n976 VGND.t340 214.456
R778 VGND.n959 VGND.t149 214.456
R779 VGND.n958 VGND.t148 214.456
R780 VGND.n936 VGND.t390 214.456
R781 VGND.n936 VGND.t389 214.456
R782 VGND.n955 VGND.t182 214.456
R783 VGND.n955 VGND.t181 214.456
R784 VGND.n619 VGND.t197 214.456
R785 VGND.n619 VGND.t196 214.456
R786 VGND.n1711 VGND.t116 214.456
R787 VGND.n1711 VGND.t115 214.456
R788 VGND.n1767 VGND.t445 214.456
R789 VGND.n1767 VGND.t444 214.456
R790 VGND.n1768 VGND.t69 214.456
R791 VGND.n1768 VGND.t68 214.456
R792 VGND.n755 VGND.t259 214.456
R793 VGND.n747 VGND.t258 214.456
R794 VGND.n755 VGND.t242 214.456
R795 VGND.n739 VGND.t241 214.456
R796 VGND.n773 VGND.t179 214.456
R797 VGND.n777 VGND.t178 214.456
R798 VGND.n1605 VGND.t90 214.456
R799 VGND.n698 VGND.t89 214.456
R800 VGND.n1623 VGND.t143 214.456
R801 VGND.n1645 VGND.t142 214.456
R802 VGND.n898 VGND.t375 214.456
R803 VGND.n1361 VGND.t374 214.456
R804 VGND.n881 VGND.t19 214.456
R805 VGND.n881 VGND.t18 214.456
R806 VGND.n894 VGND.t8 214.456
R807 VGND.n894 VGND.t7 214.456
R808 VGND.n750 VGND.t113 214.456
R809 VGND.n750 VGND.t112 214.456
R810 VGND.n751 VGND.t108 214.456
R811 VGND.n751 VGND.t107 214.456
R812 VGND.n868 VGND.t349 214.456
R813 VGND.n1375 VGND.t348 214.456
R814 VGND.n1403 VGND.t195 214.456
R815 VGND.n1401 VGND.t194 214.456
R816 VGND.n1428 VGND.t383 214.456
R817 VGND.n1430 VGND.t384 214.456
R818 VGND.n1577 VGND.t188 214.456
R819 VGND.n1575 VGND.t187 214.456
R820 VGND.n1554 VGND.t122 214.456
R821 VGND.n1552 VGND.t121 214.456
R822 VGND.n813 VGND.t11 214.456
R823 VGND.n1514 VGND.t10 214.456
R824 VGND.n1501 VGND.t440 214.456
R825 VGND.n1499 VGND.t439 214.456
R826 VGND.n1475 VGND.t310 214.456
R827 VGND.n1473 VGND.t309 214.456
R828 VGND.n1446 VGND.t408 214.456
R829 VGND.n845 VGND.t407 214.456
R830 VGND.n1682 VGND.n1681 212.317
R831 VGND VGND.t714 210.728
R832 VGND.n1704 VGND.n621 207.965
R833 VGND.n790 VGND.n720 207.965
R834 VGND.n439 VGND.n438 206.909
R835 VGND.n1304 VGND.n1303 205.971
R836 VGND.n1841 VGND.n461 205.899
R837 VGND.n1844 VGND.n1843 205.899
R838 VGND.n463 VGND.n462 205.481
R839 VGND.n1316 VGND.n986 205.481
R840 VGND.n546 VGND.n545 205.385
R841 VGND.n1824 VGND.n478 204.692
R842 VGND.n1851 VGND.n1850 204.692
R843 VGND.n1617 VGND.n694 204.457
R844 VGND.n1617 VGND.n695 204.457
R845 VGND.n708 VGND.n707 204.457
R846 VGND.n2069 VGND.n2068 204.201
R847 VGND.n1637 VGND.n675 204.201
R848 VGND.n685 VGND.n683 204.201
R849 VGND.n488 VGND.n487 202.724
R850 VGND.n523 VGND.n522 202.724
R851 VGND.n1859 VGND.n452 202.724
R852 VGND.n1288 VGND.n1269 202.724
R853 VGND.n1273 VGND.n1270 202.724
R854 VGND.t547 VGND.t782 202.299
R855 VGND VGND.t525 202.299
R856 VGND.t263 VGND.t764 202.299
R857 VGND.t715 VGND.t598 202.299
R858 VGND.n540 VGND.n508 201.458
R859 VGND.n1309 VGND.n990 201.458
R860 VGND.n1834 VGND.n465 201.129
R861 VGND.n555 VGND.n503 201.129
R862 VGND.n550 VGND.n549 201.129
R863 VGND.n988 VGND.n987 201.129
R864 VGND.n2542 VGND.n2537 200.692
R865 VGND.n1207 VGND.n1206 200.692
R866 VGND.n2229 VGND.n2228 200.692
R867 VGND.n975 VGND.n974 200.692
R868 VGND.n1539 VGND.n1538 200.692
R869 VGND.n1707 VGND.n1706 200.516
R870 VGND.n906 VGND.n905 200.516
R871 VGND.n557 VGND.n502 200.508
R872 VGND.n532 VGND.n512 200.508
R873 VGND.n510 VGND.n509 200.508
R874 VGND.n457 VGND.n456 200.508
R875 VGND.n984 VGND.n924 200.508
R876 VGND.n1298 VGND.n995 200.508
R877 VGND.n1266 VGND.n1265 200.508
R878 VGND.n1821 VGND.n482 200.231
R879 VGND.n1719 VGND.n1718 200.127
R880 VGND.n1355 VGND.n900 200.127
R881 VGND.n2565 VGND.n2564 199.739
R882 VGND.n2291 VGND.n158 199.739
R883 VGND.n2291 VGND.n159 199.739
R884 VGND.n1869 VGND.n440 199.739
R885 VGND.n1687 VGND.n1686 199.739
R886 VGND.n1001 VGND.n1000 199.739
R887 VGND.n1437 VGND.n848 199.739
R888 VGND.n1410 VGND.n858 199.739
R889 VGND.n1396 VGND.n864 199.739
R890 VGND.n866 VGND.n865 199.739
R891 VGND.n1467 VGND.n1466 199.739
R892 VGND.n1486 VGND.n1482 199.739
R893 VGND.n1509 VGND.n1508 199.739
R894 VGND.n1546 VGND.n1545 199.739
R895 VGND.n1571 VGND.n1570 199.739
R896 VGND.n1584 VGND.n1574 199.739
R897 VGND.n285 VGND.n284 199.662
R898 VGND.n230 VGND.n218 199.53
R899 VGND.n230 VGND.n220 199.53
R900 VGND.n1845 VGND.n1842 199.53
R901 VGND.n1675 VGND.n1674 199.53
R902 VGND.n1742 VGND.n607 199.53
R903 VGND.n1343 VGND.n908 199.53
R904 VGND.n1657 VGND.n657 199.53
R905 VGND.n784 VGND.n723 199.53
R906 VGND.n425 VGND.n374 197.476
R907 VGND.n2484 VGND.n61 196.831
R908 VGND.n982 VGND.n925 196.589
R909 VGND.n1750 VGND.n602 196.589
R910 VGND.n418 VGND.n377 196.442
R911 VGND.n1858 VGND.n453 196.442
R912 VGND.n992 VGND.n991 196.442
R913 VGND.n1752 VGND.n1751 196.442
R914 VGND.n1774 VGND.n1762 196.442
R915 VGND.t238 VGND.t762 193.87
R916 VGND.t419 VGND.t32 193.87
R917 VGND.t286 VGND 190.516
R918 VGND.n2544 VGND.n2543 190.399
R919 VGND.n1187 VGND.n1185 190.399
R920 VGND.n2227 VGND.n2226 190.399
R921 VGND.n930 VGND.n929 190.399
R922 VGND.n1537 VGND.n1536 190.399
R923 VGND.n672 VGND.n671 189.268
R924 VGND.n736 VGND.n735 189.201
R925 VGND.t48 VGND.t746 185.441
R926 VGND.t412 VGND.t624 185.441
R927 VGND.t797 VGND.t227 177.012
R928 VGND.t788 VGND.t416 177.012
R929 VGND.t809 VGND.t608 177.012
R930 VGND.t300 VGND.t602 168.583
R931 VGND.t664 VGND.t750 168.583
R932 VGND.n1757 VGND.t716 154.131
R933 VGND.n2060 VGND.t744 152.381
R934 VGND.n1786 VGND.t360 152.381
R935 VGND.n1766 VGND.t31 152.381
R936 VGND.n2542 VGND.n2541 152
R937 VGND.n2228 VGND.n184 152
R938 VGND.n974 VGND.n973 152
R939 VGND.n1538 VGND.n812 152
R940 VGND.n1208 VGND.n1207 152
R941 VGND.n2045 VGND.t635 150.101
R942 VGND.n1766 VGND.t354 150.101
R943 VGND.n1737 VGND.t765 144.886
R944 VGND.n1349 VGND.t798 144.886
R945 VGND VGND.t88 143.296
R946 VGND VGND.n617 143.296
R947 VGND.t274 VGND.t205 143.296
R948 VGND.t284 VGND.t229 134.867
R949 VGND.t646 VGND.t290 134.867
R950 VGND.t211 VGND.t618 134.867
R951 VGND.t676 VGND.t480 134.867
R952 VGND.t748 VGND.t682 126.438
R953 VGND.n64 VGND.t652 124.688
R954 VGND.n1763 VGND.t910 121.927
R955 VGND.n1430 VGND.t828 121.927
R956 VGND.n1554 VGND.t920 121.927
R957 VGND.n1475 VGND.t845 121.927
R958 VGND.n1446 VGND.t905 121.927
R959 VGND.t298 VGND.t611 118.008
R960 VGND.t537 VGND.t496 118.008
R961 VGND.t205 VGND 118.008
R962 VGND.t320 VGND.t571 118.008
R963 VGND.n756 VGND.t878 116.734
R964 VGND.n413 VGND.t864 116.734
R965 VGND.n660 VGND.n659 114.377
R966 VGND.n1884 VGND.n431 110.349
R967 VGND.n1012 VGND.n999 110.349
R968 VGND.t28 VGND.t812 109.579
R969 VGND.t220 VGND.t513 109.579
R970 VGND.n1264 VGND.t529 109.579
R971 VGND.t426 VGND.t730 109.579
R972 VGND.t203 VGND.t643 109.579
R973 VGND.n431 VGND.t607 108.505
R974 VGND.n999 VGND.t236 108.505
R975 VGND.n659 VGND.t734 108.505
R976 VGND.n2335 VGND.t881 102.353
R977 VGND.n2161 VGND.t852 102.353
R978 VGND.n350 VGND.t854 102.353
R979 VGND.n2068 VGND.t756 101.43
R980 VGND.n675 VGND.t805 101.43
R981 VGND.n683 VGND.t705 101.43
R982 VGND.t417 VGND.t515 101.15
R983 VGND.t633 VGND.t64 101.15
R984 VGND.n2096 VGND.t861 99.7825
R985 VGND.n748 VGND.t880 99.7825
R986 VGND VGND.t474 94.1702
R987 VGND.t811 VGND 92.7208
R988 VGND.t527 VGND 92.7208
R989 VGND.t217 VGND.t535 92.7208
R990 VGND.t219 VGND.t431 92.7208
R991 VGND.t614 VGND.t701 92.7208
R992 VGND.t686 VGND.t292 92.7208
R993 VGND VGND.t585 87.6981
R994 VGND VGND.t737 87.6981
R995 VGND VGND.t806 87.6981
R996 VGND VGND.t656 87.6981
R997 VGND VGND.t49 87.6981
R998 VGND VGND.t545 87.6981
R999 VGND.t712 VGND 87.6981
R1000 VGND.t505 VGND 87.6981
R1001 VGND.t387 VGND 87.6981
R1002 VGND.t109 VGND.t759 84.2917
R1003 VGND.t59 VGND.t491 75.8626
R1004 VGND.n218 VGND.t732 74.8666
R1005 VGND.n220 VGND.t700 74.8666
R1006 VGND.n1842 VGND.t273 74.8666
R1007 VGND.n925 VGND.t221 74.8666
R1008 VGND.n1674 VGND.t265 74.8666
R1009 VGND.n607 VGND.t420 74.8666
R1010 VGND.n602 VGND.t816 74.8666
R1011 VGND.n908 VGND.t763 74.8666
R1012 VGND.n657 VGND.t208 74.8666
R1013 VGND.n723 VGND.t502 74.8666
R1014 VGND.n694 VGND.t610 72.8576
R1015 VGND.n695 VGND.t544 72.8576
R1016 VGND.n707 VGND.t358 72.8576
R1017 VGND.t268 VGND.t20 67.4335
R1018 VGND.t278 VGND.t432 67.4335
R1019 VGND.t592 VGND.t222 67.4335
R1020 VGND.t590 VGND.t541 59.0043
R1021 VGND.n482 VGND.t767 58.5719
R1022 VGND.n374 VGND.t56 58.5719
R1023 VGND.n284 VGND.t773 52.8576
R1024 VGND VGND.t527 50.5752
R1025 VGND.t53 VGND.t662 50.5752
R1026 VGND.n641 VGND.t362 48.5719
R1027 VGND.n635 VGND.t721 47.1434
R1028 VGND.n724 VGND.t60 47.1434
R1029 VGND.n218 VGND.t719 40.0005
R1030 VGND.n220 VGND.t698 40.0005
R1031 VGND.n284 VGND.t754 40.0005
R1032 VGND.n465 VGND.t687 40.0005
R1033 VGND.n465 VGND.t691 40.0005
R1034 VGND.n503 VGND.t564 40.0005
R1035 VGND.n503 VGND.t568 40.0005
R1036 VGND.n549 VGND.t558 40.0005
R1037 VGND.n549 VGND.t562 40.0005
R1038 VGND.n502 VGND.t570 40.0005
R1039 VGND.n502 VGND.t572 40.0005
R1040 VGND.n487 VGND.t628 40.0005
R1041 VGND.n487 VGND.t43 40.0005
R1042 VGND.n522 VGND.t225 40.0005
R1043 VGND.n522 VGND.t574 40.0005
R1044 VGND.n512 VGND.t578 40.0005
R1045 VGND.n512 VGND.t582 40.0005
R1046 VGND.n509 VGND.t584 40.0005
R1047 VGND.n509 VGND.t580 40.0005
R1048 VGND.n508 VGND.t556 40.0005
R1049 VGND.n508 VGND.t560 40.0005
R1050 VGND.n545 VGND.t554 40.0005
R1051 VGND.n461 VGND.t685 40.0005
R1052 VGND.n462 VGND.t693 40.0005
R1053 VGND.n462 VGND.t665 40.0005
R1054 VGND.n478 VGND.t663 40.0005
R1055 VGND.n478 VGND.t667 40.0005
R1056 VGND.n1842 VGND.t601 40.0005
R1057 VGND.n1843 VGND.t677 40.0005
R1058 VGND.n1843 VGND.t681 40.0005
R1059 VGND.n1850 VGND.t669 40.0005
R1060 VGND.n1850 VGND.t673 40.0005
R1061 VGND.n456 VGND.t675 40.0005
R1062 VGND.n456 VGND.t679 40.0005
R1063 VGND.n452 VGND.t206 40.0005
R1064 VGND.n452 VGND.t683 40.0005
R1065 VGND.n438 VGND.t364 40.0005
R1066 VGND.n438 VGND.t632 40.0005
R1067 VGND.n924 VGND.t508 40.0005
R1068 VGND.n924 VGND.t510 40.0005
R1069 VGND.n925 VGND.t725 40.0005
R1070 VGND.n986 VGND.t512 40.0005
R1071 VGND.n986 VGND.t538 40.0005
R1072 VGND.n987 VGND.t516 40.0005
R1073 VGND.n987 VGND.t518 40.0005
R1074 VGND.n990 VGND.t524 40.0005
R1075 VGND.n1303 VGND.t528 40.0005
R1076 VGND.n1303 VGND.t532 40.0005
R1077 VGND.n995 VGND.t522 40.0005
R1078 VGND.n995 VGND.t526 40.0005
R1079 VGND.n1265 VGND.t530 40.0005
R1080 VGND.n1265 VGND.t534 40.0005
R1081 VGND.n1269 VGND.t536 40.0005
R1082 VGND.n1269 VGND.t731 40.0005
R1083 VGND.n1270 VGND.t485 40.0005
R1084 VGND.n1270 VGND.t477 40.0005
R1085 VGND.n1674 VGND.t801 40.0005
R1086 VGND.n607 VGND.t37 40.0005
R1087 VGND.n602 VGND.t792 40.0005
R1088 VGND.n908 VGND.t718 40.0005
R1089 VGND.n657 VGND.t27 40.0005
R1090 VGND.n723 VGND.t492 40.0005
R1091 VGND.n431 VGND.t595 38.7697
R1092 VGND.n1706 VGND.t437 38.7697
R1093 VGND.n905 VGND.t789 38.7697
R1094 VGND.n999 VGND.t727 38.7697
R1095 VGND.n659 VGND.t619 38.7697
R1096 VGND.n158 VGND.t636 38.5719
R1097 VGND.n158 VGND.t780 38.5719
R1098 VGND.n159 VGND.t429 38.5719
R1099 VGND.n159 VGND.t232 38.5719
R1100 VGND.n545 VGND.t566 38.5719
R1101 VGND.n461 VGND.t689 38.5719
R1102 VGND.n453 VGND.t275 38.5719
R1103 VGND.n453 VGND.t749 38.5719
R1104 VGND.n990 VGND.t520 38.5719
R1105 VGND.n991 VGND.t495 38.5719
R1106 VGND.n991 VGND.t270 38.5719
R1107 VGND.n1681 VGND.t736 38.5719
R1108 VGND.n1681 VGND.t723 38.5719
R1109 VGND.n1686 VGND.t641 38.5719
R1110 VGND.n1686 VGND.t301 38.5719
R1111 VGND.n1751 VGND.t262 38.5719
R1112 VGND.n1751 VGND.t470 38.5719
R1113 VGND.n1762 VGND.t597 38.5719
R1114 VGND.n1762 VGND.t540 38.5719
R1115 VGND.n1000 VGND.t21 38.5719
R1116 VGND.n1000 VGND.t299 38.5719
R1117 VGND.n671 VGND.t213 38.5719
R1118 VGND.n671 VGND.t277 38.5719
R1119 VGND.n735 VGND.t814 38.5719
R1120 VGND.n735 VGND.t468 38.5719
R1121 VGND.n635 VGND.t603 35.4291
R1122 VGND.n724 VGND.t591 35.4291
R1123 VGND.n1853 VGND.n1852 34.6358
R1124 VGND.n1106 VGND.n1089 34.6358
R1125 VGND.n267 VGND.n266 34.6358
R1126 VGND.n232 VGND.n231 34.6358
R1127 VGND.n232 VGND.n216 34.6358
R1128 VGND.n236 VGND.n216 34.6358
R1129 VGND.n225 VGND.n221 34.6358
R1130 VGND.n229 VGND.n221 34.6358
R1131 VGND.n1834 VGND.n466 34.6358
R1132 VGND.n1849 VGND.n459 34.6358
R1133 VGND.n1857 VGND.n454 34.6358
R1134 VGND.n1291 VGND.n1290 34.6358
R1135 VGND.n1287 VGND.n1274 34.6358
R1136 VGND.n1672 VGND.n1671 34.6358
R1137 VGND.n1679 VGND.n639 34.6358
R1138 VGND.n1680 VGND.n1679 34.6358
R1139 VGND.n1703 VGND.n622 34.6358
R1140 VGND.n1739 VGND.n1738 34.6358
R1141 VGND.n1744 VGND.n603 34.6358
R1142 VGND.n1787 VGND.n1758 34.6358
R1143 VGND.n1011 VGND.n1010 34.6358
R1144 VGND.n1023 VGND.n996 34.6358
R1145 VGND.n1020 VGND.n1019 34.6358
R1146 VGND.n1019 VGND.n656 34.6358
R1147 VGND.n1658 VGND.n656 34.6358
R1148 VGND.n1618 VGND.n692 34.6358
R1149 VGND.n1616 VGND.n1615 34.6358
R1150 VGND.n1615 VGND.n696 34.6358
R1151 VGND.n789 VGND.n721 34.6358
R1152 VGND.n785 VGND.n721 34.6358
R1153 VGND.n782 VGND.n725 34.6358
R1154 VGND.n1411 VGND.n851 34.6358
R1155 VGND.n1395 VGND.n1394 34.6358
R1156 VGND.n1468 VGND.n836 34.6358
R1157 VGND.n1485 VGND.n824 34.6358
R1158 VGND.n1547 VGND.n808 34.6358
R1159 VGND.n1589 VGND.n1588 34.6358
R1160 VGND.n1588 VGND.n1572 34.6358
R1161 VGND.n2543 VGND.t903 34.2973
R1162 VGND.n1187 VGND.t832 34.2973
R1163 VGND.n2227 VGND.t887 34.2973
R1164 VGND.n929 VGND.t842 34.2973
R1165 VGND.n1537 VGND.t872 34.2973
R1166 VGND.n1305 VGND.n992 33.8829
R1167 VGND.n1752 VGND.n600 33.8829
R1168 VGND.t726 VGND.t710 33.717
R1169 VGND.t476 VGND.t215 33.717
R1170 VGND.t482 VGND.t735 33.717
R1171 VGND.t411 VGND 33.717
R1172 VGND.t739 VGND.t359 33.717
R1173 VGND.t294 VGND.t666 33.717
R1174 VGND.n2564 VGND.t475 33.462
R1175 VGND.n2564 VGND.t622 33.462
R1176 VGND.n377 VGND.t796 33.462
R1177 VGND.n377 VGND.t356 33.462
R1178 VGND.n440 VGND.t794 33.462
R1179 VGND.n440 VGND.t803 33.462
R1180 VGND.n848 VGND.t807 33.462
R1181 VGND.n848 VGND.t297 33.462
R1182 VGND.n858 VGND.t738 33.462
R1183 VGND.n858 VGND.t661 33.462
R1184 VGND.n864 VGND.t703 33.462
R1185 VGND.n864 VGND.t287 33.462
R1186 VGND.n865 VGND.t586 33.462
R1187 VGND.n865 VGND.t58 33.462
R1188 VGND.n1466 VGND.t657 33.462
R1189 VGND.n1466 VGND.t435 33.462
R1190 VGND.n1482 VGND.t50 33.462
R1191 VGND.n1482 VGND.t709 33.462
R1192 VGND.n1508 VGND.t546 33.462
R1193 VGND.n1508 VGND.t695 33.462
R1194 VGND.n1545 VGND.t713 33.462
R1195 VGND.n1545 VGND.t52 33.462
R1196 VGND.n1570 VGND.t506 33.462
R1197 VGND.n1570 VGND.t490 33.462
R1198 VGND.n1574 VGND.t388 33.462
R1199 VGND.n1574 VGND.t410 33.462
R1200 VGND.n641 VGND.t479 32.5719
R1201 VGND.n239 VGND.n238 32.377
R1202 VGND.n1351 VGND.n902 32.377
R1203 VGND.n1014 VGND.n996 32.377
R1204 VGND.n719 VGND.n718 32.377
R1205 VGND.n1311 VGND.n1310 32.377
R1206 VGND.n1012 VGND.n1011 31.624
R1207 VGND.n238 VGND.n237 31.2476
R1208 VGND.n1721 VGND.n1720 31.2476
R1209 VGND.n1351 VGND.n1350 31.2476
R1210 VGND.n792 VGND.n719 31.2476
R1211 VGND.n230 VGND.n229 30.8711
R1212 VGND.n1675 VGND.n639 30.8711
R1213 VGND.n1343 VGND.n1342 30.8711
R1214 VGND.n1657 VGND.n1656 30.8711
R1215 VGND.n985 VGND.n984 30.4946
R1216 VGND.n1692 VGND.n622 30.4946
R1217 VGND.n1342 VGND.n910 30.4946
R1218 VGND.n1836 VGND.n1835 30.1181
R1219 VGND.n1315 VGND.n988 30.1181
R1220 VGND.n1272 VGND.n1271 30.1181
R1221 VGND.n1020 VGND.n997 30.1181
R1222 VGND.n1840 VGND.n463 29.7417
R1223 VGND.n1716 VGND.n616 29.3652
R1224 VGND.n1824 VGND.n1823 28.9887
R1225 VGND.n1860 VGND.n1859 27.8593
R1226 VGND.n1288 VGND.n1287 27.8593
R1227 VGND.n225 VGND.n224 27.4829
R1228 VGND.n1682 VGND.n1680 27.4829
R1229 VGND.n1707 VGND.n618 27.4829
R1230 VGND.n1743 VGND.n1742 27.4829
R1231 VGND.n1748 VGND.n603 27.4829
R1232 VGND.n1348 VGND.n906 27.4829
R1233 VGND.n1005 VGND.n1002 27.4829
R1234 VGND.n1652 VGND.n660 27.4829
R1235 VGND.n1652 VGND.n1651 27.4829
R1236 VGND.n1860 VGND.n439 27.1064
R1237 VGND.n1691 VGND.n636 26.7299
R1238 VGND.n2560 VGND.n1 26.6009
R1239 VGND.n1622 VGND.n692 26.314
R1240 VGND.n2068 VGND.t47 25.9346
R1241 VGND.n675 VGND.t504 25.9346
R1242 VGND.n683 VGND.t210 25.9346
R1243 VGND.n1295 VGND.n1294 25.7355
R1244 VGND.n1604 VGND.n699 25.7355
R1245 VGND.n778 VGND.n725 25.7355
R1246 VGND.n1390 VGND.n1389 25.7355
R1247 VGND.n1583 VGND.n1582 25.7355
R1248 VGND.n1106 VGND.n1105 25.6926
R1249 VGND.n1427 VGND.n851 25.6926
R1250 VGND.n1409 VGND.n860 25.6926
R1251 VGND.n1400 VGND.n862 25.6926
R1252 VGND.n1472 VGND.n836 25.6926
R1253 VGND.n1498 VGND.n824 25.6926
R1254 VGND.n1507 VGND.n822 25.6926
R1255 VGND.n1551 VGND.n808 25.6926
R1256 VGND.n266 VGND.n240 25.6005
R1257 VGND.n1310 VGND.n1309 25.6005
R1258 VGND.n482 VGND.t787 25.4291
R1259 VGND.n374 VGND.t707 25.4291
R1260 VGND.t626 VGND.t542 25.2879
R1261 VGND.t680 VGND.t600 25.2879
R1262 VGND.t165 VGND.t757 25.2879
R1263 VGND.n1316 VGND.n985 25.224
R1264 VGND.n1316 VGND.n1315 25.224
R1265 VGND.n2566 VGND.n0 24.9894
R1266 VGND.n1544 VGND.n810 24.9894
R1267 VGND.n2290 VGND.n2289 24.968
R1268 VGND.n61 VGND.t414 24.9236
R1269 VGND.n61 VGND.t386 24.9236
R1270 VGND.n214 VGND.t696 24.9236
R1271 VGND.n214 VGND.t289 24.9236
R1272 VGND.n213 VGND.t500 24.9236
R1273 VGND.n213 VGND.t39 24.9236
R1274 VGND.n479 VGND.t54 24.9236
R1275 VGND.n479 VGND.t295 24.9236
R1276 VGND.n932 VGND.t552 24.9236
R1277 VGND.n932 VGND.t752 24.9236
R1278 VGND.n1268 VGND.t218 24.9236
R1279 VGND.n1268 VGND.t427 24.9236
R1280 VGND.n621 VGND.t615 24.9236
R1281 VGND.n621 VGND.t810 24.9236
R1282 VGND.n1706 VGND.t609 24.9236
R1283 VGND.n1718 VGND.t433 24.9236
R1284 VGND.n1718 VGND.t223 24.9236
R1285 VGND.n1717 VGND.t279 24.9236
R1286 VGND.n1717 VGND.t593 24.9236
R1287 VGND.n605 VGND.t33 24.9236
R1288 VGND.n605 VGND.t645 24.9236
R1289 VGND.n900 VGND.t283 24.9236
R1290 VGND.n900 VGND.t285 24.9236
R1291 VGND.n901 VGND.t230 24.9236
R1292 VGND.n901 VGND.t291 24.9236
R1293 VGND.n905 VGND.t239 24.9236
R1294 VGND.n1013 VGND.t777 24.9236
R1295 VGND.n1013 VGND.t711 24.9236
R1296 VGND.n706 VGND.t785 24.9236
R1297 VGND.n706 VGND.t605 24.9236
R1298 VGND.n720 VGND.t548 24.9236
R1299 VGND.n720 VGND.t29 24.9236
R1300 VGND.n982 VGND.n981 24.4711
R1301 VGND.n1750 VGND.n1749 24.4711
R1302 VGND.n1704 VGND.n1703 24.4711
R1303 VGND.n1757 VGND.n600 24.4711
R1304 VGND.n1758 VGND.n1757 24.4711
R1305 VGND.n790 VGND.n789 24.4711
R1306 VGND.n1713 VGND.n1712 23.7181
R1307 VGND.n1110 VGND.n1089 23.7181
R1308 VGND.n394 VGND.n381 23.7181
R1309 VGND.n405 VGND.n381 23.7181
R1310 VGND.n1808 VGND.n485 23.7181
R1311 VGND.n1808 VGND.n1807 23.7181
R1312 VGND.n1671 VGND.n642 23.7181
R1313 VGND.n1712 VGND.n618 23.7181
R1314 VGND.n1737 VGND.n609 23.7181
R1315 VGND.n1738 VGND.n1737 23.7181
R1316 VGND.n1349 VGND.n1348 23.7181
R1317 VGND.n1611 VGND.n696 23.7181
R1318 VGND.n1441 VGND.n846 23.7181
R1319 VGND.n1436 VGND.n849 23.7181
R1320 VGND.n1465 VGND.n838 23.7181
R1321 VGND.n1481 VGND.n834 23.7181
R1322 VGND.n1513 VGND.n820 23.7181
R1323 VGND.n1569 VGND.n804 23.7181
R1324 VGND.n1785 VGND.n1784 23.4338
R1325 VGND.n457 VGND.n454 23.3417
R1326 VGND.n1291 VGND.n1266 23.3417
R1327 VGND.n2291 VGND.n157 22.9652
R1328 VGND.n224 VGND.n157 22.9652
R1329 VGND.n1682 VGND.n637 22.9652
R1330 VGND.n1687 VGND.n637 22.9652
R1331 VGND.n1721 VGND.n1719 22.9652
R1332 VGND.n1749 VGND.n1748 22.9652
R1333 VGND.n1355 VGND.n1354 22.9652
R1334 VGND.n1006 VGND.n1005 22.9652
R1335 VGND.n1006 VGND.n1001 22.9652
R1336 VGND.n1651 VGND.n1650 22.9652
R1337 VGND.n1650 VGND.n669 22.9652
R1338 VGND.n784 VGND.n783 22.9652
R1339 VGND.n1271 VGND.n642 22.5887
R1340 VGND.n694 VGND.t25 22.3257
R1341 VGND.n695 VGND.t620 22.3257
R1342 VGND.n707 VGND.t498 22.3257
R1343 VGND.n2565 VGND.n1 22.2123
R1344 VGND.n2566 VGND.n2565 22.2123
R1345 VGND.n237 VGND.n236 22.2123
R1346 VGND.n1720 VGND.n609 22.2123
R1347 VGND.n1744 VGND.n1743 22.2123
R1348 VGND.n792 VGND.n791 22.2123
R1349 VGND.n1437 VGND.n846 22.2123
R1350 VGND.n1437 VGND.n1436 22.2123
R1351 VGND.n1411 VGND.n1410 22.2123
R1352 VGND.n1410 VGND.n1409 22.2123
R1353 VGND.n1396 VGND.n862 22.2123
R1354 VGND.n1394 VGND.n866 22.2123
R1355 VGND.n1396 VGND.n1395 22.2123
R1356 VGND.n1390 VGND.n866 22.2123
R1357 VGND.n1467 VGND.n1465 22.2123
R1358 VGND.n1468 VGND.n1467 22.2123
R1359 VGND.n1486 VGND.n1481 22.2123
R1360 VGND.n1486 VGND.n1485 22.2123
R1361 VGND.n1509 VGND.n1507 22.2123
R1362 VGND.n1509 VGND.n820 22.2123
R1363 VGND.n1546 VGND.n1544 22.2123
R1364 VGND.n1547 VGND.n1546 22.2123
R1365 VGND.n1571 VGND.n1569 22.2123
R1366 VGND.n1589 VGND.n1571 22.2123
R1367 VGND.n1584 VGND.n1572 22.2123
R1368 VGND.n1584 VGND.n1583 22.2123
R1369 VGND.n2291 VGND.n2290 21.4593
R1370 VGND.n1688 VGND.n1687 21.4593
R1371 VGND.n1719 VGND.n1716 21.4593
R1372 VGND.n1010 VGND.n1001 21.4593
R1373 VGND.n1656 VGND.n660 21.4593
R1374 VGND.n977 VGND.n926 20.8482
R1375 VGND.n1836 VGND.n463 20.7064
R1376 VGND.n1824 VGND.n466 20.7064
R1377 VGND.n1137 VGND.n1136 18.2791
R1378 VGND.n2074 VGND.n2073 18.2791
R1379 VGND.n1892 VGND.n428 18.2791
R1380 VGND.n1065 VGND.n1047 17.7007
R1381 VGND.n30 VGND.n29 17.4137
R1382 VGND.n1822 VGND.n1821 17.3181
R1383 VGND.n2444 VGND.n2442 17.195
R1384 VGND.n2040 VGND.n299 16.9936
R1385 VGND.n1204 VGND.n1188 16.9545
R1386 VGND.n1707 VGND.n1705 16.9417
R1387 VGND.n1344 VGND.n906 16.9417
R1388 VGND.t503 VGND.t141 16.8587
R1389 VGND.t751 VGND.t338 16.8587
R1390 VGND.t97 VGND.t795 16.8587
R1391 VGND.n1224 VGND.n1179 16.8353
R1392 VGND.n1219 VGND.n1180 16.7924
R1393 VGND.n2476 VGND.n64 16.763
R1394 VGND.n1841 VGND.n1840 16.1887
R1395 VGND.n1823 VGND.n1822 16.1887
R1396 VGND.n981 VGND.n926 16.1887
R1397 VGND.n1111 VGND.n1110 15.3963
R1398 VGND.n1871 VGND.n1870 15.3963
R1399 VGND.n1257 VGND.n1256 15.3963
R1400 VGND.n1257 VGND.n1026 14.8179
R1401 VGND.n1611 VGND.n1610 14.8179
R1402 VGND.n249 VGND.n248 14.775
R1403 VGND.n1812 VGND.n485 14.775
R1404 VGND.n957 VGND.n956 14.775
R1405 VGND.n1362 VGND.n895 14.775
R1406 VGND.n1442 VGND.n1441 14.775
R1407 VGND.n1515 VGND.n1513 14.775
R1408 VGND.n2474 VGND.n2473 14.2735
R1409 VGND.n772 VGND.n727 14.065
R1410 VGND.n2495 VGND.n2494 14.0503
R1411 VGND.n2092 VGND.n2091 14.0503
R1412 VGND.n567 VGND.n564 14.0503
R1413 VGND.n1692 VGND.n1691 13.9299
R1414 VGND.n1002 VGND.n910 13.9299
R1415 VGND.n754 VGND.n753 13.8859
R1416 VGND.n2329 VGND.n139 12.8005
R1417 VGND.n2155 VGND.n2133 12.8005
R1418 VGND.n1927 VGND.n356 12.8005
R1419 VGND.n1771 VGND.n1770 12.8005
R1420 VGND.n1356 VGND.n1355 12.5161
R1421 VGND.n2040 VGND.n2039 12.1384
R1422 VGND.n1305 VGND.n1304 11.9309
R1423 VGND.n1294 VGND.n1266 11.2946
R1424 VGND.n1350 VGND.n1349 11.2946
R1425 VGND.n2208 VGND.n186 10.9091
R1426 VGND.n1806 VGND.n1805 10.8805
R1427 VGND.n406 VGND.n405 10.5983
R1428 VGND.n231 VGND.n230 10.5417
R1429 VGND.n1845 VGND.n1841 10.5417
R1430 VGND.n1344 VGND.n1343 10.5417
R1431 VGND.n1658 VGND.n1657 10.5417
R1432 VGND.n785 VGND.n784 10.5417
R1433 VGND.n1870 VGND.n1869 10.1652
R1434 VGND.n1869 VGND.n439 10.1652
R1435 VGND.n983 VGND.n982 10.1652
R1436 VGND.n1705 VGND.n1704 10.1652
R1437 VGND.n1753 VGND.n1750 10.1652
R1438 VGND.n791 VGND.n790 10.1652
R1439 VGND.n256 VGND.n240 9.88085
R1440 VGND.n1375 VGND.n1372 9.7205
R1441 VGND.n1169 VGND.n1168 9.7205
R1442 VGND.n24 VGND.n23 9.71789
R1443 VGND.n1577 VGND.n1576 9.71789
R1444 VGND.n1675 VGND.n1673 9.41227
R1445 VGND.n1618 VGND.n1617 9.41227
R1446 VGND.n717 VGND.n708 9.41227
R1447 VGND.n2311 VGND.n139 9.3031
R1448 VGND.n2138 VGND.n2133 9.3031
R1449 VGND.n1909 VGND.n356 9.3031
R1450 VGND.n394 VGND.n393 9.3031
R1451 VGND.n956 VGND.n954 9.3031
R1452 VGND.n895 VGND.n893 9.3031
R1453 VGND.n2496 VGND.n2495 9.3005
R1454 VGND.n2498 VGND.n2497 9.3005
R1455 VGND.n2499 VGND.n2487 9.3005
R1456 VGND.n2502 VGND.n2501 9.3005
R1457 VGND.n2503 VGND.n2485 9.3005
R1458 VGND.n2511 VGND.n2510 9.3005
R1459 VGND.n2514 VGND.n2513 9.3005
R1460 VGND.n2483 VGND.n59 9.3005
R1461 VGND.n2482 VGND.n2481 9.3005
R1462 VGND.n2480 VGND.n62 9.3005
R1463 VGND.n2479 VGND.n2478 9.3005
R1464 VGND.n2475 VGND.n63 9.3005
R1465 VGND.n2318 VGND.n139 9.3005
R1466 VGND.n2314 VGND.n139 9.3005
R1467 VGND.n2331 VGND.n2330 9.3005
R1468 VGND.n2333 VGND.n2332 9.3005
R1469 VGND.n2334 VGND.n135 9.3005
R1470 VGND.n2338 VGND.n2337 9.3005
R1471 VGND.n2341 VGND.n2340 9.3005
R1472 VGND.n2343 VGND.n132 9.3005
R1473 VGND.n2345 VGND.n2344 9.3005
R1474 VGND.n2358 VGND.n2357 9.3005
R1475 VGND.n2360 VGND.n2359 9.3005
R1476 VGND.n2362 VGND.n2361 9.3005
R1477 VGND.n2363 VGND.n121 9.3005
R1478 VGND.n2366 VGND.n2365 9.3005
R1479 VGND.n2367 VGND.n120 9.3005
R1480 VGND.n2369 VGND.n2368 9.3005
R1481 VGND.n2370 VGND.n119 9.3005
R1482 VGND.n2373 VGND.n2372 9.3005
R1483 VGND.n2375 VGND.n2374 9.3005
R1484 VGND.n2377 VGND.n2376 9.3005
R1485 VGND.n2379 VGND.n2378 9.3005
R1486 VGND.n2380 VGND.n2379 9.3005
R1487 VGND.n2389 VGND.n102 9.3005
R1488 VGND.n2389 VGND.n2388 9.3005
R1489 VGND.n2391 VGND.n101 9.3005
R1490 VGND.n2394 VGND.n2393 9.3005
R1491 VGND.n2395 VGND.n100 9.3005
R1492 VGND.n2397 VGND.n2396 9.3005
R1493 VGND.n2398 VGND.n99 9.3005
R1494 VGND.n2400 VGND.n2399 9.3005
R1495 VGND.n2402 VGND.n2401 9.3005
R1496 VGND.n2403 VGND.n97 9.3005
R1497 VGND.n2406 VGND.n2405 9.3005
R1498 VGND.n2408 VGND.n2407 9.3005
R1499 VGND.n2416 VGND.n2415 9.3005
R1500 VGND.n2413 VGND.n2412 9.3005
R1501 VGND.n2425 VGND.n83 9.3005
R1502 VGND.n2427 VGND.n2426 9.3005
R1503 VGND.n2428 VGND.n82 9.3005
R1504 VGND.n2430 VGND.n2429 9.3005
R1505 VGND.n2432 VGND.n2431 9.3005
R1506 VGND.n2433 VGND.n80 9.3005
R1507 VGND.n2436 VGND.n2435 9.3005
R1508 VGND.n2438 VGND.n2437 9.3005
R1509 VGND.n2440 VGND.n2439 9.3005
R1510 VGND.n2442 VGND.n2441 9.3005
R1511 VGND.n2445 VGND.n2444 9.3005
R1512 VGND.n2446 VGND.n76 9.3005
R1513 VGND.n2452 VGND.n2451 9.3005
R1514 VGND.n2454 VGND.n2453 9.3005
R1515 VGND.n70 VGND.n69 9.3005
R1516 VGND.n2463 VGND.n2462 9.3005
R1517 VGND.n2464 VGND.n68 9.3005
R1518 VGND.n2466 VGND.n2465 9.3005
R1519 VGND.n2468 VGND.n2467 9.3005
R1520 VGND.n2469 VGND.n66 9.3005
R1521 VGND.n2471 VGND.n2470 9.3005
R1522 VGND.n2473 VGND.n2472 9.3005
R1523 VGND.n2278 VGND.n2277 9.3005
R1524 VGND.n2275 VGND.n2274 9.3005
R1525 VGND.n2273 VGND.n163 9.3005
R1526 VGND.n2272 VGND.n2271 9.3005
R1527 VGND.n2270 VGND.n2269 9.3005
R1528 VGND.n2268 VGND.n165 9.3005
R1529 VGND.n2266 VGND.n2265 9.3005
R1530 VGND.n2276 VGND.n161 9.3005
R1531 VGND.n2283 VGND.n2282 9.3005
R1532 VGND.n2284 VGND.n160 9.3005
R1533 VGND.n2286 VGND.n2285 9.3005
R1534 VGND.n2289 VGND.n153 9.3005
R1535 VGND.n2292 VGND.n2291 9.3005
R1536 VGND.n224 VGND.n223 9.3005
R1537 VGND.n258 VGND.n240 9.3005
R1538 VGND.n252 VGND.n251 9.3005
R1539 VGND.n250 VGND.n249 9.3005
R1540 VGND.n254 VGND.n242 9.3005
R1541 VGND.n257 VGND.n256 9.3005
R1542 VGND.n266 VGND.n265 9.3005
R1543 VGND.n268 VGND.n267 9.3005
R1544 VGND.n238 VGND.n211 9.3005
R1545 VGND.n237 VGND.n215 9.3005
R1546 VGND.n236 VGND.n235 9.3005
R1547 VGND.n234 VGND.n216 9.3005
R1548 VGND.n233 VGND.n232 9.3005
R1549 VGND.n231 VGND.n217 9.3005
R1550 VGND.n230 VGND.n219 9.3005
R1551 VGND.n229 VGND.n228 9.3005
R1552 VGND.n227 VGND.n221 9.3005
R1553 VGND.n226 VGND.n225 9.3005
R1554 VGND.n222 VGND.n157 9.3005
R1555 VGND.n2290 VGND.n154 9.3005
R1556 VGND.n2264 VGND.n166 9.3005
R1557 VGND.n2253 VGND.n2252 9.3005
R1558 VGND.n2255 VGND.n2254 9.3005
R1559 VGND.n2250 VGND.n2249 9.3005
R1560 VGND.n2248 VGND.n2247 9.3005
R1561 VGND.n2143 VGND.n2133 9.3005
R1562 VGND.n2145 VGND.n2133 9.3005
R1563 VGND.n2157 VGND.n2156 9.3005
R1564 VGND.n2159 VGND.n2158 9.3005
R1565 VGND.n2160 VGND.n2129 9.3005
R1566 VGND.n2164 VGND.n2163 9.3005
R1567 VGND.n2167 VGND.n2166 9.3005
R1568 VGND.n2169 VGND.n2126 9.3005
R1569 VGND.n2171 VGND.n2170 9.3005
R1570 VGND.n2184 VGND.n2183 9.3005
R1571 VGND.n2186 VGND.n2185 9.3005
R1572 VGND.n2188 VGND.n2187 9.3005
R1573 VGND.n2189 VGND.n199 9.3005
R1574 VGND.n2192 VGND.n2191 9.3005
R1575 VGND.n2193 VGND.n198 9.3005
R1576 VGND.n2195 VGND.n2194 9.3005
R1577 VGND.n2196 VGND.n197 9.3005
R1578 VGND.n2199 VGND.n2198 9.3005
R1579 VGND.n2201 VGND.n2200 9.3005
R1580 VGND.n2204 VGND.n2203 9.3005
R1581 VGND.n2206 VGND.n2205 9.3005
R1582 VGND.n2209 VGND.n2208 9.3005
R1583 VGND.n2214 VGND.n2213 9.3005
R1584 VGND.n2224 VGND.n2223 9.3005
R1585 VGND.n2225 VGND.n183 9.3005
R1586 VGND.n2231 VGND.n2230 9.3005
R1587 VGND.n2232 VGND.n182 9.3005
R1588 VGND.n2234 VGND.n2233 9.3005
R1589 VGND.n2236 VGND.n181 9.3005
R1590 VGND.n2238 VGND.n2237 9.3005
R1591 VGND.n2240 VGND.n2239 9.3005
R1592 VGND.n2241 VGND.n179 9.3005
R1593 VGND.n2243 VGND.n2242 9.3005
R1594 VGND.n2245 VGND.n2244 9.3005
R1595 VGND.n2036 VGND.n301 9.3005
R1596 VGND.n2035 VGND.n2034 9.3005
R1597 VGND.n2031 VGND.n302 9.3005
R1598 VGND.n2030 VGND.n2029 9.3005
R1599 VGND.n2028 VGND.n2027 9.3005
R1600 VGND.n2026 VGND.n304 9.3005
R1601 VGND.n2025 VGND.n2024 9.3005
R1602 VGND.n2023 VGND.n305 9.3005
R1603 VGND.n2011 VGND.n2010 9.3005
R1604 VGND.n2014 VGND.n2013 9.3005
R1605 VGND.n2038 VGND.n2037 9.3005
R1606 VGND.n2041 VGND.n2040 9.3005
R1607 VGND.n2043 VGND.n295 9.3005
R1608 VGND.n2046 VGND.n2045 9.3005
R1609 VGND.n288 VGND.n287 9.3005
R1610 VGND.n2059 VGND.n2058 9.3005
R1611 VGND.n2061 VGND.n286 9.3005
R1612 VGND.n2065 VGND.n2064 9.3005
R1613 VGND.n2066 VGND.n285 9.3005
R1614 VGND.n2067 VGND 9.3005
R1615 VGND.n2071 VGND.n2070 9.3005
R1616 VGND.n2073 VGND.n2072 9.3005
R1617 VGND.n2074 VGND.n282 9.3005
R1618 VGND.n2077 VGND.n2076 9.3005
R1619 VGND.n2078 VGND.n281 9.3005
R1620 VGND.n2080 VGND.n2079 9.3005
R1621 VGND.n2081 VGND.n279 9.3005
R1622 VGND.n2110 VGND.n2109 9.3005
R1623 VGND.n2108 VGND.n2107 9.3005
R1624 VGND.n2100 VGND.n2083 9.3005
R1625 VGND.n2099 VGND.n2098 9.3005
R1626 VGND.n2097 VGND.n2085 9.3005
R1627 VGND.n2095 VGND.n2094 9.3005
R1628 VGND.n2093 VGND.n2092 9.3005
R1629 VGND.n1916 VGND.n356 9.3005
R1630 VGND.n1912 VGND.n356 9.3005
R1631 VGND.n1929 VGND.n1928 9.3005
R1632 VGND.n1931 VGND.n1930 9.3005
R1633 VGND.n1932 VGND.n352 9.3005
R1634 VGND.n1934 VGND.n1933 9.3005
R1635 VGND.n1939 VGND.n1938 9.3005
R1636 VGND.n1945 VGND.n1944 9.3005
R1637 VGND.n1947 VGND.n1946 9.3005
R1638 VGND.n1956 VGND.n1955 9.3005
R1639 VGND.n1958 VGND.n1957 9.3005
R1640 VGND.n1960 VGND.n1959 9.3005
R1641 VGND.n1961 VGND.n341 9.3005
R1642 VGND.n1964 VGND.n1963 9.3005
R1643 VGND.n1965 VGND.n340 9.3005
R1644 VGND.n1967 VGND.n1966 9.3005
R1645 VGND.n1968 VGND.n339 9.3005
R1646 VGND.n1971 VGND.n1970 9.3005
R1647 VGND.n1973 VGND.n1972 9.3005
R1648 VGND.n1975 VGND.n1974 9.3005
R1649 VGND.n1977 VGND.n1976 9.3005
R1650 VGND.n1978 VGND.n1977 9.3005
R1651 VGND.n1987 VGND.n323 9.3005
R1652 VGND.n1987 VGND.n1986 9.3005
R1653 VGND.n1989 VGND.n322 9.3005
R1654 VGND.n1992 VGND.n1991 9.3005
R1655 VGND.n1993 VGND.n321 9.3005
R1656 VGND.n1995 VGND.n1994 9.3005
R1657 VGND.n1996 VGND.n320 9.3005
R1658 VGND.n1998 VGND.n1997 9.3005
R1659 VGND.n2000 VGND.n1999 9.3005
R1660 VGND.n2001 VGND.n318 9.3005
R1661 VGND.n2004 VGND.n2003 9.3005
R1662 VGND.n2006 VGND.n2005 9.3005
R1663 VGND.n1869 VGND.n1868 9.3005
R1664 VGND.n1857 VGND.n1856 9.3005
R1665 VGND.n1854 VGND.n1853 9.3005
R1666 VGND.n1821 VGND.n1820 9.3005
R1667 VGND.n1812 VGND.n1811 9.3005
R1668 VGND.n489 VGND.n486 9.3005
R1669 VGND.n1803 VGND.n1802 9.3005
R1670 VGND.n521 VGND.n490 9.3005
R1671 VGND.n525 VGND.n524 9.3005
R1672 VGND.n514 VGND.n513 9.3005
R1673 VGND.n531 VGND.n530 9.3005
R1674 VGND.n533 VGND.n511 9.3005
R1675 VGND.n536 VGND.n535 9.3005
R1676 VGND.n538 VGND.n537 9.3005
R1677 VGND.n539 VGND.n507 9.3005
R1678 VGND.n542 VGND.n541 9.3005
R1679 VGND.n544 VGND.n543 9.3005
R1680 VGND.n547 VGND.n505 9.3005
R1681 VGND.n552 VGND.n551 9.3005
R1682 VGND.n553 VGND.n504 9.3005
R1683 VGND.n555 VGND.n554 9.3005
R1684 VGND.n556 VGND.n500 9.3005
R1685 VGND.n587 VGND.n586 9.3005
R1686 VGND.n585 VGND.n584 9.3005
R1687 VGND.n577 VGND.n576 9.3005
R1688 VGND.n574 VGND.n573 9.3005
R1689 VGND.n572 VGND.n571 9.3005
R1690 VGND.n570 VGND.n561 9.3005
R1691 VGND.n567 VGND.n566 9.3005
R1692 VGND.n1809 VGND.n1808 9.3005
R1693 VGND.n1810 VGND.n485 9.3005
R1694 VGND.n1816 VGND.n483 9.3005
R1695 VGND.n1818 VGND.n1817 9.3005
R1696 VGND.n1819 VGND.n481 9.3005
R1697 VGND.n1822 VGND.n480 9.3005
R1698 VGND.n1823 VGND.n477 9.3005
R1699 VGND.n1825 VGND.n1824 9.3005
R1700 VGND.n468 VGND.n466 9.3005
R1701 VGND.n1834 VGND.n1833 9.3005
R1702 VGND.n1837 VGND.n1836 9.3005
R1703 VGND.n1838 VGND.n463 9.3005
R1704 VGND.n1840 VGND.n1839 9.3005
R1705 VGND.n1841 VGND.n460 9.3005
R1706 VGND.n1846 VGND.n1845 9.3005
R1707 VGND.n1847 VGND.n459 9.3005
R1708 VGND.n1849 VGND.n1848 9.3005
R1709 VGND.n1852 VGND.n455 9.3005
R1710 VGND.n1855 VGND.n454 9.3005
R1711 VGND.n1861 VGND.n1860 9.3005
R1712 VGND.n451 VGND.n439 9.3005
R1713 VGND.n1870 VGND.n437 9.3005
R1714 VGND.n1872 VGND.n1871 9.3005
R1715 VGND.n1873 VGND.n435 9.3005
R1716 VGND.n1875 VGND.n1874 9.3005
R1717 VGND.n1876 VGND.n433 9.3005
R1718 VGND.n1879 VGND.n1878 9.3005
R1719 VGND.n1880 VGND.n432 9.3005
R1720 VGND.n1882 VGND.n1881 9.3005
R1721 VGND.n1883 VGND.n430 9.3005
R1722 VGND.n1886 VGND.n1885 9.3005
R1723 VGND.n1887 VGND.n429 9.3005
R1724 VGND.n1889 VGND.n1888 9.3005
R1725 VGND.n1893 VGND.n1892 9.3005
R1726 VGND.n394 VGND.n385 9.3005
R1727 VGND.n395 VGND.n394 9.3005
R1728 VGND.n403 VGND.n381 9.3005
R1729 VGND.n405 VGND.n404 9.3005
R1730 VGND.n408 VGND.n407 9.3005
R1731 VGND.n410 VGND.n409 9.3005
R1732 VGND.n411 VGND.n379 9.3005
R1733 VGND.n414 VGND.n413 9.3005
R1734 VGND.n415 VGND.n378 9.3005
R1735 VGND.n417 VGND.n416 9.3005
R1736 VGND.n418 VGND.n376 9.3005
R1737 VGND.n421 VGND.n420 9.3005
R1738 VGND.n422 VGND.n375 9.3005
R1739 VGND.n424 VGND.n423 9.3005
R1740 VGND.n426 VGND.n370 9.3005
R1741 VGND.n428 VGND.n371 9.3005
R1742 VGND.n956 VGND.n938 9.3005
R1743 VGND.n956 VGND.n937 9.3005
R1744 VGND.n957 VGND.n935 9.3005
R1745 VGND.n962 VGND.n961 9.3005
R1746 VGND.n965 VGND.n964 9.3005
R1747 VGND.n966 VGND.n931 9.3005
R1748 VGND.n969 VGND.n968 9.3005
R1749 VGND.n971 VGND.n970 9.3005
R1750 VGND.n928 VGND.n927 9.3005
R1751 VGND.n978 VGND.n977 9.3005
R1752 VGND.n979 VGND.n926 9.3005
R1753 VGND.n981 VGND.n980 9.3005
R1754 VGND.n983 VGND.n920 9.3005
R1755 VGND.n985 VGND.n921 9.3005
R1756 VGND.n1317 VGND.n1316 9.3005
R1757 VGND.n1315 VGND.n1314 9.3005
R1758 VGND.n1313 VGND.n1312 9.3005
R1759 VGND.n1310 VGND.n989 9.3005
R1760 VGND.n1308 VGND.n1307 9.3005
R1761 VGND.n1306 VGND.n1305 9.3005
R1762 VGND.n1302 VGND.n1301 9.3005
R1763 VGND.n1300 VGND.n1299 9.3005
R1764 VGND.n1295 VGND.n994 9.3005
R1765 VGND.n1294 VGND.n1293 9.3005
R1766 VGND.n1292 VGND.n1291 9.3005
R1767 VGND.n1290 VGND.n1267 9.3005
R1768 VGND.n1287 VGND.n1286 9.3005
R1769 VGND.n1276 VGND.n1274 9.3005
R1770 VGND.n1271 VGND.n643 9.3005
R1771 VGND.n1669 VGND.n642 9.3005
R1772 VGND.n1671 VGND.n1670 9.3005
R1773 VGND.n1672 VGND.n640 9.3005
R1774 VGND.n1676 VGND.n1675 9.3005
R1775 VGND.n1677 VGND.n639 9.3005
R1776 VGND.n1679 VGND.n1678 9.3005
R1777 VGND.n1680 VGND.n638 9.3005
R1778 VGND.n1683 VGND.n1682 9.3005
R1779 VGND.n1684 VGND.n637 9.3005
R1780 VGND.n1687 VGND.n1685 9.3005
R1781 VGND.n1689 VGND.n1688 9.3005
R1782 VGND.n1691 VGND.n1690 9.3005
R1783 VGND.n1693 VGND.n1692 9.3005
R1784 VGND.n631 VGND.n622 9.3005
R1785 VGND.n1703 VGND.n1702 9.3005
R1786 VGND.n1705 VGND.n620 9.3005
R1787 VGND.n1708 VGND.n1707 9.3005
R1788 VGND.n1709 VGND.n618 9.3005
R1789 VGND.n1714 VGND.n1713 9.3005
R1790 VGND.n1716 VGND.n1715 9.3005
R1791 VGND.n1719 VGND.n615 9.3005
R1792 VGND.n1722 VGND.n1721 9.3005
R1793 VGND.n1720 VGND.n614 9.3005
R1794 VGND.n1728 VGND.n609 9.3005
R1795 VGND.n1737 VGND.n1736 9.3005
R1796 VGND.n1738 VGND.n608 9.3005
R1797 VGND.n1740 VGND.n1739 9.3005
R1798 VGND.n1742 VGND.n1741 9.3005
R1799 VGND.n1743 VGND.n604 9.3005
R1800 VGND.n1745 VGND.n1744 9.3005
R1801 VGND.n1746 VGND.n603 9.3005
R1802 VGND.n1748 VGND.n1747 9.3005
R1803 VGND.n1749 VGND.n601 9.3005
R1804 VGND.n1754 VGND.n1753 9.3005
R1805 VGND.n1755 VGND.n600 9.3005
R1806 VGND.n1757 VGND.n1756 9.3005
R1807 VGND.n1758 VGND.n598 9.3005
R1808 VGND.n1788 VGND.n1787 9.3005
R1809 VGND.n1784 VGND.n1783 9.3005
R1810 VGND.n1776 VGND.n1775 9.3005
R1811 VGND.n1773 VGND.n1761 9.3005
R1812 VGND.n1771 VGND.n1765 9.3005
R1813 VGND.n895 VGND.n884 9.3005
R1814 VGND.n895 VGND.n883 9.3005
R1815 VGND.n1363 VGND.n1362 9.3005
R1816 VGND.n1360 VGND.n880 9.3005
R1817 VGND.n1359 VGND.n1358 9.3005
R1818 VGND.n1357 VGND.n1356 9.3005
R1819 VGND.n1355 VGND.n899 9.3005
R1820 VGND.n1354 VGND.n1353 9.3005
R1821 VGND.n1352 VGND.n1351 9.3005
R1822 VGND.n1350 VGND.n903 9.3005
R1823 VGND.n1349 VGND.n904 9.3005
R1824 VGND.n1348 VGND.n1347 9.3005
R1825 VGND.n1346 VGND.n906 9.3005
R1826 VGND.n1345 VGND.n1344 9.3005
R1827 VGND.n1343 VGND.n909 9.3005
R1828 VGND.n1342 VGND.n1341 9.3005
R1829 VGND.n912 VGND.n910 9.3005
R1830 VGND.n1003 VGND.n1002 9.3005
R1831 VGND.n1005 VGND.n1004 9.3005
R1832 VGND.n1007 VGND.n1006 9.3005
R1833 VGND.n1008 VGND.n1001 9.3005
R1834 VGND.n1010 VGND.n1009 9.3005
R1835 VGND.n1011 VGND.n998 9.3005
R1836 VGND.n1016 VGND.n1015 9.3005
R1837 VGND.n1017 VGND.n996 9.3005
R1838 VGND.n1023 VGND.n1022 9.3005
R1839 VGND.n1021 VGND.n1020 9.3005
R1840 VGND.n1019 VGND.n1018 9.3005
R1841 VGND.n656 VGND.n654 9.3005
R1842 VGND.n1659 VGND.n1658 9.3005
R1843 VGND.n1657 VGND.n658 9.3005
R1844 VGND.n1656 VGND.n1655 9.3005
R1845 VGND.n1654 VGND.n660 9.3005
R1846 VGND.n1653 VGND.n1652 9.3005
R1847 VGND.n1651 VGND.n668 9.3005
R1848 VGND.n1650 VGND.n1649 9.3005
R1849 VGND.n1648 VGND.n1647 9.3005
R1850 VGND.n1644 VGND.n670 9.3005
R1851 VGND.n1643 VGND.n1642 9.3005
R1852 VGND.n1641 VGND.n673 9.3005
R1853 VGND.n1640 VGND.n1639 9.3005
R1854 VGND.n1638 VGND.n674 9.3005
R1855 VGND.n1636 VGND.n1635 9.3005
R1856 VGND.n687 VGND.n676 9.3005
R1857 VGND.n691 VGND.n690 9.3005
R1858 VGND.n1626 VGND.n1625 9.3005
R1859 VGND.n1624 VGND.n682 9.3005
R1860 VGND.n1622 VGND.n1621 9.3005
R1861 VGND.n1620 VGND.n692 9.3005
R1862 VGND.n1619 VGND.n1618 9.3005
R1863 VGND.n1616 VGND.n693 9.3005
R1864 VGND.n1615 VGND.n1614 9.3005
R1865 VGND.n1613 VGND.n696 9.3005
R1866 VGND.n1612 VGND.n1611 9.3005
R1867 VGND.n1610 VGND.n1609 9.3005
R1868 VGND.n1608 VGND.n1607 9.3005
R1869 VGND.n1604 VGND.n1603 9.3005
R1870 VGND.n709 VGND.n699 9.3005
R1871 VGND.n717 VGND.n716 9.3005
R1872 VGND.n719 VGND.n704 9.3005
R1873 VGND.n793 VGND.n792 9.3005
R1874 VGND.n791 VGND.n705 9.3005
R1875 VGND.n789 VGND.n788 9.3005
R1876 VGND.n787 VGND.n721 9.3005
R1877 VGND.n786 VGND.n785 9.3005
R1878 VGND.n784 VGND.n722 9.3005
R1879 VGND.n782 VGND.n781 9.3005
R1880 VGND.n780 VGND.n725 9.3005
R1881 VGND.n779 VGND.n778 9.3005
R1882 VGND.n776 VGND.n726 9.3005
R1883 VGND.n772 VGND.n771 9.3005
R1884 VGND.n737 VGND.n728 9.3005
R1885 VGND.n745 VGND.n744 9.3005
R1886 VGND.n746 VGND.n733 9.3005
R1887 VGND.n762 VGND.n761 9.3005
R1888 VGND.n760 VGND.n734 9.3005
R1889 VGND.n759 VGND.n758 9.3005
R1890 VGND.n757 VGND.n756 9.3005
R1891 VGND.n754 VGND.n749 9.3005
R1892 VGND.n1580 VGND.n1579 9.3005
R1893 VGND.n1582 VGND.n1581 9.3005
R1894 VGND.n1378 VGND.n1377 9.3005
R1895 VGND.n1389 VGND.n1388 9.3005
R1896 VGND.n1391 VGND.n1390 9.3005
R1897 VGND.n1392 VGND.n866 9.3005
R1898 VGND.n1394 VGND.n1393 9.3005
R1899 VGND.n1395 VGND.n863 9.3005
R1900 VGND.n1397 VGND.n1396 9.3005
R1901 VGND.n1398 VGND.n862 9.3005
R1902 VGND.n1400 VGND.n1399 9.3005
R1903 VGND.n1402 VGND.n861 9.3005
R1904 VGND.n1406 VGND.n1405 9.3005
R1905 VGND.n1407 VGND.n860 9.3005
R1906 VGND.n1409 VGND.n1408 9.3005
R1907 VGND.n1410 VGND.n859 9.3005
R1908 VGND.n1412 VGND.n1411 9.3005
R1909 VGND.n1414 VGND.n851 9.3005
R1910 VGND.n1427 VGND.n1426 9.3005
R1911 VGND.n1429 VGND.n850 9.3005
R1912 VGND.n1433 VGND.n1432 9.3005
R1913 VGND.n1436 VGND.n1435 9.3005
R1914 VGND.n1438 VGND.n1437 9.3005
R1915 VGND.n1439 VGND.n846 9.3005
R1916 VGND.n1443 VGND.n1442 9.3005
R1917 VGND.n1445 VGND.n1444 9.3005
R1918 VGND.n1449 VGND.n1448 9.3005
R1919 VGND.n1454 VGND.n838 9.3005
R1920 VGND.n839 VGND.n838 9.3005
R1921 VGND.n1463 VGND.n838 9.3005
R1922 VGND.n1465 VGND.n1464 9.3005
R1923 VGND.n1467 VGND.n837 9.3005
R1924 VGND.n1469 VGND.n1468 9.3005
R1925 VGND.n1470 VGND.n836 9.3005
R1926 VGND.n1472 VGND.n1471 9.3005
R1927 VGND.n1474 VGND.n835 9.3005
R1928 VGND.n1478 VGND.n1477 9.3005
R1929 VGND.n1481 VGND.n1480 9.3005
R1930 VGND.n1487 VGND.n1486 9.3005
R1931 VGND.n1485 VGND.n1484 9.3005
R1932 VGND.n1496 VGND.n824 9.3005
R1933 VGND.n1498 VGND.n1497 9.3005
R1934 VGND.n1500 VGND.n823 9.3005
R1935 VGND.n1504 VGND.n1503 9.3005
R1936 VGND.n1505 VGND.n822 9.3005
R1937 VGND.n1507 VGND.n1506 9.3005
R1938 VGND.n1510 VGND.n1509 9.3005
R1939 VGND.n1511 VGND.n820 9.3005
R1940 VGND.n1513 VGND.n1512 9.3005
R1941 VGND.n1516 VGND.n1515 9.3005
R1942 VGND.n1517 VGND.n819 9.3005
R1943 VGND.n1519 VGND.n1518 9.3005
R1944 VGND.n1521 VGND.n1520 9.3005
R1945 VGND.n815 VGND.n814 9.3005
R1946 VGND.n1535 VGND.n1534 9.3005
R1947 VGND.n1541 VGND.n1540 9.3005
R1948 VGND.n1542 VGND.n810 9.3005
R1949 VGND.n1544 VGND.n1543 9.3005
R1950 VGND.n1546 VGND.n809 9.3005
R1951 VGND.n1548 VGND.n1547 9.3005
R1952 VGND.n1549 VGND.n808 9.3005
R1953 VGND.n1551 VGND.n1550 9.3005
R1954 VGND.n1553 VGND.n807 9.3005
R1955 VGND.n1557 VGND.n1556 9.3005
R1956 VGND.n1560 VGND.n804 9.3005
R1957 VGND.n1569 VGND.n1568 9.3005
R1958 VGND.n1571 VGND.n803 9.3005
R1959 VGND.n1590 VGND.n1589 9.3005
R1960 VGND.n1588 VGND.n1587 9.3005
R1961 VGND.n1586 VGND.n1572 9.3005
R1962 VGND.n1585 VGND.n1584 9.3005
R1963 VGND.n1583 VGND.n1573 9.3005
R1964 VGND.n1441 VGND.n1440 9.3005
R1965 VGND.n1166 VGND.n1164 9.3005
R1966 VGND.n1179 VGND.n1178 9.3005
R1967 VGND.n1225 VGND.n1224 9.3005
R1968 VGND.n1222 VGND.n1162 9.3005
R1969 VGND.n1219 VGND.n1218 9.3005
R1970 VGND.n1217 VGND.n1180 9.3005
R1971 VGND.n1216 VGND.n1215 9.3005
R1972 VGND.n1214 VGND.n1181 9.3005
R1973 VGND.n1213 VGND.n1212 9.3005
R1974 VGND.n1211 VGND.n1183 9.3005
R1975 VGND.n1210 VGND.n1209 9.3005
R1976 VGND.n1186 VGND.n1184 9.3005
R1977 VGND.n1204 VGND.n1203 9.3005
R1978 VGND.n1202 VGND.n1188 9.3005
R1979 VGND.n1200 VGND.n1199 9.3005
R1980 VGND.n1198 VGND.n1197 9.3005
R1981 VGND.n1192 VGND.n1033 9.3005
R1982 VGND.n1244 VGND.n1032 9.3005
R1983 VGND.n1246 VGND.n1245 9.3005
R1984 VGND.n1247 VGND.n1031 9.3005
R1985 VGND.n1249 VGND.n1248 9.3005
R1986 VGND.n1251 VGND.n1250 9.3005
R1987 VGND.n1252 VGND.n1029 9.3005
R1988 VGND.n1254 VGND.n1253 9.3005
R1989 VGND.n1256 VGND.n1255 9.3005
R1990 VGND.n1257 VGND.n1027 9.3005
R1991 VGND.n1050 VGND.n1026 9.3005
R1992 VGND.n1055 VGND.n1054 9.3005
R1993 VGND.n1057 VGND.n1047 9.3005
R1994 VGND.n1065 VGND.n1064 9.3005
R1995 VGND.n1067 VGND.n1045 9.3005
R1996 VGND.n1153 VGND.n1152 9.3005
R1997 VGND.n1151 VGND.n1046 9.3005
R1998 VGND.n1150 VGND.n1149 9.3005
R1999 VGND.n1148 VGND.n1068 9.3005
R2000 VGND.n1147 VGND.n1146 9.3005
R2001 VGND.n1145 VGND.n1069 9.3005
R2002 VGND.n1143 VGND.n1142 9.3005
R2003 VGND.n1141 VGND.n1070 9.3005
R2004 VGND.n1140 VGND.n1139 9.3005
R2005 VGND.n1137 VGND 9.3005
R2006 VGND.n1136 VGND.n1135 9.3005
R2007 VGND.n1134 VGND.n1133 9.3005
R2008 VGND.n1132 VGND.n1131 9.3005
R2009 VGND.n1075 VGND.n1073 9.3005
R2010 VGND.n1123 VGND.n1122 9.3005
R2011 VGND.n1121 VGND.n1084 9.3005
R2012 VGND.n1120 VGND.n1119 9.3005
R2013 VGND.n1118 VGND.n1085 9.3005
R2014 VGND.n1117 VGND.n1116 9.3005
R2015 VGND.n1115 VGND.n1086 9.3005
R2016 VGND.n1114 VGND.n1113 9.3005
R2017 VGND.n1112 VGND.n1111 9.3005
R2018 VGND.n1110 VGND.n1109 9.3005
R2019 VGND.n1108 VGND.n1089 9.3005
R2020 VGND.n1107 VGND.n1106 9.3005
R2021 VGND.n1105 VGND.n1104 9.3005
R2022 VGND.n1100 VGND.n47 9.3005
R2023 VGND.n2533 VGND.n2532 9.3005
R2024 VGND.n2534 VGND.n45 9.3005
R2025 VGND.n2546 VGND.n2545 9.3005
R2026 VGND.n2535 VGND.n46 9.3005
R2027 VGND.n2540 VGND.n2539 9.3005
R2028 VGND.n2538 VGND.n0 9.3005
R2029 VGND.n2567 VGND.n2566 9.3005
R2030 VGND.n2565 VGND.n2563 9.3005
R2031 VGND.n2562 VGND.n1 9.3005
R2032 VGND.n2561 VGND.n2560 9.3005
R2033 VGND.n2558 VGND.n2 9.3005
R2034 VGND.n2557 VGND.n2556 9.3005
R2035 VGND.n2555 VGND.n3 9.3005
R2036 VGND.n12 VGND.n4 9.3005
R2037 VGND.n18 VGND.n17 9.3005
R2038 VGND.n19 VGND.n10 9.3005
R2039 VGND.n38 VGND.n37 9.3005
R2040 VGND.n35 VGND.n11 9.3005
R2041 VGND.n34 VGND.n33 9.3005
R2042 VGND.n32 VGND.n20 9.3005
R2043 VGND.n31 VGND.n30 9.3005
R2044 VGND.n29 VGND.n28 9.3005
R2045 VGND.n27 VGND.n26 9.3005
R2046 VGND.n1821 VGND.n481 9.12791
R2047 VGND.n1852 VGND.n1851 9.03579
R2048 VGND.n458 VGND.n457 9.03579
R2049 VGND.n1309 VGND.n1308 9.03579
R2050 VGND.n547 VGND.n546 8.9684
R2051 VGND.t183 VGND.t521 8.42962
R2052 VGND.t365 VGND.t793 8.42962
R2053 VGND.t802 VGND.t363 8.42962
R2054 VGND.n1742 VGND.n606 8.28285
R2055 VGND.n2558 VGND.n2557 8.23546
R2056 VGND.n2557 VGND.n3 8.23546
R2057 VGND.n12 VGND.n3 8.23546
R2058 VGND.n18 VGND.n12 8.23546
R2059 VGND.n19 VGND.n18 8.23546
R2060 VGND.n37 VGND.n19 8.23546
R2061 VGND.n35 VGND.n34 8.23546
R2062 VGND.n34 VGND.n20 8.23546
R2063 VGND.n1133 VGND.n1132 8.23546
R2064 VGND.n1132 VGND.n1073 8.23546
R2065 VGND.n1122 VGND.n1073 8.23546
R2066 VGND.n1122 VGND.n1121 8.23546
R2067 VGND.n1121 VGND.n1120 8.23546
R2068 VGND.n1120 VGND.n1085 8.23546
R2069 VGND.n1116 VGND.n1115 8.23546
R2070 VGND.n1115 VGND.n1114 8.23546
R2071 VGND.n1152 VGND.n1067 8.23546
R2072 VGND.n1152 VGND.n1151 8.23546
R2073 VGND.n1151 VGND.n1150 8.23546
R2074 VGND.n1150 VGND.n1068 8.23546
R2075 VGND.n1146 VGND.n1068 8.23546
R2076 VGND.n1146 VGND.n1145 8.23546
R2077 VGND.n1143 VGND.n1070 8.23546
R2078 VGND.n1139 VGND.n1070 8.23546
R2079 VGND.n2376 VGND.n2375 8.23546
R2080 VGND.n2478 VGND.n62 8.23546
R2081 VGND.n2482 VGND.n62 8.23546
R2082 VGND.n2483 VGND.n2482 8.23546
R2083 VGND.n2511 VGND.n2485 8.23546
R2084 VGND.n2076 VGND.n281 8.23546
R2085 VGND.n2080 VGND.n281 8.23546
R2086 VGND.n2045 VGND.n287 8.23546
R2087 VGND.n2059 VGND.n287 8.23546
R2088 VGND.n2067 VGND.n285 8.23546
R2089 VGND.n2070 VGND.n2067 8.23546
R2090 VGND.n1974 VGND.n1973 8.23546
R2091 VGND.n555 VGND.n504 8.23546
R2092 VGND.n556 VGND.n555 8.23546
R2093 VGND.n586 VGND.n585 8.23546
R2094 VGND.n524 VGND.n521 8.23546
R2095 VGND.n531 VGND.n513 8.23546
R2096 VGND.n535 VGND.n533 8.23546
R2097 VGND.n539 VGND.n538 8.23546
R2098 VGND.n418 VGND.n417 8.23546
R2099 VGND.n420 VGND.n418 8.23546
R2100 VGND.n424 VGND.n375 8.23546
R2101 VGND.n1889 VGND.n429 8.23546
R2102 VGND.n1885 VGND.n429 8.23546
R2103 VGND.n1883 VGND.n1882 8.23546
R2104 VGND.n1882 VGND.n432 8.23546
R2105 VGND.n1878 VGND.n432 8.23546
R2106 VGND.n1876 VGND.n1875 8.23546
R2107 VGND.n1875 VGND.n435 8.23546
R2108 VGND.n1644 VGND.n1643 8.23546
R2109 VGND.n1643 VGND.n673 8.23546
R2110 VGND.n1639 VGND.n673 8.23546
R2111 VGND.n1639 VGND.n1638 8.23546
R2112 VGND.n1636 VGND.n676 8.23546
R2113 VGND.n1625 VGND.n691 8.23546
R2114 VGND.n1625 VGND.n1624 8.23546
R2115 VGND.n1199 VGND.n1198 8.23546
R2116 VGND.n1198 VGND.n1192 8.23546
R2117 VGND.n1192 VGND.n1032 8.23546
R2118 VGND.n1246 VGND.n1032 8.23546
R2119 VGND.n1247 VGND.n1246 8.23546
R2120 VGND.n1248 VGND.n1247 8.23546
R2121 VGND.n1252 VGND.n1251 8.23546
R2122 VGND.n1253 VGND.n1252 8.23546
R2123 VGND.n2061 VGND.n2060 8.14595
R2124 VGND.n2513 VGND.n2484 8.05644
R2125 VGND.n1845 VGND.n1844 7.90638
R2126 VGND.n1688 VGND.n636 7.90638
R2127 VGND.n783 VGND.n782 7.90638
R2128 VGND.n426 VGND.n425 7.78791
R2129 VGND.n1646 VGND.n672 7.72113
R2130 VGND.n2559 VGND.n2558 7.6984
R2131 VGND.n21 VGND.n20 7.6984
R2132 VGND.n1133 VGND.n1071 7.6984
R2133 VGND.n1114 VGND.n1088 7.6984
R2134 VGND.n1067 VGND.n1066 7.6984
R2135 VGND.n1139 VGND.n1138 7.6984
R2136 VGND.n2439 VGND.n77 7.6984
R2137 VGND.n2478 VGND.n2477 7.6984
R2138 VGND.n2076 VGND.n2075 7.6984
R2139 VGND.n2064 VGND.n2062 7.6984
R2140 VGND.n551 VGND.n548 7.6984
R2141 VGND.n1804 VGND.n1803 7.6984
R2142 VGND.n1803 VGND.n488 7.6984
R2143 VGND.n541 VGND.n506 7.6984
R2144 VGND.n427 VGND.n426 7.6984
R2145 VGND.n436 VGND.n435 7.6984
R2146 VGND.n1645 VGND.n1644 7.6984
R2147 VGND.n1624 VGND.n1623 7.6984
R2148 VGND.n1199 VGND.n1191 7.6984
R2149 VGND.n1253 VGND.n1028 7.6984
R2150 VGND.n738 VGND.n736 7.6005
R2151 VGND.n1884 VGND.n1883 7.51938
R2152 VGND.n2070 VGND.n2069 7.34036
R2153 VGND.n1637 VGND.n1636 7.34036
R2154 VGND.n557 VGND.n556 7.25085
R2155 VGND.n1891 VGND.n1890 7.25085
R2156 VGND.n550 VGND.n504 7.16134
R2157 VGND.n2439 VGND.n2438 7.11268
R2158 VGND.n2038 VGND.n301 7.11268
R2159 VGND.n2513 VGND.n2512 6.98232
R2160 VGND.n2081 VGND.n2080 6.88949
R2161 VGND.n417 VGND.n378 6.88949
R2162 VGND.n524 VGND.n523 6.62428
R2163 VGND.n2389 VGND.n104 6.61527
R2164 VGND.n1987 VGND.n325 6.61527
R2165 VGND.n2379 VGND.n104 6.57117
R2166 VGND.n1977 VGND.n325 6.57117
R2167 VGND.n934 VGND.n933 6.57117
R2168 VGND.n960 VGND.n934 6.57117
R2169 VGND.n585 VGND.n558 6.53477
R2170 VGND.n1617 VGND.n1616 6.4005
R2171 VGND.n708 VGND.n699 6.4005
R2172 VGND.n2533 VGND.n47 6.26433
R2173 VGND.n2534 VGND.n2533 6.26433
R2174 VGND.n1817 VGND.n1816 6.26433
R2175 VGND.n966 VGND.n965 6.26433
R2176 VGND.n1360 VGND.n1359 6.26433
R2177 VGND.n1432 VGND.n1429 6.26433
R2178 VGND.n1405 VGND.n1402 6.26433
R2179 VGND.n1448 VGND.n1445 6.26433
R2180 VGND.n1477 VGND.n1474 6.26433
R2181 VGND.n1503 VGND.n1500 6.26433
R2182 VGND.n1519 VGND.n819 6.26433
R2183 VGND.n1520 VGND.n1519 6.26433
R2184 VGND.n1556 VGND.n1553 6.26433
R2185 VGND.n1215 VGND.n1214 6.26433
R2186 VGND.n1214 VGND.n1213 6.26433
R2187 VGND.n1774 VGND.n1773 6.12816
R2188 VGND.n254 VGND.n253 6.06007
R2189 VGND.n2359 VGND.n2358 6.02861
R2190 VGND.n2185 VGND.n2184 6.02861
R2191 VGND.n2247 VGND.n2245 6.02861
R2192 VGND.n2266 VGND.n166 6.02861
R2193 VGND.n1957 VGND.n1956 6.02861
R2194 VGND.n1851 VGND.n1849 6.02403
R2195 VGND.n1859 VGND.n1858 6.02403
R2196 VGND.n26 VGND.n22 5.98311
R2197 VGND.n1054 VGND.n1051 5.98311
R2198 VGND.n1299 VGND.n993 5.98311
R2199 VGND.n1607 VGND.n698 5.98311
R2200 VGND.n777 VGND.n776 5.98311
R2201 VGND.n1377 VGND.n868 5.98311
R2202 VGND.n1579 VGND.n1575 5.98311
R2203 VGND.n1223 VGND.n1222 5.98311
R2204 VGND.n1166 VGND.n1163 5.98311
R2205 VGND.n1099 VGND.n47 5.85582
R2206 VGND.n255 VGND.n254 5.85582
R2207 VGND.n1817 VGND.n484 5.85582
R2208 VGND.n961 VGND.n958 5.85582
R2209 VGND.n1775 VGND.n1759 5.85582
R2210 VGND.n1361 VGND.n1360 5.85582
R2211 VGND.n745 VGND.n739 5.85582
R2212 VGND.n1429 VGND.n1428 5.85582
R2213 VGND.n1402 VGND.n1401 5.85582
R2214 VGND.n1445 VGND.n845 5.85582
R2215 VGND.n1474 VGND.n1473 5.85582
R2216 VGND.n1500 VGND.n1499 5.85582
R2217 VGND.n1514 VGND.n819 5.85582
R2218 VGND.n1553 VGND.n1552 5.85582
R2219 VGND.n1215 VGND.n1182 5.85582
R2220 VGND.n2545 VGND.n2534 5.65809
R2221 VGND.n1520 VGND.n814 5.65809
R2222 VGND.n1213 VGND.n1183 5.65809
R2223 VGND.n2376 VGND.n116 5.63966
R2224 VGND.n2045 VGND.n2044 5.63966
R2225 VGND.n2039 VGND.n2038 5.63966
R2226 VGND.n1974 VGND.n336 5.63966
R2227 VGND.n2279 VGND.n161 5.5878
R2228 VGND.n532 VGND.n531 5.55015
R2229 VGND.n2202 VGND.n2201 5.48621
R2230 VGND.n2234 VGND.n182 5.48128
R2231 VGND.n746 VGND.n745 5.37524
R2232 VGND.n1713 VGND.n616 5.27109
R2233 VGND.n968 VGND.n967 5.24958
R2234 VGND.n139 VGND.n137 5.13108
R2235 VGND.n139 VGND.n138 5.13108
R2236 VGND.n2329 VGND.n140 5.13108
R2237 VGND.n2329 VGND.n2328 5.13108
R2238 VGND.n2494 VGND.n2491 5.13108
R2239 VGND.n2494 VGND.n2492 5.13108
R2240 VGND.n248 VGND.n245 5.13108
R2241 VGND.n248 VGND.n247 5.13108
R2242 VGND.n2133 VGND.n2131 5.13108
R2243 VGND.n2133 VGND.n2132 5.13108
R2244 VGND.n2155 VGND.n2134 5.13108
R2245 VGND.n2155 VGND.n2154 5.13108
R2246 VGND.n2091 VGND.n2088 5.13108
R2247 VGND.n2091 VGND.n2090 5.13108
R2248 VGND.n356 VGND.n354 5.13108
R2249 VGND.n356 VGND.n355 5.13108
R2250 VGND.n1927 VGND.n357 5.13108
R2251 VGND.n1927 VGND.n1926 5.13108
R2252 VGND.n394 VGND.n387 5.13108
R2253 VGND.n394 VGND.n388 5.13108
R2254 VGND.n564 VGND.n562 5.13108
R2255 VGND.n564 VGND.n563 5.13108
R2256 VGND.n956 VGND.n936 5.13108
R2257 VGND.n956 VGND.n955 5.13108
R2258 VGND.n1770 VGND.n1767 5.13108
R2259 VGND.n1770 VGND.n1768 5.13108
R2260 VGND.n895 VGND.n881 5.13108
R2261 VGND.n895 VGND.n894 5.13108
R2262 VGND.n753 VGND.n750 5.13108
R2263 VGND.n753 VGND.n751 5.13108
R2264 VGND.n541 VGND.n540 4.92358
R2265 VGND.n2543 VGND.n2542 4.85762
R2266 VGND.n1207 VGND.n1187 4.85762
R2267 VGND.n2228 VGND.n2227 4.85762
R2268 VGND.n974 VGND.n929 4.85762
R2269 VGND.n1538 VGND.n1537 4.85762
R2270 VGND.n26 VGND.n25 4.8005
R2271 VGND.n1054 VGND.n1053 4.8005
R2272 VGND.n1607 VGND.n1606 4.8005
R2273 VGND.n1377 VGND.n1376 4.8005
R2274 VGND.n1579 VGND.n1578 4.8005
R2275 VGND.n1222 VGND.n1221 4.8005
R2276 VGND.n1167 VGND.n1166 4.8005
R2277 VGND.n2410 VGND.n2409 4.72533
R2278 VGND.n2008 VGND.n2007 4.72533
R2279 VGND.n2344 VGND.n2343 4.67352
R2280 VGND.n2363 VGND.n2362 4.67352
R2281 VGND.n2365 VGND.n2363 4.67352
R2282 VGND.n2369 VGND.n120 4.67352
R2283 VGND.n2370 VGND.n2369 4.67352
R2284 VGND.n2393 VGND.n100 4.67352
R2285 VGND.n2397 VGND.n100 4.67352
R2286 VGND.n2398 VGND.n2397 4.67352
R2287 VGND.n2399 VGND.n2398 4.67352
R2288 VGND.n2403 VGND.n2402 4.67352
R2289 VGND.n2413 VGND.n83 4.67352
R2290 VGND.n2427 VGND.n83 4.67352
R2291 VGND.n2428 VGND.n2427 4.67352
R2292 VGND.n2429 VGND.n2428 4.67352
R2293 VGND.n2433 VGND.n2432 4.67352
R2294 VGND.n2452 VGND.n76 4.67352
R2295 VGND.n2453 VGND.n2452 4.67352
R2296 VGND.n2453 VGND.n69 4.67352
R2297 VGND.n2463 VGND.n69 4.67352
R2298 VGND.n2464 VGND.n2463 4.67352
R2299 VGND.n2465 VGND.n2464 4.67352
R2300 VGND.n2469 VGND.n2468 4.67352
R2301 VGND.n2470 VGND.n2469 4.67352
R2302 VGND.n2170 VGND.n2169 4.67352
R2303 VGND.n2189 VGND.n2188 4.67352
R2304 VGND.n2191 VGND.n2189 4.67352
R2305 VGND.n2195 VGND.n198 4.67352
R2306 VGND.n2196 VGND.n2195 4.67352
R2307 VGND.n2237 VGND.n2236 4.67352
R2308 VGND.n2241 VGND.n2240 4.67352
R2309 VGND.n2242 VGND.n2241 4.67352
R2310 VGND.n2254 VGND.n2250 4.67352
R2311 VGND.n2254 VGND.n2253 4.67352
R2312 VGND.n2269 VGND.n2268 4.67352
R2313 VGND.n2273 VGND.n2272 4.67352
R2314 VGND.n2274 VGND.n2273 4.67352
R2315 VGND.n1946 VGND.n1945 4.67352
R2316 VGND.n1961 VGND.n1960 4.67352
R2317 VGND.n1963 VGND.n1961 4.67352
R2318 VGND.n1967 VGND.n340 4.67352
R2319 VGND.n1968 VGND.n1967 4.67352
R2320 VGND.n1991 VGND.n321 4.67352
R2321 VGND.n1995 VGND.n321 4.67352
R2322 VGND.n1996 VGND.n1995 4.67352
R2323 VGND.n1997 VGND.n1996 4.67352
R2324 VGND.n2001 VGND.n2000 4.67352
R2325 VGND.n2011 VGND.n305 4.67352
R2326 VGND.n2025 VGND.n305 4.67352
R2327 VGND.n2026 VGND.n2025 4.67352
R2328 VGND.n2027 VGND.n2026 4.67352
R2329 VGND.n2031 VGND.n2030 4.67352
R2330 VGND.n2390 VGND.n2389 4.63943
R2331 VGND.n2411 VGND.n2410 4.63943
R2332 VGND.n1988 VGND.n1987 4.63943
R2333 VGND.n2009 VGND.n2008 4.63943
R2334 VGND.n1771 VGND.n1764 4.62124
R2335 VGND.n1558 VGND.n804 4.62124
R2336 VGND.n2410 VGND.n95 4.62124
R2337 VGND.n2043 VGND.n2042 4.62124
R2338 VGND.n2008 VGND.n316 4.62124
R2339 VGND.n963 VGND.n934 4.62124
R2340 VGND.n2379 VGND.n116 4.6085
R2341 VGND.n1977 VGND.n336 4.6085
R2342 VGND.n2409 VGND.n2408 4.60638
R2343 VGND.n2007 VGND.n2006 4.60638
R2344 VGND.n2391 VGND.n2390 4.55559
R2345 VGND.n2415 VGND.n2411 4.55559
R2346 VGND.n1989 VGND.n1988 4.55559
R2347 VGND.n2013 VGND.n2009 4.55559
R2348 VGND.n1835 VGND.n1834 4.51815
R2349 VGND.n1844 VGND.n459 4.51815
R2350 VGND.n1312 VGND.n988 4.51815
R2351 VGND.n1289 VGND.n1288 4.51815
R2352 VGND.n1023 VGND.n997 4.51815
R2353 VGND.n1381 VGND.n1372 4.51401
R2354 VGND.n1385 VGND.n867 4.51401
R2355 VGND.n1725 VGND.n1723 4.51401
R2356 VGND.n1735 VGND.n1734 4.51401
R2357 VGND.n1079 VGND.n1072 4.51401
R2358 VGND.n1125 VGND.n1124 4.51401
R2359 VGND.n1103 VGND.n1102 4.51401
R2360 VGND.n2548 VGND.n2547 4.51401
R2361 VGND.n2554 VGND.n2553 4.51401
R2362 VGND.n40 VGND.n39 4.51401
R2363 VGND.n1056 VGND.n1049 4.51401
R2364 VGND.n1155 VGND.n1154 4.51401
R2365 VGND.n1201 VGND.n1037 4.51401
R2366 VGND.n1243 VGND.n1242 4.51401
R2367 VGND.n1169 VGND.n1165 4.51401
R2368 VGND.n1227 VGND.n1226 4.51401
R2369 VGND.n2450 VGND.n2449 4.51401
R2370 VGND.n2461 VGND.n2460 4.51401
R2371 VGND.n2383 VGND.n111 4.51401
R2372 VGND VGND.n2387 4.51401
R2373 VGND.n2351 VGND.n130 4.51401
R2374 VGND.n2356 VGND.n2355 4.51401
R2375 VGND.n2321 VGND.n2311 4.51401
R2376 VGND.n2326 VGND.n2325 4.51401
R2377 VGND.n2517 VGND.n57 4.51401
R2378 VGND.n2509 VGND.n2508 4.51401
R2379 VGND.n2419 VGND.n90 4.51401
R2380 VGND.n2424 VGND.n2423 4.51401
R2381 VGND.n2177 VGND.n2124 4.51401
R2382 VGND.n2182 VGND.n2181 4.51401
R2383 VGND.n2140 VGND.n2138 4.51401
R2384 VGND.n2152 VGND.n2151 4.51401
R2385 VGND.n271 VGND.n209 4.51401
R2386 VGND.n264 VGND.n263 4.51401
R2387 VGND.n2301 VGND.n151 4.51401
R2388 VGND.n156 VGND.n155 4.51401
R2389 VGND.n2217 VGND.n192 4.51401
R2390 VGND.n2222 VGND.n2221 4.51401
R2391 VGND.n2258 VGND.n172 4.51401
R2392 VGND.n2263 VGND.n2262 4.51401
R2393 VGND.n1943 VGND.n1942 4.51401
R2394 VGND.n1954 VGND.n1953 4.51401
R2395 VGND.n1919 VGND.n1909 4.51401
R2396 VGND.n1924 VGND.n1923 4.51401
R2397 VGND.n2113 VGND.n277 4.51401
R2398 VGND.n2106 VGND.n2105 4.51401
R2399 VGND.n2052 VGND.n293 4.51401
R2400 VGND.n2057 VGND.n2056 4.51401
R2401 VGND.n1981 VGND.n331 4.51401
R2402 VGND VGND.n1985 4.51401
R2403 VGND.n2017 VGND.n311 4.51401
R2404 VGND.n2022 VGND.n2021 4.51401
R2405 VGND.n393 VGND.n392 4.51401
R2406 VGND.n402 VGND.n401 4.51401
R2407 VGND.n590 VGND.n498 4.51401
R2408 VGND.n583 VGND.n582 4.51401
R2409 VGND.n1801 VGND.n1800 4.51401
R2410 VGND.n529 VGND.n528 4.51401
R2411 VGND.n448 VGND.n446 4.51401
R2412 VGND.n1862 VGND 4.51401
R2413 VGND.n1902 VGND.n368 4.51401
R2414 VGND.n373 VGND.n372 4.51401
R2415 VGND.n473 VGND.n464 4.51401
R2416 VGND.n1827 VGND.n1826 4.51401
R2417 VGND.n1696 VGND.n629 4.51401
R2418 VGND.n1701 VGND.n1700 4.51401
R2419 VGND.n1634 VGND.n1633 4.51401
R2420 VGND.n1628 VGND.n1627 4.51401
R2421 VGND.n1490 VGND.n829 4.51401
R2422 VGND.n1495 VGND.n1494 4.51401
R2423 VGND.n1662 VGND.n652 4.51401
R2424 VGND.n667 VGND.n666 4.51401
R2425 VGND.n1457 VGND.n843 4.51401
R2426 VGND.n1462 VGND.n1461 4.51401
R2427 VGND.n1277 VGND.n1275 4.51401
R2428 VGND.n1668 VGND.n1667 4.51401
R2429 VGND.n954 VGND.n953 4.51401
R2430 VGND.n948 VGND.n947 4.51401
R2431 VGND.n1791 VGND.n596 4.51401
R2432 VGND.n1782 VGND.n1781 4.51401
R2433 VGND.n1326 VGND.n918 4.51401
R2434 VGND.n923 VGND.n922 4.51401
R2435 VGND.n1334 VGND.n907 4.51401
R2436 VGND.n1338 VGND.n914 4.51401
R2437 VGND.n1420 VGND.n856 4.51401
R2438 VGND.n1425 VGND.n1424 4.51401
R2439 VGND.n893 VGND.n892 4.51401
R2440 VGND.n1365 VGND.n1364 4.51401
R2441 VGND.n770 VGND.n769 4.51401
R2442 VGND.n764 VGND.n763 4.51401
R2443 VGND.n1602 VGND.n1601 4.51401
R2444 VGND.n795 VGND.n794 4.51401
R2445 VGND.n1526 VGND.n818 4.51401
R2446 VGND.n1531 VGND.n811 4.51401
R2447 VGND.n1559 VGND.n806 4.51401
R2448 VGND.n1592 VGND.n1591 4.51401
R2449 VGND.n2516 VGND.n2515 4.5005
R2450 VGND.n2504 VGND.n60 4.5005
R2451 VGND.n2507 VGND.n2486 4.5005
R2452 VGND.n2320 VGND.n2319 4.5005
R2453 VGND.n2317 VGND.n2316 4.5005
R2454 VGND.n2313 VGND.n141 4.5005
R2455 VGND.n2350 VGND.n2349 4.5005
R2456 VGND.n2348 VGND.n2347 4.5005
R2457 VGND.n125 VGND.n124 4.5005
R2458 VGND.n2382 VGND.n2381 4.5005
R2459 VGND.n114 VGND.n113 4.5005
R2460 VGND.n106 VGND.n105 4.5005
R2461 VGND.n2447 VGND.n74 4.5005
R2462 VGND.n2456 VGND.n2455 4.5005
R2463 VGND.n75 VGND.n71 4.5005
R2464 VGND.n2418 VGND.n2417 4.5005
R2465 VGND.n94 VGND.n93 4.5005
R2466 VGND.n85 VGND.n84 4.5005
R2467 VGND.n188 VGND.n187 4.5005
R2468 VGND.n2300 VGND.n2299 4.5005
R2469 VGND.n2298 VGND.n2297 4.5005
R2470 VGND.n2294 VGND.n2293 4.5005
R2471 VGND.n270 VGND.n269 4.5005
R2472 VGND.n259 VGND.n212 4.5005
R2473 VGND.n262 VGND.n241 4.5005
R2474 VGND.n2142 VGND.n2141 4.5005
R2475 VGND.n2147 VGND.n2146 4.5005
R2476 VGND.n2144 VGND.n2135 4.5005
R2477 VGND.n2176 VGND.n2175 4.5005
R2478 VGND.n2174 VGND.n2173 4.5005
R2479 VGND.n203 VGND.n202 4.5005
R2480 VGND.n2216 VGND.n2215 4.5005
R2481 VGND.n2212 VGND.n2211 4.5005
R2482 VGND.n2257 VGND.n2256 4.5005
R2483 VGND.n176 VGND.n175 4.5005
R2484 VGND.n168 VGND.n167 4.5005
R2485 VGND.n327 VGND.n326 4.5005
R2486 VGND.n2051 VGND.n2050 4.5005
R2487 VGND.n2049 VGND.n2048 4.5005
R2488 VGND.n296 VGND.n289 4.5005
R2489 VGND.n2112 VGND.n2111 4.5005
R2490 VGND.n2101 VGND.n280 4.5005
R2491 VGND.n2104 VGND.n2084 4.5005
R2492 VGND.n1918 VGND.n1917 4.5005
R2493 VGND.n1915 VGND.n1914 4.5005
R2494 VGND.n1911 VGND.n358 4.5005
R2495 VGND.n1940 VGND.n348 4.5005
R2496 VGND.n1949 VGND.n1948 4.5005
R2497 VGND.n345 VGND.n344 4.5005
R2498 VGND.n1980 VGND.n1979 4.5005
R2499 VGND.n334 VGND.n333 4.5005
R2500 VGND.n2016 VGND.n2015 4.5005
R2501 VGND.n315 VGND.n314 4.5005
R2502 VGND.n307 VGND.n306 4.5005
R2503 VGND.n447 VGND.n441 4.5005
R2504 VGND.n1867 VGND.n1866 4.5005
R2505 VGND.n444 VGND.n442 4.5005
R2506 VGND.n517 VGND.n491 4.5005
R2507 VGND.n520 VGND.n519 4.5005
R2508 VGND.n527 VGND.n526 4.5005
R2509 VGND.n589 VGND.n588 4.5005
R2510 VGND.n578 VGND.n501 4.5005
R2511 VGND.n581 VGND.n559 4.5005
R2512 VGND.n390 VGND.n389 4.5005
R2513 VGND.n397 VGND.n396 4.5005
R2514 VGND.n386 VGND.n382 4.5005
R2515 VGND.n1901 VGND.n1900 4.5005
R2516 VGND.n1899 VGND.n1898 4.5005
R2517 VGND.n1895 VGND.n1894 4.5005
R2518 VGND.n472 VGND.n467 4.5005
R2519 VGND.n1832 VGND.n1831 4.5005
R2520 VGND.n476 VGND.n470 4.5005
R2521 VGND.n1780 VGND.n1760 4.5005
R2522 VGND.n940 VGND.n939 4.5005
R2523 VGND.n943 VGND.n942 4.5005
R2524 VGND.n946 VGND.n945 4.5005
R2525 VGND.n1285 VGND.n1284 4.5005
R2526 VGND.n1281 VGND.n1280 4.5005
R2527 VGND.n1279 VGND.n644 4.5005
R2528 VGND.n1695 VGND.n1694 4.5005
R2529 VGND.n634 VGND.n633 4.5005
R2530 VGND.n624 VGND.n623 4.5005
R2531 VGND.n1727 VGND.n1726 4.5005
R2532 VGND.n1730 VGND.n1729 4.5005
R2533 VGND.n611 VGND.n610 4.5005
R2534 VGND.n1790 VGND.n1789 4.5005
R2535 VGND.n1777 VGND.n599 4.5005
R2536 VGND.n1325 VGND.n1324 4.5005
R2537 VGND.n1323 VGND.n1322 4.5005
R2538 VGND.n1319 VGND.n1318 4.5005
R2539 VGND.n741 VGND.n732 4.5005
R2540 VGND.n891 VGND.n890 4.5005
R2541 VGND.n887 VGND.n886 4.5005
R2542 VGND.n882 VGND.n879 4.5005
R2543 VGND.n1333 VGND.n1332 4.5005
R2544 VGND.n1330 VGND.n911 4.5005
R2545 VGND.n1340 VGND.n1339 4.5005
R2546 VGND.n1661 VGND.n1660 4.5005
R2547 VGND.n661 VGND.n655 4.5005
R2548 VGND.n665 VGND.n664 4.5005
R2549 VGND.n686 VGND.n677 4.5005
R2550 VGND.n689 VGND.n688 4.5005
R2551 VGND.n681 VGND.n680 4.5005
R2552 VGND.n740 VGND.n729 4.5005
R2553 VGND.n743 VGND.n742 4.5005
R2554 VGND.n710 VGND.n700 4.5005
R2555 VGND.n714 VGND.n713 4.5005
R2556 VGND.n715 VGND.n703 4.5005
R2557 VGND.n805 VGND.n802 4.5005
R2558 VGND.n1380 VGND.n1379 4.5005
R2559 VGND.n1373 VGND.n869 4.5005
R2560 VGND.n1387 VGND.n1386 4.5005
R2561 VGND.n1419 VGND.n1418 4.5005
R2562 VGND.n1417 VGND.n1416 4.5005
R2563 VGND.n1413 VGND.n852 4.5005
R2564 VGND.n1456 VGND.n1455 4.5005
R2565 VGND.n1453 VGND.n1452 4.5005
R2566 VGND.n1450 VGND.n840 4.5005
R2567 VGND.n1489 VGND.n1488 4.5005
R2568 VGND.n833 VGND.n832 4.5005
R2569 VGND.n1483 VGND.n825 4.5005
R2570 VGND.n1525 VGND.n1524 4.5005
R2571 VGND.n1523 VGND.n1522 4.5005
R2572 VGND.n1533 VGND.n1532 4.5005
R2573 VGND.n1562 VGND.n1561 4.5005
R2574 VGND.n1567 VGND.n1566 4.5005
R2575 VGND.n14 VGND.n9 4.5005
R2576 VGND.n1171 VGND.n1170 4.5005
R2577 VGND.n1176 VGND.n1175 4.5005
R2578 VGND.n1177 VGND.n1161 4.5005
R2579 VGND.n1190 VGND.n1189 4.5005
R2580 VGND.n1195 VGND.n1194 4.5005
R2581 VGND.n1196 VGND.n1034 4.5005
R2582 VGND.n1059 VGND.n1058 4.5005
R2583 VGND.n1063 VGND.n1062 4.5005
R2584 VGND.n1048 VGND.n1044 4.5005
R2585 VGND.n1078 VGND.n1074 4.5005
R2586 VGND.n1130 VGND.n1129 4.5005
R2587 VGND.n1083 VGND.n1077 4.5005
R2588 VGND.n1101 VGND.n48 4.5005
R2589 VGND.n2530 VGND.n2529 4.5005
R2590 VGND.n2531 VGND.n44 4.5005
R2591 VGND.n13 VGND.n5 4.5005
R2592 VGND.n16 VGND.n15 4.5005
R2593 VGND.n775 VGND.n774 4.38311
R2594 VGND.n2343 VGND.n2342 4.36875
R2595 VGND.n2344 VGND.n123 4.36875
R2596 VGND.n2362 VGND.n122 4.36875
R2597 VGND.n2371 VGND.n2370 4.36875
R2598 VGND.n2393 VGND.n2392 4.36875
R2599 VGND.n2405 VGND.n96 4.36875
R2600 VGND.n2414 VGND.n2413 4.36875
R2601 VGND.n2435 VGND.n79 4.36875
R2602 VGND.n2443 VGND.n76 4.36875
R2603 VGND.n2470 VGND.n65 4.36875
R2604 VGND.n2169 VGND.n2168 4.36875
R2605 VGND.n2170 VGND.n201 4.36875
R2606 VGND.n2188 VGND.n200 4.36875
R2607 VGND.n2197 VGND.n2196 4.36875
R2608 VGND.n2236 VGND.n2235 4.36875
R2609 VGND.n2242 VGND.n178 4.36875
R2610 VGND.n2253 VGND.n2251 4.36875
R2611 VGND.n2268 VGND.n2267 4.36875
R2612 VGND.n2274 VGND.n162 4.36875
R2613 VGND.n1945 VGND.n349 4.36875
R2614 VGND.n1946 VGND.n343 4.36875
R2615 VGND.n1960 VGND.n342 4.36875
R2616 VGND.n1969 VGND.n1968 4.36875
R2617 VGND.n1991 VGND.n1990 4.36875
R2618 VGND.n2003 VGND.n317 4.36875
R2619 VGND.n2012 VGND.n2011 4.36875
R2620 VGND.n2034 VGND.n2033 4.36875
R2621 VGND.n961 VGND.n960 4.28986
R2622 VGND.n965 VGND.n933 4.28986
R2623 VGND.n1773 VGND.n1772 4.28986
R2624 VGND.n1432 VGND.n1431 4.28986
R2625 VGND.n1448 VGND.n1447 4.28986
R2626 VGND.n1477 VGND.n1476 4.28986
R2627 VGND.n1556 VGND.n1555 4.28986
R2628 VGND.n984 VGND.n983 4.14168
R2629 VGND.n37 VGND.n36 4.11798
R2630 VGND.n36 VGND.n35 4.11798
R2631 VGND.n1087 VGND.n1085 4.11798
R2632 VGND.n1116 VGND.n1087 4.11798
R2633 VGND.n1145 VGND.n1144 4.11798
R2634 VGND.n1144 VGND.n1143 4.11798
R2635 VGND.n2064 VGND.n2063 4.11798
R2636 VGND.n2063 VGND.n285 4.11798
R2637 VGND.n535 VGND.n534 4.11798
R2638 VGND.n420 VGND.n419 4.11798
R2639 VGND.n419 VGND.n375 4.11798
R2640 VGND.n1878 VGND.n1877 4.11798
R2641 VGND.n1877 VGND.n1876 4.11798
R2642 VGND.n684 VGND.n676 4.11798
R2643 VGND.n1248 VGND.n1030 4.11798
R2644 VGND.n1251 VGND.n1030 4.11798
R2645 VGND.n2043 VGND.n298 4.09013
R2646 VGND.n1772 VGND.n1771 4.07323
R2647 VGND.n1431 VGND.n849 4.07323
R2648 VGND.n1447 VGND.n838 4.07323
R2649 VGND.n1476 VGND.n834 4.07323
R2650 VGND.n1555 VGND.n804 4.07323
R2651 VGND.n2488 VGND.n2485 4.03876
R2652 VGND.n576 VGND.n575 4.03876
R2653 VGND.n2375 VGND.n118 3.97459
R2654 VGND.n1973 VGND.n338 3.97459
R2655 VGND.n2334 VGND.n2333 3.96548
R2656 VGND.n2337 VGND.n2334 3.96548
R2657 VGND.n2499 VGND.n2498 3.96548
R2658 VGND.n2286 VGND.n160 3.96548
R2659 VGND.n2160 VGND.n2159 3.96548
R2660 VGND.n2163 VGND.n2160 3.96548
R2661 VGND.n2109 VGND.n2108 3.96548
R2662 VGND.n2108 VGND.n2083 3.96548
R2663 VGND.n2098 VGND.n2097 3.96548
R2664 VGND.n1932 VGND.n1931 3.96548
R2665 VGND.n1933 VGND.n1932 3.96548
R2666 VGND.n571 VGND.n570 3.96548
R2667 VGND.n411 VGND.n410 3.96548
R2668 VGND.n413 VGND.n411 3.96548
R2669 VGND.n1712 VGND.n619 3.90948
R2670 VGND.n1712 VGND.n1711 3.90948
R2671 VGND.n538 VGND.n510 3.75994
R2672 VGND.n2333 VGND.n136 3.7069
R2673 VGND.n2500 VGND.n2499 3.7069
R2674 VGND.n2281 VGND.n160 3.7069
R2675 VGND.n2159 VGND.n2130 3.7069
R2676 VGND.n2206 VGND.n194 3.7069
R2677 VGND.n2207 VGND.n2206 3.7069
R2678 VGND.n2109 VGND.n2082 3.7069
R2679 VGND.n2095 VGND.n2087 3.7069
R2680 VGND.n1931 VGND.n353 3.7069
R2681 VGND.n571 VGND.n560 3.7069
R2682 VGND.n410 VGND.n380 3.7069
R2683 VGND.n413 VGND.n412 3.7069
R2684 VGND.n2544 VGND.n2535 3.50735
R2685 VGND.n971 VGND.n930 3.50735
R2686 VGND.n1536 VGND.n1535 3.50735
R2687 VGND.n1209 VGND.n1185 3.50735
R2688 VGND.n761 VGND.n760 3.44377
R2689 VGND.n760 VGND.n759 3.44377
R2690 VGND.n1385 VGND.n1384 3.43925
R2691 VGND.n1382 VGND.n1381 3.43925
R2692 VGND.n1734 VGND.n1733 3.43925
R2693 VGND.n1725 VGND.n1724 3.43925
R2694 VGND.n2460 VGND.n2459 3.43925
R2695 VGND.n2449 VGND.n2448 3.43925
R2696 VGND.n2387 VGND.n2386 3.43925
R2697 VGND.n2384 VGND.n2383 3.43925
R2698 VGND.n2355 VGND.n2354 3.43925
R2699 VGND.n2352 VGND.n2351 3.43925
R2700 VGND.n2325 VGND.n2324 3.43925
R2701 VGND.n2322 VGND.n2321 3.43925
R2702 VGND.n2508 VGND.n54 3.43925
R2703 VGND.n2518 VGND.n2517 3.43925
R2704 VGND.n2423 VGND.n2422 3.43925
R2705 VGND.n2420 VGND.n2419 3.43925
R2706 VGND.n2181 VGND.n2180 3.43925
R2707 VGND.n2178 VGND.n2177 3.43925
R2708 VGND.n2151 VGND.n2150 3.43925
R2709 VGND.n2140 VGND.n2139 3.43925
R2710 VGND.n263 VGND.n207 3.43925
R2711 VGND.n272 VGND.n271 3.43925
R2712 VGND.n155 VGND.n148 3.43925
R2713 VGND.n2302 VGND.n2301 3.43925
R2714 VGND.n2221 VGND.n2220 3.43925
R2715 VGND.n2218 VGND.n2217 3.43925
R2716 VGND.n2262 VGND.n2261 3.43925
R2717 VGND.n2259 VGND.n2258 3.43925
R2718 VGND.n1953 VGND.n1952 3.43925
R2719 VGND.n1942 VGND.n1941 3.43925
R2720 VGND.n1923 VGND.n1922 3.43925
R2721 VGND.n1920 VGND.n1919 3.43925
R2722 VGND.n2105 VGND.n274 3.43925
R2723 VGND.n2114 VGND.n2113 3.43925
R2724 VGND.n2056 VGND.n2055 3.43925
R2725 VGND.n2053 VGND.n2052 3.43925
R2726 VGND.n1985 VGND.n1984 3.43925
R2727 VGND.n1982 VGND.n1981 3.43925
R2728 VGND.n2021 VGND.n2020 3.43925
R2729 VGND.n2018 VGND.n2017 3.43925
R2730 VGND.n401 VGND.n400 3.43925
R2731 VGND.n392 VGND.n391 3.43925
R2732 VGND.n582 VGND.n496 3.43925
R2733 VGND.n591 VGND.n590 3.43925
R2734 VGND.n528 VGND.n493 3.43925
R2735 VGND.n1800 VGND.n1799 3.43925
R2736 VGND.n1863 VGND.n1862 3.43925
R2737 VGND.n449 VGND.n448 3.43925
R2738 VGND.n372 VGND.n365 3.43925
R2739 VGND.n1903 VGND.n1902 3.43925
R2740 VGND.n1828 VGND.n1827 3.43925
R2741 VGND.n474 VGND.n473 3.43925
R2742 VGND.n1700 VGND.n1699 3.43925
R2743 VGND.n1697 VGND.n1696 3.43925
R2744 VGND.n1629 VGND.n1628 3.43925
R2745 VGND.n1633 VGND.n1632 3.43925
R2746 VGND.n1494 VGND.n1493 3.43925
R2747 VGND.n1491 VGND.n1490 3.43925
R2748 VGND.n666 VGND.n649 3.43925
R2749 VGND.n1663 VGND.n1662 3.43925
R2750 VGND.n1461 VGND.n1460 3.43925
R2751 VGND.n1458 VGND.n1457 3.43925
R2752 VGND.n949 VGND.n948 3.43925
R2753 VGND.n953 VGND.n952 3.43925
R2754 VGND.n1781 VGND.n593 3.43925
R2755 VGND.n1792 VGND.n1791 3.43925
R2756 VGND.n922 VGND.n916 3.43925
R2757 VGND.n1327 VGND.n1326 3.43925
R2758 VGND.n1338 VGND.n1337 3.43925
R2759 VGND.n1335 VGND.n1334 3.43925
R2760 VGND.n1424 VGND.n1423 3.43925
R2761 VGND.n1421 VGND.n1420 3.43925
R2762 VGND.n765 VGND.n764 3.43925
R2763 VGND.n769 VGND.n768 3.43925
R2764 VGND.n796 VGND.n795 3.43925
R2765 VGND.n1601 VGND.n1600 3.43925
R2766 VGND.n1531 VGND.n1530 3.43925
R2767 VGND.n1527 VGND.n1526 3.43925
R2768 VGND.n41 VGND.n40 3.41902
R2769 VGND.n2553 VGND.n2552 3.41902
R2770 VGND.n1228 VGND.n1227 3.41646
R2771 VGND.n1165 VGND.n1159 3.41646
R2772 VGND.n1242 VGND.n1241 3.41636
R2773 VGND.n1239 VGND.n1037 3.41636
R2774 VGND.n1156 VGND.n1155 3.41624
R2775 VGND.n1049 VGND.n1043 3.41624
R2776 VGND.n1126 VGND.n1125 3.41605
R2777 VGND.n1081 VGND.n1079 3.41605
R2778 VGND.n1374 VGND.n1371 3.4105
R2779 VGND.n871 VGND.n870 3.4105
R2780 VGND.n613 VGND.n612 3.4105
R2781 VGND.n1732 VGND.n1731 3.4105
R2782 VGND.n2551 VGND.n7 3.4105
R2783 VGND.n42 VGND.n8 3.4105
R2784 VGND.n2549 VGND.n2548 3.4105
R2785 VGND.n1102 VGND.n50 3.4105
R2786 VGND.n2526 VGND.n49 3.4105
R2787 VGND.n2528 VGND.n2527 3.4105
R2788 VGND.n1060 VGND.n1040 3.4105
R2789 VGND.n1061 VGND.n1041 3.4105
R2790 VGND.n1238 VGND.n1038 3.4105
R2791 VGND.n1193 VGND.n1035 3.4105
R2792 VGND.n1173 VGND.n1172 3.4105
R2793 VGND.n1174 VGND.n1160 3.4105
R2794 VGND.n1080 VGND.n1076 3.4105
R2795 VGND.n1128 VGND.n1127 3.4105
R2796 VGND.n73 VGND.n72 3.4105
R2797 VGND.n2458 VGND.n2457 3.4105
R2798 VGND.n115 VGND.n110 3.4105
R2799 VGND.n112 VGND.n107 3.4105
R2800 VGND.n131 VGND.n129 3.4105
R2801 VGND.n2346 VGND.n126 3.4105
R2802 VGND.n2312 VGND.n2310 3.4105
R2803 VGND.n2315 VGND.n142 3.4105
R2804 VGND.n58 VGND.n56 3.4105
R2805 VGND.n2506 VGND.n2505 3.4105
R2806 VGND.n91 VGND.n89 3.4105
R2807 VGND.n92 VGND.n86 3.4105
R2808 VGND.n2125 VGND.n2123 3.4105
R2809 VGND.n2172 VGND.n204 3.4105
R2810 VGND.n2137 VGND.n2136 3.4105
R2811 VGND.n2149 VGND.n2148 3.4105
R2812 VGND.n210 VGND.n208 3.4105
R2813 VGND.n261 VGND.n260 3.4105
R2814 VGND.n152 VGND.n150 3.4105
R2815 VGND.n2296 VGND.n2295 3.4105
R2816 VGND.n193 VGND.n191 3.4105
R2817 VGND.n2210 VGND.n189 3.4105
R2818 VGND.n173 VGND.n171 3.4105
R2819 VGND.n174 VGND.n169 3.4105
R2820 VGND.n347 VGND.n346 3.4105
R2821 VGND.n1951 VGND.n1950 3.4105
R2822 VGND.n1910 VGND.n1908 3.4105
R2823 VGND.n1913 VGND.n359 3.4105
R2824 VGND.n278 VGND.n276 3.4105
R2825 VGND.n2103 VGND.n2102 3.4105
R2826 VGND.n294 VGND.n292 3.4105
R2827 VGND.n2047 VGND.n290 3.4105
R2828 VGND.n335 VGND.n330 3.4105
R2829 VGND.n332 VGND.n328 3.4105
R2830 VGND.n312 VGND.n310 3.4105
R2831 VGND.n313 VGND.n308 3.4105
R2832 VGND.n384 VGND.n383 3.4105
R2833 VGND.n399 VGND.n398 3.4105
R2834 VGND.n499 VGND.n497 3.4105
R2835 VGND.n580 VGND.n579 3.4105
R2836 VGND.n518 VGND.n492 3.4105
R2837 VGND.n516 VGND.n515 3.4105
R2838 VGND.n445 VGND.n443 3.4105
R2839 VGND.n1865 VGND.n1864 3.4105
R2840 VGND.n369 VGND.n367 3.4105
R2841 VGND.n1897 VGND.n1896 3.4105
R2842 VGND.n471 VGND.n469 3.4105
R2843 VGND.n1830 VGND.n1829 3.4105
R2844 VGND.n630 VGND.n628 3.4105
R2845 VGND.n632 VGND.n625 3.4105
R2846 VGND.n1631 VGND.n678 3.4105
R2847 VGND.n1630 VGND.n679 3.4105
R2848 VGND.n830 VGND.n828 3.4105
R2849 VGND.n831 VGND.n826 3.4105
R2850 VGND.n653 VGND.n651 3.4105
R2851 VGND.n663 VGND.n662 3.4105
R2852 VGND.n844 VGND.n842 3.4105
R2853 VGND.n1451 VGND.n841 3.4105
R2854 VGND.n1666 VGND.n1665 3.4105
R2855 VGND.n1665 VGND.n648 3.4105
R2856 VGND.n1667 VGND.n1666 3.4105
R2857 VGND.n1277 VGND.n648 3.4105
R2858 VGND.n1283 VGND.n1282 3.4105
R2859 VGND.n1278 VGND.n645 3.4105
R2860 VGND.n951 VGND.n941 3.4105
R2861 VGND.n950 VGND.n944 3.4105
R2862 VGND.n597 VGND.n595 3.4105
R2863 VGND.n1779 VGND.n1778 3.4105
R2864 VGND.n919 VGND.n917 3.4105
R2865 VGND.n1321 VGND.n1320 3.4105
R2866 VGND.n1331 VGND.n1329 3.4105
R2867 VGND.n915 VGND.n913 3.4105
R2868 VGND.n857 VGND.n855 3.4105
R2869 VGND.n1415 VGND.n853 3.4105
R2870 VGND.n1367 VGND.n1366 3.4105
R2871 VGND.n1367 VGND.n877 3.4105
R2872 VGND.n1366 VGND.n1365 3.4105
R2873 VGND.n892 VGND.n877 3.4105
R2874 VGND.n889 VGND.n888 3.4105
R2875 VGND.n885 VGND.n878 3.4105
R2876 VGND.n767 VGND.n730 3.4105
R2877 VGND.n766 VGND.n731 3.4105
R2878 VGND.n711 VGND.n701 3.4105
R2879 VGND.n712 VGND.n702 3.4105
R2880 VGND.n1528 VGND.n817 3.4105
R2881 VGND.n1529 VGND.n816 3.4105
R2882 VGND.n1594 VGND.n1593 3.4105
R2883 VGND.n1594 VGND.n800 3.4105
R2884 VGND.n1593 VGND.n1592 3.4105
R2885 VGND.n806 VGND.n800 3.4105
R2886 VGND.n1564 VGND.n1563 3.4105
R2887 VGND.n1565 VGND.n801 3.4105
R2888 VGND.n540 VGND.n539 3.31239
R2889 VGND.n685 VGND.n684 3.22288
R2890 VGND.n761 VGND.n747 3.21921
R2891 VGND.n756 VGND.n755 3.21921
R2892 VGND.n2541 VGND.n2540 3.2005
R2893 VGND.n973 VGND.n928 3.2005
R2894 VGND.n1540 VGND.n812 3.2005
R2895 VGND.n1208 VGND.n1186 3.2005
R2896 VGND.n252 VGND.n243 3.13241
R2897 VGND.n1816 VGND.n1815 3.13241
R2898 VGND.n1405 VGND.n1404 3.13241
R2899 VGND.n1503 VGND.n1502 3.13241
R2900 VGND.n2213 VGND.n186 3.09945
R2901 VGND.n2372 VGND.n118 3.05276
R2902 VGND.n1970 VGND.n338 3.05276
R2903 VGND.n2494 VGND.n2493 3.04861
R2904 VGND.n2329 VGND.n2327 3.04861
R2905 VGND.n248 VGND.n246 3.04861
R2906 VGND.n2155 VGND.n2153 3.04861
R2907 VGND.n2091 VGND.n2089 3.04861
R2908 VGND.n1927 VGND.n1925 3.04861
R2909 VGND.n565 VGND.n564 3.04861
R2910 VGND.n1770 VGND.n1769 3.04861
R2911 VGND.n753 VGND.n752 3.04861
R2912 VGND.n1479 VGND.n834 3.04861
R2913 VGND.n1434 VGND.n849 3.04861
R2914 VGND.n1015 VGND.n1012 3.01226
R2915 VGND.n1299 VGND.n1298 2.92224
R2916 VGND.n2044 VGND.n2043 2.92166
R2917 VGND.n2337 VGND.n2336 2.88804
R2918 VGND.n2163 VGND.n2162 2.88804
R2919 VGND.n1933 VGND.n351 2.88804
R2920 VGND.n2336 VGND.n2335 2.79323
R2921 VGND.n2162 VGND.n2161 2.79323
R2922 VGND.n351 VGND.n350 2.79323
R2923 VGND.n2501 VGND.n2488 2.77203
R2924 VGND.n575 VGND.n574 2.77203
R2925 VGND.n244 VGND.n243 2.7239
R2926 VGND.n1815 VGND.n1814 2.7239
R2927 VGND.n898 VGND.n897 2.7239
R2928 VGND.n1404 VGND.n1403 2.7239
R2929 VGND.n1502 VGND.n1501 2.7239
R2930 VGND.n533 VGND.n532 2.68581
R2931 VGND.n2537 VGND.n2536 2.63064
R2932 VGND.n976 VGND.n975 2.63064
R2933 VGND.n1539 VGND.n813 2.63064
R2934 VGND.n1206 VGND.n1205 2.63064
R2935 VGND.n2226 VGND.n2225 2.55412
R2936 VGND.n2475 VGND.n2474 2.50679
R2937 VGND.n1807 VGND.n486 2.50679
R2938 VGND.n1647 VGND.n669 2.50679
R2939 VGND.n299 VGND.n298 2.38348
R2940 VGND.n2365 VGND.n2364 2.33701
R2941 VGND.n2364 VGND.n120 2.33701
R2942 VGND.n2399 VGND.n98 2.33701
R2943 VGND.n2402 VGND.n98 2.33701
R2944 VGND.n2404 VGND.n2403 2.33701
R2945 VGND.n2405 VGND.n2404 2.33701
R2946 VGND.n2429 VGND.n81 2.33701
R2947 VGND.n2432 VGND.n81 2.33701
R2948 VGND.n2434 VGND.n2433 2.33701
R2949 VGND.n2435 VGND.n2434 2.33701
R2950 VGND.n2465 VGND.n67 2.33701
R2951 VGND.n2468 VGND.n67 2.33701
R2952 VGND.n2191 VGND.n2190 2.33701
R2953 VGND.n2190 VGND.n198 2.33701
R2954 VGND.n2237 VGND.n180 2.33701
R2955 VGND.n2240 VGND.n180 2.33701
R2956 VGND.n2250 VGND.n177 2.33701
R2957 VGND.n2269 VGND.n164 2.33701
R2958 VGND.n2272 VGND.n164 2.33701
R2959 VGND.n1963 VGND.n1962 2.33701
R2960 VGND.n1962 VGND.n340 2.33701
R2961 VGND.n1997 VGND.n319 2.33701
R2962 VGND.n2000 VGND.n319 2.33701
R2963 VGND.n2002 VGND.n2001 2.33701
R2964 VGND.n2003 VGND.n2002 2.33701
R2965 VGND.n2027 VGND.n303 2.33701
R2966 VGND.n2030 VGND.n303 2.33701
R2967 VGND.n2032 VGND.n2031 2.33701
R2968 VGND.n2034 VGND.n2032 2.33701
R2969 VGND.n2230 VGND.n184 2.33067
R2970 VGND.n267 VGND.n239 2.25932
R2971 VGND.n1853 VGND.n458 2.25932
R2972 VGND.n1312 VGND.n1311 2.25932
R2973 VGND.n1290 VGND.n1289 2.25932
R2974 VGND.n1274 VGND.n1273 2.25932
R2975 VGND.n1273 VGND.n1272 2.25932
R2976 VGND.n1739 VGND.n606 2.25932
R2977 VGND.n1354 VGND.n902 2.25932
R2978 VGND.n1015 VGND.n1014 2.25932
R2979 VGND.n718 VGND.n717 2.25932
R2980 VGND.n2339 VGND.n134 2.25312
R2981 VGND.n2165 VGND.n2128 2.25312
R2982 VGND.n1936 VGND.n1935 2.25312
R2983 VGND.n1712 VGND.n1710 2.25293
R2984 VGND.n134 VGND.n133 2.2228
R2985 VGND.n2128 VGND.n2127 2.2228
R2986 VGND.n1937 VGND.n1936 2.2228
R2987 VGND.n897 VGND.n896 2.17922
R2988 VGND.n960 VGND.n959 2.13383
R2989 VGND.n104 VGND.n103 2.11085
R2990 VGND.n325 VGND.n324 2.11085
R2991 VGND.n2097 VGND.n2096 2.06919
R2992 VGND.n2246 VGND.n177 2.03225
R2993 VGND.n2498 VGND.n2489 1.98299
R2994 VGND.n2287 VGND.n2286 1.98299
R2995 VGND.n2086 VGND.n2083 1.98299
R2996 VGND.n2098 VGND.n2086 1.98299
R2997 VGND.n570 VGND.n569 1.98299
R2998 VGND.n737 VGND.n727 1.97497
R2999 VGND.n2229 VGND.n185 1.91571
R3000 VGND.n2096 VGND.n2095 1.8968
R3001 VGND.n1786 VGND.n1785 1.88285
R3002 VGND.n1298 VGND.n1297 1.87876
R3003 VGND.n759 VGND.n748 1.79699
R3004 VGND.n546 VGND.n544 1.75824
R3005 VGND.n1304 VGND.n1302 1.7528
R3006 VGND.n2490 VGND.n2489 1.72441
R3007 VGND.n2288 VGND.n2287 1.72441
R3008 VGND.n569 VGND.n568 1.72441
R3009 VGND.n2524 VGND.n43 1.70468
R3010 VGND.n2525 VGND.n2524 1.70468
R3011 VGND.n1126 VGND.n1082 1.70348
R3012 VGND.n1082 VGND.n1081 1.70348
R3013 VGND.n1157 VGND.n1156 1.70338
R3014 VGND.n1157 VGND.n1043 1.70338
R3015 VGND.n1241 VGND.n1240 1.70332
R3016 VGND.n1240 VGND.n1239 1.70332
R3017 VGND.n1229 VGND.n1228 1.70327
R3018 VGND.n1229 VGND.n1159 1.70327
R3019 VGND.n41 VGND.n6 1.70199
R3020 VGND.n2552 VGND.n6 1.70199
R3021 VGND.n576 VGND.n558 1.7012
R3022 VGND.n1493 VGND.n1492 1.69188
R3023 VGND.n1492 VGND.n1491 1.69188
R3024 VGND.n1629 VGND.n627 1.69188
R3025 VGND.n1632 VGND.n627 1.69188
R3026 VGND.n1699 VGND.n1698 1.69188
R3027 VGND.n1698 VGND.n1697 1.69188
R3028 VGND.n1828 VGND.n475 1.69188
R3029 VGND.n475 VGND.n474 1.69188
R3030 VGND.n2020 VGND.n2019 1.69188
R3031 VGND.n2019 VGND.n2018 1.69188
R3032 VGND.n2261 VGND.n2260 1.69188
R3033 VGND.n2260 VGND.n2259 1.69188
R3034 VGND.n2422 VGND.n2421 1.69188
R3035 VGND.n2421 VGND.n2420 1.69188
R3036 VGND.n1460 VGND.n1459 1.69188
R3037 VGND.n1459 VGND.n1458 1.69188
R3038 VGND.n1664 VGND.n649 1.69188
R3039 VGND.n1664 VGND.n1663 1.69188
R3040 VGND.n1863 VGND.n450 1.69188
R3041 VGND.n450 VGND.n449 1.69188
R3042 VGND.n1984 VGND.n1983 1.69188
R3043 VGND.n1983 VGND.n1982 1.69188
R3044 VGND.n2220 VGND.n2219 1.69188
R3045 VGND.n2219 VGND.n2218 1.69188
R3046 VGND.n2386 VGND.n2385 1.69188
R3047 VGND.n2385 VGND.n2384 1.69188
R3048 VGND.n1665 VGND.n647 1.69188
R3049 VGND.n1423 VGND.n1422 1.69188
R3050 VGND.n1422 VGND.n1421 1.69188
R3051 VGND.n1337 VGND.n1336 1.69188
R3052 VGND.n1336 VGND.n1335 1.69188
R3053 VGND.n1328 VGND.n916 1.69188
R3054 VGND.n1328 VGND.n1327 1.69188
R3055 VGND.n1904 VGND.n365 1.69188
R3056 VGND.n1904 VGND.n1903 1.69188
R3057 VGND.n1952 VGND.n205 1.69188
R3058 VGND.n1941 VGND.n205 1.69188
R3059 VGND.n2180 VGND.n2179 1.69188
R3060 VGND.n2179 VGND.n2178 1.69188
R3061 VGND.n2354 VGND.n2353 1.69188
R3062 VGND.n2353 VGND.n2352 1.69188
R3063 VGND.n1384 VGND.n1383 1.69188
R3064 VGND.n1383 VGND.n1382 1.69188
R3065 VGND.n949 VGND.n875 1.69188
R3066 VGND.n952 VGND.n875 1.69188
R3067 VGND.n400 VGND.n360 1.69188
R3068 VGND.n391 VGND.n360 1.69188
R3069 VGND.n1922 VGND.n1921 1.69188
R3070 VGND.n1921 VGND.n1920 1.69188
R3071 VGND.n2150 VGND.n146 1.69188
R3072 VGND.n2139 VGND.n146 1.69188
R3073 VGND.n2324 VGND.n2323 1.69188
R3074 VGND.n2323 VGND.n2322 1.69188
R3075 VGND.n1367 VGND.n876 1.69188
R3076 VGND.n1530 VGND.n797 1.69188
R3077 VGND.n1527 VGND.n797 1.69188
R3078 VGND.n1599 VGND.n796 1.69188
R3079 VGND.n1600 VGND.n1599 1.69188
R3080 VGND.n1733 VGND.n494 1.69188
R3081 VGND.n1724 VGND.n494 1.69188
R3082 VGND.n1798 VGND.n493 1.69188
R3083 VGND.n1799 VGND.n1798 1.69188
R3084 VGND.n2055 VGND.n2054 1.69188
R3085 VGND.n2054 VGND.n2053 1.69188
R3086 VGND.n2303 VGND.n148 1.69188
R3087 VGND.n2303 VGND.n2302 1.69188
R3088 VGND.n2459 VGND.n52 1.69188
R3089 VGND.n2448 VGND.n52 1.69188
R3090 VGND.n765 VGND.n594 1.69188
R3091 VGND.n768 VGND.n594 1.69188
R3092 VGND.n1793 VGND.n593 1.69188
R3093 VGND.n1793 VGND.n1792 1.69188
R3094 VGND.n592 VGND.n496 1.69188
R3095 VGND.n592 VGND.n591 1.69188
R3096 VGND.n2115 VGND.n274 1.69188
R3097 VGND.n2115 VGND.n2114 1.69188
R3098 VGND.n273 VGND.n207 1.69188
R3099 VGND.n273 VGND.n272 1.69188
R3100 VGND.n2519 VGND.n54 1.69188
R3101 VGND.n2519 VGND.n2518 1.69188
R3102 VGND.n1594 VGND.n799 1.69188
R3103 VGND.n756 VGND.n748 1.64728
R3104 VGND.n523 VGND.n513 1.61169
R3105 VGND.n2279 VGND.n2278 1.47352
R3106 VGND.n2198 VGND.n195 1.34658
R3107 VGND.n298 VGND.n297 1.3283
R3108 VGND.n2341 VGND.n133 1.29527
R3109 VGND.n2167 VGND.n2127 1.29527
R3110 VGND.n1938 VGND.n1937 1.29527
R3111 VGND.n2512 VGND.n2511 1.25365
R3112 VGND.n2203 VGND.n2202 1.25033
R3113 VGND.n407 VGND.n406 1.20723
R3114 VGND.n25 VGND.n24 1.18311
R3115 VGND.n1053 VGND.n1052 1.18311
R3116 VGND.n1297 VGND.n1296 1.18311
R3117 VGND.n1606 VGND.n1605 1.18311
R3118 VGND.n774 VGND.n773 1.18311
R3119 VGND.n1376 VGND.n1375 1.18311
R3120 VGND.n1578 VGND.n1577 1.18311
R3121 VGND.n1221 VGND.n1220 1.18311
R3122 VGND.n1168 VGND.n1167 1.18311
R3123 VGND.n2540 VGND.n2537 1.14023
R3124 VGND.n975 VGND.n928 1.14023
R3125 VGND.n1540 VGND.n1539 1.14023
R3126 VGND.n1206 VGND.n1186 1.14023
R3127 VGND.n1673 VGND.n1672 1.12991
R3128 VGND.n2282 VGND.n2280 1.12954
R3129 VGND.n1036 VGND 1.12383
R3130 VGND.n1158 VGND 1.11689
R3131 VGND.n1232 VGND 1.11689
R3132 VGND.n51 VGND 1.07702
R3133 VGND.n551 VGND.n550 1.07463
R3134 VGND.n586 VGND.n557 0.985115
R3135 VGND.n1359 VGND.n896 0.953691
R3136 VGND.n1772 VGND.n1763 0.952566
R3137 VGND.n1431 VGND.n1430 0.952566
R3138 VGND.n1447 VGND.n1446 0.952566
R3139 VGND.n1476 VGND.n1475 0.952566
R3140 VGND.n1555 VGND.n1554 0.952566
R3141 VGND.n1771 VGND.n1766 0.899674
R3142 VGND.n1638 VGND.n1637 0.895605
R3143 VGND.n691 VGND.n685 0.895605
R3144 VGND.n2336 VGND.n134 0.892621
R3145 VGND.n2162 VGND.n2128 0.892621
R3146 VGND.n1936 VGND.n351 0.892621
R3147 VGND.n2541 VGND.n2535 0.833377
R3148 VGND.n1535 VGND.n812 0.833377
R3149 VGND.n1209 VGND.n1208 0.833377
R3150 VGND.n2230 VGND.n2229 0.830425
R3151 VGND.n2224 VGND.n186 0.798505
R3152 VGND.n1858 VGND.n1857 0.753441
R3153 VGND.n1308 VGND.n992 0.753441
R3154 VGND.n1753 VGND.n1752 0.753441
R3155 VGND.n1885 VGND.n1884 0.716584
R3156 VGND.n2225 VGND.n184 0.606984
R3157 VGND.n2560 VGND.n2559 0.537563
R3158 VGND.n30 VGND.n21 0.537563
R3159 VGND.n1136 VGND.n1071 0.537563
R3160 VGND.n1111 VGND.n1088 0.537563
R3161 VGND.n1066 VGND.n1065 0.537563
R3162 VGND.n1138 VGND.n1137 0.537563
R3163 VGND.n2442 VGND.n77 0.537563
R3164 VGND.n2075 VGND.n2074 0.537563
R3165 VGND.n2062 VGND.n2061 0.537563
R3166 VGND.n2073 VGND.n283 0.537563
R3167 VGND.n548 VGND.n547 0.537563
R3168 VGND.n521 VGND.n488 0.537563
R3169 VGND.n544 VGND.n506 0.537563
R3170 VGND.n428 VGND.n427 0.537563
R3171 VGND.n1892 VGND.n1891 0.537563
R3172 VGND.n1871 VGND.n436 0.537563
R3173 VGND.n1623 VGND.n1622 0.537563
R3174 VGND.n1191 VGND.n1188 0.537563
R3175 VGND.n1256 VGND.n1028 0.537563
R3176 VGND.n2545 VGND.n2544 0.526527
R3177 VGND.n968 VGND.n930 0.526527
R3178 VGND.n972 VGND.n971 0.526527
R3179 VGND.n1536 VGND.n814 0.526527
R3180 VGND.n1185 VGND.n1183 0.526527
R3181 VGND.n874 VGND.n873 0.500125
R3182 VGND.n1370 VGND.n1369 0.500125
R3183 VGND.n2309 VGND.n2308 0.500125
R3184 VGND.n2121 VGND.n206 0.500125
R3185 VGND.n1907 VGND.n1906 0.500125
R3186 VGND.n145 VGND.n144 0.500125
R3187 VGND.n2477 VGND.n2476 0.448052
R3188 VGND.n425 VGND.n424 0.448052
R3189 VGND.n1890 VGND.n1889 0.448052
R3190 VGND.n29 VGND.n22 0.417891
R3191 VGND.n1051 VGND.n1026 0.417891
R3192 VGND.n1052 VGND.n1047 0.417891
R3193 VGND.n1302 VGND.n993 0.417891
R3194 VGND.n1296 VGND.n1295 0.417891
R3195 VGND.n1610 VGND.n698 0.417891
R3196 VGND.n1605 VGND.n1604 0.417891
R3197 VGND.n778 VGND.n777 0.417891
R3198 VGND.n776 VGND.n775 0.417891
R3199 VGND.n773 VGND.n772 0.417891
R3200 VGND.n1389 VGND.n868 0.417891
R3201 VGND.n1582 VGND.n1575 0.417891
R3202 VGND.n1224 VGND.n1223 0.417891
R3203 VGND.n1220 VGND.n1219 0.417891
R3204 VGND.n1179 VGND.n1163 0.417891
R3205 VGND.n1105 VGND.n1099 0.409011
R3206 VGND.n256 VGND.n255 0.409011
R3207 VGND.n249 VGND.n244 0.409011
R3208 VGND.n484 VGND.n481 0.409011
R3209 VGND.n958 VGND.n957 0.409011
R3210 VGND.n967 VGND.n966 0.409011
R3211 VGND.n1784 VGND.n1759 0.409011
R3212 VGND.n1362 VGND.n1361 0.409011
R3213 VGND.n1356 VGND.n898 0.409011
R3214 VGND.n1428 VGND.n1427 0.409011
R3215 VGND.n1401 VGND.n1400 0.409011
R3216 VGND.n1403 VGND.n860 0.409011
R3217 VGND.n1442 VGND.n845 0.409011
R3218 VGND.n1473 VGND.n1472 0.409011
R3219 VGND.n1499 VGND.n1498 0.409011
R3220 VGND.n1501 VGND.n822 0.409011
R3221 VGND.n1515 VGND.n1514 0.409011
R3222 VGND.n1552 VGND.n1551 0.409011
R3223 VGND.n1182 VGND.n1180 0.409011
R3224 VGND.n2226 VGND.n2224 0.383542
R3225 VGND.n363 VGND.n309 0.3805
R3226 VGND.n2119 VGND.n170 0.3805
R3227 VGND.n2306 VGND.n88 0.3805
R3228 VGND.n827 VGND.n798 0.3805
R3229 VGND.n626 VGND.n495 0.3805
R3230 VGND.n87 VGND.n53 0.3805
R3231 VGND.n143 VGND.n108 0.3805
R3232 VGND.n2307 VGND.n109 0.3805
R3233 VGND.n2120 VGND.n190 0.3805
R3234 VGND.n364 VGND.n329 0.3805
R3235 VGND.n872 VGND.n646 0.3805
R3236 VGND.n1368 VGND.n650 0.3805
R3237 VGND.n144 VGND.n127 0.3805
R3238 VGND.n2308 VGND.n128 0.3805
R3239 VGND.n2122 VGND.n2121 0.3805
R3240 VGND.n1906 VGND.n1905 0.3805
R3241 VGND.n873 VGND.n366 0.3805
R3242 VGND.n1369 VGND.n854 0.3805
R3243 VGND.n2523 VGND.n2522 0.3805
R3244 VGND.n2305 VGND.n2304 0.3805
R3245 VGND.n2118 VGND.n149 0.3805
R3246 VGND.n362 VGND.n291 0.3805
R3247 VGND.n1797 VGND.n1796 0.3805
R3248 VGND.n1598 VGND.n1597 0.3805
R3249 VGND.n361 VGND.n275 0.3805
R3250 VGND.n2117 VGND.n2116 0.3805
R3251 VGND.n147 VGND.n55 0.3805
R3252 VGND.n2521 VGND.n2520 0.3805
R3253 VGND.n1596 VGND.n1595 0.3805
R3254 VGND.n1795 VGND.n1794 0.3805
R3255 VGND.n1787 VGND.n1786 0.376971
R3256 VGND.n2069 VGND.n283 0.358542
R3257 VGND.n1805 VGND.n1804 0.358542
R3258 VGND.n534 VGND.n510 0.358542
R3259 VGND.n1647 VGND.n1646 0.358542
R3260 VGND.n1813 VGND.n1812 0.340926
R3261 VGND.n973 VGND.n972 0.307349
R3262 VGND.n2342 VGND.n2341 0.305262
R3263 VGND.n2358 VGND.n123 0.305262
R3264 VGND.n2359 VGND.n122 0.305262
R3265 VGND.n2372 VGND.n2371 0.305262
R3266 VGND.n2392 VGND.n2391 0.305262
R3267 VGND.n2408 VGND.n96 0.305262
R3268 VGND.n2415 VGND.n2414 0.305262
R3269 VGND.n2438 VGND.n79 0.305262
R3270 VGND.n2444 VGND.n2443 0.305262
R3271 VGND.n2473 VGND.n65 0.305262
R3272 VGND.n2168 VGND.n2167 0.305262
R3273 VGND.n2184 VGND.n201 0.305262
R3274 VGND.n2185 VGND.n200 0.305262
R3275 VGND.n2198 VGND.n2197 0.305262
R3276 VGND.n2235 VGND.n2234 0.305262
R3277 VGND.n2245 VGND.n178 0.305262
R3278 VGND.n2247 VGND.n2246 0.305262
R3279 VGND.n2251 VGND.n166 0.305262
R3280 VGND.n2267 VGND.n2266 0.305262
R3281 VGND.n2278 VGND.n162 0.305262
R3282 VGND.n1938 VGND.n349 0.305262
R3283 VGND.n1956 VGND.n343 0.305262
R3284 VGND.n1957 VGND.n342 0.305262
R3285 VGND.n1970 VGND.n1969 0.305262
R3286 VGND.n1990 VGND.n1989 0.305262
R3287 VGND.n2006 VGND.n317 0.305262
R3288 VGND.n2013 VGND.n2012 0.305262
R3289 VGND.n2033 VGND.n301 0.305262
R3290 VGND.n2339 VGND.n2338 0.298074
R3291 VGND.n2165 VGND.n2164 0.298074
R3292 VGND.n1935 VGND.n1934 0.298074
R3293 VGND.n1234 VGND.n1233 0.278782
R3294 VGND.n2536 VGND.n0 0.263514
R3295 VGND.n977 VGND.n976 0.263514
R3296 VGND.n813 VGND.n810 0.263514
R3297 VGND.n1205 VGND.n1204 0.263514
R3298 VGND.n2330 VGND.n136 0.259086
R3299 VGND.n2501 VGND.n2500 0.259086
R3300 VGND.n2495 VGND.n2490 0.259086
R3301 VGND.n2282 VGND.n2281 0.259086
R3302 VGND.n2289 VGND.n2288 0.259086
R3303 VGND.n2156 VGND.n2130 0.259086
R3304 VGND.n2203 VGND.n194 0.259086
R3305 VGND.n2208 VGND.n2207 0.259086
R3306 VGND.n2082 VGND.n2081 0.259086
R3307 VGND.n2092 VGND.n2087 0.259086
R3308 VGND.n1928 VGND.n353 0.259086
R3309 VGND.n574 VGND.n560 0.259086
R3310 VGND.n568 VGND.n567 0.259086
R3311 VGND.n407 VGND.n380 0.259086
R3312 VGND.n412 VGND.n378 0.259086
R3313 VGND.n1434 VGND.n1433 0.239726
R3314 VGND.n1479 VGND.n1478 0.239381
R3315 VGND.n1710 VGND 0.237784
R3316 VGND.n747 VGND.n746 0.225061
R3317 VGND.n755 VGND.n754 0.225061
R3318 VGND.n1230 VGND.n1229 0.218753
R3319 VGND.n253 VGND.n252 0.204755
R3320 VGND.n738 VGND.n737 0.204755
R3321 VGND.n739 VGND.n738 0.204755
R3322 VGND.n1710 VGND 0.200023
R3323 VGND VGND.n2339 0.199635
R3324 VGND VGND.n2165 0.199635
R3325 VGND.n1935 VGND 0.199635
R3326 VGND.n1237 VGND.n1236 0.196532
R3327 VGND.n1231 VGND.n1230 0.196532
R3328 VGND.n1237 VGND.n1039 0.196234
R3329 VGND.n1233 VGND.n1232 0.195539
R3330 VGND.n185 VGND.n182 0.192021
R3331 VGND.n1558 VGND.n1557 0.180304
R3332 VGND.n1769 VGND 0.17983
R3333 VGND.n752 VGND 0.17983
R3334 VGND.n2484 VGND.n2483 0.179521
R3335 VGND.n1805 VGND.n486 0.179521
R3336 VGND.n1646 VGND.n1645 0.179521
R3337 VGND.n2493 VGND 0.179485
R3338 VGND.n246 VGND 0.179485
R3339 VGND.n2089 VGND 0.179485
R3340 VGND VGND.n565 0.179485
R3341 VGND.n2550 VGND.n2549 0.178787
R3342 VGND.n1042 VGND.n50 0.175416
R3343 VGND.n1698 VGND.n627 0.1603
R3344 VGND.n1665 VGND.n1664 0.1603
R3345 VGND.n1336 VGND.n1328 0.1603
R3346 VGND.n1367 VGND.n875 0.1603
R3347 VGND.n1599 VGND.n494 0.1603
R3348 VGND.n1793 VGND.n594 0.1603
R3349 VGND.n626 VGND.n475 0.159712
R3350 VGND.n646 VGND.n450 0.159712
R3351 VGND.n1904 VGND.n366 0.159712
R3352 VGND.n874 VGND.n360 0.159712
R3353 VGND.n1798 VGND.n1797 0.159712
R3354 VGND.n1794 VGND.n592 0.159712
R3355 VGND VGND.n95 0.158169
R3356 VGND VGND.n316 0.158169
R3357 VGND.n2042 VGND 0.158169
R3358 VGND VGND.n1764 0.156867
R3359 VGND.n1559 VGND.n1558 0.151658
R3360 VGND.n2327 VGND.n2326 0.143027
R3361 VGND.n2153 VGND.n2152 0.143027
R3362 VGND.n1925 VGND.n1924 0.143027
R3363 VGND.n2327 VGND 0.14207
R3364 VGND.n2493 VGND 0.14207
R3365 VGND.n2153 VGND 0.14207
R3366 VGND.n246 VGND 0.14207
R3367 VGND.n1925 VGND 0.14207
R3368 VGND.n2089 VGND 0.14207
R3369 VGND.n565 VGND 0.14207
R3370 VGND VGND.n1479 0.14207
R3371 VGND.n1769 VGND 0.141725
R3372 VGND.n752 VGND 0.141725
R3373 VGND VGND.n1434 0.141725
R3374 VGND.n2421 VGND.n87 0.137387
R3375 VGND.n2385 VGND.n108 0.137387
R3376 VGND.n2353 VGND.n127 0.137387
R3377 VGND.n2323 VGND.n145 0.137387
R3378 VGND.n2523 VGND.n52 0.137387
R3379 VGND.n2520 VGND.n2519 0.137387
R3380 VGND.n1775 VGND.n1774 0.13667
R3381 VGND.n1492 VGND.n827 0.126812
R3382 VGND.n1459 VGND.n650 0.126812
R3383 VGND.n1422 VGND.n854 0.126812
R3384 VGND.n1383 VGND.n1370 0.126812
R3385 VGND.n1598 VGND.n797 0.126812
R3386 VGND.n1595 VGND.n1594 0.126812
R3387 VGND.n2202 VGND.n195 0.126617
R3388 VGND.n2019 VGND.n309 0.125637
R3389 VGND.n1983 VGND.n329 0.125637
R3390 VGND.n1905 VGND.n205 0.125637
R3391 VGND.n1921 VGND.n1907 0.125637
R3392 VGND.n2054 VGND.n291 0.125637
R3393 VGND.n2115 VGND.n275 0.125637
R3394 VGND.n2280 VGND.n2279 0.120632
R3395 VGND.n963 VGND 0.120408
R3396 VGND.n2332 VGND.n2331 0.120292
R3397 VGND.n2332 VGND.n135 0.120292
R3398 VGND.n2338 VGND.n135 0.120292
R3399 VGND.n2361 VGND.n2360 0.120292
R3400 VGND.n2361 VGND.n121 0.120292
R3401 VGND.n2366 VGND.n121 0.120292
R3402 VGND.n2367 VGND.n2366 0.120292
R3403 VGND.n2368 VGND.n2367 0.120292
R3404 VGND.n2368 VGND.n119 0.120292
R3405 VGND.n2373 VGND.n119 0.120292
R3406 VGND.n2394 VGND.n101 0.120292
R3407 VGND.n2395 VGND.n2394 0.120292
R3408 VGND.n2396 VGND.n2395 0.120292
R3409 VGND.n2396 VGND.n99 0.120292
R3410 VGND.n2400 VGND.n99 0.120292
R3411 VGND.n2401 VGND.n2400 0.120292
R3412 VGND.n2401 VGND.n97 0.120292
R3413 VGND.n2406 VGND.n97 0.120292
R3414 VGND.n2407 VGND.n2406 0.120292
R3415 VGND.n2426 VGND.n2425 0.120292
R3416 VGND.n2426 VGND.n82 0.120292
R3417 VGND.n2430 VGND.n82 0.120292
R3418 VGND.n2431 VGND.n2430 0.120292
R3419 VGND.n2431 VGND.n80 0.120292
R3420 VGND.n2436 VGND.n80 0.120292
R3421 VGND.n2437 VGND.n2436 0.120292
R3422 VGND.n2446 VGND.n2445 0.120292
R3423 VGND.n2462 VGND.n68 0.120292
R3424 VGND.n2466 VGND.n68 0.120292
R3425 VGND.n2467 VGND.n2466 0.120292
R3426 VGND.n2467 VGND.n66 0.120292
R3427 VGND.n2471 VGND.n66 0.120292
R3428 VGND.n2472 VGND.n2471 0.120292
R3429 VGND.n2479 VGND.n63 0.120292
R3430 VGND.n2480 VGND.n2479 0.120292
R3431 VGND.n2481 VGND.n2480 0.120292
R3432 VGND.n2502 VGND.n2487 0.120292
R3433 VGND.n2497 VGND.n2487 0.120292
R3434 VGND.n2497 VGND.n2496 0.120292
R3435 VGND.n2158 VGND.n2157 0.120292
R3436 VGND.n2158 VGND.n2129 0.120292
R3437 VGND.n2164 VGND.n2129 0.120292
R3438 VGND.n2187 VGND.n2186 0.120292
R3439 VGND.n2187 VGND.n199 0.120292
R3440 VGND.n2192 VGND.n199 0.120292
R3441 VGND.n2193 VGND.n2192 0.120292
R3442 VGND.n2194 VGND.n2193 0.120292
R3443 VGND.n2194 VGND.n197 0.120292
R3444 VGND.n2199 VGND.n197 0.120292
R3445 VGND.n2205 VGND.n2204 0.120292
R3446 VGND.n2231 VGND.n183 0.120292
R3447 VGND.n2232 VGND.n2231 0.120292
R3448 VGND.n2233 VGND.n181 0.120292
R3449 VGND.n2238 VGND.n181 0.120292
R3450 VGND.n2239 VGND.n2238 0.120292
R3451 VGND.n2239 VGND.n179 0.120292
R3452 VGND.n2243 VGND.n179 0.120292
R3453 VGND.n2244 VGND.n2243 0.120292
R3454 VGND.n2249 VGND.n2248 0.120292
R3455 VGND.n2265 VGND.n165 0.120292
R3456 VGND.n2270 VGND.n165 0.120292
R3457 VGND.n2271 VGND.n2270 0.120292
R3458 VGND.n2271 VGND.n163 0.120292
R3459 VGND.n2275 VGND.n163 0.120292
R3460 VGND.n2277 VGND.n2275 0.120292
R3461 VGND.n2284 VGND.n2283 0.120292
R3462 VGND.n2285 VGND.n2284 0.120292
R3463 VGND.n223 VGND.n222 0.120292
R3464 VGND.n226 VGND.n223 0.120292
R3465 VGND.n227 VGND.n226 0.120292
R3466 VGND.n228 VGND.n227 0.120292
R3467 VGND.n228 VGND.n219 0.120292
R3468 VGND.n219 VGND.n217 0.120292
R3469 VGND.n233 VGND.n217 0.120292
R3470 VGND.n234 VGND.n233 0.120292
R3471 VGND.n235 VGND.n234 0.120292
R3472 VGND.n235 VGND.n215 0.120292
R3473 VGND.n257 VGND.n242 0.120292
R3474 VGND.n251 VGND.n242 0.120292
R3475 VGND.n1930 VGND.n1929 0.120292
R3476 VGND.n1930 VGND.n352 0.120292
R3477 VGND.n1934 VGND.n352 0.120292
R3478 VGND.n1959 VGND.n1958 0.120292
R3479 VGND.n1959 VGND.n341 0.120292
R3480 VGND.n1964 VGND.n341 0.120292
R3481 VGND.n1965 VGND.n1964 0.120292
R3482 VGND.n1966 VGND.n1965 0.120292
R3483 VGND.n1966 VGND.n339 0.120292
R3484 VGND.n1971 VGND.n339 0.120292
R3485 VGND.n1992 VGND.n322 0.120292
R3486 VGND.n1993 VGND.n1992 0.120292
R3487 VGND.n1994 VGND.n1993 0.120292
R3488 VGND.n1994 VGND.n320 0.120292
R3489 VGND.n1998 VGND.n320 0.120292
R3490 VGND.n1999 VGND.n1998 0.120292
R3491 VGND.n1999 VGND.n318 0.120292
R3492 VGND.n2004 VGND.n318 0.120292
R3493 VGND.n2005 VGND.n2004 0.120292
R3494 VGND.n2024 VGND.n2023 0.120292
R3495 VGND.n2024 VGND.n304 0.120292
R3496 VGND.n2028 VGND.n304 0.120292
R3497 VGND.n2029 VGND.n2028 0.120292
R3498 VGND.n2029 VGND.n302 0.120292
R3499 VGND.n2035 VGND.n302 0.120292
R3500 VGND.n2036 VGND.n2035 0.120292
R3501 VGND.n2065 VGND.n286 0.120292
R3502 VGND.n2066 VGND.n2065 0.120292
R3503 VGND VGND.n2066 0.120292
R3504 VGND.n2072 VGND.n2071 0.120292
R3505 VGND.n2077 VGND.n282 0.120292
R3506 VGND.n2078 VGND.n2077 0.120292
R3507 VGND.n2100 VGND.n2099 0.120292
R3508 VGND.n2099 VGND.n2085 0.120292
R3509 VGND.n2094 VGND.n2085 0.120292
R3510 VGND.n2094 VGND.n2093 0.120292
R3511 VGND.n409 VGND.n408 0.120292
R3512 VGND.n409 VGND.n379 0.120292
R3513 VGND.n414 VGND.n379 0.120292
R3514 VGND.n415 VGND.n414 0.120292
R3515 VGND.n421 VGND.n376 0.120292
R3516 VGND.n423 VGND.n422 0.120292
R3517 VGND.n1887 VGND.n1886 0.120292
R3518 VGND.n1886 VGND.n430 0.120292
R3519 VGND.n1881 VGND.n430 0.120292
R3520 VGND.n1881 VGND.n1880 0.120292
R3521 VGND.n1880 VGND.n1879 0.120292
R3522 VGND.n1879 VGND.n433 0.120292
R3523 VGND.n1873 VGND.n1872 0.120292
R3524 VGND.n1856 VGND.n1855 0.120292
R3525 VGND.n1855 VGND.n1854 0.120292
R3526 VGND.n1854 VGND.n455 0.120292
R3527 VGND.n1848 VGND.n455 0.120292
R3528 VGND.n1848 VGND.n1847 0.120292
R3529 VGND.n1847 VGND.n1846 0.120292
R3530 VGND.n1846 VGND.n460 0.120292
R3531 VGND.n1839 VGND.n460 0.120292
R3532 VGND.n1839 VGND.n1838 0.120292
R3533 VGND.n1838 VGND.n1837 0.120292
R3534 VGND.n1825 VGND.n477 0.120292
R3535 VGND.n1819 VGND.n1818 0.120292
R3536 VGND.n1818 VGND.n483 0.120292
R3537 VGND.n1811 VGND.n483 0.120292
R3538 VGND.n530 VGND.n511 0.120292
R3539 VGND.n536 VGND.n511 0.120292
R3540 VGND.n537 VGND.n536 0.120292
R3541 VGND.n537 VGND.n507 0.120292
R3542 VGND.n542 VGND.n507 0.120292
R3543 VGND.n543 VGND.n542 0.120292
R3544 VGND.n552 VGND.n505 0.120292
R3545 VGND.n553 VGND.n552 0.120292
R3546 VGND.n554 VGND.n553 0.120292
R3547 VGND.n573 VGND.n572 0.120292
R3548 VGND.n572 VGND.n561 0.120292
R3549 VGND.n566 VGND.n561 0.120292
R3550 VGND.n962 VGND.n935 0.120292
R3551 VGND.n964 VGND.n931 0.120292
R3552 VGND.n969 VGND.n931 0.120292
R3553 VGND.n970 VGND.n969 0.120292
R3554 VGND.n970 VGND.n927 0.120292
R3555 VGND.n978 VGND.n927 0.120292
R3556 VGND.n980 VGND.n979 0.120292
R3557 VGND.n1314 VGND.n1313 0.120292
R3558 VGND.n1313 VGND.n989 0.120292
R3559 VGND.n1307 VGND.n989 0.120292
R3560 VGND.n1307 VGND.n1306 0.120292
R3561 VGND.n1301 VGND.n1300 0.120292
R3562 VGND.n1300 VGND.n994 0.120292
R3563 VGND.n1292 VGND.n1267 0.120292
R3564 VGND.n1676 VGND.n640 0.120292
R3565 VGND.n1677 VGND.n1676 0.120292
R3566 VGND.n1678 VGND.n1677 0.120292
R3567 VGND.n1678 VGND.n638 0.120292
R3568 VGND.n1683 VGND.n638 0.120292
R3569 VGND.n1684 VGND.n1683 0.120292
R3570 VGND.n1702 VGND.n620 0.120292
R3571 VGND.n1708 VGND.n620 0.120292
R3572 VGND.n1715 VGND.n615 0.120292
R3573 VGND.n1722 VGND.n615 0.120292
R3574 VGND.n1740 VGND.n608 0.120292
R3575 VGND.n1741 VGND.n1740 0.120292
R3576 VGND.n1741 VGND.n604 0.120292
R3577 VGND.n1745 VGND.n604 0.120292
R3578 VGND.n1746 VGND.n1745 0.120292
R3579 VGND.n1747 VGND.n1746 0.120292
R3580 VGND.n1747 VGND.n601 0.120292
R3581 VGND.n1754 VGND.n601 0.120292
R3582 VGND.n1755 VGND.n1754 0.120292
R3583 VGND.n1776 VGND.n1761 0.120292
R3584 VGND.n1363 VGND.n880 0.120292
R3585 VGND.n1353 VGND.n899 0.120292
R3586 VGND.n1353 VGND.n1352 0.120292
R3587 VGND.n1352 VGND.n903 0.120292
R3588 VGND.n904 VGND.n903 0.120292
R3589 VGND.n1346 VGND.n1345 0.120292
R3590 VGND.n1008 VGND.n1007 0.120292
R3591 VGND.n1009 VGND.n1008 0.120292
R3592 VGND.n1016 VGND.n998 0.120292
R3593 VGND.n1017 VGND.n1016 0.120292
R3594 VGND.n1655 VGND.n1654 0.120292
R3595 VGND.n1654 VGND.n1653 0.120292
R3596 VGND.n1649 VGND.n668 0.120292
R3597 VGND.n1648 VGND.n670 0.120292
R3598 VGND.n1641 VGND.n1640 0.120292
R3599 VGND.n1640 VGND.n674 0.120292
R3600 VGND.n1635 VGND.n674 0.120292
R3601 VGND.n1626 VGND.n682 0.120292
R3602 VGND.n1621 VGND.n682 0.120292
R3603 VGND.n1620 VGND.n1619 0.120292
R3604 VGND.n1619 VGND.n693 0.120292
R3605 VGND.n1614 VGND.n693 0.120292
R3606 VGND.n1614 VGND.n1613 0.120292
R3607 VGND.n793 VGND.n705 0.120292
R3608 VGND.n788 VGND.n705 0.120292
R3609 VGND.n788 VGND.n787 0.120292
R3610 VGND.n787 VGND.n786 0.120292
R3611 VGND.n786 VGND.n722 0.120292
R3612 VGND.n781 VGND.n722 0.120292
R3613 VGND.n781 VGND.n780 0.120292
R3614 VGND.n779 VGND.n726 0.120292
R3615 VGND.n771 VGND.n726 0.120292
R3616 VGND.n762 VGND.n734 0.120292
R3617 VGND.n758 VGND.n734 0.120292
R3618 VGND.n758 VGND.n757 0.120292
R3619 VGND.n757 VGND.n749 0.120292
R3620 VGND.n1393 VGND.n1392 0.120292
R3621 VGND.n1397 VGND.n863 0.120292
R3622 VGND.n1398 VGND.n1397 0.120292
R3623 VGND.n1399 VGND.n861 0.120292
R3624 VGND.n1406 VGND.n861 0.120292
R3625 VGND.n1407 VGND.n1406 0.120292
R3626 VGND.n1433 VGND.n850 0.120292
R3627 VGND.n1439 VGND.n1438 0.120292
R3628 VGND.n1444 VGND.n1443 0.120292
R3629 VGND.n1469 VGND.n837 0.120292
R3630 VGND.n1471 VGND.n835 0.120292
R3631 VGND.n1478 VGND.n835 0.120292
R3632 VGND.n1497 VGND.n823 0.120292
R3633 VGND.n1504 VGND.n823 0.120292
R3634 VGND.n1505 VGND.n1504 0.120292
R3635 VGND.n1511 VGND.n1510 0.120292
R3636 VGND.n1517 VGND.n1516 0.120292
R3637 VGND.n1518 VGND.n1517 0.120292
R3638 VGND.n1542 VGND.n1541 0.120292
R3639 VGND.n1548 VGND.n809 0.120292
R3640 VGND.n1550 VGND.n807 0.120292
R3641 VGND.n1557 VGND.n807 0.120292
R3642 VGND.n1585 VGND.n1573 0.120292
R3643 VGND.n1581 VGND.n1580 0.120292
R3644 VGND.n1580 VGND.n1576 0.120292
R3645 VGND.n1225 VGND.n1162 0.120292
R3646 VGND.n1218 VGND.n1162 0.120292
R3647 VGND.n1217 VGND.n1216 0.120292
R3648 VGND.n1216 VGND.n1181 0.120292
R3649 VGND.n1212 VGND.n1181 0.120292
R3650 VGND.n1212 VGND.n1211 0.120292
R3651 VGND.n1211 VGND.n1210 0.120292
R3652 VGND.n1210 VGND.n1184 0.120292
R3653 VGND.n1203 VGND.n1184 0.120292
R3654 VGND.n1245 VGND.n1244 0.120292
R3655 VGND.n1245 VGND.n1031 0.120292
R3656 VGND.n1249 VGND.n1031 0.120292
R3657 VGND.n1250 VGND.n1249 0.120292
R3658 VGND.n1250 VGND.n1029 0.120292
R3659 VGND.n1254 VGND.n1029 0.120292
R3660 VGND.n1255 VGND.n1254 0.120292
R3661 VGND.n1055 VGND.n1050 0.120292
R3662 VGND.n1153 VGND.n1046 0.120292
R3663 VGND.n1149 VGND.n1046 0.120292
R3664 VGND.n1149 VGND.n1148 0.120292
R3665 VGND.n1148 VGND.n1147 0.120292
R3666 VGND.n1147 VGND.n1069 0.120292
R3667 VGND.n1142 VGND.n1069 0.120292
R3668 VGND.n1142 VGND.n1141 0.120292
R3669 VGND.n1141 VGND.n1140 0.120292
R3670 VGND.n1140 VGND 0.120292
R3671 VGND.n1135 VGND.n1134 0.120292
R3672 VGND.n1123 VGND.n1084 0.120292
R3673 VGND.n1119 VGND.n1084 0.120292
R3674 VGND.n1119 VGND.n1118 0.120292
R3675 VGND.n1118 VGND.n1117 0.120292
R3676 VGND.n1117 VGND.n1086 0.120292
R3677 VGND.n1113 VGND.n1086 0.120292
R3678 VGND.n1113 VGND.n1112 0.120292
R3679 VGND.n1108 VGND.n1107 0.120292
R3680 VGND.n2546 VGND.n46 0.120292
R3681 VGND.n2539 VGND.n46 0.120292
R3682 VGND.n2539 VGND.n2538 0.120292
R3683 VGND.n2563 VGND.n2562 0.120292
R3684 VGND.n2561 VGND.n2 0.120292
R3685 VGND.n2556 VGND.n2 0.120292
R3686 VGND.n2556 VGND.n2555 0.120292
R3687 VGND.n38 VGND.n11 0.120292
R3688 VGND.n33 VGND.n11 0.120292
R3689 VGND.n33 VGND.n32 0.120292
R3690 VGND.n32 VGND.n31 0.120292
R3691 VGND.n28 VGND.n27 0.120292
R3692 VGND.n27 VGND.n23 0.120292
R3693 VGND.n873 VGND.n872 0.120125
R3694 VGND.n872 VGND.n495 0.120125
R3695 VGND.n1796 VGND.n495 0.120125
R3696 VGND.n1796 VGND.n1795 0.120125
R3697 VGND.n1369 VGND.n1368 0.120125
R3698 VGND.n1368 VGND.n798 0.120125
R3699 VGND.n1597 VGND.n798 0.120125
R3700 VGND.n1597 VGND.n1596 0.120125
R3701 VGND.n2308 VGND.n2307 0.120125
R3702 VGND.n2307 VGND.n2306 0.120125
R3703 VGND.n2306 VGND.n2305 0.120125
R3704 VGND.n2305 VGND.n147 0.120125
R3705 VGND.n2121 VGND.n2120 0.120125
R3706 VGND.n2120 VGND.n2119 0.120125
R3707 VGND.n2119 VGND.n2118 0.120125
R3708 VGND.n2118 VGND.n2117 0.120125
R3709 VGND.n1906 VGND.n364 0.120125
R3710 VGND.n364 VGND.n363 0.120125
R3711 VGND.n363 VGND.n362 0.120125
R3712 VGND.n362 VGND.n361 0.120125
R3713 VGND.n144 VGND.n143 0.120125
R3714 VGND.n143 VGND.n53 0.120125
R3715 VGND.n2522 VGND.n53 0.120125
R3716 VGND.n2522 VGND.n2521 0.120125
R3717 VGND.n2042 VGND.n293 0.109992
R3718 VGND.n1235 VGND.n1042 0.10744
R3719 VGND.n2260 VGND.n88 0.103312
R3720 VGND.n2219 VGND.n109 0.103312
R3721 VGND.n2179 VGND.n128 0.103312
R3722 VGND.n2309 VGND.n146 0.103312
R3723 VGND.n2304 VGND.n2303 0.103312
R3724 VGND.n273 VGND.n55 0.103312
R3725 VGND.n1888 VGND.n373 0.102062
R3726 VGND.n1314 VGND.n923 0.102062
R3727 VGND.n1003 VGND.n914 0.102062
R3728 VGND.n1425 VGND.n850 0.102062
R3729 VGND.n1244 VGND.n1243 0.102062
R3730 VGND.n2360 VGND 0.0981562
R3731 VGND.n2374 VGND 0.0981562
R3732 VGND.n2440 VGND 0.0981562
R3733 VGND VGND.n63 0.0981562
R3734 VGND.n2186 VGND 0.0981562
R3735 VGND.n2200 VGND 0.0981562
R3736 VGND.n2248 VGND 0.0981562
R3737 VGND.n2265 VGND 0.0981562
R3738 VGND VGND.n2276 0.0981562
R3739 VGND.n1958 VGND 0.0981562
R3740 VGND.n1972 VGND 0.0981562
R3741 VGND.n2037 VGND 0.0981562
R3742 VGND VGND.n282 0.0981562
R3743 VGND VGND.n376 0.0981562
R3744 VGND.n1856 VGND 0.0981562
R3745 VGND.n1802 VGND 0.0981562
R3746 VGND VGND.n505 0.0981562
R3747 VGND.n1689 VGND 0.0981562
R3748 VGND VGND.n1357 0.0981562
R3749 VGND.n1007 VGND 0.0981562
R3750 VGND VGND.n1641 0.0981562
R3751 VGND.n1603 VGND 0.0981562
R3752 VGND VGND.n1027 0.0981562
R3753 VGND.n1135 VGND 0.0981562
R3754 VGND.n1109 VGND 0.0981562
R3755 VGND.n28 VGND 0.0981562
R3756 VGND.n2462 VGND.n2461 0.0968542
R3757 VGND.n222 VGND.n156 0.0968542
R3758 VGND.n2058 VGND.n2057 0.0968542
R3759 VGND.n530 VGND.n529 0.0968542
R3760 VGND VGND.n640 0.0968542
R3761 VGND VGND.n1346 0.0968542
R3762 VGND.n1541 VGND.n811 0.0968542
R3763 VGND.n2547 VGND.n2546 0.0968542
R3764 VGND.n1392 VGND 0.0955521
R3765 VGND VGND.n859 0.0955521
R3766 VGND.n1438 VGND 0.0955521
R3767 VGND VGND.n837 0.0955521
R3768 VGND.n1510 VGND 0.0955521
R3769 VGND VGND.n809 0.0955521
R3770 VGND VGND.n1585 0.0955521
R3771 VGND.n2563 VGND 0.0955521
R3772 VGND.n1381 VGND.n1380 0.0950946
R3773 VGND.n1386 VGND.n1385 0.0950946
R3774 VGND.n1726 VGND.n1725 0.0950946
R3775 VGND.n1734 VGND.n611 0.0950946
R3776 VGND.n1079 VGND.n1078 0.0950946
R3777 VGND.n1125 VGND.n1077 0.0950946
R3778 VGND.n1102 VGND.n1101 0.0950946
R3779 VGND.n2548 VGND.n44 0.0950946
R3780 VGND.n2553 VGND.n5 0.0950946
R3781 VGND.n40 VGND.n9 0.0950946
R3782 VGND.n1059 VGND.n1049 0.0950946
R3783 VGND.n1155 VGND.n1044 0.0950946
R3784 VGND.n1189 VGND.n1037 0.0950946
R3785 VGND.n1242 VGND.n1034 0.0950946
R3786 VGND.n1171 VGND.n1165 0.0950946
R3787 VGND.n1227 VGND.n1161 0.0950946
R3788 VGND.n2449 VGND.n2447 0.0950946
R3789 VGND.n2460 VGND.n71 0.0950946
R3790 VGND.n2383 VGND.n2382 0.0950946
R3791 VGND.n2387 VGND.n106 0.0950946
R3792 VGND.n2351 VGND.n2350 0.0950946
R3793 VGND.n2355 VGND.n125 0.0950946
R3794 VGND.n2321 VGND.n2320 0.0950946
R3795 VGND.n2325 VGND.n141 0.0950946
R3796 VGND.n2517 VGND.n2516 0.0950946
R3797 VGND.n2508 VGND.n2507 0.0950946
R3798 VGND.n2419 VGND.n2418 0.0950946
R3799 VGND.n2423 VGND.n85 0.0950946
R3800 VGND.n2177 VGND.n2176 0.0950946
R3801 VGND.n2181 VGND.n203 0.0950946
R3802 VGND.n2141 VGND.n2140 0.0950946
R3803 VGND.n2151 VGND.n2135 0.0950946
R3804 VGND.n271 VGND.n270 0.0950946
R3805 VGND.n263 VGND.n262 0.0950946
R3806 VGND.n2301 VGND.n2300 0.0950946
R3807 VGND.n2294 VGND.n155 0.0950946
R3808 VGND.n2217 VGND.n2216 0.0950946
R3809 VGND.n2221 VGND.n188 0.0950946
R3810 VGND.n2258 VGND.n2257 0.0950946
R3811 VGND.n2262 VGND.n168 0.0950946
R3812 VGND.n1942 VGND.n1940 0.0950946
R3813 VGND.n1953 VGND.n345 0.0950946
R3814 VGND.n1919 VGND.n1918 0.0950946
R3815 VGND.n1923 VGND.n358 0.0950946
R3816 VGND.n2113 VGND.n2112 0.0950946
R3817 VGND.n2105 VGND.n2104 0.0950946
R3818 VGND.n2052 VGND.n2051 0.0950946
R3819 VGND.n2056 VGND.n289 0.0950946
R3820 VGND.n1981 VGND.n1980 0.0950946
R3821 VGND.n1985 VGND.n327 0.0950946
R3822 VGND.n2017 VGND.n2016 0.0950946
R3823 VGND.n2021 VGND.n307 0.0950946
R3824 VGND.n392 VGND.n390 0.0950946
R3825 VGND.n401 VGND.n382 0.0950946
R3826 VGND.n590 VGND.n589 0.0950946
R3827 VGND.n582 VGND.n581 0.0950946
R3828 VGND.n1800 VGND.n491 0.0950946
R3829 VGND.n528 VGND.n527 0.0950946
R3830 VGND.n448 VGND.n447 0.0950946
R3831 VGND.n1862 VGND.n444 0.0950946
R3832 VGND.n1902 VGND.n1901 0.0950946
R3833 VGND.n1895 VGND.n372 0.0950946
R3834 VGND.n473 VGND.n472 0.0950946
R3835 VGND.n1827 VGND.n470 0.0950946
R3836 VGND.n1696 VGND.n1695 0.0950946
R3837 VGND.n1700 VGND.n624 0.0950946
R3838 VGND.n1633 VGND.n677 0.0950946
R3839 VGND.n1628 VGND.n680 0.0950946
R3840 VGND.n1490 VGND.n1489 0.0950946
R3841 VGND.n1494 VGND.n825 0.0950946
R3842 VGND.n1662 VGND.n1661 0.0950946
R3843 VGND.n666 VGND.n665 0.0950946
R3844 VGND.n1457 VGND.n1456 0.0950946
R3845 VGND.n1461 VGND.n840 0.0950946
R3846 VGND.n1284 VGND.n1277 0.0950946
R3847 VGND.n1667 VGND.n644 0.0950946
R3848 VGND.n953 VGND.n940 0.0950946
R3849 VGND.n948 VGND.n945 0.0950946
R3850 VGND.n1791 VGND.n1790 0.0950946
R3851 VGND.n1781 VGND.n1780 0.0950946
R3852 VGND.n1326 VGND.n1325 0.0950946
R3853 VGND.n1319 VGND.n922 0.0950946
R3854 VGND.n1334 VGND.n1333 0.0950946
R3855 VGND.n1339 VGND.n1338 0.0950946
R3856 VGND.n1420 VGND.n1419 0.0950946
R3857 VGND.n1424 VGND.n852 0.0950946
R3858 VGND.n892 VGND.n891 0.0950946
R3859 VGND.n1365 VGND.n879 0.0950946
R3860 VGND.n769 VGND.n729 0.0950946
R3861 VGND.n764 VGND.n732 0.0950946
R3862 VGND.n1601 VGND.n700 0.0950946
R3863 VGND.n795 VGND.n703 0.0950946
R3864 VGND.n1526 VGND.n1525 0.0950946
R3865 VGND.n1532 VGND.n1531 0.0950946
R3866 VGND.n1562 VGND.n806 0.0950946
R3867 VGND.n1592 VGND.n802 0.0950946
R3868 VGND.n2481 VGND.n57 0.0916458
R3869 VGND.n215 VGND.n209 0.0916458
R3870 VGND.n554 VGND.n498 0.0916458
R3871 VGND.n1756 VGND.n596 0.0916458
R3872 VGND.n2555 VGND.n2554 0.0916458
R3873 VGND.n2260 VGND.n170 0.0915625
R3874 VGND.n2219 VGND.n190 0.0915625
R3875 VGND.n2179 VGND.n2122 0.0915625
R3876 VGND.n206 VGND.n146 0.0915625
R3877 VGND.n2303 VGND.n149 0.0915625
R3878 VGND.n2116 VGND.n273 0.0915625
R3879 VGND.n2476 VGND.n2475 0.0900105
R3880 VGND.n2060 VGND.n2059 0.0900105
R3881 VGND.n1236 VGND.n1235 0.0898892
R3882 VGND.n1234 VGND.n1231 0.0898892
R3883 VGND.n2378 VGND.n111 0.0864375
R3884 VGND.n2205 VGND.n192 0.0864375
R3885 VGND.n1976 VGND.n331 0.0864375
R3886 VGND.n1275 VGND.n1267 0.0864375
R3887 VGND.n1444 VGND.n843 0.0864375
R3888 VGND.n1056 VGND.n1055 0.0864375
R3889 VGND.n2349 VGND.n2348 0.0838333
R3890 VGND.n113 VGND.n105 0.0838333
R3891 VGND.n2424 VGND.n84 0.0838333
R3892 VGND.n2455 VGND.n74 0.0838333
R3893 VGND.n2486 VGND.n60 0.0838333
R3894 VGND.n2175 VGND.n2174 0.0838333
R3895 VGND.n2212 VGND.n187 0.0838333
R3896 VGND.n2256 VGND.n172 0.0838333
R3897 VGND.n2263 VGND.n167 0.0838333
R3898 VGND.n241 VGND.n212 0.0838333
R3899 VGND.n1948 VGND.n348 0.0838333
R3900 VGND.n333 VGND.n326 0.0838333
R3901 VGND.n2022 VGND.n306 0.0838333
R3902 VGND.n2084 VGND.n280 0.0838333
R3903 VGND.n1900 VGND.n1899 0.0838333
R3904 VGND.n1867 VGND.n442 0.0838333
R3905 VGND.n467 VGND.n464 0.0838333
R3906 VGND.n1826 VGND.n476 0.0838333
R3907 VGND.n520 VGND.n517 0.0838333
R3908 VGND.n559 VGND.n501 0.0838333
R3909 VGND.n1324 VGND.n1323 0.0838333
R3910 VGND.n1280 VGND.n1279 0.0838333
R3911 VGND.n1694 VGND.n629 0.0838333
R3912 VGND.n1701 VGND.n623 0.0838333
R3913 VGND.n1729 VGND.n1727 0.0838333
R3914 VGND.n1332 VGND.n911 0.0838333
R3915 VGND.n664 VGND.n655 0.0838333
R3916 VGND.n1627 VGND.n681 0.0838333
R3917 VGND.n714 VGND.n710 0.0838333
R3918 VGND.n1453 VGND.n1450 0.0838333
R3919 VGND.n1524 VGND.n1523 0.0838333
R3920 VGND.n1195 VGND.n1190 0.0838333
R3921 VGND.n1063 VGND.n1048 0.0838333
R3922 VGND.n1074 VGND.n1072 0.0838333
R3923 VGND.n1124 VGND.n1083 0.0838333
R3924 VGND.n2530 VGND.n48 0.0838333
R3925 VGND.n16 VGND.n14 0.0838333
R3926 VGND.n1795 VGND 0.0827875
R3927 VGND.n1596 VGND 0.0827875
R3928 VGND.n147 VGND 0.0827875
R3929 VGND.n2117 VGND 0.0827875
R3930 VGND.n361 VGND 0.0827875
R3931 VGND.n2521 VGND 0.0827875
R3932 VGND VGND.n1764 0.082648
R3933 VGND VGND.n963 0.082648
R3934 VGND VGND.n805 0.0773229
R3935 VGND.n132 VGND.n130 0.0760208
R3936 VGND.n2126 VGND.n2124 0.0760208
R3937 VGND.n1944 VGND.n1943 0.0760208
R3938 VGND.n370 VGND.n368 0.0760208
R3939 VGND.n920 VGND.n918 0.0760208
R3940 VGND.n909 VGND.n907 0.0760208
R3941 VGND.n1412 VGND.n856 0.0760208
R3942 VGND.n1201 VGND.n1200 0.0760208
R3943 VGND.n2317 VGND.n2314 0.0708125
R3944 VGND.n2381 VGND.n102 0.0708125
R3945 VGND.n2451 VGND.n2450 0.0708125
R3946 VGND.n2146 VGND.n2145 0.0708125
R3947 VGND.n2215 VGND.n2214 0.0708125
R3948 VGND.n153 VGND.n151 0.0708125
R3949 VGND.n1915 VGND.n1912 0.0708125
R3950 VGND.n1979 VGND.n323 0.0708125
R3951 VGND.n295 VGND.n293 0.0708125
R3952 VGND.n396 VGND.n395 0.0708125
R3953 VGND.n1868 VGND.n441 0.0708125
R3954 VGND.n1801 VGND.n490 0.0708125
R3955 VGND.n942 VGND.n937 0.0708125
R3956 VGND.n1285 VGND.n1276 0.0708125
R3957 VGND.n1723 VGND.n614 0.0708125
R3958 VGND.n886 VGND.n883 0.0708125
R3959 VGND.n1660 VGND.n1659 0.0708125
R3960 VGND.n1388 VGND.n869 0.0708125
R3961 VGND.n1455 VGND.n1454 0.0708125
R3962 VGND.n1521 VGND.n818 0.0708125
R3963 VGND.n1178 VGND.n1176 0.0708125
R3964 VGND.n1103 VGND.n1100 0.0708125
R3965 VGND.n2417 VGND 0.0695104
R3966 VGND.n2015 VGND 0.0695104
R3967 VGND.n2019 VGND.n170 0.0692375
R3968 VGND.n1983 VGND.n190 0.0692375
R3969 VGND.n2122 VGND.n205 0.0692375
R3970 VGND.n1921 VGND.n206 0.0692375
R3971 VGND.n2054 VGND.n149 0.0692375
R3972 VGND.n2116 VGND.n2115 0.0692375
R3973 VGND.n1814 VGND.n1813 0.0685851
R3974 VGND.n95 VGND.n90 0.068325
R3975 VGND.n316 VGND.n311 0.068325
R3976 VGND.n1374 VGND.n1373 0.0680676
R3977 VGND.n1373 VGND.n870 0.0680676
R3978 VGND.n1730 VGND.n613 0.0680676
R3979 VGND.n1731 VGND.n1730 0.0680676
R3980 VGND.n1129 VGND.n1076 0.0680676
R3981 VGND.n1129 VGND.n1128 0.0680676
R3982 VGND.n2529 VGND.n49 0.0680676
R3983 VGND.n2529 VGND.n2528 0.0680676
R3984 VGND.n15 VGND.n7 0.0680676
R3985 VGND.n15 VGND.n8 0.0680676
R3986 VGND.n1062 VGND.n1060 0.0680676
R3987 VGND.n1062 VGND.n1061 0.0680676
R3988 VGND.n1194 VGND.n1038 0.0680676
R3989 VGND.n1194 VGND.n1193 0.0680676
R3990 VGND.n1175 VGND.n1173 0.0680676
R3991 VGND.n1175 VGND.n1174 0.0680676
R3992 VGND.n2456 VGND.n73 0.0680676
R3993 VGND.n2457 VGND.n2456 0.0680676
R3994 VGND.n115 VGND.n114 0.0680676
R3995 VGND.n114 VGND.n112 0.0680676
R3996 VGND.n2347 VGND.n131 0.0680676
R3997 VGND.n2347 VGND.n2346 0.0680676
R3998 VGND.n2316 VGND.n2312 0.0680676
R3999 VGND.n2316 VGND.n2315 0.0680676
R4000 VGND.n2504 VGND.n58 0.0680676
R4001 VGND.n2506 VGND.n2504 0.0680676
R4002 VGND.n93 VGND.n91 0.0680676
R4003 VGND.n93 VGND.n92 0.0680676
R4004 VGND.n2173 VGND.n2125 0.0680676
R4005 VGND.n2173 VGND.n2172 0.0680676
R4006 VGND.n2147 VGND.n2137 0.0680676
R4007 VGND.n2148 VGND.n2147 0.0680676
R4008 VGND.n259 VGND.n210 0.0680676
R4009 VGND.n261 VGND.n259 0.0680676
R4010 VGND.n2297 VGND.n152 0.0680676
R4011 VGND.n2297 VGND.n2296 0.0680676
R4012 VGND.n2211 VGND.n193 0.0680676
R4013 VGND.n2211 VGND.n2210 0.0680676
R4014 VGND.n175 VGND.n173 0.0680676
R4015 VGND.n175 VGND.n174 0.0680676
R4016 VGND.n1949 VGND.n347 0.0680676
R4017 VGND.n1950 VGND.n1949 0.0680676
R4018 VGND.n1914 VGND.n1910 0.0680676
R4019 VGND.n1914 VGND.n1913 0.0680676
R4020 VGND.n2101 VGND.n278 0.0680676
R4021 VGND.n2103 VGND.n2101 0.0680676
R4022 VGND.n2048 VGND.n294 0.0680676
R4023 VGND.n2048 VGND.n2047 0.0680676
R4024 VGND.n335 VGND.n334 0.0680676
R4025 VGND.n334 VGND.n332 0.0680676
R4026 VGND.n314 VGND.n312 0.0680676
R4027 VGND.n314 VGND.n313 0.0680676
R4028 VGND.n397 VGND.n384 0.0680676
R4029 VGND.n398 VGND.n397 0.0680676
R4030 VGND.n578 VGND.n499 0.0680676
R4031 VGND.n580 VGND.n578 0.0680676
R4032 VGND.n519 VGND.n518 0.0680676
R4033 VGND.n519 VGND.n516 0.0680676
R4034 VGND.n1866 VGND.n443 0.0680676
R4035 VGND.n1866 VGND.n1865 0.0680676
R4036 VGND.n1898 VGND.n369 0.0680676
R4037 VGND.n1898 VGND.n1897 0.0680676
R4038 VGND.n1831 VGND.n469 0.0680676
R4039 VGND.n1831 VGND.n1830 0.0680676
R4040 VGND.n633 VGND.n630 0.0680676
R4041 VGND.n633 VGND.n632 0.0680676
R4042 VGND.n688 VGND.n678 0.0680676
R4043 VGND.n688 VGND.n679 0.0680676
R4044 VGND.n832 VGND.n830 0.0680676
R4045 VGND.n832 VGND.n831 0.0680676
R4046 VGND.n661 VGND.n653 0.0680676
R4047 VGND.n663 VGND.n661 0.0680676
R4048 VGND.n1452 VGND.n844 0.0680676
R4049 VGND.n1452 VGND.n1451 0.0680676
R4050 VGND.n1283 VGND.n1281 0.0680676
R4051 VGND.n1281 VGND.n1278 0.0680676
R4052 VGND.n943 VGND.n941 0.0680676
R4053 VGND.n944 VGND.n943 0.0680676
R4054 VGND.n1777 VGND.n597 0.0680676
R4055 VGND.n1779 VGND.n1777 0.0680676
R4056 VGND.n1322 VGND.n919 0.0680676
R4057 VGND.n1322 VGND.n1321 0.0680676
R4058 VGND.n1331 VGND.n1330 0.0680676
R4059 VGND.n1330 VGND.n913 0.0680676
R4060 VGND.n1416 VGND.n857 0.0680676
R4061 VGND.n1416 VGND.n1415 0.0680676
R4062 VGND.n889 VGND.n887 0.0680676
R4063 VGND.n887 VGND.n885 0.0680676
R4064 VGND.n742 VGND.n730 0.0680676
R4065 VGND.n742 VGND.n731 0.0680676
R4066 VGND.n713 VGND.n711 0.0680676
R4067 VGND.n713 VGND.n712 0.0680676
R4068 VGND.n1522 VGND.n817 0.0680676
R4069 VGND.n1522 VGND.n816 0.0680676
R4070 VGND.n1566 VGND.n1564 0.0680676
R4071 VGND.n1566 VGND.n1565 0.0680676
R4072 VGND.n1488 VGND 0.0669062
R4073 VGND.n2357 VGND.n124 0.0656042
R4074 VGND.n2412 VGND.n94 0.0656042
R4075 VGND.n2515 VGND.n2514 0.0656042
R4076 VGND.n2183 VGND.n202 0.0656042
R4077 VGND.n2252 VGND.n176 0.0656042
R4078 VGND.n269 VGND.n268 0.0656042
R4079 VGND.n1955 VGND.n344 0.0656042
R4080 VGND.n2010 VGND.n315 0.0656042
R4081 VGND.n2111 VGND.n2110 0.0656042
R4082 VGND.n2107 VGND.n2106 0.0656042
R4083 VGND.n1894 VGND.n1893 0.0656042
R4084 VGND.n1832 VGND.n468 0.0656042
R4085 VGND.n588 VGND.n587 0.0656042
R4086 VGND.n584 VGND.n583 0.0656042
R4087 VGND.n1318 VGND.n1317 0.0656042
R4088 VGND.n634 VGND.n631 0.0656042
R4089 VGND.n1789 VGND.n1788 0.0656042
R4090 VGND.n1783 VGND.n1782 0.0656042
R4091 VGND.n1340 VGND.n912 0.0656042
R4092 VGND.n690 VGND.n689 0.0656042
R4093 VGND.n744 VGND.n740 0.0656042
R4094 VGND.n763 VGND.n733 0.0656042
R4095 VGND.n1484 VGND.n833 0.0656042
R4096 VGND.n1591 VGND.n803 0.0656042
R4097 VGND.n1196 VGND.n1033 0.0656042
R4098 VGND.n1130 VGND.n1075 0.0656042
R4099 VGND.n17 VGND.n13 0.0656042
R4100 VGND.n39 VGND.n10 0.0656042
R4101 VGND.n2319 VGND 0.0643021
R4102 VGND.n2142 VGND 0.0643021
R4103 VGND.n1917 VGND 0.0643021
R4104 VGND.n389 VGND 0.0643021
R4105 VGND.n939 VGND 0.0643021
R4106 VGND.n890 VGND 0.0643021
R4107 VGND VGND.n652 0.0643021
R4108 VGND.n1379 VGND 0.0643021
R4109 VGND.n1170 VGND 0.0643021
R4110 VGND.n2331 VGND 0.0603958
R4111 VGND.n2340 VGND 0.0603958
R4112 VGND.n2377 VGND 0.0603958
R4113 VGND.n2378 VGND 0.0603958
R4114 VGND VGND.n101 0.0603958
R4115 VGND.n2441 VGND 0.0603958
R4116 VGND.n2445 VGND 0.0603958
R4117 VGND.n2454 VGND.n75 0.0603958
R4118 VGND.n75 VGND.n70 0.0603958
R4119 VGND VGND.n2502 0.0603958
R4120 VGND.n2157 VGND 0.0603958
R4121 VGND.n2166 VGND 0.0603958
R4122 VGND.n2204 VGND 0.0603958
R4123 VGND.n2223 VGND.n2222 0.0603958
R4124 VGND.n2222 VGND.n183 0.0603958
R4125 VGND.n2233 VGND 0.0603958
R4126 VGND.n2283 VGND 0.0603958
R4127 VGND.n2293 VGND.n2292 0.0603958
R4128 VGND.n265 VGND 0.0603958
R4129 VGND VGND.n257 0.0603958
R4130 VGND.n251 VGND 0.0603958
R4131 VGND VGND.n250 0.0603958
R4132 VGND.n1929 VGND 0.0603958
R4133 VGND.n1939 VGND 0.0603958
R4134 VGND.n1975 VGND 0.0603958
R4135 VGND.n1976 VGND 0.0603958
R4136 VGND VGND.n322 0.0603958
R4137 VGND.n2041 VGND 0.0603958
R4138 VGND.n2046 VGND.n296 0.0603958
R4139 VGND.n296 VGND.n288 0.0603958
R4140 VGND VGND.n286 0.0603958
R4141 VGND.n2071 VGND 0.0603958
R4142 VGND.n2079 VGND 0.0603958
R4143 VGND.n404 VGND 0.0603958
R4144 VGND.n408 VGND 0.0603958
R4145 VGND.n416 VGND 0.0603958
R4146 VGND VGND.n421 0.0603958
R4147 VGND.n422 VGND 0.0603958
R4148 VGND VGND.n1887 0.0603958
R4149 VGND.n1874 VGND 0.0603958
R4150 VGND VGND.n1873 0.0603958
R4151 VGND VGND.n451 0.0603958
R4152 VGND VGND.n1861 0.0603958
R4153 VGND VGND.n477 0.0603958
R4154 VGND.n480 VGND 0.0603958
R4155 VGND VGND.n480 0.0603958
R4156 VGND.n1820 VGND 0.0603958
R4157 VGND VGND.n1819 0.0603958
R4158 VGND VGND.n1810 0.0603958
R4159 VGND VGND.n1809 0.0603958
R4160 VGND.n489 VGND 0.0603958
R4161 VGND.n526 VGND.n525 0.0603958
R4162 VGND.n526 VGND.n514 0.0603958
R4163 VGND.n577 VGND 0.0603958
R4164 VGND.n573 VGND 0.0603958
R4165 VGND.n964 VGND 0.0603958
R4166 VGND.n979 VGND 0.0603958
R4167 VGND.n1301 VGND 0.0603958
R4168 VGND.n1293 VGND 0.0603958
R4169 VGND VGND.n1292 0.0603958
R4170 VGND.n1668 VGND.n643 0.0603958
R4171 VGND.n1669 VGND.n1668 0.0603958
R4172 VGND.n1670 VGND 0.0603958
R4173 VGND VGND.n1684 0.0603958
R4174 VGND.n1685 VGND 0.0603958
R4175 VGND.n1690 VGND 0.0603958
R4176 VGND VGND.n1708 0.0603958
R4177 VGND.n1709 VGND 0.0603958
R4178 VGND.n1714 VGND 0.0603958
R4179 VGND.n1715 VGND 0.0603958
R4180 VGND.n1728 VGND.n610 0.0603958
R4181 VGND.n1736 VGND.n610 0.0603958
R4182 VGND VGND.n608 0.0603958
R4183 VGND.n1756 VGND 0.0603958
R4184 VGND.n1765 VGND 0.0603958
R4185 VGND.n1358 VGND 0.0603958
R4186 VGND.n899 VGND 0.0603958
R4187 VGND VGND.n904 0.0603958
R4188 VGND.n1347 VGND 0.0603958
R4189 VGND VGND.n1003 0.0603958
R4190 VGND.n1004 VGND 0.0603958
R4191 VGND VGND.n998 0.0603958
R4192 VGND VGND.n1017 0.0603958
R4193 VGND.n1022 VGND 0.0603958
R4194 VGND VGND.n1021 0.0603958
R4195 VGND.n1018 VGND 0.0603958
R4196 VGND.n667 VGND.n658 0.0603958
R4197 VGND.n1655 VGND.n667 0.0603958
R4198 VGND.n1653 VGND 0.0603958
R4199 VGND.n668 VGND 0.0603958
R4200 VGND VGND.n1648 0.0603958
R4201 VGND.n1642 VGND 0.0603958
R4202 VGND VGND.n1620 0.0603958
R4203 VGND VGND.n1612 0.0603958
R4204 VGND.n1609 VGND 0.0603958
R4205 VGND VGND.n1608 0.0603958
R4206 VGND.n709 VGND 0.0603958
R4207 VGND.n716 VGND.n715 0.0603958
R4208 VGND.n715 VGND.n704 0.0603958
R4209 VGND VGND.n793 0.0603958
R4210 VGND VGND.n779 0.0603958
R4211 VGND.n1393 VGND 0.0603958
R4212 VGND VGND.n863 0.0603958
R4213 VGND.n1399 VGND 0.0603958
R4214 VGND.n1408 VGND 0.0603958
R4215 VGND.n1426 VGND 0.0603958
R4216 VGND.n1435 VGND 0.0603958
R4217 VGND VGND.n1439 0.0603958
R4218 VGND.n1440 VGND 0.0603958
R4219 VGND.n1443 VGND 0.0603958
R4220 VGND.n1462 VGND.n839 0.0603958
R4221 VGND.n1463 VGND.n1462 0.0603958
R4222 VGND.n1464 VGND 0.0603958
R4223 VGND VGND.n1469 0.0603958
R4224 VGND.n1470 VGND 0.0603958
R4225 VGND.n1471 VGND 0.0603958
R4226 VGND.n1480 VGND 0.0603958
R4227 VGND.n1497 VGND 0.0603958
R4228 VGND.n1506 VGND 0.0603958
R4229 VGND VGND.n1511 0.0603958
R4230 VGND.n1512 VGND 0.0603958
R4231 VGND.n1516 VGND 0.0603958
R4232 VGND.n1533 VGND.n815 0.0603958
R4233 VGND.n1534 VGND.n1533 0.0603958
R4234 VGND.n1543 VGND 0.0603958
R4235 VGND VGND.n1548 0.0603958
R4236 VGND.n1549 VGND 0.0603958
R4237 VGND.n1550 VGND 0.0603958
R4238 VGND.n1568 VGND 0.0603958
R4239 VGND.n1590 VGND 0.0603958
R4240 VGND.n1587 VGND 0.0603958
R4241 VGND VGND.n1586 0.0603958
R4242 VGND VGND.n1573 0.0603958
R4243 VGND.n1581 VGND 0.0603958
R4244 VGND VGND.n1217 0.0603958
R4245 VGND VGND.n1202 0.0603958
R4246 VGND.n1050 VGND 0.0603958
R4247 VGND.n1064 VGND 0.0603958
R4248 VGND.n1154 VGND.n1045 0.0603958
R4249 VGND.n1154 VGND.n1153 0.0603958
R4250 VGND VGND.n1108 0.0603958
R4251 VGND.n1104 VGND 0.0603958
R4252 VGND.n2532 VGND.n2531 0.0603958
R4253 VGND.n2531 VGND.n45 0.0603958
R4254 VGND VGND.n2567 0.0603958
R4255 VGND.n2562 VGND 0.0603958
R4256 VGND VGND.n2561 0.0603958
R4257 VGND.n2421 VGND.n88 0.0574875
R4258 VGND.n2385 VGND.n109 0.0574875
R4259 VGND.n2353 VGND.n128 0.0574875
R4260 VGND.n2323 VGND.n2309 0.0574875
R4261 VGND.n2304 VGND.n52 0.0574875
R4262 VGND.n2519 VGND.n55 0.0574875
R4263 VGND.n1371 VGND.n871 0.0574697
R4264 VGND.n1732 VGND.n612 0.0574697
R4265 VGND.n2458 VGND.n72 0.0574697
R4266 VGND.n110 VGND.n107 0.0574697
R4267 VGND.n129 VGND.n126 0.0574697
R4268 VGND.n2310 VGND.n142 0.0574697
R4269 VGND.n2505 VGND.n56 0.0574697
R4270 VGND.n89 VGND.n86 0.0574697
R4271 VGND.n2123 VGND.n204 0.0574697
R4272 VGND.n2149 VGND.n2136 0.0574697
R4273 VGND.n260 VGND.n208 0.0574697
R4274 VGND.n2295 VGND.n150 0.0574697
R4275 VGND.n191 VGND.n189 0.0574697
R4276 VGND.n171 VGND.n169 0.0574697
R4277 VGND.n1951 VGND.n346 0.0574697
R4278 VGND.n1908 VGND.n359 0.0574697
R4279 VGND.n2102 VGND.n276 0.0574697
R4280 VGND.n292 VGND.n290 0.0574697
R4281 VGND.n330 VGND.n328 0.0574697
R4282 VGND.n310 VGND.n308 0.0574697
R4283 VGND.n399 VGND.n383 0.0574697
R4284 VGND.n579 VGND.n497 0.0574697
R4285 VGND.n515 VGND.n492 0.0574697
R4286 VGND.n1864 VGND.n445 0.0574697
R4287 VGND.n1896 VGND.n367 0.0574697
R4288 VGND.n1829 VGND.n471 0.0574697
R4289 VGND.n628 VGND.n625 0.0574697
R4290 VGND.n1631 VGND.n1630 0.0574697
R4291 VGND.n828 VGND.n826 0.0574697
R4292 VGND.n662 VGND.n651 0.0574697
R4293 VGND.n842 VGND.n841 0.0574697
R4294 VGND.n1282 VGND.n648 0.0574697
R4295 VGND.n1666 VGND.n645 0.0574697
R4296 VGND.n951 VGND.n950 0.0574697
R4297 VGND.n1778 VGND.n595 0.0574697
R4298 VGND.n1320 VGND.n917 0.0574697
R4299 VGND.n1329 VGND.n915 0.0574697
R4300 VGND.n855 VGND.n853 0.0574697
R4301 VGND.n888 VGND.n877 0.0574697
R4302 VGND.n1366 VGND.n878 0.0574697
R4303 VGND.n767 VGND.n766 0.0574697
R4304 VGND.n702 VGND.n701 0.0574697
R4305 VGND.n1529 VGND.n1528 0.0574697
R4306 VGND.n1563 VGND.n800 0.0574697
R4307 VGND.n1593 VGND.n801 0.0574697
R4308 VGND.n2345 VGND.n124 0.0551875
R4309 VGND.n2416 VGND.n94 0.0551875
R4310 VGND.n2515 VGND.n59 0.0551875
R4311 VGND.n2509 VGND.n2503 0.0551875
R4312 VGND.n2171 VGND.n202 0.0551875
R4313 VGND.n2255 VGND.n176 0.0551875
R4314 VGND.n269 VGND.n211 0.0551875
R4315 VGND.n264 VGND.n258 0.0551875
R4316 VGND.n1947 VGND.n344 0.0551875
R4317 VGND.n2014 VGND.n315 0.0551875
R4318 VGND.n2111 VGND.n279 0.0551875
R4319 VGND.n2106 VGND.n2100 0.0551875
R4320 VGND.n1833 VGND.n1832 0.0551875
R4321 VGND.n588 VGND.n500 0.0551875
R4322 VGND.n583 VGND.n577 0.0551875
R4323 VGND.n1318 VGND.n921 0.0551875
R4324 VGND.n1693 VGND.n634 0.0551875
R4325 VGND.n1789 VGND.n598 0.0551875
R4326 VGND.n1782 VGND.n1776 0.0551875
R4327 VGND.n1341 VGND.n1340 0.0551875
R4328 VGND.n689 VGND.n687 0.0551875
R4329 VGND.n740 VGND.n728 0.0551875
R4330 VGND.n763 VGND.n762 0.0551875
R4331 VGND.n1487 VGND.n833 0.0551875
R4332 VGND.n1591 VGND.n1590 0.0551875
R4333 VGND.n1197 VGND.n1196 0.0551875
R4334 VGND.n1131 VGND.n1130 0.0551875
R4335 VGND.n13 VGND.n4 0.0551875
R4336 VGND.n39 VGND.n38 0.0551875
R4337 VGND.n1634 VGND 0.0525833
R4338 VGND.n1418 VGND 0.0525833
R4339 VGND.n2318 VGND.n2317 0.0499792
R4340 VGND.n2450 VGND.n2446 0.0499792
R4341 VGND.n2146 VGND.n2143 0.0499792
R4342 VGND.n2285 VGND.n151 0.0499792
R4343 VGND.n1916 VGND.n1915 0.0499792
R4344 VGND.n396 VGND.n385 0.0499792
R4345 VGND.n1802 VGND.n1801 0.0499792
R4346 VGND.n942 VGND.n938 0.0499792
R4347 VGND.n1286 VGND.n1285 0.0499792
R4348 VGND.n1723 VGND.n1722 0.0499792
R4349 VGND.n886 VGND.n884 0.0499792
R4350 VGND.n1660 VGND.n654 0.0499792
R4351 VGND.n1378 VGND.n869 0.0499792
R4352 VGND.n1455 VGND.n1449 0.0499792
R4353 VGND.n1518 VGND.n818 0.0499792
R4354 VGND.n1176 VGND.n1164 0.0499792
R4355 VGND.n1104 VGND.n1103 0.0499792
R4356 VGND.n2313 VGND 0.047375
R4357 VGND.n2144 VGND 0.047375
R4358 VGND.n1911 VGND 0.047375
R4359 VGND.n386 VGND 0.047375
R4360 VGND VGND.n946 0.047375
R4361 VGND.n882 VGND 0.047375
R4362 VGND.n1387 VGND 0.047375
R4363 VGND.n1177 VGND 0.047375
R4364 VGND.n2340 VGND.n130 0.0447708
R4365 VGND.n2166 VGND.n2124 0.0447708
R4366 VGND.n1943 VGND.n1939 0.0447708
R4367 VGND.n423 VGND.n368 0.0447708
R4368 VGND.n980 VGND.n918 0.0447708
R4369 VGND.n1345 VGND.n907 0.0447708
R4370 VGND.n859 VGND.n856 0.0447708
R4371 VGND.n1202 VGND.n1201 0.0447708
R4372 VGND.n1760 VGND 0.0421667
R4373 VGND VGND.n741 0.0421667
R4374 VGND.n1483 VGND 0.0421667
R4375 VGND.n1495 VGND 0.0421667
R4376 VGND.n1380 VGND.n1374 0.0410405
R4377 VGND.n1386 VGND.n870 0.0410405
R4378 VGND.n1726 VGND.n613 0.0410405
R4379 VGND.n1731 VGND.n611 0.0410405
R4380 VGND.n1078 VGND.n1076 0.0410405
R4381 VGND.n1128 VGND.n1077 0.0410405
R4382 VGND.n1101 VGND.n49 0.0410405
R4383 VGND.n2528 VGND.n44 0.0410405
R4384 VGND.n7 VGND.n5 0.0410405
R4385 VGND.n9 VGND.n8 0.0410405
R4386 VGND.n1060 VGND.n1059 0.0410405
R4387 VGND.n1061 VGND.n1044 0.0410405
R4388 VGND.n1189 VGND.n1038 0.0410405
R4389 VGND.n1193 VGND.n1034 0.0410405
R4390 VGND.n1173 VGND.n1171 0.0410405
R4391 VGND.n1174 VGND.n1161 0.0410405
R4392 VGND.n2447 VGND.n73 0.0410405
R4393 VGND.n2457 VGND.n71 0.0410405
R4394 VGND.n2382 VGND.n115 0.0410405
R4395 VGND.n112 VGND.n106 0.0410405
R4396 VGND.n2350 VGND.n131 0.0410405
R4397 VGND.n2346 VGND.n125 0.0410405
R4398 VGND.n2320 VGND.n2312 0.0410405
R4399 VGND.n2315 VGND.n141 0.0410405
R4400 VGND.n2516 VGND.n58 0.0410405
R4401 VGND.n2507 VGND.n2506 0.0410405
R4402 VGND.n2418 VGND.n91 0.0410405
R4403 VGND.n92 VGND.n85 0.0410405
R4404 VGND.n2176 VGND.n2125 0.0410405
R4405 VGND.n2172 VGND.n203 0.0410405
R4406 VGND.n2141 VGND.n2137 0.0410405
R4407 VGND.n2148 VGND.n2135 0.0410405
R4408 VGND.n270 VGND.n210 0.0410405
R4409 VGND.n262 VGND.n261 0.0410405
R4410 VGND.n2300 VGND.n152 0.0410405
R4411 VGND.n2296 VGND.n2294 0.0410405
R4412 VGND.n2216 VGND.n193 0.0410405
R4413 VGND.n2210 VGND.n188 0.0410405
R4414 VGND.n2257 VGND.n173 0.0410405
R4415 VGND.n174 VGND.n168 0.0410405
R4416 VGND.n1940 VGND.n347 0.0410405
R4417 VGND.n1950 VGND.n345 0.0410405
R4418 VGND.n1918 VGND.n1910 0.0410405
R4419 VGND.n1913 VGND.n358 0.0410405
R4420 VGND.n2112 VGND.n278 0.0410405
R4421 VGND.n2104 VGND.n2103 0.0410405
R4422 VGND.n2051 VGND.n294 0.0410405
R4423 VGND.n2047 VGND.n289 0.0410405
R4424 VGND.n1980 VGND.n335 0.0410405
R4425 VGND.n332 VGND.n327 0.0410405
R4426 VGND.n2016 VGND.n312 0.0410405
R4427 VGND.n313 VGND.n307 0.0410405
R4428 VGND.n390 VGND.n384 0.0410405
R4429 VGND.n398 VGND.n382 0.0410405
R4430 VGND.n589 VGND.n499 0.0410405
R4431 VGND.n581 VGND.n580 0.0410405
R4432 VGND.n518 VGND.n491 0.0410405
R4433 VGND.n527 VGND.n516 0.0410405
R4434 VGND.n447 VGND.n443 0.0410405
R4435 VGND.n1865 VGND.n444 0.0410405
R4436 VGND.n1901 VGND.n369 0.0410405
R4437 VGND.n1897 VGND.n1895 0.0410405
R4438 VGND.n472 VGND.n469 0.0410405
R4439 VGND.n1830 VGND.n470 0.0410405
R4440 VGND.n1695 VGND.n630 0.0410405
R4441 VGND.n632 VGND.n624 0.0410405
R4442 VGND.n678 VGND.n677 0.0410405
R4443 VGND.n680 VGND.n679 0.0410405
R4444 VGND.n1489 VGND.n830 0.0410405
R4445 VGND.n831 VGND.n825 0.0410405
R4446 VGND.n1661 VGND.n653 0.0410405
R4447 VGND.n665 VGND.n663 0.0410405
R4448 VGND.n1456 VGND.n844 0.0410405
R4449 VGND.n1451 VGND.n840 0.0410405
R4450 VGND.n1284 VGND.n1283 0.0410405
R4451 VGND.n1278 VGND.n644 0.0410405
R4452 VGND.n941 VGND.n940 0.0410405
R4453 VGND.n945 VGND.n944 0.0410405
R4454 VGND.n1790 VGND.n597 0.0410405
R4455 VGND.n1780 VGND.n1779 0.0410405
R4456 VGND.n1325 VGND.n919 0.0410405
R4457 VGND.n1321 VGND.n1319 0.0410405
R4458 VGND.n1333 VGND.n1331 0.0410405
R4459 VGND.n1339 VGND.n913 0.0410405
R4460 VGND.n1419 VGND.n857 0.0410405
R4461 VGND.n1415 VGND.n852 0.0410405
R4462 VGND.n891 VGND.n889 0.0410405
R4463 VGND.n885 VGND.n879 0.0410405
R4464 VGND.n730 VGND.n729 0.0410405
R4465 VGND.n732 VGND.n731 0.0410405
R4466 VGND.n711 VGND.n700 0.0410405
R4467 VGND.n712 VGND.n703 0.0410405
R4468 VGND.n1525 VGND.n817 0.0410405
R4469 VGND.n1532 VGND.n816 0.0410405
R4470 VGND.n1564 VGND.n1562 0.0410405
R4471 VGND.n1565 VGND.n802 0.0410405
R4472 VGND.n1233 VGND.n51 0.0393869
R4473 VGND.n2293 VGND 0.0382604
R4474 VGND.n2326 VGND 0.0369583
R4475 VGND.n2152 VGND 0.0369583
R4476 VGND VGND.n2298 0.0369583
R4477 VGND.n1924 VGND 0.0369583
R4478 VGND VGND.n2049 0.0369583
R4479 VGND.n402 VGND 0.0369583
R4480 VGND.n947 VGND 0.0369583
R4481 VGND.n1735 VGND 0.0369583
R4482 VGND.n1364 VGND 0.0369583
R4483 VGND.n794 VGND 0.0369583
R4484 VGND VGND.n867 0.0369583
R4485 VGND.n1226 VGND 0.0369583
R4486 VGND.n475 VGND.n309 0.0351625
R4487 VGND.n450 VGND.n329 0.0351625
R4488 VGND.n1905 VGND.n1904 0.0351625
R4489 VGND.n1907 VGND.n360 0.0351625
R4490 VGND.n1798 VGND.n291 0.0351625
R4491 VGND.n592 VGND.n275 0.0351625
R4492 VGND.n2319 VGND.n2318 0.0343542
R4493 VGND.n2380 VGND.n111 0.0343542
R4494 VGND.n2143 VGND.n2142 0.0343542
R4495 VGND.n2209 VGND.n192 0.0343542
R4496 VGND.n1917 VGND.n1916 0.0343542
R4497 VGND.n1978 VGND.n331 0.0343542
R4498 VGND.n389 VGND.n385 0.0343542
R4499 VGND.n404 VGND 0.0343542
R4500 VGND.n446 VGND.n437 0.0343542
R4501 VGND.n939 VGND.n938 0.0343542
R4502 VGND VGND.n962 0.0343542
R4503 VGND.n1286 VGND.n1275 0.0343542
R4504 VGND.n890 VGND.n884 0.0343542
R4505 VGND VGND.n880 0.0343542
R4506 VGND.n654 VGND.n652 0.0343542
R4507 VGND.n1649 VGND 0.0343542
R4508 VGND.n1609 VGND 0.0343542
R4509 VGND.n1379 VGND.n1378 0.0343542
R4510 VGND.n1449 VGND.n843 0.0343542
R4511 VGND.n1170 VGND.n1164 0.0343542
R4512 VGND.n1057 VGND.n1056 0.0343542
R4513 VGND.n1107 VGND 0.0343542
R4514 VGND.n827 VGND.n627 0.0339875
R4515 VGND.n1664 VGND.n650 0.0339875
R4516 VGND.n1336 VGND.n854 0.0339875
R4517 VGND.n1370 VGND.n1367 0.0339875
R4518 VGND.n1599 VGND.n1598 0.0339875
R4519 VGND.n1595 VGND.n594 0.0339875
R4520 VGND.n2374 VGND 0.0330521
R4521 VGND VGND.n2440 0.0330521
R4522 VGND.n2200 VGND 0.0330521
R4523 VGND.n2276 VGND 0.0330521
R4524 VGND.n1972 VGND 0.0330521
R4525 VGND.n2037 VGND 0.0330521
R4526 VGND.n1894 VGND 0.0330521
R4527 VGND.n1874 VGND 0.0330521
R4528 VGND.n1810 VGND 0.0330521
R4529 VGND.n1293 VGND 0.0330521
R4530 VGND.n1022 VGND 0.0330521
R4531 VGND.n1612 VGND 0.0330521
R4532 VGND.n1440 VGND 0.0330521
R4533 VGND.n1512 VGND 0.0330521
R4534 VGND.n1561 VGND 0.0330521
R4535 VGND VGND.n1027 0.0330521
R4536 VGND.n1109 VGND 0.0330521
R4537 VGND VGND.n2377 0.03175
R4538 VGND.n2503 VGND 0.03175
R4539 VGND VGND.n1975 0.03175
R4540 VGND.n2079 VGND 0.03175
R4541 VGND VGND.n277 0.03175
R4542 VGND VGND.n403 0.03175
R4543 VGND.n1820 VGND 0.03175
R4544 VGND.n1809 VGND 0.03175
R4545 VGND.n1021 VGND 0.03175
R4546 VGND.n686 VGND 0.03175
R4547 VGND VGND.n770 0.03175
R4548 VGND VGND.n1417 0.03175
R4549 VGND.n1414 VGND 0.03175
R4550 VGND VGND.n1470 0.03175
R4551 VGND VGND.n1496 0.03175
R4552 VGND VGND.n1549 0.03175
R4553 VGND.n1587 VGND 0.03175
R4554 VGND.n1491 VGND.n828 0.0292489
R4555 VGND.n1493 VGND.n826 0.0292489
R4556 VGND.n1632 VGND.n1631 0.0292489
R4557 VGND.n1630 VGND.n1629 0.0292489
R4558 VGND.n1697 VGND.n628 0.0292489
R4559 VGND.n1699 VGND.n625 0.0292489
R4560 VGND.n474 VGND.n471 0.0292489
R4561 VGND.n1829 VGND.n1828 0.0292489
R4562 VGND.n2018 VGND.n310 0.0292489
R4563 VGND.n2020 VGND.n308 0.0292489
R4564 VGND.n2259 VGND.n171 0.0292489
R4565 VGND.n2261 VGND.n169 0.0292489
R4566 VGND.n2420 VGND.n89 0.0292489
R4567 VGND.n2422 VGND.n86 0.0292489
R4568 VGND.n1458 VGND.n842 0.0292489
R4569 VGND.n1460 VGND.n841 0.0292489
R4570 VGND.n1663 VGND.n651 0.0292489
R4571 VGND.n662 VGND.n649 0.0292489
R4572 VGND.n449 VGND.n445 0.0292489
R4573 VGND.n1864 VGND.n1863 0.0292489
R4574 VGND.n1982 VGND.n330 0.0292489
R4575 VGND.n1984 VGND.n328 0.0292489
R4576 VGND.n2218 VGND.n191 0.0292489
R4577 VGND.n2220 VGND.n189 0.0292489
R4578 VGND.n2384 VGND.n110 0.0292489
R4579 VGND.n2386 VGND.n107 0.0292489
R4580 VGND.n647 VGND.n645 0.0292489
R4581 VGND.n1282 VGND.n647 0.0292489
R4582 VGND.n1421 VGND.n855 0.0292489
R4583 VGND.n1423 VGND.n853 0.0292489
R4584 VGND.n1335 VGND.n1329 0.0292489
R4585 VGND.n1337 VGND.n915 0.0292489
R4586 VGND.n1327 VGND.n917 0.0292489
R4587 VGND.n1320 VGND.n916 0.0292489
R4588 VGND.n1903 VGND.n367 0.0292489
R4589 VGND.n1896 VGND.n365 0.0292489
R4590 VGND.n1941 VGND.n346 0.0292489
R4591 VGND.n1952 VGND.n1951 0.0292489
R4592 VGND.n2178 VGND.n2123 0.0292489
R4593 VGND.n2180 VGND.n204 0.0292489
R4594 VGND.n2352 VGND.n129 0.0292489
R4595 VGND.n2354 VGND.n126 0.0292489
R4596 VGND.n1382 VGND.n1371 0.0292489
R4597 VGND.n1384 VGND.n871 0.0292489
R4598 VGND.n952 VGND.n951 0.0292489
R4599 VGND.n950 VGND.n949 0.0292489
R4600 VGND.n391 VGND.n383 0.0292489
R4601 VGND.n400 VGND.n399 0.0292489
R4602 VGND.n1920 VGND.n1908 0.0292489
R4603 VGND.n1922 VGND.n359 0.0292489
R4604 VGND.n2139 VGND.n2136 0.0292489
R4605 VGND.n2150 VGND.n2149 0.0292489
R4606 VGND.n2322 VGND.n2310 0.0292489
R4607 VGND.n2324 VGND.n142 0.0292489
R4608 VGND.n878 VGND.n876 0.0292489
R4609 VGND.n888 VGND.n876 0.0292489
R4610 VGND.n1528 VGND.n1527 0.0292489
R4611 VGND.n1530 VGND.n1529 0.0292489
R4612 VGND.n1600 VGND.n701 0.0292489
R4613 VGND.n796 VGND.n702 0.0292489
R4614 VGND.n1724 VGND.n612 0.0292489
R4615 VGND.n1733 VGND.n1732 0.0292489
R4616 VGND.n1799 VGND.n492 0.0292489
R4617 VGND.n515 VGND.n493 0.0292489
R4618 VGND.n2053 VGND.n292 0.0292489
R4619 VGND.n2055 VGND.n290 0.0292489
R4620 VGND.n2302 VGND.n150 0.0292489
R4621 VGND.n2295 VGND.n148 0.0292489
R4622 VGND.n2448 VGND.n72 0.0292489
R4623 VGND.n2459 VGND.n2458 0.0292489
R4624 VGND.n768 VGND.n767 0.0292489
R4625 VGND.n766 VGND.n765 0.0292489
R4626 VGND.n1792 VGND.n595 0.0292489
R4627 VGND.n1778 VGND.n593 0.0292489
R4628 VGND.n591 VGND.n497 0.0292489
R4629 VGND.n579 VGND.n496 0.0292489
R4630 VGND.n2114 VGND.n276 0.0292489
R4631 VGND.n2102 VGND.n274 0.0292489
R4632 VGND.n272 VGND.n208 0.0292489
R4633 VGND.n260 VGND.n207 0.0292489
R4634 VGND.n2518 VGND.n56 0.0292489
R4635 VGND.n2505 VGND.n54 0.0292489
R4636 VGND.n801 VGND.n799 0.0292489
R4637 VGND.n1563 VGND.n799 0.0292489
R4638 VGND.n2348 VGND.n2345 0.0291458
R4639 VGND.n2417 VGND.n2416 0.0291458
R4640 VGND.n59 VGND.n57 0.0291458
R4641 VGND.n2174 VGND.n2171 0.0291458
R4642 VGND.n2256 VGND.n2255 0.0291458
R4643 VGND.n211 VGND.n209 0.0291458
R4644 VGND.n1948 VGND.n1947 0.0291458
R4645 VGND.n2015 VGND.n2014 0.0291458
R4646 VGND.n279 VGND.n277 0.0291458
R4647 VGND.n1899 VGND.n371 0.0291458
R4648 VGND.n1833 VGND.n467 0.0291458
R4649 VGND.n500 VGND.n498 0.0291458
R4650 VGND.n1323 VGND.n921 0.0291458
R4651 VGND.n1694 VGND.n1693 0.0291458
R4652 VGND.n598 VGND.n596 0.0291458
R4653 VGND.n1341 VGND.n911 0.0291458
R4654 VGND.n687 VGND.n686 0.0291458
R4655 VGND.n770 VGND.n728 0.0291458
R4656 VGND.n1417 VGND.n1414 0.0291458
R4657 VGND.n1488 VGND.n1487 0.0291458
R4658 VGND.n1560 VGND.n1559 0.0291458
R4659 VGND.n1197 VGND.n1195 0.0291458
R4660 VGND.n1131 VGND.n1074 0.0291458
R4661 VGND.n2554 VGND.n4 0.0291458
R4662 VGND.n2381 VGND 0.0278438
R4663 VGND.n2215 VGND 0.0278438
R4664 VGND.n1979 VGND 0.0278438
R4665 VGND.n441 VGND 0.0278438
R4666 VGND VGND.n1602 0.0278438
R4667 VGND.n1058 VGND 0.0278438
R4668 VGND.n446 VGND 0.0265417
R4669 VGND VGND.n1391 0.0252396
R4670 VGND.n1408 VGND 0.0252396
R4671 VGND.n1435 VGND 0.0252396
R4672 VGND.n1464 VGND 0.0252396
R4673 VGND.n1506 VGND 0.0252396
R4674 VGND.n1543 VGND 0.0252396
R4675 VGND.n1586 VGND 0.0252396
R4676 VGND.n2567 VGND 0.0252396
R4677 VGND.n2388 VGND.n105 0.0239375
R4678 VGND.n2455 VGND.n2454 0.0239375
R4679 VGND.n2461 VGND.n70 0.0239375
R4680 VGND.n2223 VGND.n187 0.0239375
R4681 VGND.n2298 VGND.n154 0.0239375
R4682 VGND.n2292 VGND.n156 0.0239375
R4683 VGND.n1986 VGND.n326 0.0239375
R4684 VGND.n2049 VGND.n2046 0.0239375
R4685 VGND.n2057 VGND.n288 0.0239375
R4686 VGND.n403 VGND.n402 0.0239375
R4687 VGND.n451 VGND.n442 0.0239375
R4688 VGND.n525 VGND.n520 0.0239375
R4689 VGND.n529 VGND.n514 0.0239375
R4690 VGND.n947 VGND.n935 0.0239375
R4691 VGND.n1279 VGND.n643 0.0239375
R4692 VGND.n1670 VGND 0.0239375
R4693 VGND.n1729 VGND.n1728 0.0239375
R4694 VGND.n1736 VGND.n1735 0.0239375
R4695 VGND.n1765 VGND 0.0239375
R4696 VGND.n1364 VGND.n1363 0.0239375
R4697 VGND.n1347 VGND 0.0239375
R4698 VGND.n664 VGND.n658 0.0239375
R4699 VGND.n716 VGND.n714 0.0239375
R4700 VGND.n794 VGND.n704 0.0239375
R4701 VGND.n1391 VGND.n867 0.0239375
R4702 VGND VGND.n1413 0.0239375
R4703 VGND.n1450 VGND.n839 0.0239375
R4704 VGND.n1523 VGND.n815 0.0239375
R4705 VGND.n1534 VGND.n811 0.0239375
R4706 VGND.n1226 VGND.n1225 0.0239375
R4707 VGND.n1048 VGND.n1045 0.0239375
R4708 VGND.n2532 VGND.n2530 0.0239375
R4709 VGND.n2547 VGND.n45 0.0239375
R4710 VGND.n1082 VGND.n87 0.0234125
R4711 VGND.n1157 VGND.n108 0.0234125
R4712 VGND.n1240 VGND.n127 0.0234125
R4713 VGND.n1229 VGND.n145 0.0234125
R4714 VGND.n2524 VGND.n2523 0.0234125
R4715 VGND.n2520 VGND.n6 0.0234125
R4716 VGND VGND.n2373 0.0226354
R4717 VGND VGND.n2380 0.0226354
R4718 VGND.n2388 VGND 0.0226354
R4719 VGND.n2407 VGND 0.0226354
R4720 VGND.n2437 VGND 0.0226354
R4721 VGND.n2441 VGND 0.0226354
R4722 VGND.n2472 VGND 0.0226354
R4723 VGND.n2510 VGND 0.0226354
R4724 VGND.n2496 VGND 0.0226354
R4725 VGND VGND.n2199 0.0226354
R4726 VGND VGND.n2209 0.0226354
R4727 VGND VGND.n2232 0.0226354
R4728 VGND.n2244 VGND 0.0226354
R4729 VGND VGND.n2264 0.0226354
R4730 VGND.n2277 VGND 0.0226354
R4731 VGND VGND.n154 0.0226354
R4732 VGND.n258 VGND 0.0226354
R4733 VGND.n250 VGND 0.0226354
R4734 VGND VGND.n1971 0.0226354
R4735 VGND VGND.n1978 0.0226354
R4736 VGND.n1986 VGND 0.0226354
R4737 VGND.n2005 VGND 0.0226354
R4738 VGND VGND.n2036 0.0226354
R4739 VGND VGND.n2041 0.0226354
R4740 VGND.n2072 VGND 0.0226354
R4741 VGND VGND.n2078 0.0226354
R4742 VGND.n2093 VGND 0.0226354
R4743 VGND VGND.n415 0.0226354
R4744 VGND.n416 VGND 0.0226354
R4745 VGND VGND.n371 0.0226354
R4746 VGND.n1888 VGND 0.0226354
R4747 VGND VGND.n433 0.0226354
R4748 VGND.n1872 VGND 0.0226354
R4749 VGND VGND.n437 0.0226354
R4750 VGND.n1861 VGND 0.0226354
R4751 VGND.n1811 VGND 0.0226354
R4752 VGND VGND.n489 0.0226354
R4753 VGND.n543 VGND 0.0226354
R4754 VGND.n566 VGND 0.0226354
R4755 VGND VGND.n978 0.0226354
R4756 VGND.n1306 VGND 0.0226354
R4757 VGND VGND.n994 0.0226354
R4758 VGND VGND.n1669 0.0226354
R4759 VGND.n1685 VGND 0.0226354
R4760 VGND VGND.n1689 0.0226354
R4761 VGND VGND.n1714 0.0226354
R4762 VGND VGND.n1755 0.0226354
R4763 VGND VGND.n1761 0.0226354
R4764 VGND.n1358 VGND 0.0226354
R4765 VGND.n1357 VGND 0.0226354
R4766 VGND.n1004 VGND 0.0226354
R4767 VGND.n1009 VGND 0.0226354
R4768 VGND.n1018 VGND 0.0226354
R4769 VGND VGND.n670 0.0226354
R4770 VGND.n1642 VGND 0.0226354
R4771 VGND.n1621 VGND 0.0226354
R4772 VGND.n1613 VGND 0.0226354
R4773 VGND.n1608 VGND 0.0226354
R4774 VGND.n1603 VGND 0.0226354
R4775 VGND.n780 VGND 0.0226354
R4776 VGND.n771 VGND 0.0226354
R4777 VGND VGND.n749 0.0226354
R4778 VGND VGND.n1407 0.0226354
R4779 VGND VGND.n1463 0.0226354
R4780 VGND VGND.n1505 0.0226354
R4781 VGND VGND.n1542 0.0226354
R4782 VGND VGND.n1560 0.0226354
R4783 VGND.n1576 VGND 0.0226354
R4784 VGND.n1218 VGND 0.0226354
R4785 VGND.n1203 VGND 0.0226354
R4786 VGND.n1255 VGND 0.0226354
R4787 VGND VGND.n1057 0.0226354
R4788 VGND.n1112 VGND 0.0226354
R4789 VGND.n2538 VGND 0.0226354
R4790 VGND.n31 VGND 0.0226354
R4791 VGND.n23 VGND 0.0226354
R4792 VGND.n1235 VGND.n1234 0.0218125
R4793 VGND.n2058 VGND 0.0213333
R4794 VGND VGND.n1709 0.0213333
R4795 VGND VGND.n2311 0.0200312
R4796 VGND.n2138 VGND 0.0200312
R4797 VGND VGND.n1909 0.0200312
R4798 VGND.n393 VGND 0.0200312
R4799 VGND.n954 VGND 0.0200312
R4800 VGND.n893 VGND 0.0200312
R4801 VGND VGND.n1372 0.0200312
R4802 VGND VGND.n1398 0.0200312
R4803 VGND VGND.n1169 0.0200312
R4804 VGND.n2357 VGND.n2356 0.0187292
R4805 VGND.n2412 VGND.n84 0.0187292
R4806 VGND.n2425 VGND.n2424 0.0187292
R4807 VGND.n2514 VGND.n60 0.0187292
R4808 VGND.n2510 VGND.n2486 0.0187292
R4809 VGND.n2183 VGND.n2182 0.0187292
R4810 VGND.n2252 VGND.n167 0.0187292
R4811 VGND.n2264 VGND.n2263 0.0187292
R4812 VGND.n268 VGND.n212 0.0187292
R4813 VGND.n265 VGND.n241 0.0187292
R4814 VGND.n1955 VGND.n1954 0.0187292
R4815 VGND.n2010 VGND.n306 0.0187292
R4816 VGND.n2023 VGND.n2022 0.0187292
R4817 VGND.n2110 VGND.n280 0.0187292
R4818 VGND.n2107 VGND.n2084 0.0187292
R4819 VGND.n1893 VGND.n373 0.0187292
R4820 VGND.n476 VGND.n468 0.0187292
R4821 VGND.n1826 VGND.n1825 0.0187292
R4822 VGND.n587 VGND.n501 0.0187292
R4823 VGND.n584 VGND.n559 0.0187292
R4824 VGND.n1317 VGND.n923 0.0187292
R4825 VGND.n631 VGND.n623 0.0187292
R4826 VGND.n1702 VGND.n1701 0.0187292
R4827 VGND.n1788 VGND.n599 0.0187292
R4828 VGND.n1783 VGND.n1760 0.0187292
R4829 VGND.n914 VGND.n912 0.0187292
R4830 VGND.n690 VGND.n681 0.0187292
R4831 VGND.n1627 VGND.n1626 0.0187292
R4832 VGND.n744 VGND.n743 0.0187292
R4833 VGND.n741 VGND.n733 0.0187292
R4834 VGND.n1426 VGND.n1425 0.0187292
R4835 VGND.n1484 VGND.n1483 0.0187292
R4836 VGND.n1496 VGND.n1495 0.0187292
R4837 VGND.n1568 VGND.n1567 0.0187292
R4838 VGND.n805 VGND.n803 0.0187292
R4839 VGND.n1243 VGND.n1033 0.0187292
R4840 VGND.n1083 VGND.n1075 0.0187292
R4841 VGND.n1124 VGND.n1123 0.0187292
R4842 VGND.n17 VGND.n16 0.0187292
R4843 VGND.n14 VGND.n10 0.0187292
R4844 VGND.n1230 VGND.n1036 0.0183038
R4845 VGND.n1231 VGND.n1158 0.0182893
R4846 VGND VGND.n829 0.0174271
R4847 VGND VGND.n90 0.0148229
R4848 VGND VGND.n311 0.0148229
R4849 VGND.n2314 VGND.n2313 0.0135208
R4850 VGND.n113 VGND.n102 0.0135208
R4851 VGND.n2451 VGND.n74 0.0135208
R4852 VGND.n2145 VGND.n2144 0.0135208
R4853 VGND.n2214 VGND.n2212 0.0135208
R4854 VGND.n2299 VGND.n153 0.0135208
R4855 VGND.n1912 VGND.n1911 0.0135208
R4856 VGND.n333 VGND.n323 0.0135208
R4857 VGND.n2050 VGND.n295 0.0135208
R4858 VGND.n395 VGND.n386 0.0135208
R4859 VGND.n1868 VGND.n1867 0.0135208
R4860 VGND.n517 VGND.n490 0.0135208
R4861 VGND.n946 VGND.n937 0.0135208
R4862 VGND.n1280 VGND.n1276 0.0135208
R4863 VGND.n1727 VGND.n614 0.0135208
R4864 VGND.n883 VGND.n882 0.0135208
R4865 VGND.n1659 VGND.n655 0.0135208
R4866 VGND.n710 VGND.n709 0.0135208
R4867 VGND.n1388 VGND.n1387 0.0135208
R4868 VGND.n1454 VGND.n1453 0.0135208
R4869 VGND.n1524 VGND.n1521 0.0135208
R4870 VGND.n1178 VGND.n1177 0.0135208
R4871 VGND.n1064 VGND.n1063 0.0135208
R4872 VGND.n1100 VGND.n48 0.0135208
R4873 VGND.n2551 VGND.n2550 0.012953
R4874 VGND.n1602 VGND 0.0109167
R4875 VGND.n1058 VGND 0.0109167
R4876 VGND.n2299 VGND 0.00961458
R4877 VGND.n2050 VGND 0.00961458
R4878 VGND.n2552 VGND.n2551 0.0090153
R4879 VGND.n42 VGND.n41 0.0090153
R4880 VGND.n2349 VGND.n132 0.0083125
R4881 VGND.n2175 VGND.n2126 0.0083125
R4882 VGND.n2249 VGND.n172 0.0083125
R4883 VGND.n1944 VGND.n348 0.0083125
R4884 VGND.n1900 VGND.n370 0.0083125
R4885 VGND.n1837 VGND.n464 0.0083125
R4886 VGND.n1324 VGND.n920 0.0083125
R4887 VGND.n1690 VGND.n629 0.0083125
R4888 VGND.n1332 VGND.n909 0.0083125
R4889 VGND.n1635 VGND.n1634 0.0083125
R4890 VGND.n1418 VGND.n1412 0.0083125
R4891 VGND.n1480 VGND.n829 0.0083125
R4892 VGND.n1200 VGND.n1190 0.0083125
R4893 VGND.n1134 VGND.n1072 0.0083125
R4894 VGND.n1492 VGND 0.00755
R4895 VGND.n1459 VGND 0.00755
R4896 VGND.n1422 VGND 0.00755
R4897 VGND.n1383 VGND 0.00755
R4898 VGND.n797 VGND 0.00755
R4899 VGND.n1594 VGND 0.00755
R4900 VGND.n1567 VGND 0.00701042
R4901 VGND.n1236 VGND.n1041 0.00653911
R4902 VGND.n1172 VGND.n1159 0.00645637
R4903 VGND.n1228 VGND.n1160 0.00645637
R4904 VGND.n1237 VGND.n1035 0.00640857
R4905 VGND.n1239 VGND.n1238 0.00636298
R4906 VGND.n1241 VGND.n1035 0.00636298
R4907 VGND.n1127 VGND.n1042 0.00631183
R4908 VGND.n1043 VGND.n1040 0.00624332
R4909 VGND.n1156 VGND.n1041 0.00624332
R4910 VGND.n1081 VGND.n1080 0.00604629
R4911 VGND.n1127 VGND.n1126 0.00604629
R4912 VGND.n1172 VGND.n1039 0.00596512
R4913 VGND.n1160 VGND.n1039 0.00596512
R4914 VGND.n2527 VGND.n2526 0.00579577
R4915 VGND VGND.n2509 0.00570833
R4916 VGND VGND.n264 0.00570833
R4917 VGND.n1413 VGND 0.00570833
R4918 VGND.n1561 VGND 0.00570833
R4919 VGND.n1238 VGND.n1237 0.00533429
R4920 VGND.n1158 VGND.n1157 0.0052
R4921 VGND.n1240 VGND.n1036 0.0052
R4922 VGND.n2524 VGND.n51 0.0052
R4923 VGND.n1232 VGND.n6 0.0052
R4924 VGND.n1236 VGND.n1040 0.00496369
R4925 VGND.n1080 VGND.n1042 0.0047957
R4926 VGND.n2356 VGND 0.00440625
R4927 VGND.n2182 VGND 0.00440625
R4928 VGND.n1954 VGND 0.00440625
R4929 VGND.n743 VGND 0.00440625
R4930 VGND.n2550 VGND.n42 0.00411538
R4931 VGND.n2526 VGND.n2525 0.00364583
R4932 VGND.n2549 VGND.n43 0.00364583
R4933 VGND.n2527 VGND.n43 0.00364583
R4934 VGND.n2525 VGND.n50 0.00364583
R4935 VGND VGND.n599 0.00310417
R4936 VGND.n1698 VGND.n626 0.0010875
R4937 VGND.n1665 VGND.n646 0.0010875
R4938 VGND.n1328 VGND.n366 0.0010875
R4939 VGND.n875 VGND.n874 0.0010875
R4940 VGND.n1797 VGND.n494 0.0010875
R4941 VGND.n1794 VGND.n1793 0.0010875
R4942 clknet_0_clk.n12 clknet_0_clk.n10 333.392
R4943 clknet_0_clk.n12 clknet_0_clk.n11 301.392
R4944 clknet_0_clk.n14 clknet_0_clk.n13 301.392
R4945 clknet_0_clk.n16 clknet_0_clk.n15 301.392
R4946 clknet_0_clk.n18 clknet_0_clk.n17 301.392
R4947 clknet_0_clk.n20 clknet_0_clk.n19 301.392
R4948 clknet_0_clk.n22 clknet_0_clk.n21 301.392
R4949 clknet_0_clk.n24 clknet_0_clk.n23 297.863
R4950 clknet_0_clk.n31 clknet_0_clk.n29 248.638
R4951 clknet_0_clk.n31 clknet_0_clk.n30 203.463
R4952 clknet_0_clk.n33 clknet_0_clk.n32 203.463
R4953 clknet_0_clk.n28 clknet_0_clk.n27 203.463
R4954 clknet_0_clk.n37 clknet_0_clk.n36 203.463
R4955 clknet_0_clk.n35 clknet_0_clk.n34 202.456
R4956 clknet_0_clk clknet_0_clk.n25 199.607
R4957 clknet_0_clk.n40 clknet_0_clk.n39 188.201
R4958 clknet_0_clk.n8 clknet_0_clk.t45 184.768
R4959 clknet_0_clk.n7 clknet_0_clk.t33 184.768
R4960 clknet_0_clk.n6 clknet_0_clk.t43 184.768
R4961 clknet_0_clk.n5 clknet_0_clk.t46 184.768
R4962 clknet_0_clk.n0 clknet_0_clk.t42 184.768
R4963 clknet_0_clk.n1 clknet_0_clk.t36 184.768
R4964 clknet_0_clk.n2 clknet_0_clk.t40 184.768
R4965 clknet_0_clk.n3 clknet_0_clk.t38 184.768
R4966 clknet_0_clk clknet_0_clk.n8 173.609
R4967 clknet_0_clk.n4 clknet_0_clk.n3 171.375
R4968 clknet_0_clk.n8 clknet_0_clk.t37 146.208
R4969 clknet_0_clk.n7 clknet_0_clk.t41 146.208
R4970 clknet_0_clk.n6 clknet_0_clk.t35 146.208
R4971 clknet_0_clk.n5 clknet_0_clk.t39 146.208
R4972 clknet_0_clk.n0 clknet_0_clk.t34 146.208
R4973 clknet_0_clk.n1 clknet_0_clk.t44 146.208
R4974 clknet_0_clk.n2 clknet_0_clk.t32 146.208
R4975 clknet_0_clk.n3 clknet_0_clk.t47 146.208
R4976 clknet_0_clk.n33 clknet_0_clk.n31 45.177
R4977 clknet_0_clk.n38 clknet_0_clk.n28 45.177
R4978 clknet_0_clk.n38 clknet_0_clk.n37 45.177
R4979 clknet_0_clk.n35 clknet_0_clk.n33 44.0476
R4980 clknet_0_clk.n37 clknet_0_clk.n35 44.0476
R4981 clknet_0_clk.n8 clknet_0_clk.n7 40.6397
R4982 clknet_0_clk.n7 clknet_0_clk.n6 40.6397
R4983 clknet_0_clk.n6 clknet_0_clk.n5 40.6397
R4984 clknet_0_clk.n1 clknet_0_clk.n0 40.6397
R4985 clknet_0_clk.n2 clknet_0_clk.n1 40.6397
R4986 clknet_0_clk.n3 clknet_0_clk.n2 40.6397
R4987 clknet_0_clk.n29 clknet_0_clk.t26 40.0005
R4988 clknet_0_clk.n29 clknet_0_clk.t22 40.0005
R4989 clknet_0_clk.n30 clknet_0_clk.t24 40.0005
R4990 clknet_0_clk.n30 clknet_0_clk.t19 40.0005
R4991 clknet_0_clk.n32 clknet_0_clk.t21 40.0005
R4992 clknet_0_clk.n32 clknet_0_clk.t23 40.0005
R4993 clknet_0_clk.n34 clknet_0_clk.t25 40.0005
R4994 clknet_0_clk.n34 clknet_0_clk.t27 40.0005
R4995 clknet_0_clk.n25 clknet_0_clk.t18 40.0005
R4996 clknet_0_clk.n25 clknet_0_clk.t20 40.0005
R4997 clknet_0_clk.n27 clknet_0_clk.t30 40.0005
R4998 clknet_0_clk.n27 clknet_0_clk.t16 40.0005
R4999 clknet_0_clk.n39 clknet_0_clk.t17 40.0005
R5000 clknet_0_clk.n39 clknet_0_clk.t28 40.0005
R5001 clknet_0_clk.n36 clknet_0_clk.t29 40.0005
R5002 clknet_0_clk.n36 clknet_0_clk.t31 40.0005
R5003 clknet_0_clk.n14 clknet_0_clk.n12 32.0005
R5004 clknet_0_clk.n16 clknet_0_clk.n14 32.0005
R5005 clknet_0_clk.n20 clknet_0_clk.n18 32.0005
R5006 clknet_0_clk.n22 clknet_0_clk.n20 32.0005
R5007 clknet_0_clk.n18 clknet_0_clk.n16 31.2005
R5008 clknet_0_clk.n21 clknet_0_clk.t12 27.5805
R5009 clknet_0_clk.n21 clknet_0_clk.t5 27.5805
R5010 clknet_0_clk.n10 clknet_0_clk.t15 27.5805
R5011 clknet_0_clk.n10 clknet_0_clk.t2 27.5805
R5012 clknet_0_clk.n11 clknet_0_clk.t13 27.5805
R5013 clknet_0_clk.n11 clknet_0_clk.t8 27.5805
R5014 clknet_0_clk.n13 clknet_0_clk.t1 27.5805
R5015 clknet_0_clk.n13 clknet_0_clk.t3 27.5805
R5016 clknet_0_clk.n15 clknet_0_clk.t14 27.5805
R5017 clknet_0_clk.n15 clknet_0_clk.t9 27.5805
R5018 clknet_0_clk.n17 clknet_0_clk.t11 27.5805
R5019 clknet_0_clk.n17 clknet_0_clk.t4 27.5805
R5020 clknet_0_clk.n19 clknet_0_clk.t6 27.5805
R5021 clknet_0_clk.n19 clknet_0_clk.t10 27.5805
R5022 clknet_0_clk.n23 clknet_0_clk.t7 27.5805
R5023 clknet_0_clk.n23 clknet_0_clk.t0 27.5805
R5024 clknet_0_clk clknet_0_clk.n4 25.9814
R5025 clknet_0_clk.n40 clknet_0_clk.n38 15.262
R5026 clknet_0_clk.n41 clknet_0_clk.n9 14.7771
R5027 clknet_0_clk.n28 clknet_0_clk.n26 13.177
R5028 clknet_0_clk.n24 clknet_0_clk.n22 10.4484
R5029 clknet_0_clk.n9 clknet_0_clk 10.3624
R5030 clknet_0_clk.n41 clknet_0_clk.n40 9.3005
R5031 clknet_0_clk.n9 clknet_0_clk 3.45447
R5032 clknet_0_clk.n26 clknet_0_clk 3.13183
R5033 clknet_0_clk.n4 clknet_0_clk 2.23542
R5034 clknet_0_clk clknet_0_clk.n24 1.75844
R5035 clknet_0_clk clknet_0_clk.n41 1.5927
R5036 clknet_0_clk.n26 clknet_0_clk 0.604792
R5037 VPWR.n234 VPWR.n216 2296.22
R5038 VPWR.n2075 VPWR.n2074 2296.22
R5039 VPWR.n293 VPWR.n275 2296.22
R5040 VPWR.n1758 VPWR.n1757 2291.62
R5041 VPWR.n1757 VPWR.n1754 1418.92
R5042 VPWR.n234 VPWR.n233 1408
R5043 VPWR.n2074 VPWR.n2073 1408
R5044 VPWR.n293 VPWR.n292 1408
R5045 VPWR VPWR.t446 975.178
R5046 VPWR VPWR.t510 975.178
R5047 VPWR VPWR.t481 975.178
R5048 VPWR.t446 VPWR 877.827
R5049 VPWR.t510 VPWR 877.827
R5050 VPWR.t481 VPWR 877.827
R5051 VPWR.n958 VPWR.t340 843.261
R5052 VPWR.n91 VPWR.t745 842.073
R5053 VPWR.n1647 VPWR.t90 842.073
R5054 VPWR.n2224 VPWR.t775 832.876
R5055 VPWR.n2306 VPWR.t603 812.014
R5056 VPWR.n1146 VPWR.t664 811.918
R5057 VPWR.n1236 VPWR.t553 811.793
R5058 VPWR.n1515 VPWR.t52 808.141
R5059 VPWR.n560 VPWR.t636 807.567
R5060 VPWR.n1766 VPWR.t457 807.548
R5061 VPWR.n577 VPWR.t608 807.481
R5062 VPWR.n602 VPWR.t408 807.481
R5063 VPWR.n608 VPWR.t418 807.462
R5064 VPWR.n38 VPWR.t500 806.484
R5065 VPWR.n186 VPWR.t412 806.423
R5066 VPWR.n337 VPWR.t619 806.423
R5067 VPWR.n860 VPWR.t320 804.845
R5068 VPWR.n70 VPWR.t501 804.731
R5069 VPWR.t599 VPWR.n33 804.731
R5070 VPWR.n561 VPWR.t602 804.731
R5071 VPWR.n26 VPWR.t609 804.731
R5072 VPWR.n542 VPWR.t635 804.731
R5073 VPWR.n582 VPWR.t409 804.731
R5074 VPWR.n607 VPWR.t423 804.731
R5075 VPWR.n538 VPWR.t489 804.731
R5076 VPWR.n627 VPWR.t417 804.731
R5077 VPWR.n243 VPWR.t488 804.731
R5078 VPWR.n632 VPWR.t454 804.731
R5079 VPWR.n217 VPWR.t453 804.731
R5080 VPWR.n220 VPWR.t486 804.731
R5081 VPWR.n223 VPWR.t586 804.731
R5082 VPWR.n227 VPWR.t442 804.731
R5083 VPWR.n232 VPWR.t550 804.731
R5084 VPWR.n58 VPWR.t477 804.731
R5085 VPWR.n61 VPWR.t573 804.731
R5086 VPWR.n65 VPWR.t655 804.731
R5087 VPWR.n115 VPWR.t474 804.731
R5088 VPWR.n2054 VPWR.t438 804.731
R5089 VPWR.n2098 VPWR.t567 804.731
R5090 VPWR.n202 VPWR.t439 804.731
R5091 VPWR.n189 VPWR.t568 804.731
R5092 VPWR.n2106 VPWR.t411 804.731
R5093 VPWR.t497 VPWR.n2134 804.731
R5094 VPWR.n184 VPWR.t402 804.731
R5095 VPWR.n2151 VPWR.t680 804.731
R5096 VPWR.n171 VPWR.t403 804.731
R5097 VPWR.n168 VPWR.t681 804.731
R5098 VPWR.n170 VPWR.t605 804.731
R5099 VPWR.n2185 VPWR.t581 804.731
R5100 VPWR.n2193 VPWR.t606 804.731
R5101 VPWR.n153 VPWR.t582 804.731
R5102 VPWR.n2058 VPWR.t533 804.731
R5103 VPWR.n2064 VPWR.t548 804.731
R5104 VPWR.n2067 VPWR.t565 804.731
R5105 VPWR.n2071 VPWR.t584 804.731
R5106 VPWR.n2253 VPWR.t570 804.731
R5107 VPWR.n134 VPWR.t427 804.731
R5108 VPWR.n2273 VPWR.t468 804.731
R5109 VPWR.n1137 VPWR.t556 804.731
R5110 VPWR.n1140 VPWR.t667 804.731
R5111 VPWR.n2004 VPWR.t546 804.731
R5112 VPWR.n675 VPWR.t545 804.731
R5113 VPWR.n674 VPWR.t576 804.731
R5114 VPWR.n1258 VPWR.t575 804.731
R5115 VPWR.n1290 VPWR.t678 804.731
R5116 VPWR.n1092 VPWR.t677 804.731
R5117 VPWR.n1088 VPWR.t406 804.731
R5118 VPWR.n1211 VPWR.t405 804.731
R5119 VPWR.n1235 VPWR.t520 804.731
R5120 VPWR.n1191 VPWR.t559 804.731
R5121 VPWR.n1180 VPWR.t552 804.731
R5122 VPWR.n1175 VPWR.t558 804.731
R5123 VPWR.n1119 VPWR.t665 804.731
R5124 VPWR.n1133 VPWR.t526 804.731
R5125 VPWR.n690 VPWR.t421 804.731
R5126 VPWR.n693 VPWR.t543 804.731
R5127 VPWR.n1378 VPWR.t660 804.731
R5128 VPWR.n1381 VPWR.t463 804.731
R5129 VPWR.n767 VPWR.t641 804.731
R5130 VPWR.n805 VPWR.t640 804.731
R5131 VPWR.n746 VPWR.t672 804.731
R5132 VPWR.n730 VPWR.t671 804.731
R5133 VPWR.t562 VPWR.n1373 804.731
R5134 VPWR.n1375 VPWR.t621 804.731
R5135 VPWR.n1390 VPWR.t561 804.731
R5136 VPWR.n771 VPWR.t536 804.731
R5137 VPWR.n774 VPWR.t633 804.731
R5138 VPWR.n1006 VPWR.t436 804.731
R5139 VPWR.n1009 VPWR.t538 804.731
R5140 VPWR.n999 VPWR.t579 804.731
R5141 VPWR.n1002 VPWR.t669 804.731
R5142 VPWR.n1031 VPWR.t433 804.731
R5143 VPWR.n1625 VPWR.t687 804.731
R5144 VPWR.n1900 VPWR.t624 804.731
R5145 VPWR.n1903 VPWR.t415 804.731
R5146 VPWR.n867 VPWR.t675 804.731
R5147 VPWR.n973 VPWR.t530 804.731
R5148 VPWR.n977 VPWR.t631 804.731
R5149 VPWR.n1781 VPWR.t649 804.731
R5150 VPWR.n1802 VPWR.t456 804.731
R5151 VPWR.n886 VPWR.t397 804.731
R5152 VPWR.n889 VPWR.t506 804.731
R5153 VPWR.n423 VPWR.t611 804.731
R5154 VPWR.n470 VPWR.t610 804.731
R5155 VPWR.n423 VPWR.t483 804.731
R5156 VPWR.n470 VPWR.t482 804.731
R5157 VPWR.n413 VPWR.t509 804.731
R5158 VPWR.n398 VPWR.t508 804.731
R5159 VPWR.n385 VPWR.t638 804.731
R5160 VPWR.n349 VPWR.t637 804.731
R5161 VPWR.n385 VPWR.t512 804.731
R5162 VPWR.n349 VPWR.t511 804.731
R5163 VPWR.n350 VPWR.t448 804.731
R5164 VPWR.n2341 VPWR.t447 804.731
R5165 VPWR.n350 VPWR.t616 804.731
R5166 VPWR.n2341 VPWR.t615 804.731
R5167 VPWR.n2 VPWR.t460 804.731
R5168 VPWR.n509 VPWR.t629 804.731
R5169 VPWR.n328 VPWR.t618 804.731
R5170 VPWR.n320 VPWR.t628 804.731
R5171 VPWR.n261 VPWR.t644 804.731
R5172 VPWR.n276 VPWR.t643 804.731
R5173 VPWR.n279 VPWR.t626 804.731
R5174 VPWR.n282 VPWR.t492 804.731
R5175 VPWR.n286 VPWR.t591 804.731
R5176 VPWR.n291 VPWR.t466 804.731
R5177 VPWR.n434 VPWR.t504 804.731
R5178 VPWR.n440 VPWR.t662 804.731
R5179 VPWR.n1364 VPWR.t226 783.403
R5180 VPWR.n1095 VPWR.t374 779.372
R5181 VPWR.n684 VPWR.t248 779.372
R5182 VPWR.t401 VPWR.t679 772.086
R5183 VPWR.t604 VPWR.t580 772.086
R5184 VPWR.n34 VPWR.t599 751.692
R5185 VPWR.t423 VPWR.n606 751.692
R5186 VPWR.t477 VPWR.n57 751.692
R5187 VPWR.t573 VPWR.n60 751.692
R5188 VPWR.n2135 VPWR.t497 751.692
R5189 VPWR.t570 VPWR.n2252 751.692
R5190 VPWR.t520 VPWR.n1234 751.692
R5191 VPWR.n1387 VPWR.t562 751.692
R5192 VPWR.t621 VPWR.n1374 751.692
R5193 VPWR.t561 VPWR.n1389 751.692
R5194 VPWR.t579 VPWR.n998 751.692
R5195 VPWR.t669 VPWR.n1001 751.692
R5196 VPWR.t649 VPWR.n1780 751.692
R5197 VPWR.t486 VPWR.n219 725.173
R5198 VPWR.t586 VPWR.n222 725.173
R5199 VPWR.t442 VPWR.n226 725.173
R5200 VPWR.t550 VPWR.n231 725.173
R5201 VPWR.t655 VPWR.n64 725.173
R5202 VPWR.t474 VPWR.n114 725.173
R5203 VPWR.t533 VPWR.n2057 725.173
R5204 VPWR.t548 VPWR.n2063 725.173
R5205 VPWR.t565 VPWR.n2066 725.173
R5206 VPWR.t584 VPWR.n2070 725.173
R5207 VPWR.t427 VPWR.n133 725.173
R5208 VPWR.t468 VPWR.n2272 725.173
R5209 VPWR.t556 VPWR.n1136 725.173
R5210 VPWR.t667 VPWR.n1139 725.173
R5211 VPWR.t526 VPWR.n1132 725.173
R5212 VPWR.t421 VPWR.n689 725.173
R5213 VPWR.t543 VPWR.n692 725.173
R5214 VPWR.t660 VPWR.n1377 725.173
R5215 VPWR.t463 VPWR.n1380 725.173
R5216 VPWR.t536 VPWR.n770 725.173
R5217 VPWR.t633 VPWR.n773 725.173
R5218 VPWR.t436 VPWR.n1005 725.173
R5219 VPWR.t538 VPWR.n1008 725.173
R5220 VPWR.t433 VPWR.n1030 725.173
R5221 VPWR.t687 VPWR.n1624 725.173
R5222 VPWR.t624 VPWR.n1899 725.173
R5223 VPWR.t415 VPWR.n1902 725.173
R5224 VPWR.t675 VPWR.n866 725.173
R5225 VPWR.t530 VPWR.n972 725.173
R5226 VPWR.t631 VPWR.n976 725.173
R5227 VPWR.t397 VPWR.n885 725.173
R5228 VPWR.t506 VPWR.n888 725.173
R5229 VPWR.t460 VPWR.n1 725.173
R5230 VPWR.t626 VPWR.n278 725.173
R5231 VPWR.t492 VPWR.n281 725.173
R5232 VPWR.t591 VPWR.n285 725.173
R5233 VPWR.t466 VPWR.n290 725.173
R5234 VPWR.t504 VPWR.n433 725.173
R5235 VPWR.t662 VPWR.n439 725.173
R5236 VPWR.n1592 VPWR.n1059 717.729
R5237 VPWR.n1587 VPWR.n1062 717.729
R5238 VPWR.n143 VPWR.n142 713.462
R5239 VPWR.n1610 VPWR.t326 671.408
R5240 VPWR.n842 VPWR.t710 671.408
R5241 VPWR.n1872 VPWR.t708 671.408
R5242 VPWR.n1492 VPWR.t718 669.655
R5243 VPWR.n92 VPWR.t21 667.734
R5244 VPWR.n138 VPWR.t108 667.734
R5245 VPWR.n1516 VPWR.t116 667.734
R5246 VPWR.n1017 VPWR.t239 667.734
R5247 VPWR.n1017 VPWR.t60 667.734
R5248 VPWR.n1641 VPWR.t791 667.734
R5249 VPWR.n1636 VPWR.t11 667.734
R5250 VPWR.n1484 VPWR.t332 666.677
R5251 VPWR.n1568 VPWR.t773 666.677
R5252 VPWR.n1668 VPWR.t144 666.677
R5253 VPWR.n1668 VPWR.t721 666.677
R5254 VPWR.n1932 VPWR.t23 666.677
R5255 VPWR.n1927 VPWR.t730 666.677
R5256 VPWR.t513 VPWR 666.343
R5257 VPWR VPWR.t407 666.343
R5258 VPWR VPWR.t607 666.343
R5259 VPWR.t592 VPWR 666.343
R5260 VPWR.t587 VPWR 666.343
R5261 VPWR.t645 VPWR 666.343
R5262 VPWR VPWR.t449 664.664
R5263 VPWR.n1585 VPWR.t174 664.37
R5264 VPWR.n1968 VPWR.t100 664.279
R5265 VPWR.n1559 VPWR.t48 664.279
R5266 VPWR.n1045 VPWR.t781 664.279
R5267 VPWR.n751 VPWR.t318 663.024
R5268 VPWR.n42 VPWR.t732 662.571
R5269 VPWR.n2222 VPWR.t808 662.571
R5270 VPWR.n1448 VPWR.t136 659.593
R5271 VPWR.n1729 VPWR.t274 659.593
R5272 VPWR.n1746 VPWR.t80 659.593
R5273 VPWR.n1346 VPWR.n1345 642.188
R5274 VPWR.t416 VPWR.t487 617.668
R5275 VPWR.t410 VPWR.t566 617.668
R5276 VPWR.t617 VPWR.t627 617.668
R5277 VPWR.n923 VPWR.n922 614.562
R5278 VPWR.n1494 VPWR.n1493 613.71
R5279 VPWR.n2248 VPWR.n141 611.178
R5280 VPWR.n1595 VPWR.n1594 611.178
R5281 VPWR.n1585 VPWR.n1066 611.178
R5282 VPWR.n1431 VPWR.n1430 610.861
R5283 VPWR.n1422 VPWR.n1421 609.847
R5284 VPWR.n1362 VPWR.n1361 609.717
R5285 VPWR.n2027 VPWR.n2026 609.303
R5286 VPWR.n1087 VPWR.n1086 606.42
R5287 VPWR.n1319 VPWR.n1084 606.42
R5288 VPWR.n1090 VPWR.n1089 606.42
R5289 VPWR.n680 VPWR.n679 606.42
R5290 VPWR.n2021 VPWR.n678 606.42
R5291 VPWR.n1434 VPWR.n1433 606.42
R5292 VPWR.n1309 VPWR.n1093 605.581
R5293 VPWR.n2015 VPWR.n683 605.581
R5294 VPWR.n1081 VPWR.n1080 605.186
R5295 VPWR.n1079 VPWR.n1078 605.186
R5296 VPWR.n1220 VPWR.n1215 605.186
R5297 VPWR.n1270 VPWR.n1268 605.186
R5298 VPWR.n1267 VPWR.n1266 605.186
R5299 VPWR.n1277 VPWR.n1264 605.186
R5300 VPWR.n1445 VPWR.n1358 605.186
R5301 VPWR.n1449 VPWR.n1447 605.186
R5302 VPWR.n1464 VPWR.n1349 605.186
R5303 VPWR.n152 VPWR.n151 604.394
R5304 VPWR.n1480 VPWR.n1479 604.394
R5305 VPWR.n1586 VPWR.n1063 604.394
R5306 VPWR.n1068 VPWR.n1067 604.394
R5307 VPWR.n1666 VPWR.n1026 604.394
R5308 VPWR.n1666 VPWR.n1028 604.394
R5309 VPWR.n825 VPWR.n824 604.394
R5310 VPWR.n1593 VPWR.n1057 603.231
R5311 VPWR.n952 VPWR.n951 603.231
R5312 VPWR.n2258 VPWR.n136 603.052
R5313 VPWR.n1426 VPWR.n1425 602.456
R5314 VPWR.n2299 VPWR.n39 601.097
R5315 VPWR.n803 VPWR.n752 601.097
R5316 VPWR.n1922 VPWR.n828 601.097
R5317 VPWR.n719 VPWR.n718 599.159
R5318 VPWR.n1446 VPWR.n1357 596.442
R5319 VPWR.n1733 VPWR.n1731 596.442
R5320 VPWR.n1817 VPWR.n1748 596.442
R5321 VPWR.n1420 VPWR.n1419 589.481
R5322 VPWR.n1503 VPWR.n1502 588.318
R5323 VPWR.n1487 VPWR.n1486 585
R5324 VPWR.n1501 VPWR.n1500 585
R5325 VPWR.n1418 VPWR.n1417 585
R5326 VPWR.t634 VPWR 568.994
R5327 VPWR.t601 VPWR 568.994
R5328 VPWR.t496 VPWR 568.994
R5329 VPWR.t577 VPWR.t434 540.46
R5330 VPWR.t557 VPWR 511.926
R5331 VPWR VPWR.t612 510.248
R5332 VPWR.t247 VPWR.t651 496.82
R5333 VPWR.n188 VPWR 491.784
R5334 VPWR.t440 VPWR.t484 463.252
R5335 VPWR.t531 VPWR.t563 463.252
R5336 VPWR.t525 VPWR.t554 463.252
R5337 VPWR.t551 VPWR.t557 463.252
R5338 VPWR.t639 VPWR.t428 463.252
R5339 VPWR.t464 VPWR.t490 463.252
R5340 VPWR.t186 VPWR.t233 458.216
R5341 VPWR VPWR.t663 414.577
R5342 VPWR VPWR.t551 414.577
R5343 VPWR.t428 VPWR 414.577
R5344 VPWR.t612 VPWR 414.577
R5345 VPWR.t507 VPWR 414.577
R5346 VPWR.n911 VPWR.t400 390.875
R5347 VPWR.n604 VPWR.t424 389.526
R5348 VPWR.n1778 VPWR.t650 389.361
R5349 VPWR.n36 VPWR.t600 388.721
R5350 VPWR.n217 VPWR.t514 388.656
R5351 VPWR.n242 VPWR.t515 388.656
R5352 VPWR.n2144 VPWR.t498 388.656
R5353 VPWR.n2054 VPWR.t593 388.656
R5354 VPWR.n2092 VPWR.t594 388.656
R5355 VPWR.n1129 VPWR.t588 388.656
R5356 VPWR.n1121 VPWR.t589 388.656
R5357 VPWR.n1227 VPWR.t521 388.656
R5358 VPWR.n1605 VPWR.t470 388.656
R5359 VPWR.n1609 VPWR.t471 388.656
R5360 VPWR.n882 VPWR.t518 388.656
R5361 VPWR.n276 VPWR.t646 388.656
R5362 VPWR.n314 VPWR.t647 388.656
R5363 VPWR.n496 VPWR.t450 388.656
R5364 VPWR.n402 VPWR.t451 388.656
R5365 VPWR.n2210 VPWR.t596 388.656
R5366 VPWR.n153 VPWR.t597 388.656
R5367 VPWR.n2260 VPWR.t571 388.656
R5368 VPWR.n1244 VPWR.t683 388.656
R5369 VPWR.n1253 VPWR.t684 388.656
R5370 VPWR.n685 VPWR.t652 388.656
R5371 VPWR.n2004 VPWR.t653 388.656
R5372 VPWR.n1504 VPWR.t479 388.656
R5373 VPWR.n724 VPWR.t480 388.656
R5374 VPWR.n1411 VPWR.t622 388.656
R5375 VPWR.n757 VPWR.t429 388.656
R5376 VPWR.n767 VPWR.t430 388.656
R5377 VPWR.n826 VPWR.t523 388.656
R5378 VPWR.n1896 VPWR.t524 388.656
R5379 VPWR.n1723 VPWR.t657 388.656
R5380 VPWR.n1732 VPWR.t658 388.656
R5381 VPWR.n1710 VPWR.t494 388.656
R5382 VPWR.n956 VPWR.t495 388.656
R5383 VPWR.n1823 VPWR.t444 388.656
R5384 VPWR.n1749 VPWR.t445 388.656
R5385 VPWR.n1802 VPWR.t613 388.656
R5386 VPWR.n1763 VPWR.t614 388.656
R5387 VPWR.n845 VPWR.t540 388.656
R5388 VPWR.n851 VPWR.t541 388.656
R5389 VPWR.n862 VPWR.t399 388.656
R5390 VPWR.n56 VPWR.t476 387.682
R5391 VPWR.n59 VPWR.t572 387.682
R5392 VPWR.n997 VPWR.t578 387.682
R5393 VPWR.n1000 VPWR.t668 387.682
R5394 VPWR.n187 VPWR.t595 386.043
R5395 VPWR.n869 VPWR.t517 385.026
R5396 VPWR.n1130 VPWR.t527 383.42
R5397 VPWR VPWR.t277 381.007
R5398 VPWR.n218 VPWR.t485 380.193
R5399 VPWR.n221 VPWR.t585 380.193
R5400 VPWR.n225 VPWR.t441 380.193
R5401 VPWR.n230 VPWR.t549 380.193
R5402 VPWR.n63 VPWR.t654 380.193
R5403 VPWR.n113 VPWR.t473 380.193
R5404 VPWR.n2056 VPWR.t532 380.193
R5405 VPWR.n2062 VPWR.t547 380.193
R5406 VPWR.n2065 VPWR.t564 380.193
R5407 VPWR.n2069 VPWR.t583 380.193
R5408 VPWR.n132 VPWR.t426 380.193
R5409 VPWR.n2271 VPWR.t467 380.193
R5410 VPWR.n1135 VPWR.t555 380.193
R5411 VPWR.n1138 VPWR.t666 380.193
R5412 VPWR.n688 VPWR.t420 380.193
R5413 VPWR.n691 VPWR.t542 380.193
R5414 VPWR.n1376 VPWR.t659 380.193
R5415 VPWR.n1379 VPWR.t462 380.193
R5416 VPWR.n769 VPWR.t535 380.193
R5417 VPWR.n772 VPWR.t632 380.193
R5418 VPWR.n1004 VPWR.t435 380.193
R5419 VPWR.n1007 VPWR.t537 380.193
R5420 VPWR.n1029 VPWR.t432 380.193
R5421 VPWR.n1623 VPWR.t686 380.193
R5422 VPWR.n1898 VPWR.t623 380.193
R5423 VPWR.n1901 VPWR.t414 380.193
R5424 VPWR.n865 VPWR.t674 380.193
R5425 VPWR.n971 VPWR.t529 380.193
R5426 VPWR.n975 VPWR.t630 380.193
R5427 VPWR.n884 VPWR.t396 380.193
R5428 VPWR.n887 VPWR.t505 380.193
R5429 VPWR.n0 VPWR.t459 380.193
R5430 VPWR.n277 VPWR.t625 380.193
R5431 VPWR.n280 VPWR.t491 380.193
R5432 VPWR.n284 VPWR.t590 380.193
R5433 VPWR.n289 VPWR.t465 380.193
R5434 VPWR.n432 VPWR.t503 380.193
R5435 VPWR.n438 VPWR.t661 380.193
R5436 VPWR VPWR.t475 360.866
R5437 VPWR.t487 VPWR 357.51
R5438 VPWR.t566 VPWR 357.51
R5439 VPWR.t627 VPWR 357.51
R5440 VPWR.t560 VPWR 355.83
R5441 VPWR.t280 VPWR.t99 352.474
R5442 VPWR.t59 VPWR.t111 352.474
R5443 VPWR.n1478 VPWR.t765 340.212
R5444 VPWR VPWR.t528 337.368
R5445 VPWR.n1208 VPWR.t72 336.524
R5446 VPWR.n1257 VPWR.t757 336.524
R5447 VPWR.n1033 VPWR.n1032 334.247
R5448 VPWR VPWR.t461 334.012
R5449 VPWR.n2254 VPWR.n139 333.99
R5450 VPWR.n95 VPWR.n94 333.348
R5451 VPWR.n731 VPWR.n729 333.348
R5452 VPWR.n1692 VPWR.n1016 333.348
R5453 VPWR.n1628 VPWR.n1627 333.348
R5454 VPWR.n1514 VPWR.n1497 333.346
R5455 VPWR.n1553 VPWR.n1552 333.346
R5456 VPWR.n1692 VPWR.n1015 333.346
R5457 VPWR.n1631 VPWR.n1630 333.346
R5458 VPWR.n985 VPWR.n965 328.036
R5459 VPWR.n245 VPWR.t901 328.005
R5460 VPWR.n326 VPWR.t931 328.005
R5461 VPWR.n2104 VPWR.t869 328.005
R5462 VPWR.n1777 VPWR.n1768 326.202
R5463 VPWR.n1648 VPWR.n1621 325.639
R5464 VPWR.n96 VPWR.n93 324.74
R5465 VPWR.n1606 VPWR.n1053 322.329
R5466 VPWR.n849 VPWR.n848 322.329
R5467 VPWR.t292 VPWR.t12 322.262
R5468 VPWR.n1260 VPWR.t863 321.911
R5469 VPWR.n72 VPWR.n71 320.976
R5470 VPWR.n735 VPWR.n734 320.976
R5471 VPWR.n1560 VPWR.n1548 320.976
R5472 VPWR.n1023 VPWR.n1022 320.976
R5473 VPWR.n1634 VPWR.n1633 320.976
R5474 VPWR.n2235 VPWR.n2234 320.976
R5475 VPWR.n1491 VPWR.n1490 320.976
R5476 VPWR.n1567 VPWR.n1545 320.976
R5477 VPWR.n1023 VPWR.n1021 320.976
R5478 VPWR.n822 VPWR.n821 320.976
R5479 VPWR.t1 VPWR.t143 315.548
R5480 VPWR.t806 VPWR.t339 315.548
R5481 VPWR.n1466 VPWR.n1465 315.089
R5482 VPWR.n1474 VPWR.n1473 314.447
R5483 VPWR.t115 VPWR.t51 313.87
R5484 VPWR.n149 VPWR.n148 312.829
R5485 VPWR.n1718 VPWR.n953 312.053
R5486 VPWR.n985 VPWR.n967 312.053
R5487 VPWR.n980 VPWR.n970 312.053
R5488 VPWR.n1811 VPWR.n1753 312.053
R5489 VPWR.n1474 VPWR.n1472 312.051
R5490 VPWR.n1227 VPWR.n1210 311.151
R5491 VPWR.n1284 VPWR.n1259 311.151
R5492 VPWR.n1214 VPWR.n1213 310.904
R5493 VPWR.n1263 VPWR.n1262 310.904
R5494 VPWR.n1812 VPWR.n1750 310.5
R5495 VPWR.n907 VPWR.n906 309.533
R5496 VPWR.t452 VPWR.t513 308.834
R5497 VPWR.t407 VPWR.t634 308.834
R5498 VPWR.t607 VPWR.t601 308.834
R5499 VPWR.t437 VPWR.t592 308.834
R5500 VPWR.t682 VPWR.t676 308.834
R5501 VPWR.t620 VPWR.t560 308.834
R5502 VPWR.t642 VPWR.t645 308.834
R5503 VPWR.n504 VPWR.t458 308.834
R5504 VPWR.n873 VPWR.n872 308.755
R5505 VPWR.n853 VPWR.n852 308.755
R5506 VPWR.n1770 VPWR.n1769 308.755
R5507 VPWR.n1765 VPWR.n1764 308.755
R5508 VPWR.n1829 VPWR.n946 308.755
R5509 VPWR.n1410 VPWR.n1366 308.755
R5510 VPWR.n404 VPWR.n403 308.755
R5511 VPWR.n1435 VPWR.n1432 307.204
R5512 VPWR.n1743 VPWR.n947 307.204
R5513 VPWR.n240 VPWR.t926 306.735
R5514 VPWR.n527 VPWR.t832 306.735
R5515 VPWR.n544 VPWR.t847 306.735
R5516 VPWR.n597 VPWR.t835 306.735
R5517 VPWR.n563 VPWR.t854 306.735
R5518 VPWR.n572 VPWR.t866 306.735
R5519 VPWR.n2300 VPWR.t895 306.735
R5520 VPWR.n2191 VPWR.t862 306.735
R5521 VPWR.n2179 VPWR.t840 306.735
R5522 VPWR.n2168 VPWR.t830 306.735
R5523 VPWR.n2145 VPWR.t906 306.735
R5524 VPWR.n2112 VPWR.t903 306.735
R5525 VPWR.n206 VPWR.t894 306.735
R5526 VPWR.n1156 VPWR.t925 306.735
R5527 VPWR.n1118 VPWR.t873 306.735
R5528 VPWR.n1116 VPWR.t851 306.735
R5529 VPWR.n1217 VPWR.t928 306.735
R5530 VPWR.n1094 VPWR.t833 306.735
R5531 VPWR.n682 VPWR.t876 306.735
R5532 VPWR.n732 VPWR.t838 306.735
R5533 VPWR.n756 VPWR.t848 306.735
R5534 VPWR.n1795 VPWR.t891 306.735
R5535 VPWR.n7 VPWR.t858 306.735
R5536 VPWR.n7 VPWR.t888 306.735
R5537 VPWR.n347 VPWR.t898 306.735
R5538 VPWR.n347 VPWR.t927 306.735
R5539 VPWR.n265 VPWR.t849 306.735
R5540 VPWR.n334 VPWR.t856 306.735
R5541 VPWR.n399 VPWR.t900 306.735
R5542 VPWR.n420 VPWR.t908 306.735
R5543 VPWR.n420 VPWR.t834 306.735
R5544 VPWR VPWR.t373 290.372
R5545 VPWR VPWR.t472 280.3
R5546 VPWR.t109 VPWR 280.3
R5547 VPWR VPWR.t425 280.3
R5548 VPWR VPWR.t419 280.3
R5549 VPWR VPWR.t534 280.3
R5550 VPWR VPWR.t413 280.3
R5551 VPWR VPWR.t395 280.3
R5552 VPWR VPWR.t502 280.3
R5553 VPWR.t192 VPWR.t348 278.623
R5554 VPWR.t748 VPWR 261.837
R5555 VPWR VPWR.t452 260.159
R5556 VPWR VPWR.t416 260.159
R5557 VPWR.t422 VPWR 260.159
R5558 VPWR.t598 VPWR 260.159
R5559 VPWR.t475 VPWR 260.159
R5560 VPWR VPWR.t437 260.159
R5561 VPWR VPWR.t410 260.159
R5562 VPWR.t595 VPWR 260.159
R5563 VPWR VPWR.t682 260.159
R5564 VPWR.t651 VPWR 260.159
R5565 VPWR VPWR.t577 260.159
R5566 VPWR VPWR.t493 260.159
R5567 VPWR.t163 VPWR 260.159
R5568 VPWR.t699 VPWR 260.159
R5569 VPWR.t28 VPWR 260.159
R5570 VPWR VPWR.t642 260.159
R5571 VPWR VPWR.t617 260.159
R5572 VPWR.n1132 VPWR.t881 246.71
R5573 VPWR.n219 VPWR.t902 245.667
R5574 VPWR.n222 VPWR.t875 245.667
R5575 VPWR.n226 VPWR.t911 245.667
R5576 VPWR.n231 VPWR.t886 245.667
R5577 VPWR.n64 VPWR.t841 245.667
R5578 VPWR.n114 VPWR.t921 245.667
R5579 VPWR.n2057 VPWR.t880 245.667
R5580 VPWR.n2063 VPWR.t853 245.667
R5581 VPWR.n2066 VPWR.t870 245.667
R5582 VPWR.n2070 VPWR.t846 245.667
R5583 VPWR.n133 VPWR.t914 245.667
R5584 VPWR.n2272 VPWR.t890 245.667
R5585 VPWR.n1136 VPWR.t874 245.667
R5586 VPWR.n1139 VPWR.t924 245.667
R5587 VPWR.n689 VPWR.t916 245.667
R5588 VPWR.n692 VPWR.t855 245.667
R5589 VPWR.n1377 VPWR.t844 245.667
R5590 VPWR.n1380 VPWR.t893 245.667
R5591 VPWR.n770 VPWR.t885 245.667
R5592 VPWR.n773 VPWR.t831 245.667
R5593 VPWR.n1005 VPWR.t919 245.667
R5594 VPWR.n1008 VPWR.t864 245.667
R5595 VPWR.n1030 VPWR.t920 245.667
R5596 VPWR.n1624 VPWR.t922 245.667
R5597 VPWR.n1899 VPWR.t852 245.667
R5598 VPWR.n1902 VPWR.t909 245.667
R5599 VPWR.n866 VPWR.t918 245.667
R5600 VPWR.n972 VPWR.t860 245.667
R5601 VPWR.n976 VPWR.t839 245.667
R5602 VPWR.n885 VPWR.t907 245.667
R5603 VPWR.n888 VPWR.t879 245.667
R5604 VPWR.n1 VPWR.t884 245.667
R5605 VPWR.n278 VPWR.t932 245.667
R5606 VPWR.n281 VPWR.t904 245.667
R5607 VPWR.n285 VPWR.t837 245.667
R5608 VPWR.n290 VPWR.t917 245.667
R5609 VPWR.n433 VPWR.t867 245.667
R5610 VPWR.n439 VPWR.t845 245.667
R5611 VPWR.n1499 VPWR.t814 245.064
R5612 VPWR.n2217 VPWR.t127 243.512
R5613 VPWR.n850 VPWR.t234 241.767
R5614 VPWR.n755 VPWR.t704 240.215
R5615 VPWR.n1896 VPWR.t123 240.214
R5616 VPWR.n34 VPWR.t868 235.319
R5617 VPWR.n1744 VPWR.t117 234.982
R5618 VPWR VPWR.t703 233.304
R5619 VPWR.t648 VPWR.t311 231.625
R5620 VPWR.t813 VPWR.t792 229.947
R5621 VPWR.n1717 VPWR.n954 223.868
R5622 VPWR.t57 VPWR 223.233
R5623 VPWR.t778 VPWR 223.233
R5624 VPWR.t713 VPWR.t722 221.555
R5625 VPWR.t145 VPWR.t16 221.555
R5626 VPWR.t711 VPWR.t53 221.555
R5627 VPWR.n1595 VPWR.n1056 221.314
R5628 VPWR.n606 VPWR.t915 215.827
R5629 VPWR.n1780 VPWR.t829 215.827
R5630 VPWR VPWR.t73 213.163
R5631 VPWR VPWR.t284 213.163
R5632 VPWR.n57 VPWR.t905 213.148
R5633 VPWR.n60 VPWR.t878 213.148
R5634 VPWR.n998 VPWR.t872 213.148
R5635 VPWR.n1001 VPWR.t930 213.148
R5636 VPWR.n1975 VPWR.n726 213.119
R5637 VPWR.n1650 VPWR.n1649 213.119
R5638 VPWR.n1877 VPWR.n844 213.119
R5639 VPWR.n1233 VPWR.t889 211.263
R5640 VPWR.n2211 VPWR.t842 210.964
R5641 VPWR.n1245 VPWR.t913 210.964
R5642 VPWR.n687 VPWR.t929 210.964
R5643 VPWR.n717 VPWR.t883 210.964
R5644 VPWR.n1607 VPWR.t910 210.964
R5645 VPWR.n1711 VPWR.t882 210.964
R5646 VPWR.n2307 VPWR.n31 209.368
R5647 VPWR.n613 VPWR.n539 209.368
R5648 VPWR.n187 VPWR.n155 209.368
R5649 VPWR.n2130 VPWR.n188 209.368
R5650 VPWR.n1291 VPWR.n1243 209.368
R5651 VPWR.n1242 VPWR.n1241 209.368
R5652 VPWR.n1463 VPWR.n1462 209.368
R5653 VPWR.n1652 VPWR.n1651 209.368
R5654 VPWR.n505 VPWR.n504 209.368
R5655 VPWR.t697 VPWR 206.45
R5656 VPWR VPWR.t598 203.093
R5657 VPWR VPWR.t496 203.093
R5658 VPWR VPWR.t401 203.093
R5659 VPWR VPWR.t604 203.093
R5660 VPWR VPWR.t398 203.093
R5661 VPWR VPWR.t807 201.413
R5662 VPWR VPWR.t391 199.736
R5663 VPWR VPWR.t770 199.736
R5664 VPWR.t89 VPWR.t788 198.058
R5665 VPWR.n2137 VPWR.n2136 197.508
R5666 VPWR.t179 VPWR.t20 191.344
R5667 VPWR.t99 VPWR.t151 191.344
R5668 VPWR.t142 VPWR.t59 191.344
R5669 VPWR.t37 VPWR.t278 189.665
R5670 VPWR.n726 VPWR 184.63
R5671 VPWR.n844 VPWR 184.63
R5672 VPWR VPWR.t440 182.952
R5673 VPWR.n31 VPWR 182.952
R5674 VPWR.t472 VPWR 182.952
R5675 VPWR VPWR.t531 182.952
R5676 VPWR.t425 VPWR 182.952
R5677 VPWR.t419 VPWR 182.952
R5678 VPWR.t534 VPWR 182.952
R5679 VPWR.t413 VPWR 182.952
R5680 VPWR.t673 VPWR 182.952
R5681 VPWR.t395 VPWR 182.952
R5682 VPWR VPWR.t464 182.952
R5683 VPWR.t458 VPWR 182.952
R5684 VPWR.t502 VPWR 182.952
R5685 VPWR.t4 VPWR.t300 181.273
R5686 VPWR.n539 VPWR 179.595
R5687 VPWR VPWR.n1242 179.595
R5688 VPWR.n1243 VPWR 179.595
R5689 VPWR.n1744 VPWR 179.595
R5690 VPWR.n503 VPWR 179.595
R5691 VPWR.t302 VPWR.t119 174.559
R5692 VPWR.t351 VPWR.t819 174.559
R5693 VPWR.t784 VPWR.t713 172.881
R5694 VPWR.t16 VPWR.t75 172.881
R5695 VPWR.t0 VPWR.t711 172.881
R5696 VPWR.t809 VPWR.t45 172.881
R5697 VPWR.t325 VPWR 169.524
R5698 VPWR.t119 VPWR.t273 167.845
R5699 VPWR.t782 VPWR.t499 164.488
R5700 VPWR.t169 VPWR.t87 162.81
R5701 VPWR.t190 VPWR.t139 162.81
R5702 VPWR.t22 VPWR.t287 161.131
R5703 VPWR.t83 VPWR.t298 161.131
R5704 VPWR.n1502 VPWR.n1501 159.476
R5705 VPWR.n1419 VPWR.n1418 159.476
R5706 VPWR.t180 VPWR.t784 159.452
R5707 VPWR.t171 VPWR.t736 159.452
R5708 VPWR.t91 VPWR.t739 159.452
R5709 VPWR.t75 VPWR.t152 159.452
R5710 VPWR.t53 VPWR.t3 159.452
R5711 VPWR.t141 VPWR.t0 159.452
R5712 VPWR.t43 VPWR.t39 159.452
R5713 VPWR.t181 VPWR.t516 157.774
R5714 VPWR.t776 VPWR.t61 154.417
R5715 VPWR.t663 VPWR.t587 154.417
R5716 VPWR.t287 VPWR.t821 154.417
R5717 VPWR.t449 VPWR.t507 154.417
R5718 VPWR VPWR.t235 152.739
R5719 VPWR.t499 VPWR.t731 151.06
R5720 VPWR.t478 VPWR.t306 151.06
R5721 VPWR.t79 VPWR.t443 151.06
R5722 VPWR.t393 VPWR.t24 149.382
R5723 VPWR.t157 VPWR.t748 149.382
R5724 VPWR.t124 VPWR.t804 147.703
R5725 VPWR.t770 VPWR.t55 147.703
R5726 VPWR.t117 VPWR.t815 147.703
R5727 VPWR.t349 VPWR.t163 147.703
R5728 VPWR.t26 VPWR.t699 147.703
R5729 VPWR.t95 VPWR.t181 147.703
R5730 VPWR.t133 VPWR.t137 147.703
R5731 VPWR.t167 VPWR.t313 147.703
R5732 VPWR.t194 VPWR.t157 144.346
R5733 VPWR.t321 VPWR.t71 144.346
R5734 VPWR.t750 VPWR.t14 144.346
R5735 VPWR.t385 VPWR.t750 144.346
R5736 VPWR.t377 VPWR.t385 144.346
R5737 VPWR.t381 VPWR.t377 144.346
R5738 VPWR.t371 VPWR.t381 144.346
R5739 VPWR.t375 VPWR.t371 144.346
R5740 VPWR.t383 VPWR.t379 144.346
R5741 VPWR.t355 VPWR.t383 144.346
R5742 VPWR.t363 VPWR.t359 144.346
R5743 VPWR.t367 VPWR.t363 144.346
R5744 VPWR.t361 VPWR.t357 144.346
R5745 VPWR.t365 VPWR.t361 144.346
R5746 VPWR.t369 VPWR.t365 144.346
R5747 VPWR.t373 VPWR.t369 144.346
R5748 VPWR.t756 VPWR.t768 144.346
R5749 VPWR.t768 VPWR.t758 144.346
R5750 VPWR.t758 VPWR.t754 144.346
R5751 VPWR.t754 VPWR.t245 144.346
R5752 VPWR.t245 VPWR.t249 144.346
R5753 VPWR.t253 VPWR.t255 144.346
R5754 VPWR.t255 VPWR.t251 144.346
R5755 VPWR.t251 VPWR.t259 144.346
R5756 VPWR.t259 VPWR.t263 144.346
R5757 VPWR.t263 VPWR.t257 144.346
R5758 VPWR.t269 VPWR.t261 144.346
R5759 VPWR.t261 VPWR.t265 144.346
R5760 VPWR.t265 VPWR.t267 144.346
R5761 VPWR.t267 VPWR.t271 144.346
R5762 VPWR.t271 VPWR.t241 144.346
R5763 VPWR.t241 VPWR.t243 144.346
R5764 VPWR.t219 VPWR.t225 144.346
R5765 VPWR.t217 VPWR.t223 144.346
R5766 VPWR.t197 VPWR.t227 144.346
R5767 VPWR.t213 VPWR.t215 144.346
R5768 VPWR.t762 VPWR.t764 144.346
R5769 VPWR.t819 VPWR.t725 144.346
R5770 VPWR.t731 VPWR.t180 142.668
R5771 VPWR.t359 VPWR.t355 142.668
R5772 VPWR.t203 VPWR.t199 142.668
R5773 VPWR.t152 VPWR.t317 142.668
R5774 VPWR.t143 VPWR.t141 142.668
R5775 VPWR.t772 VPWR.t809 142.668
R5776 VPWR.t155 VPWR.t782 140.989
R5777 VPWR.t744 VPWR.t159 140.989
R5778 VPWR.t391 VPWR.t109 140.989
R5779 VPWR.t97 VPWR.t280 140.989
R5780 VPWR.t151 VPWR.t76 140.989
R5781 VPWR.t73 VPWR.t229 140.989
R5782 VPWR.t111 VPWR.t57 140.989
R5783 VPWR.t3 VPWR.t142 140.989
R5784 VPWR.t93 VPWR.t1 140.989
R5785 VPWR.t45 VPWR.t128 140.989
R5786 VPWR.t161 VPWR.t346 140.989
R5787 VPWR.t36 VPWR.t329 140.989
R5788 VPWR.t232 VPWR.t824 140.989
R5789 VPWR.t284 VPWR.t131 140.989
R5790 VPWR.t103 VPWR.t338 140.989
R5791 VPWR.t101 VPWR.t103 140.989
R5792 VPWR.t707 VPWR.t692 140.989
R5793 VPWR.t87 VPWR.t331 139.311
R5794 VPWR.t159 VPWR.t188 137.633
R5795 VPWR.t798 VPWR.t18 137.633
R5796 VPWR.t774 VPWR.t390 135.954
R5797 VPWR.t766 VPWR.t811 135.954
R5798 VPWR.t786 VPWR.t288 135.954
R5799 VPWR.t333 VPWR.t817 135.954
R5800 VPWR.t140 VPWR.t177 135.954
R5801 VPWR.t122 VPWR 135.954
R5802 VPWR.n1486 VPWR.t787 135.268
R5803 VPWR.t353 VPWR.t67 134.276
R5804 VPWR.t824 VPWR.t10 130.919
R5805 VPWR.t231 VPWR.t800 130.919
R5806 VPWR.n793 VPWR.t896 129.344
R5807 VPWR.n1923 VPWR.t871 129.344
R5808 VPWR.n917 VPWR.t912 129.344
R5809 VPWR.n1822 VPWR.t899 129.344
R5810 VPWR.n950 VPWR.t933 129.344
R5811 VPWR VPWR.t785 129.24
R5812 VPWR.n1758 VPWR.t843 127.695
R5813 VPWR.t315 VPWR.t221 127.562
R5814 VPWR.n1651 VPWR.t780 127.562
R5815 VPWR.t294 VPWR.t304 127.562
R5816 VPWR VPWR.t4 127.562
R5817 VPWR.t484 VPWR 125.883
R5818 VPWR.n539 VPWR 125.883
R5819 VPWR VPWR.n31 125.883
R5820 VPWR.t563 VPWR 125.883
R5821 VPWR.n188 VPWR 125.883
R5822 VPWR VPWR.n187 125.883
R5823 VPWR.t554 VPWR 125.883
R5824 VPWR.n1242 VPWR 125.883
R5825 VPWR.n1243 VPWR 125.883
R5826 VPWR.t461 VPWR 125.883
R5827 VPWR.t172 VPWR.t715 125.883
R5828 VPWR VPWR.n726 125.883
R5829 VPWR.t434 VPWR 125.883
R5830 VPWR.n1651 VPWR 125.883
R5831 VPWR.t39 VPWR.t47 125.883
R5832 VPWR.t695 VPWR.t147 125.883
R5833 VPWR VPWR.n1650 125.883
R5834 VPWR.t528 VPWR 125.883
R5835 VPWR VPWR.n844 125.883
R5836 VPWR.t490 VPWR 125.883
R5837 VPWR.n504 VPWR 125.883
R5838 VPWR VPWR.n503 125.883
R5839 VPWR.n1388 VPWR.t877 124.953
R5840 VPWR.t32 VPWR.t219 124.206
R5841 VPWR.t780 VPWR.t49 124.206
R5842 VPWR.t41 VPWR.t327 124.206
R5843 VPWR.t743 VPWR 122.526
R5844 VPWR.t207 VPWR.t296 122.526
R5845 VPWR.t211 VPWR.t690 122.526
R5846 VPWR.n1462 VPWR.t213 122.526
R5847 VPWR.t30 VPWR.t308 122.526
R5848 VPWR.t544 VPWR.t247 120.849
R5849 VPWR.t724 VPWR.t717 120.849
R5850 VPWR.t703 VPWR.t121 120.849
R5851 VPWR.t9 VPWR.t122 120.849
R5852 VPWR.n870 VPWR.t865 120.76
R5853 VPWR.n1374 VPWR.t836 119.007
R5854 VPWR.n2252 VPWR.t850 118.853
R5855 VPWR.n1486 VPWR.t66 118.549
R5856 VPWR.t788 VPWR.t753 117.492
R5857 VPWR.n1432 VPWR.t297 117.451
R5858 VPWR.n947 VPWR.t70 117.451
R5859 VPWR.n1750 VPWR.t726 117.451
R5860 VPWR.n1155 VPWR.t859 117.294
R5861 VPWR.n1871 VPWR.t861 117.294
R5862 VPWR.n494 VPWR.t887 117.294
R5863 VPWR.n1768 VPWR.t236 116.343
R5864 VPWR.n1053 VPWR.t301 116.341
R5865 VPWR.n848 VPWR.t693 116.341
R5866 VPWR.t81 VPWR 115.814
R5867 VPWR.n1493 VPWR.t716 114.918
R5868 VPWR.n922 VPWR.t38 114.918
R5869 VPWR.n216 VPWR.t892 114.546
R5870 VPWR.n2075 VPWR.t857 114.546
R5871 VPWR.n275 VPWR.t923 114.546
R5872 VPWR.t126 VPWR.t62 114.135
R5873 VPWR.t199 VPWR.t282 114.135
R5874 VPWR.n71 VPWR.t714 113.98
R5875 VPWR.n2234 VPWR.t394 113.98
R5876 VPWR.n1490 VPWR.t289 113.98
R5877 VPWR.n734 VPWR.t17 113.98
R5878 VPWR.n1545 VPWR.t810 113.98
R5879 VPWR.n1548 VPWR.t7 113.98
R5880 VPWR.n1022 VPWR.t712 113.98
R5881 VPWR.n1021 VPWR.t719 113.98
R5882 VPWR.n821 VPWR.t801 113.98
R5883 VPWR.n1633 VPWR.t184 113.98
R5884 VPWR VPWR.t707 112.457
R5885 VPWR.t741 VPWR 110.778
R5886 VPWR VPWR.t321 110.778
R5887 VPWR.t790 VPWR.t336 110.778
R5888 VPWR VPWR.t124 109.1
R5889 VPWR VPWR.t341 109.1
R5890 VPWR.t306 VPWR 109.1
R5891 VPWR.t149 VPWR 109.1
R5892 VPWR.t165 VPWR 109.1
R5893 VPWR VPWR.t34 109.1
R5894 VPWR VPWR.t105 109.1
R5895 VPWR.t387 VPWR 109.1
R5896 VPWR.t278 VPWR 109.1
R5897 VPWR.t137 VPWR 109.1
R5898 VPWR.t313 VPWR 109.1
R5899 VPWR.t733 VPWR 107.421
R5900 VPWR.t796 VPWR.t107 107.421
R5901 VPWR.t121 VPWR 107.421
R5902 VPWR.t522 VPWR 107.421
R5903 VPWR.n503 VPWR.n502 106.561
R5904 VPWR.n1745 VPWR.n1744 106.559
R5905 VPWR.t679 VPWR 105.743
R5906 VPWR.t580 VPWR 105.743
R5907 VPWR VPWR.t620 105.743
R5908 VPWR.t455 VPWR 105.743
R5909 VPWR.t319 VPWR.t28 105.743
R5910 VPWR.t209 VPWR 104.064
R5911 VPWR.t827 VPWR 104.064
R5912 VPWR VPWR.t275 104.064
R5913 VPWR.t692 VPWR.t539 104.064
R5914 VPWR.t113 VPWR.t813 102.385
R5915 VPWR.t317 VPWR 102.385
R5916 VPWR.t173 VPWR 102.385
R5917 VPWR.t516 VPWR 102.385
R5918 VPWR.n2136 VPWR.n2135 101.591
R5919 VPWR VPWR.t794 100.707
R5920 VPWR.t574 VPWR.t253 99.0288
R5921 VPWR.t792 VPWR 99.0288
R5922 VPWR VPWR.t701 99.0288
R5923 VPWR.t65 VPWR.t171 97.3503
R5924 VPWR.n1345 VPWR.t88 96.1553
R5925 VPWR.n718 VPWR.t56 96.1553
R5926 VPWR.n1425 VPWR.t316 96.1553
R5927 VPWR.t47 VPWR.t6 95.6719
R5928 VPWR.t6 VPWR.t323 95.6719
R5929 VPWR.t335 VPWR.t735 95.6719
R5930 VPWR.n142 VPWR.t747 93.81
R5931 VPWR.n1059 VPWR.t696 93.81
R5932 VPWR.n1062 VPWR.t818 93.81
R5933 VPWR.t201 VPWR.t344 92.315
R5934 VPWR.t785 VPWR.t343 90.6365
R5935 VPWR.t469 VPWR.t325 90.6365
R5936 VPWR.t286 VPWR.t823 90.6365
R5937 VPWR.t825 VPWR.t231 90.6365
R5938 VPWR VPWR.t367 88.9581
R5939 VPWR.t688 VPWR.t746 87.2797
R5940 VPWR.t237 VPWR.t709 87.2797
R5941 VPWR VPWR.t8 87.2797
R5942 VPWR.n1502 VPWR.t771 86.7743
R5943 VPWR.n1419 VPWR.t33 86.7743
R5944 VPWR.n1357 VPWR.t691 86.7743
R5945 VPWR.n1357 VPWR.t345 86.7743
R5946 VPWR.n1731 VPWR.t120 86.7743
R5947 VPWR.n1731 VPWR.t303 86.7743
R5948 VPWR.n1748 VPWR.t352 86.7743
R5949 VPWR.n1748 VPWR.t820 86.7743
R5950 VPWR VPWR.t269 85.6012
R5951 VPWR.t277 VPWR 85.6012
R5952 VPWR.t64 VPWR.t195 83.9228
R5953 VPWR.t389 VPWR.t796 83.9228
R5954 VPWR.t701 VPWR.t431 83.9228
R5955 VPWR.t764 VPWR 82.2443
R5956 VPWR.t183 VPWR.t286 82.2443
R5957 VPWR.t760 VPWR 80.5659
R5958 VPWR.t76 VPWR.t670 80.5659
R5959 VPWR.t229 VPWR 80.5659
R5960 VPWR VPWR.t93 80.5659
R5961 VPWR.t85 VPWR 80.5659
R5962 VPWR.t336 VPWR.t232 80.5659
R5963 VPWR.t131 VPWR 80.5659
R5964 VPWR.t717 VPWR.t91 78.8874
R5965 VPWR.t670 VPWR.t145 78.8874
R5966 VPWR.t77 VPWR.t772 78.8874
R5967 VPWR VPWR.t69 78.8874
R5968 VPWR.t725 VPWR 78.8874
R5969 VPWR.t323 VPWR.t44 77.209
R5970 VPWR.t539 VPWR.t186 77.209
R5971 VPWR.t398 VPWR.t673 77.209
R5972 VPWR.t404 VPWR.t375 75.5305
R5973 VPWR.t135 VPWR.t201 75.5305
R5974 VPWR VPWR.t83 75.5305
R5975 VPWR.t69 VPWR 75.5305
R5976 VPWR.t20 VPWR.t744 73.8521
R5977 VPWR.t734 VPWR.t153 73.8521
R5978 VPWR.t329 VPWR.t685 73.8521
R5979 VPWR.t729 VPWR 73.8521
R5980 VPWR.t24 VPWR.t688 72.1736
R5981 VPWR.t746 VPWR.t64 72.1736
R5982 VPWR.t215 VPWR 72.1736
R5983 VPWR VPWR.t760 72.1736
R5984 VPWR.t379 VPWR.t404 68.8168
R5985 VPWR.t205 VPWR.t135 68.8168
R5986 VPWR.t823 VPWR.t825 68.8168
R5987 VPWR VPWR.t302 68.8168
R5988 VPWR VPWR.t97 67.1383
R5989 VPWR.t49 VPWR.t734 67.1383
R5990 VPWR.t153 VPWR.t43 67.1383
R5991 VPWR.t685 VPWR.t81 67.1383
R5992 VPWR.t8 VPWR 67.1383
R5993 VPWR.n1501 VPWR.t793 66.8398
R5994 VPWR.n1418 VPWR.t698 66.8398
R5995 VPWR.t715 VPWR.t115 65.4599
R5996 VPWR VPWR.t36 65.4599
R5997 VPWR.t338 VPWR 65.4599
R5998 VPWR.t290 VPWR.t172 63.7814
R5999 VPWR.t44 VPWR.t335 63.7814
R6000 VPWR.t735 VPWR.t77 63.7814
R6001 VPWR.n141 VPWR.t196 63.3219
R6002 VPWR.n141 VPWR.t797 63.3219
R6003 VPWR.n718 VPWR.t307 63.3219
R6004 VPWR.n1425 VPWR.t342 63.3219
R6005 VPWR.n1594 VPWR.t295 63.3219
R6006 VPWR.n1594 VPWR.t150 63.3219
R6007 VPWR.n1066 VPWR.t162 63.3219
R6008 VPWR.n1066 VPWR.t347 63.3219
R6009 VPWR.t324 VPWR 62.103
R6010 VPWR.t709 VPWR.t387 60.4245
R6011 VPWR.t139 VPWR.t183 58.7461
R6012 VPWR VPWR.t393 57.0676
R6013 VPWR.t195 VPWR.t389 57.0676
R6014 VPWR.t257 VPWR 57.0676
R6015 VPWR.t431 VPWR.t778 57.0676
R6016 VPWR.t357 VPWR 55.3892
R6017 VPWR VPWR.t756 53.7107
R6018 VPWR VPWR.t155 52.0323
R6019 VPWR VPWR.t175 52.0323
R6020 VPWR.t676 VPWR 52.0323
R6021 VPWR.t804 VPWR 52.0323
R6022 VPWR.t344 VPWR.t211 52.0323
R6023 VPWR VPWR.t802 52.0323
R6024 VPWR VPWR.t827 52.0323
R6025 VPWR VPWR.t290 52.0323
R6026 VPWR VPWR.t173 52.0323
R6027 VPWR VPWR.t161 52.0323
R6028 VPWR.t275 VPWR 52.0323
R6029 VPWR.t794 VPWR 52.0323
R6030 VPWR.t727 VPWR 52.0323
R6031 VPWR.t815 VPWR 52.0323
R6032 VPWR VPWR.t79 52.0323
R6033 VPWR VPWR.t26 52.0323
R6034 VPWR VPWR.t237 52.0323
R6035 VPWR VPWR.t705 52.0323
R6036 VPWR VPWR.t95 52.0323
R6037 VPWR VPWR.t133 52.0323
R6038 VPWR VPWR.t167 52.0323
R6039 VPWR.n2136 VPWR.t897 50.5057
R6040 VPWR.t343 VPWR.t179 50.3539
R6041 VPWR VPWR.t639 50.3539
R6042 VPWR.t300 VPWR.t469 50.3539
R6043 VPWR VPWR.t9 50.3539
R6044 VPWR VPWR.t422 48.6754
R6045 VPWR VPWR.t569 48.6754
R6046 VPWR.t519 VPWR 48.6754
R6047 VPWR VPWR.t522 48.6754
R6048 VPWR.t656 VPWR 48.6754
R6049 VPWR VPWR.t455 48.6754
R6050 VPWR VPWR.t648 48.6754
R6051 VPWR.n2137 VPWR.n185 46.0805
R6052 VPWR.t249 VPWR.t574 45.3185
R6053 VPWR.t331 VPWR.t65 45.3185
R6054 VPWR VPWR.t192 45.3185
R6055 VPWR VPWR.t309 45.3185
R6056 VPWR VPWR.t165 43.6401
R6057 VPWR.t34 VPWR 43.6401
R6058 VPWR.n1432 VPWR.t283 42.3555
R6059 VPWR.n947 VPWR.t720 42.3555
R6060 VPWR.n1750 VPWR.t310 42.3555
R6061 VPWR.t705 VPWR.t319 41.9616
R6062 VPWR.n39 VPWR.t156 41.5552
R6063 VPWR.n39 VPWR.t783 41.5552
R6064 VPWR.n151 VPWR.t176 41.5552
R6065 VPWR.n151 VPWR.t63 41.5552
R6066 VPWR.n1479 VPWR.t828 41.5552
R6067 VPWR.n1479 VPWR.t738 41.5552
R6068 VPWR.n752 VPWR.t74 41.5552
R6069 VPWR.n752 VPWR.t230 41.5552
R6070 VPWR.n1063 VPWR.t334 41.5552
R6071 VPWR.n1063 VPWR.t86 41.5552
R6072 VPWR.n1067 VPWR.t46 41.5552
R6073 VPWR.n1067 VPWR.t129 41.5552
R6074 VPWR.n1026 VPWR.t185 41.5552
R6075 VPWR.n1026 VPWR.t94 41.5552
R6076 VPWR.n1028 VPWR.t2 41.5552
R6077 VPWR.n1028 VPWR.t130 41.5552
R6078 VPWR.n824 VPWR.t822 41.5552
R6079 VPWR.n824 VPWR.t178 41.5552
R6080 VPWR.n828 VPWR.t285 41.5552
R6081 VPWR.n828 VPWR.t132 41.5552
R6082 VPWR VPWR.t205 40.2832
R6083 VPWR.t51 VPWR.t30 38.6047
R6084 VPWR VPWR.t737 36.9263
R6085 VPWR.t736 VPWR.t786 36.9263
R6086 VPWR.t348 VPWR.t41 36.9263
R6087 VPWR.n148 VPWR.t777 36.4455
R6088 VPWR.n1366 VPWR.t805 36.1587
R6089 VPWR.n1366 VPWR.t125 36.1587
R6090 VPWR.n1472 VPWR.t803 36.1587
R6091 VPWR.n1472 VPWR.t812 36.1587
R6092 VPWR.n872 VPWR.t134 36.1587
R6093 VPWR.n872 VPWR.t138 36.1587
R6094 VPWR.n852 VPWR.t706 36.1587
R6095 VPWR.n852 VPWR.t29 36.1587
R6096 VPWR.n1769 VPWR.t238 36.1587
R6097 VPWR.n1769 VPWR.t388 36.1587
R6098 VPWR.n1764 VPWR.t27 36.1587
R6099 VPWR.n1764 VPWR.t700 36.1587
R6100 VPWR.n946 VPWR.t816 36.1587
R6101 VPWR.n946 VPWR.t118 36.1587
R6102 VPWR.n953 VPWR.t728 36.1587
R6103 VPWR.n953 VPWR.t354 36.1587
R6104 VPWR.n967 VPWR.t694 36.1587
R6105 VPWR.n967 VPWR.t106 36.1587
R6106 VPWR.n970 VPWR.t276 36.1587
R6107 VPWR.n970 VPWR.t35 36.1587
R6108 VPWR.n1753 VPWR.t350 36.1587
R6109 VPWR.n1753 VPWR.t164 36.1587
R6110 VPWR.n906 VPWR.t96 36.1587
R6111 VPWR.n906 VPWR.t182 36.1587
R6112 VPWR.n403 VPWR.t168 36.1587
R6113 VPWR.n403 VPWR.t314 36.1587
R6114 VPWR.n71 VPWR.t723 35.4605
R6115 VPWR.n2234 VPWR.t689 35.4605
R6116 VPWR.n1490 VPWR.t92 35.4605
R6117 VPWR.n734 VPWR.t146 35.4605
R6118 VPWR.n1545 VPWR.t78 35.4605
R6119 VPWR.n1548 VPWR.t40 35.4605
R6120 VPWR.n1022 VPWR.t752 35.4605
R6121 VPWR.n1021 VPWR.t54 35.4605
R6122 VPWR.n821 VPWR.t826 35.4605
R6123 VPWR.n1633 VPWR.t191 35.4605
R6124 VPWR.t327 VPWR.t695 35.2479
R6125 VPWR.n2247 VPWR.n2246 34.6358
R6126 VPWR.n1829 VPWR.n1828 34.6358
R6127 VPWR.n1776 VPWR.n1770 34.6358
R6128 VPWR.n1860 VPWR.n853 34.6358
R6129 VPWR.n86 VPWR.n68 34.6358
R6130 VPWR.n90 VPWR.n68 34.6358
R6131 VPWR.n101 VPWR.n66 34.6358
R6132 VPWR.n102 VPWR.n101 34.6358
R6133 VPWR.n2248 VPWR.n2247 34.6358
R6134 VPWR.n2236 VPWR.n2233 34.6358
R6135 VPWR.n1532 VPWR.n1488 34.6358
R6136 VPWR.n1522 VPWR.n1521 34.6358
R6137 VPWR.n1513 VPWR.n1498 34.6358
R6138 VPWR.n1591 VPWR.n1060 34.6358
R6139 VPWR.n1558 VPWR.n1549 34.6358
R6140 VPWR.n1562 VPWR.n1561 34.6358
R6141 VPWR.n1562 VPWR.n1546 34.6358
R6142 VPWR.n1566 VPWR.n1546 34.6358
R6143 VPWR.n1554 VPWR.n1551 34.6358
R6144 VPWR.n1693 VPWR.n1014 34.6358
R6145 VPWR.n1680 VPWR.n1679 34.6358
R6146 VPWR.n1679 VPWR.n1678 34.6358
R6147 VPWR.n1678 VPWR.n1019 34.6358
R6148 VPWR.n1674 VPWR.n1673 34.6358
R6149 VPWR.n1673 VPWR.n1672 34.6358
R6150 VPWR.n1672 VPWR.n1024 34.6358
R6151 VPWR.n1646 VPWR.n1626 34.6358
R6152 VPWR.n1937 VPWR.n820 34.6358
R6153 VPWR.n1937 VPWR.n1936 34.6358
R6154 VPWR.n984 VPWR.n968 34.6358
R6155 VPWR.n1810 VPWR.n1754 34.6358
R6156 VPWR.n924 VPWR.n861 34.6358
R6157 VPWR.n1056 VPWR.t305 34.4755
R6158 VPWR.n954 VPWR.t68 34.4755
R6159 VPWR.n1444 VPWR.n1359 33.6462
R6160 VPWR.n1451 VPWR.n1450 33.6462
R6161 VPWR.n1463 VPWR.n1350 33.6462
R6162 VPWR.t14 VPWR 33.5694
R6163 VPWR.t233 VPWR 33.5694
R6164 VPWR.n1493 VPWR.t291 33.4905
R6165 VPWR.n1056 VPWR.t166 33.4905
R6166 VPWR.n954 VPWR.t795 33.4905
R6167 VPWR.n922 VPWR.t279 33.4905
R6168 VPWR.n1345 VPWR.t170 32.7439
R6169 VPWR.n1057 VPWR.t328 32.5055
R6170 VPWR.n1057 VPWR.t148 32.5055
R6171 VPWR.n951 VPWR.t299 32.5055
R6172 VPWR.n951 VPWR.t84 32.5055
R6173 VPWR.n2225 VPWR.n2224 32.377
R6174 VPWR.n1533 VPWR.n1532 32.2581
R6175 VPWR.n2222 VPWR.n2221 32.0005
R6176 VPWR.t227 VPWR 31.891
R6177 VPWR.n1553 VPWR.n1549 31.624
R6178 VPWR.n1692 VPWR.n1691 31.624
R6179 VPWR.n1642 VPWR.n1628 31.624
R6180 VPWR.n1637 VPWR.n1631 31.624
R6181 VPWR.n96 VPWR.n95 30.8711
R6182 VPWR.n1515 VPWR.n1514 30.8711
R6183 VPWR.n1467 VPWR.n1466 30.7205
R6184 VPWR.n136 VPWR.t749 30.5355
R6185 VPWR.n97 VPWR.n92 30.4946
R6186 VPWR.n1691 VPWR.n1017 30.4946
R6187 VPWR.n1642 VPWR.n1641 30.4946
R6188 VPWR.n1637 VPWR.n1636 30.4946
R6189 VPWR.t722 VPWR 30.2125
R6190 VPWR VPWR.t525 30.2125
R6191 VPWR.t225 VPWR.t697 30.2125
R6192 VPWR.t282 VPWR.t197 30.2125
R6193 VPWR.t147 VPWR.t294 30.2125
R6194 VPWR.t12 VPWR.t790 30.2125
R6195 VPWR.n1743 VPWR.n1742 29.3652
R6196 VPWR.n1436 VPWR.n1431 29.2576
R6197 VPWR.n1509 VPWR.n1508 29.1064
R6198 VPWR.n1650 VPWR 28.5341
R6199 VPWR.t10 VPWR.t190 28.5341
R6200 VPWR.t311 VPWR 28.5341
R6201 VPWR.n1053 VPWR.t5 28.4453
R6202 VPWR.n848 VPWR.t187 28.4453
R6203 VPWR.n1768 VPWR.t312 28.4433
R6204 VPWR.n148 VPWR.t742 27.5805
R6205 VPWR.n136 VPWR.t158 27.5805
R6206 VPWR.n2026 VPWR.t258 27.5805
R6207 VPWR.n1210 VPWR.t322 27.5805
R6208 VPWR.n1210 VPWR.t15 27.5805
R6209 VPWR.n1086 VPWR.t364 27.5805
R6210 VPWR.n1086 VPWR.t368 27.5805
R6211 VPWR.n1084 VPWR.t356 27.5805
R6212 VPWR.n1080 VPWR.t380 27.5805
R6213 VPWR.n1080 VPWR.t384 27.5805
R6214 VPWR.n1078 VPWR.t372 27.5805
R6215 VPWR.n1078 VPWR.t376 27.5805
R6216 VPWR.n1215 VPWR.t378 27.5805
R6217 VPWR.n1215 VPWR.t382 27.5805
R6218 VPWR.n1213 VPWR.t751 27.5805
R6219 VPWR.n1213 VPWR.t386 27.5805
R6220 VPWR.n1093 VPWR.t366 27.5805
R6221 VPWR.n1093 VPWR.t370 27.5805
R6222 VPWR.n1089 VPWR.t358 27.5805
R6223 VPWR.n1089 VPWR.t362 27.5805
R6224 VPWR.n1259 VPWR.t769 27.5805
R6225 VPWR.n1259 VPWR.t759 27.5805
R6226 VPWR.n1268 VPWR.t260 27.5805
R6227 VPWR.n1268 VPWR.t264 27.5805
R6228 VPWR.n1266 VPWR.t256 27.5805
R6229 VPWR.n1266 VPWR.t252 27.5805
R6230 VPWR.n1264 VPWR.t250 27.5805
R6231 VPWR.n1264 VPWR.t254 27.5805
R6232 VPWR.n1262 VPWR.t755 27.5805
R6233 VPWR.n1262 VPWR.t246 27.5805
R6234 VPWR.n683 VPWR.t242 27.5805
R6235 VPWR.n683 VPWR.t244 27.5805
R6236 VPWR.n679 VPWR.t268 27.5805
R6237 VPWR.n679 VPWR.t272 27.5805
R6238 VPWR.n678 VPWR.t262 27.5805
R6239 VPWR.n678 VPWR.t266 27.5805
R6240 VPWR.n1473 VPWR.t767 27.5805
R6241 VPWR.n1473 VPWR.t763 27.5805
R6242 VPWR.n1465 VPWR.t216 27.5805
R6243 VPWR.n1465 VPWR.t761 27.5805
R6244 VPWR.n1421 VPWR.t220 27.5805
R6245 VPWR.n1421 VPWR.t222 27.5805
R6246 VPWR.n1361 VPWR.t224 27.5805
R6247 VPWR.n1361 VPWR.t218 27.5805
R6248 VPWR.n1430 VPWR.t228 27.5805
R6249 VPWR.n1430 VPWR.t198 27.5805
R6250 VPWR.n1433 VPWR.t204 27.5805
R6251 VPWR.n1358 VPWR.t208 27.5805
R6252 VPWR.n1358 VPWR.t212 27.5805
R6253 VPWR.n1447 VPWR.t202 27.5805
R6254 VPWR.n1447 VPWR.t206 27.5805
R6255 VPWR.n1349 VPWR.t210 27.5805
R6256 VPWR.n1349 VPWR.t214 27.5805
R6257 VPWR.n1485 VPWR.n1484 27.4829
R6258 VPWR.n1521 VPWR.n1494 27.4829
R6259 VPWR.n1595 VPWR.n1593 27.4829
R6260 VPWR.n1668 VPWR.n1024 27.4829
R6261 VPWR.n1933 VPWR.n1932 27.4829
R6262 VPWR.n1974 VPWR.n727 27.0566
R6263 VPWR.n501 VPWR.n396 27.0566
R6264 VPWR.n142 VPWR.t25 26.9729
R6265 VPWR.n1059 VPWR.t42 26.9729
R6266 VPWR.n1062 VPWR.t193 26.9729
R6267 VPWR.t175 VPWR.t126 26.8556
R6268 VPWR.n86 VPWR.n85 26.7859
R6269 VPWR.n1551 VPWR.n1045 26.7299
R6270 VPWR.n93 VPWR.t160 26.5955
R6271 VPWR.n93 VPWR.t799 26.5955
R6272 VPWR.n94 VPWR.t189 26.5955
R6273 VPWR.n94 VPWR.t19 26.5955
R6274 VPWR.n139 VPWR.t392 26.5955
R6275 VPWR.n139 VPWR.t110 26.5955
R6276 VPWR.n2026 VPWR.t270 26.5955
R6277 VPWR.n1084 VPWR.t360 26.5955
R6278 VPWR.n1497 VPWR.t31 26.5955
R6279 VPWR.n1497 VPWR.t114 26.5955
R6280 VPWR.n1433 VPWR.t200 26.5955
R6281 VPWR.n729 VPWR.t98 26.5955
R6282 VPWR.n729 VPWR.t281 26.5955
R6283 VPWR.n1552 VPWR.t50 26.5955
R6284 VPWR.n1552 VPWR.t154 26.5955
R6285 VPWR.n1016 VPWR.t58 26.5955
R6286 VPWR.n1016 VPWR.t112 26.5955
R6287 VPWR.n1015 VPWR.t240 26.5955
R6288 VPWR.n1015 VPWR.t740 26.5955
R6289 VPWR.n1032 VPWR.t779 26.5955
R6290 VPWR.n1032 VPWR.t702 26.5955
R6291 VPWR.n1621 VPWR.t330 26.5955
R6292 VPWR.n1621 VPWR.t82 26.5955
R6293 VPWR.n1627 VPWR.t789 26.5955
R6294 VPWR.n1627 VPWR.t293 26.5955
R6295 VPWR.n1630 VPWR.t13 26.5955
R6296 VPWR.n1630 VPWR.t337 26.5955
R6297 VPWR.n965 VPWR.t104 26.5955
R6298 VPWR.n965 VPWR.t102 26.5955
R6299 VPWR.n910 VPWR.n869 26.3341
R6300 VPWR.n1604 VPWR.n1054 25.1912
R6301 VPWR.n1742 VPWR.n948 25.1912
R6302 VPWR.n1724 VPWR.n1722 25.1912
R6303 VPWR.n1861 VPWR.n1860 25.1912
R6304 VPWR.t739 VPWR 25.1772
R6305 VPWR VPWR.t89 25.1772
R6306 VPWR.t339 VPWR 25.1772
R6307 VPWR.n986 VPWR.n958 24.0841
R6308 VPWR.n1234 VPWR.n1233 24.0557
R6309 VPWR.n1652 VPWR.n1033 23.7181
R6310 VPWR.n102 VPWR.n62 23.7181
R6311 VPWR.n1385 VPWR.n1382 23.7181
R6312 VPWR.n1391 VPWR.n1385 23.7181
R6313 VPWR.n1975 VPWR.n1974 23.7181
R6314 VPWR.n1595 VPWR.n1054 23.7181
R6315 VPWR.n1585 VPWR.n1584 23.7181
R6316 VPWR.n1014 VPWR.n1003 23.7181
R6317 VPWR.n1665 VPWR.n1033 23.7181
R6318 VPWR.n1828 VPWR.n1745 23.7181
R6319 VPWR.n979 VPWR.n978 23.7181
R6320 VPWR.n1878 VPWR.n1877 23.7181
R6321 VPWR.n502 VPWR.n501 23.7181
R6322 VPWR.t243 VPWR.t544 23.4987
R6323 VPWR.t753 VPWR.t292 23.4987
R6324 VPWR.t298 VPWR.t353 23.4987
R6325 VPWR.n861 VPWR.n860 22.9652
R6326 VPWR.n2221 VPWR.n152 22.9652
R6327 VPWR.n1586 VPWR.n1585 22.9652
R6328 VPWR.n1569 VPWR.n1068 22.9652
R6329 VPWR.n1667 VPWR.n1666 22.9652
R6330 VPWR.n1931 VPWR.n825 22.9652
R6331 VPWR.n1467 VPWR.n1464 22.6748
R6332 VPWR.n1478 VPWR.n1347 22.5887
R6333 VPWR.n1587 VPWR.n1060 22.5887
R6334 VPWR.n1592 VPWR.n1591 22.5887
R6335 VPWR.n1423 VPWR.n1362 22.3091
R6336 VPWR.n2233 VPWR.n149 22.2123
R6337 VPWR.n2225 VPWR.n149 22.2123
R6338 VPWR.n1474 VPWR.n1471 22.2123
R6339 VPWR.n1474 VPWR.n1347 22.2123
R6340 VPWR.n986 VPWR.n985 22.2123
R6341 VPWR.n980 VPWR.n968 22.2123
R6342 VPWR.n985 VPWR.n984 22.2123
R6343 VPWR.n1811 VPWR.n1810 22.2123
R6344 VPWR.n1569 VPWR.n1568 21.8358
R6345 VPWR.n1668 VPWR.n1667 21.8358
R6346 VPWR.n1932 VPWR.n1931 21.8358
R6347 VPWR.t296 VPWR.t203 21.8203
R6348 VPWR.t690 VPWR.t207 21.8203
R6349 VPWR.n1462 VPWR.t209 21.8203
R6350 VPWR.t288 VPWR.t724 21.8203
R6351 VPWR.n1584 VPWR.n1068 21.4593
R6352 VPWR.n1666 VPWR.n1665 21.4593
R6353 VPWR.n1412 VPWR.n1364 21.05
R6354 VPWR.n1145 VPWR.n1130 20.912
R6355 VPWR.n1429 VPWR.n1362 20.8462
R6356 VPWR.n911 VPWR.n910 20.4852
R6357 VPWR.n1423 VPWR.n1422 20.4805
R6358 VPWR.t221 VPWR.t32 20.1418
R6359 VPWR.t346 VPWR.t333 20.1418
R6360 VPWR.n1431 VPWR.n1429 20.1148
R6361 VPWR.n2139 VPWR.n185 20.0749
R6362 VPWR.n1770 VPWR.n842 19.9534
R6363 VPWR.n1389 VPWR.n1388 19.9237
R6364 VPWR.n1435 VPWR.n1434 19.7491
R6365 VPWR.n1445 VPWR.n1444 19.7491
R6366 VPWR.n2254 VPWR.n138 19.577
R6367 VPWR.n1289 VPWR.n1255 19.2067
R6368 VPWR.n1314 VPWR.n1313 18.7808
R6369 VPWR.n35 VPWR.n33 18.7591
R6370 VPWR.t308 VPWR.t113 18.4634
R6371 VPWR.t128 VPWR.t324 18.4634
R6372 VPWR.n2236 VPWR.n2235 18.4476
R6373 VPWR.n1491 VPWR.n1488 18.4476
R6374 VPWR.n1561 VPWR.n1560 18.4476
R6375 VPWR.n1674 VPWR.n1023 18.4476
R6376 VPWR.n1634 VPWR.n820 18.4476
R6377 VPWR.n1933 VPWR.n822 18.4476
R6378 VPWR.n1471 VPWR.n1348 18.0711
R6379 VPWR.n1717 VPWR.n1716 18.0382
R6380 VPWR.n471 VPWR.n417 17.9678
R6381 VPWR.n1226 VPWR.n1225 17.612
R6382 VPWR.n1648 VPWR.n1647 16.9417
R6383 VPWR.n1722 VPWR.n952 16.9417
R6384 VPWR.t223 VPWR.t315 16.785
R6385 VPWR.t493 VPWR.t806 16.785
R6386 VPWR.t443 VPWR.t351 16.785
R6387 VPWR.n2305 VPWR.n33 16.7729
R6388 VPWR.n1237 VPWR.n1235 16.7729
R6389 VPWR.n364 VPWR.n363 16.6847
R6390 VPWR.n806 VPWR.n751 16.5825
R6391 VPWR.n1449 VPWR.n1448 16.4576
R6392 VPWR.n1567 VPWR.n1566 16.1887
R6393 VPWR.n1023 VPWR.n1019 16.1887
R6394 VPWR.n1635 VPWR.n1634 16.1887
R6395 VPWR.n1936 VPWR.n822 16.1887
R6396 VPWR.n980 VPWR 15.8123
R6397 VPWR.n1450 VPWR.n1449 15.3605
R6398 VPWR.n1234 VPWR.n1207 15.2281
R6399 VPWR.n36 VPWR.n35 15.101
R6400 VPWR.n1517 VPWR.n1516 15.0593
R6401 VPWR.n1680 VPWR.n1017 15.0593
R6402 VPWR.n1641 VPWR.n1640 15.0593
R6403 VPWR.n1636 VPWR.n1635 15.0593
R6404 VPWR.n1718 VPWR.n952 15.0593
R6405 VPWR.n1812 VPWR.n1811 15.0593
R6406 VPWR.n2342 VPWR.n3 14.9
R6407 VPWR.n1878 VPWR.n842 14.6829
R6408 VPWR.n2217 VPWR.n2216 14.6484
R6409 VPWR.n502 VPWR.n338 14.5851
R6410 VPWR.n441 VPWR.n431 14.5851
R6411 VPWR.n1492 VPWR.n1491 14.3064
R6412 VPWR.n1587 VPWR.n1586 14.3064
R6413 VPWR.n1927 VPWR.n825 14.3064
R6414 VPWR.n2274 VPWR.n131 14.2735
R6415 VPWR.n1975 VPWR.n725 14.2735
R6416 VPWR.n1649 VPWR.n1046 14.2735
R6417 VPWR.n1909 VPWR.n1897 14.2735
R6418 VPWR.n1824 VPWR.n1745 14.2735
R6419 VPWR.n1877 VPWR.n1876 14.2735
R6420 VPWR.n892 VPWR.n883 14.2735
R6421 VPWR.n2235 VPWR.n143 13.9299
R6422 VPWR.n2003 VPWR.n694 13.8955
R6423 VPWR.n780 VPWR.n768 13.8955
R6424 VPWR.t737 VPWR.t169 13.4281
R6425 VPWR.t55 VPWR.t478 13.4281
R6426 VPWR.t304 VPWR.t149 13.4281
R6427 VPWR.t67 VPWR.t727 13.4281
R6428 VPWR VPWR.t37 13.4281
R6429 VPWR.n1416 VPWR.n1364 12.9181
R6430 VPWR.n233 VPWR.n224 12.8005
R6431 VPWR.n116 VPWR.n62 12.8005
R6432 VPWR.n2073 VPWR.n2072 12.8005
R6433 VPWR.n1141 VPWR.n1134 12.8005
R6434 VPWR.n1010 VPWR.n1003 12.8005
R6435 VPWR.n1649 VPWR.n1648 12.8005
R6436 VPWR.n292 VPWR.n283 12.8005
R6437 VPWR.n1487 VPWR.n1485 12.3976
R6438 VPWR.n1927 VPWR.n1926 12.3912
R6439 VPWR.t802 VPWR.t766 11.7496
R6440 VPWR.t800 VPWR.t22 11.7496
R6441 VPWR.n924 VPWR.n923 11.6993
R6442 VPWR.n860 VPWR.n853 11.6711
R6443 VPWR.n1480 VPWR.n1478 11.2946
R6444 VPWR.n1568 VPWR.n1567 11.2946
R6445 VPWR.n1464 VPWR.n1463 10.9719
R6446 VPWR.n1517 VPWR.n1494 10.9181
R6447 VPWR.n2138 VPWR.n2137 10.912
R6448 VPWR.n1391 VPWR.n1390 10.5744
R6449 VPWR.n1718 VPWR.n1717 10.5417
R6450 VPWR.n1484 VPWR.n1346 10.1652
R6451 VPWR.t569 VPWR.t194 10.0712
R6452 VPWR.n1146 VPWR.n1145 9.8812
R6453 VPWR.n1480 VPWR.n1346 9.78874
R6454 VPWR.n1593 VPWR.n1592 9.78874
R6455 VPWR.n613 VPWR.n540 9.73273
R6456 VPWR.n2298 VPWR.n40 9.73273
R6457 VPWR.n2294 VPWR.n2293 9.73273
R6458 VPWR.n2293 VPWR.n2292 9.73273
R6459 VPWR.n2292 VPWR.n43 9.73273
R6460 VPWR.n73 VPWR.n43 9.73273
R6461 VPWR.n1241 VPWR.n1104 9.73273
R6462 VPWR.n1304 VPWR.n1303 9.73273
R6463 VPWR.n1283 VPWR.n1282 9.73273
R6464 VPWR.n1970 VPWR.n1969 9.73273
R6465 VPWR.n1964 VPWR.n1963 9.73273
R6466 VPWR.n1963 VPWR.n1962 9.73273
R6467 VPWR.n1959 VPWR.n1958 9.73273
R6468 VPWR.n1958 VPWR.n1957 9.73273
R6469 VPWR.n1957 VPWR.n737 9.73273
R6470 VPWR.n802 VPWR.n753 9.73273
R6471 VPWR.n798 VPWR.n797 9.73273
R6472 VPWR.n1790 VPWR.n1765 9.73273
R6473 VPWR.n1786 VPWR.n1765 9.73273
R6474 VPWR.n1786 VPWR.n1785 9.73273
R6475 VPWR.n483 VPWR.n404 9.73273
R6476 VPWR.n1308 VPWR.n1307 9.71972
R6477 VPWR.n2014 VPWR.n2013 9.71972
R6478 VPWR.n1237 VPWR.n1236 9.71084
R6479 VPWR.n1222 VPWR.n1221 9.65296
R6480 VPWR.n1331 VPWR.n1330 9.65296
R6481 VPWR.n1321 VPWR.n1320 9.65296
R6482 VPWR.n1318 VPWR.n1085 9.65296
R6483 VPWR.n1279 VPWR.n1278 9.65296
R6484 VPWR.n1276 VPWR.n1265 9.65296
R6485 VPWR.n1272 VPWR.n1271 9.65296
R6486 VPWR.n2020 VPWR.n2019 9.65296
R6487 VPWR.n1389 VPWR.n1386 9.6005
R6488 VPWR.n1431 VPWR.n1360 9.56172
R6489 VPWR.n803 VPWR.n802 9.52116
R6490 VPWR.n2306 VPWR.n2305 9.49016
R6491 VPWR.n2027 VPWR.n2025 9.35121
R6492 VPWR.n117 VPWR.n116 9.3005
R6493 VPWR.n116 VPWR.n55 9.3005
R6494 VPWR.n116 VPWR.n112 9.3005
R6495 VPWR.n236 VPWR.n235 9.3005
R6496 VPWR.n238 VPWR.n237 9.3005
R6497 VPWR.n655 VPWR.n654 9.3005
R6498 VPWR.n653 VPWR.n652 9.3005
R6499 VPWR.n644 VPWR.n643 9.3005
R6500 VPWR.n642 VPWR.n241 9.3005
R6501 VPWR.n641 VPWR.n640 9.3005
R6502 VPWR.n639 VPWR.n638 9.3005
R6503 VPWR.n637 VPWR.n636 9.3005
R6504 VPWR.n635 VPWR.n634 9.3005
R6505 VPWR.n633 VPWR.n244 9.3005
R6506 VPWR.n631 VPWR.n630 9.3005
R6507 VPWR.n629 VPWR.n628 9.3005
R6508 VPWR.n626 VPWR.n246 9.3005
R6509 VPWR.n625 VPWR.n624 9.3005
R6510 VPWR.n623 VPWR.n247 9.3005
R6511 VPWR.n528 VPWR.n248 9.3005
R6512 VPWR.n536 VPWR.n535 9.3005
R6513 VPWR.n537 VPWR.n526 9.3005
R6514 VPWR.n615 VPWR.n614 9.3005
R6515 VPWR.n613 VPWR.n612 9.3005
R6516 VPWR.n611 VPWR.n540 9.3005
R6517 VPWR.n601 VPWR.n600 9.3005
R6518 VPWR.n599 VPWR.n598 9.3005
R6519 VPWR.n596 VPWR.n543 9.3005
R6520 VPWR.n595 VPWR.n594 9.3005
R6521 VPWR.n552 VPWR.n545 9.3005
R6522 VPWR.n558 VPWR.n557 9.3005
R6523 VPWR.n559 VPWR.n550 9.3005
R6524 VPWR.n585 VPWR.n584 9.3005
R6525 VPWR.n583 VPWR.n551 9.3005
R6526 VPWR.n581 VPWR.n580 9.3005
R6527 VPWR.n576 VPWR.n575 9.3005
R6528 VPWR.n574 VPWR.n573 9.3005
R6529 VPWR.n571 VPWR.n562 9.3005
R6530 VPWR.n570 VPWR.n569 9.3005
R6531 VPWR.n568 VPWR.n567 9.3005
R6532 VPWR.n566 VPWR.n565 9.3005
R6533 VPWR.n564 VPWR.n25 9.3005
R6534 VPWR.n2316 VPWR.n2315 9.3005
R6535 VPWR.n2314 VPWR.n2313 9.3005
R6536 VPWR.n32 VPWR.n27 9.3005
R6537 VPWR.n2308 VPWR.n2307 9.3005
R6538 VPWR.n2305 VPWR.n2304 9.3005
R6539 VPWR.n2302 VPWR.n2301 9.3005
R6540 VPWR.n2298 VPWR.n2297 9.3005
R6541 VPWR.n2296 VPWR.n40 9.3005
R6542 VPWR.n2295 VPWR.n2294 9.3005
R6543 VPWR.n2293 VPWR.n41 9.3005
R6544 VPWR.n2292 VPWR.n2291 9.3005
R6545 VPWR.n44 VPWR.n43 9.3005
R6546 VPWR.n74 VPWR.n73 9.3005
R6547 VPWR.n85 VPWR.n84 9.3005
R6548 VPWR.n87 VPWR.n86 9.3005
R6549 VPWR.n88 VPWR.n68 9.3005
R6550 VPWR.n90 VPWR.n89 9.3005
R6551 VPWR.n92 VPWR.n67 9.3005
R6552 VPWR.n98 VPWR.n97 9.3005
R6553 VPWR.n99 VPWR.n66 9.3005
R6554 VPWR.n101 VPWR.n100 9.3005
R6555 VPWR.n103 VPWR.n102 9.3005
R6556 VPWR.n105 VPWR.n62 9.3005
R6557 VPWR.n2275 VPWR.n2274 9.3005
R6558 VPWR.n2274 VPWR.n130 9.3005
R6559 VPWR.n2274 VPWR.n2270 9.3005
R6560 VPWR.n2060 VPWR.n2055 9.3005
R6561 VPWR.n2059 VPWR.n2053 9.3005
R6562 VPWR.n2080 VPWR.n2079 9.3005
R6563 VPWR.n2078 VPWR.n2077 9.3005
R6564 VPWR.n2090 VPWR.n2089 9.3005
R6565 VPWR.n2091 VPWR.n205 9.3005
R6566 VPWR.n2094 VPWR.n2093 9.3005
R6567 VPWR.n2095 VPWR.n204 9.3005
R6568 VPWR.n2097 VPWR.n2096 9.3005
R6569 VPWR.n2099 VPWR.n203 9.3005
R6570 VPWR.n2101 VPWR.n2100 9.3005
R6571 VPWR.n2103 VPWR.n2102 9.3005
R6572 VPWR.n2105 VPWR.n201 9.3005
R6573 VPWR.n2108 VPWR.n2107 9.3005
R6574 VPWR.n2109 VPWR.n200 9.3005
R6575 VPWR.n2111 VPWR.n2110 9.3005
R6576 VPWR.n2113 VPWR.n198 9.3005
R6577 VPWR.n2116 VPWR.n2115 9.3005
R6578 VPWR.n2114 VPWR.n190 9.3005
R6579 VPWR.n2129 VPWR.n2128 9.3005
R6580 VPWR.n2131 VPWR.n2130 9.3005
R6581 VPWR.n2140 VPWR.n2139 9.3005
R6582 VPWR.n2142 VPWR.n2141 9.3005
R6583 VPWR.n2143 VPWR.n183 9.3005
R6584 VPWR.n2147 VPWR.n2146 9.3005
R6585 VPWR.n2148 VPWR.n182 9.3005
R6586 VPWR.n2150 VPWR.n2149 9.3005
R6587 VPWR.n2153 VPWR.n2152 9.3005
R6588 VPWR.n2157 VPWR.n173 9.3005
R6589 VPWR.n2167 VPWR.n2166 9.3005
R6590 VPWR.n2169 VPWR.n172 9.3005
R6591 VPWR.n2171 VPWR.n2170 9.3005
R6592 VPWR.n2173 VPWR.n2172 9.3005
R6593 VPWR.n2175 VPWR.n2174 9.3005
R6594 VPWR.n2177 VPWR.n2176 9.3005
R6595 VPWR.n2178 VPWR.n169 9.3005
R6596 VPWR.n2181 VPWR.n2180 9.3005
R6597 VPWR.n2183 VPWR.n2182 9.3005
R6598 VPWR.n2184 VPWR.n167 9.3005
R6599 VPWR.n2187 VPWR.n2186 9.3005
R6600 VPWR.n2188 VPWR.n166 9.3005
R6601 VPWR.n2190 VPWR.n2189 9.3005
R6602 VPWR.n2198 VPWR.n2197 9.3005
R6603 VPWR.n2196 VPWR.n2195 9.3005
R6604 VPWR.n2192 VPWR.n156 9.3005
R6605 VPWR.n2207 VPWR.n155 9.3005
R6606 VPWR.n2209 VPWR.n2208 9.3005
R6607 VPWR.n2212 VPWR.n154 9.3005
R6608 VPWR.n2214 VPWR.n2213 9.3005
R6609 VPWR.n2216 VPWR.n2215 9.3005
R6610 VPWR.n2218 VPWR.n2217 9.3005
R6611 VPWR.n2219 VPWR.n152 9.3005
R6612 VPWR.n2221 VPWR.n2220 9.3005
R6613 VPWR.n2223 VPWR.n150 9.3005
R6614 VPWR.n2226 VPWR.n2225 9.3005
R6615 VPWR.n2227 VPWR.n149 9.3005
R6616 VPWR.n2233 VPWR 9.3005
R6617 VPWR.n2237 VPWR.n2236 9.3005
R6618 VPWR.n2246 VPWR.n2245 9.3005
R6619 VPWR.n2247 VPWR.n140 9.3005
R6620 VPWR.n2250 VPWR.n138 9.3005
R6621 VPWR.n2255 VPWR.n2254 9.3005
R6622 VPWR.n2257 VPWR.n2256 9.3005
R6623 VPWR.n2259 VPWR.n135 9.3005
R6624 VPWR.n2262 VPWR.n2261 9.3005
R6625 VPWR.n2263 VPWR.n131 9.3005
R6626 VPWR.n705 VPWR.n694 9.3005
R6627 VPWR.n703 VPWR.n694 9.3005
R6628 VPWR.n696 VPWR.n694 9.3005
R6629 VPWR.n1145 VPWR.n1144 9.3005
R6630 VPWR.n1148 VPWR.n1147 9.3005
R6631 VPWR.n1154 VPWR.n1153 9.3005
R6632 VPWR.n1158 VPWR.n1157 9.3005
R6633 VPWR.n1159 VPWR.n1123 9.3005
R6634 VPWR.n1168 VPWR.n1167 9.3005
R6635 VPWR.n1169 VPWR.n1122 9.3005
R6636 VPWR.n1171 VPWR.n1170 9.3005
R6637 VPWR.n1173 VPWR.n1172 9.3005
R6638 VPWR.n1174 VPWR.n1120 9.3005
R6639 VPWR.n1177 VPWR.n1176 9.3005
R6640 VPWR.n1179 VPWR.n1178 9.3005
R6641 VPWR.n1182 VPWR.n1181 9.3005
R6642 VPWR.n1184 VPWR.n1183 9.3005
R6643 VPWR.n1185 VPWR.n1117 9.3005
R6644 VPWR.n1187 VPWR.n1186 9.3005
R6645 VPWR.n1189 VPWR.n1188 9.3005
R6646 VPWR.n1190 VPWR.n1114 9.3005
R6647 VPWR.n1194 VPWR.n1193 9.3005
R6648 VPWR.n1192 VPWR.n1105 9.3005
R6649 VPWR.n1206 VPWR.n1103 9.3005
R6650 VPWR.n1241 VPWR.n1240 9.3005
R6651 VPWR.n1239 VPWR.n1104 9.3005
R6652 VPWR.n1238 VPWR.n1237 9.3005
R6653 VPWR.n1231 VPWR.n1230 9.3005
R6654 VPWR.n1229 VPWR.n1228 9.3005
R6655 VPWR.n1226 VPWR.n1209 9.3005
R6656 VPWR.n1225 VPWR.n1224 9.3005
R6657 VPWR.n1223 VPWR.n1222 9.3005
R6658 VPWR.n1221 VPWR.n1212 9.3005
R6659 VPWR.n1219 VPWR.n1218 9.3005
R6660 VPWR.n1216 VPWR.n1076 9.3005
R6661 VPWR.n1332 VPWR.n1331 9.3005
R6662 VPWR.n1330 VPWR.n1329 9.3005
R6663 VPWR.n1322 VPWR.n1321 9.3005
R6664 VPWR.n1320 VPWR.n1083 9.3005
R6665 VPWR.n1318 VPWR.n1317 9.3005
R6666 VPWR.n1316 VPWR.n1085 9.3005
R6667 VPWR.n1315 VPWR.n1314 9.3005
R6668 VPWR.n1313 VPWR.n1312 9.3005
R6669 VPWR.n1311 VPWR.n1310 9.3005
R6670 VPWR.n1308 VPWR.n1091 9.3005
R6671 VPWR.n1307 VPWR.n1306 9.3005
R6672 VPWR.n1305 VPWR.n1304 9.3005
R6673 VPWR.n1303 VPWR.n1302 9.3005
R6674 VPWR.n1301 VPWR.n1096 9.3005
R6675 VPWR.n1247 VPWR.n1246 9.3005
R6676 VPWR.n1252 VPWR.n1251 9.3005
R6677 VPWR.n1254 VPWR.n1102 9.3005
R6678 VPWR.n1292 VPWR.n1291 9.3005
R6679 VPWR.n1289 VPWR.n1288 9.3005
R6680 VPWR.n1287 VPWR.n1255 9.3005
R6681 VPWR.n1286 VPWR.n1285 9.3005
R6682 VPWR.n1283 VPWR.n1256 9.3005
R6683 VPWR.n1282 VPWR.n1281 9.3005
R6684 VPWR.n1280 VPWR.n1279 9.3005
R6685 VPWR.n1278 VPWR.n1261 9.3005
R6686 VPWR.n1276 VPWR.n1275 9.3005
R6687 VPWR.n1274 VPWR.n1265 9.3005
R6688 VPWR.n1273 VPWR.n1272 9.3005
R6689 VPWR.n1271 VPWR.n671 9.3005
R6690 VPWR.n1269 VPWR.n672 9.3005
R6691 VPWR.n2029 VPWR.n2028 9.3005
R6692 VPWR.n2025 VPWR.n2024 9.3005
R6693 VPWR.n2023 VPWR.n2022 9.3005
R6694 VPWR.n2020 VPWR.n677 9.3005
R6695 VPWR.n2019 VPWR.n2018 9.3005
R6696 VPWR.n2017 VPWR.n2016 9.3005
R6697 VPWR.n2014 VPWR.n681 9.3005
R6698 VPWR.n2013 VPWR.n2012 9.3005
R6699 VPWR.n2011 VPWR.n2010 9.3005
R6700 VPWR.n2009 VPWR.n2008 9.3005
R6701 VPWR.n2007 VPWR.n2006 9.3005
R6702 VPWR.n2005 VPWR.n686 9.3005
R6703 VPWR.n2003 VPWR.n2002 9.3005
R6704 VPWR.n780 VPWR.n779 9.3005
R6705 VPWR.n781 VPWR.n780 9.3005
R6706 VPWR.n780 VPWR.n765 9.3005
R6707 VPWR.n1385 VPWR.n1384 9.3005
R6708 VPWR.n1392 VPWR.n1391 9.3005
R6709 VPWR.n1399 VPWR.n1371 9.3005
R6710 VPWR.n1400 VPWR.n1399 9.3005
R6711 VPWR.n1409 VPWR.n1408 9.3005
R6712 VPWR.n1410 VPWR.n1365 9.3005
R6713 VPWR.n1413 VPWR.n1412 9.3005
R6714 VPWR.n1414 VPWR.n1364 9.3005
R6715 VPWR.n1416 VPWR.n1415 9.3005
R6716 VPWR.n1420 VPWR.n1363 9.3005
R6717 VPWR.n1424 VPWR.n1423 9.3005
R6718 VPWR.n1427 VPWR.n1426 9.3005
R6719 VPWR.n1429 VPWR.n1428 9.3005
R6720 VPWR.n1437 VPWR.n1436 9.3005
R6721 VPWR.n1438 VPWR.n1359 9.3005
R6722 VPWR.n1444 VPWR.n1443 9.3005
R6723 VPWR.n1452 VPWR.n1451 9.3005
R6724 VPWR.n1450 VPWR.n1351 9.3005
R6725 VPWR.n1460 VPWR.n1350 9.3005
R6726 VPWR.n1463 VPWR.n1461 9.3005
R6727 VPWR.n1468 VPWR.n1467 9.3005
R6728 VPWR.n1469 VPWR.n1348 9.3005
R6729 VPWR.n1471 VPWR.n1470 9.3005
R6730 VPWR.n1475 VPWR.n1474 9.3005
R6731 VPWR.n1476 VPWR.n1347 9.3005
R6732 VPWR.n1478 VPWR.n1477 9.3005
R6733 VPWR.n1481 VPWR.n1480 9.3005
R6734 VPWR.n1482 VPWR.n1346 9.3005
R6735 VPWR.n1484 VPWR.n1483 9.3005
R6736 VPWR.n1485 VPWR.n1343 9.3005
R6737 VPWR.n1534 VPWR.n1533 9.3005
R6738 VPWR.n1532 VPWR.n1531 9.3005
R6739 VPWR.n1524 VPWR.n1488 9.3005
R6740 VPWR.n1523 VPWR.n1522 9.3005
R6741 VPWR.n1521 VPWR.n1520 9.3005
R6742 VPWR.n1519 VPWR.n1494 9.3005
R6743 VPWR.n1518 VPWR.n1517 9.3005
R6744 VPWR.n1516 VPWR.n1495 9.3005
R6745 VPWR.n1515 VPWR.n1496 9.3005
R6746 VPWR.n1513 VPWR.n1512 9.3005
R6747 VPWR.n1511 VPWR.n1498 9.3005
R6748 VPWR.n1510 VPWR.n1509 9.3005
R6749 VPWR.n1508 VPWR.n1507 9.3005
R6750 VPWR.n1506 VPWR.n1505 9.3005
R6751 VPWR.n1984 VPWR.n1983 9.3005
R6752 VPWR.n1982 VPWR.n1981 9.3005
R6753 VPWR.n725 VPWR.n720 9.3005
R6754 VPWR.n1976 VPWR.n1975 9.3005
R6755 VPWR.n1974 VPWR.n1973 9.3005
R6756 VPWR.n1972 VPWR.n727 9.3005
R6757 VPWR.n1971 VPWR.n1970 9.3005
R6758 VPWR.n1969 VPWR.n728 9.3005
R6759 VPWR.n1967 VPWR.n1966 9.3005
R6760 VPWR.n1965 VPWR.n1964 9.3005
R6761 VPWR.n1963 VPWR.n733 9.3005
R6762 VPWR.n1962 VPWR.n1961 9.3005
R6763 VPWR.n1960 VPWR.n1959 9.3005
R6764 VPWR.n1958 VPWR.n736 9.3005
R6765 VPWR.n1957 VPWR.n1956 9.3005
R6766 VPWR.n747 VPWR.n737 9.3005
R6767 VPWR.n750 VPWR.n749 9.3005
R6768 VPWR.n807 VPWR.n806 9.3005
R6769 VPWR.n804 VPWR.n745 9.3005
R6770 VPWR.n802 VPWR.n801 9.3005
R6771 VPWR.n800 VPWR.n753 9.3005
R6772 VPWR.n799 VPWR.n798 9.3005
R6773 VPWR.n797 VPWR.n754 9.3005
R6774 VPWR.n796 VPWR.n795 9.3005
R6775 VPWR.n794 VPWR.n793 9.3005
R6776 VPWR.n792 VPWR.n758 9.3005
R6777 VPWR.n791 VPWR.n790 9.3005
R6778 VPWR.n789 VPWR.n759 9.3005
R6779 VPWR.n768 VPWR.n760 9.3005
R6780 VPWR.n1909 VPWR.n1908 9.3005
R6781 VPWR.n1910 VPWR.n1909 9.3005
R6782 VPWR.n1909 VPWR.n1894 9.3005
R6783 VPWR.n1014 VPWR.n1013 9.3005
R6784 VPWR.n1694 VPWR.n1693 9.3005
R6785 VPWR.n1691 VPWR.n1690 9.3005
R6786 VPWR.n1682 VPWR.n1017 9.3005
R6787 VPWR.n1681 VPWR.n1680 9.3005
R6788 VPWR.n1679 VPWR.n1018 9.3005
R6789 VPWR.n1678 VPWR.n1677 9.3005
R6790 VPWR.n1676 VPWR.n1019 9.3005
R6791 VPWR.n1675 VPWR.n1674 9.3005
R6792 VPWR.n1673 VPWR.n1020 9.3005
R6793 VPWR.n1672 VPWR.n1671 9.3005
R6794 VPWR.n1670 VPWR.n1024 9.3005
R6795 VPWR.n1669 VPWR.n1668 9.3005
R6796 VPWR.n1667 VPWR.n1025 9.3005
R6797 VPWR.n1666 VPWR.n1027 9.3005
R6798 VPWR.n1665 VPWR.n1664 9.3005
R6799 VPWR.n1042 VPWR.n1033 9.3005
R6800 VPWR.n1044 VPWR.n1033 9.3005
R6801 VPWR.n1654 VPWR.n1033 9.3005
R6802 VPWR.n1653 VPWR.n1652 9.3005
R6803 VPWR.n1551 VPWR.n1550 9.3005
R6804 VPWR.n1555 VPWR.n1554 9.3005
R6805 VPWR.n1556 VPWR.n1549 9.3005
R6806 VPWR.n1558 VPWR.n1557 9.3005
R6807 VPWR.n1561 VPWR.n1547 9.3005
R6808 VPWR.n1563 VPWR.n1562 9.3005
R6809 VPWR.n1564 VPWR.n1546 9.3005
R6810 VPWR.n1566 VPWR.n1565 9.3005
R6811 VPWR.n1568 VPWR.n1544 9.3005
R6812 VPWR.n1570 VPWR.n1569 9.3005
R6813 VPWR.n1574 VPWR.n1068 9.3005
R6814 VPWR.n1584 VPWR.n1583 9.3005
R6815 VPWR.n1585 VPWR.n1065 9.3005
R6816 VPWR.n1585 VPWR.n1064 9.3005
R6817 VPWR.n1586 VPWR.n1061 9.3005
R6818 VPWR.n1588 VPWR.n1587 9.3005
R6819 VPWR.n1589 VPWR.n1060 9.3005
R6820 VPWR.n1591 VPWR.n1590 9.3005
R6821 VPWR.n1592 VPWR.n1058 9.3005
R6822 VPWR.n1593 VPWR.n1055 9.3005
R6823 VPWR.n1597 VPWR.n1054 9.3005
R6824 VPWR.n1604 VPWR.n1603 9.3005
R6825 VPWR.n1608 VPWR.n1051 9.3005
R6826 VPWR.n1612 VPWR.n1611 9.3005
R6827 VPWR.n1047 VPWR.n1046 9.3005
R6828 VPWR.n1649 VPWR.n1620 9.3005
R6829 VPWR.n1646 VPWR.n1645 9.3005
R6830 VPWR.n1644 VPWR.n1626 9.3005
R6831 VPWR.n1643 VPWR.n1642 9.3005
R6832 VPWR.n1641 VPWR.n1629 9.3005
R6833 VPWR.n1640 VPWR.n1639 9.3005
R6834 VPWR.n1638 VPWR.n1637 9.3005
R6835 VPWR.n1636 VPWR.n1632 9.3005
R6836 VPWR.n1635 VPWR.n816 9.3005
R6837 VPWR.n820 VPWR.n817 9.3005
R6838 VPWR.n1938 VPWR.n1937 9.3005
R6839 VPWR.n1936 VPWR.n1935 9.3005
R6840 VPWR.n1934 VPWR.n1933 9.3005
R6841 VPWR.n1932 VPWR.n823 9.3005
R6842 VPWR.n1931 VPWR.n1930 9.3005
R6843 VPWR.n1929 VPWR.n825 9.3005
R6844 VPWR.n1928 VPWR.n1927 9.3005
R6845 VPWR.n1926 VPWR.n1925 9.3005
R6846 VPWR.n1924 VPWR.n1923 9.3005
R6847 VPWR.n1921 VPWR.n827 9.3005
R6848 VPWR.n1920 VPWR.n1919 9.3005
R6849 VPWR.n1918 VPWR.n829 9.3005
R6850 VPWR.n1897 VPWR.n830 9.3005
R6851 VPWR.n892 VPWR.n891 9.3005
R6852 VPWR.n893 VPWR.n892 9.3005
R6853 VPWR.n892 VPWR.n879 9.3005
R6854 VPWR.n979 VPWR.n969 9.3005
R6855 VPWR.n981 VPWR.n980 9.3005
R6856 VPWR.n982 VPWR.n968 9.3005
R6857 VPWR.n984 VPWR.n983 9.3005
R6858 VPWR.n985 VPWR.n966 9.3005
R6859 VPWR.n987 VPWR.n986 9.3005
R6860 VPWR.n1709 VPWR.n1708 9.3005
R6861 VPWR.n1712 VPWR.n957 9.3005
R6862 VPWR.n1714 VPWR.n1713 9.3005
R6863 VPWR.n1716 VPWR.n1715 9.3005
R6864 VPWR.n1717 VPWR.n955 9.3005
R6865 VPWR.n1719 VPWR.n1718 9.3005
R6866 VPWR.n1720 VPWR.n952 9.3005
R6867 VPWR.n1722 VPWR.n1721 9.3005
R6868 VPWR.n1725 VPWR.n1724 9.3005
R6869 VPWR.n1726 VPWR.n950 9.3005
R6870 VPWR.n1728 VPWR.n1727 9.3005
R6871 VPWR.n1730 VPWR.n949 9.3005
R6872 VPWR.n1735 VPWR.n1734 9.3005
R6873 VPWR.n1737 VPWR.n948 9.3005
R6874 VPWR.n1742 VPWR.n1741 9.3005
R6875 VPWR.n1830 VPWR.n1829 9.3005
R6876 VPWR.n1828 VPWR.n1827 9.3005
R6877 VPWR.n1826 VPWR.n1745 9.3005
R6878 VPWR.n1825 VPWR.n1824 9.3005
R6879 VPWR.n1822 VPWR.n1821 9.3005
R6880 VPWR.n1820 VPWR.n1819 9.3005
R6881 VPWR.n1818 VPWR.n1747 9.3005
R6882 VPWR.n1816 VPWR.n1815 9.3005
R6883 VPWR.n1814 VPWR.n1813 9.3005
R6884 VPWR.n1812 VPWR.n1751 9.3005
R6885 VPWR.n1811 VPWR.n1752 9.3005
R6886 VPWR.n1810 VPWR.n1809 9.3005
R6887 VPWR.n1807 VPWR.n1754 9.3005
R6888 VPWR.n1804 VPWR.n1803 9.3005
R6889 VPWR.n1801 VPWR.n1800 9.3005
R6890 VPWR.n1798 VPWR.n1797 9.3005
R6891 VPWR.n1796 VPWR.n1762 9.3005
R6892 VPWR.n1794 VPWR.n1793 9.3005
R6893 VPWR.n1792 VPWR.n1791 9.3005
R6894 VPWR.n1790 VPWR.n1789 9.3005
R6895 VPWR.n1788 VPWR.n1765 9.3005
R6896 VPWR.n1787 VPWR.n1786 9.3005
R6897 VPWR.n1785 VPWR.n1784 9.3005
R6898 VPWR.n1776 VPWR.n1775 9.3005
R6899 VPWR.n1770 VPWR.n840 9.3005
R6900 VPWR.n1879 VPWR.n1878 9.3005
R6901 VPWR.n1877 VPWR.n843 9.3005
R6902 VPWR.n1876 VPWR.n1875 9.3005
R6903 VPWR.n1874 VPWR.n1873 9.3005
R6904 VPWR.n1870 VPWR.n1869 9.3005
R6905 VPWR.n1868 VPWR.n846 9.3005
R6906 VPWR.n1867 VPWR.n1866 9.3005
R6907 VPWR.n1865 VPWR.n847 9.3005
R6908 VPWR.n1864 VPWR.n1863 9.3005
R6909 VPWR.n1862 VPWR.n1861 9.3005
R6910 VPWR.n1860 VPWR.n1859 9.3005
R6911 VPWR.n1858 VPWR.n853 9.3005
R6912 VPWR.n861 VPWR.n854 9.3005
R6913 VPWR.n925 VPWR.n924 9.3005
R6914 VPWR.n921 VPWR.n920 9.3005
R6915 VPWR.n918 VPWR.n917 9.3005
R6916 VPWR.n916 VPWR.n915 9.3005
R6917 VPWR.n914 VPWR.n868 9.3005
R6918 VPWR.n913 VPWR.n912 9.3005
R6919 VPWR.n910 VPWR.n909 9.3005
R6920 VPWR.n908 VPWR.n907 9.3005
R6921 VPWR.n904 VPWR.n903 9.3005
R6922 VPWR.n902 VPWR.n901 9.3005
R6923 VPWR.n900 VPWR.n873 9.3005
R6924 VPWR.n883 VPWR.n874 9.3005
R6925 VPWR.n442 VPWR.n441 9.3005
R6926 VPWR.n441 VPWR.n430 9.3005
R6927 VPWR.n441 VPWR.n437 9.3005
R6928 VPWR.n295 VPWR.n294 9.3005
R6929 VPWR.n297 VPWR.n296 9.3005
R6930 VPWR.n302 VPWR.n301 9.3005
R6931 VPWR.n300 VPWR.n299 9.3005
R6932 VPWR.n312 VPWR.n311 9.3005
R6933 VPWR.n313 VPWR.n264 9.3005
R6934 VPWR.n316 VPWR.n315 9.3005
R6935 VPWR.n317 VPWR.n263 9.3005
R6936 VPWR.n319 VPWR.n318 9.3005
R6937 VPWR.n321 VPWR.n262 9.3005
R6938 VPWR.n323 VPWR.n322 9.3005
R6939 VPWR.n325 VPWR.n324 9.3005
R6940 VPWR.n327 VPWR.n260 9.3005
R6941 VPWR.n330 VPWR.n329 9.3005
R6942 VPWR.n331 VPWR.n259 9.3005
R6943 VPWR.n333 VPWR.n332 9.3005
R6944 VPWR.n335 VPWR.n255 9.3005
R6945 VPWR.n336 VPWR.n256 9.3005
R6946 VPWR.n511 VPWR.n510 9.3005
R6947 VPWR.n508 VPWR.n507 9.3005
R6948 VPWR.n506 VPWR.n505 9.3005
R6949 VPWR.n2343 VPWR.n2342 9.3005
R6950 VPWR.n2340 VPWR.n4 9.3005
R6951 VPWR.n2339 VPWR.n2338 9.3005
R6952 VPWR.n2337 VPWR.n5 9.3005
R6953 VPWR.n2336 VPWR.n2335 9.3005
R6954 VPWR.n2334 VPWR.n6 9.3005
R6955 VPWR.n2333 VPWR.n2332 9.3005
R6956 VPWR.n10 VPWR.n8 9.3005
R6957 VPWR.n359 VPWR.n358 9.3005
R6958 VPWR.n360 VPWR.n351 9.3005
R6959 VPWR.n362 VPWR.n361 9.3005
R6960 VPWR.n363 VPWR 9.3005
R6961 VPWR.n365 VPWR.n364 9.3005
R6962 VPWR.n367 VPWR.n366 9.3005
R6963 VPWR.n368 VPWR.n348 9.3005
R6964 VPWR.n370 VPWR.n369 9.3005
R6965 VPWR.n372 VPWR.n371 9.3005
R6966 VPWR.n373 VPWR.n346 9.3005
R6967 VPWR.n375 VPWR.n374 9.3005
R6968 VPWR.n376 VPWR.n345 9.3005
R6969 VPWR.n383 VPWR.n382 9.3005
R6970 VPWR.n384 VPWR.n343 9.3005
R6971 VPWR.n387 VPWR.n386 9.3005
R6972 VPWR.n339 VPWR.n338 9.3005
R6973 VPWR.n502 VPWR.n395 9.3005
R6974 VPWR.n501 VPWR.n500 9.3005
R6975 VPWR.n499 VPWR.n396 9.3005
R6976 VPWR.n498 VPWR.n497 9.3005
R6977 VPWR.n495 VPWR.n397 9.3005
R6978 VPWR.n493 VPWR.n492 9.3005
R6979 VPWR.n491 VPWR.n490 9.3005
R6980 VPWR.n489 VPWR.n400 9.3005
R6981 VPWR.n488 VPWR.n487 9.3005
R6982 VPWR.n486 VPWR.n401 9.3005
R6983 VPWR.n485 VPWR.n484 9.3005
R6984 VPWR.n483 VPWR.n482 9.3005
R6985 VPWR.n414 VPWR.n404 9.3005
R6986 VPWR.n417 VPWR.n416 9.3005
R6987 VPWR.n472 VPWR.n471 9.3005
R6988 VPWR.n469 VPWR.n412 9.3005
R6989 VPWR.n468 VPWR.n467 9.3005
R6990 VPWR.n466 VPWR.n418 9.3005
R6991 VPWR.n465 VPWR.n464 9.3005
R6992 VPWR.n463 VPWR.n419 9.3005
R6993 VPWR.n462 VPWR.n461 9.3005
R6994 VPWR.n460 VPWR.n421 9.3005
R6995 VPWR.n459 VPWR.n458 9.3005
R6996 VPWR.n457 VPWR.n422 9.3005
R6997 VPWR.n456 VPWR.n455 9.3005
R6998 VPWR.n431 VPWR.n424 9.3005
R6999 VPWR.n1291 VPWR.n1290 9.09802
R7000 VPWR.n1285 VPWR.n1258 9.09802
R7001 VPWR.n1285 VPWR.n1284 9.09802
R7002 VPWR.n746 VPWR.n737 9.09802
R7003 VPWR.n805 VPWR.n804 9.09802
R7004 VPWR.n413 VPWR.n404 9.09802
R7005 VPWR.n1310 VPWR.n1092 9.02345
R7006 VPWR.n1269 VPWR.n674 9.02345
R7007 VPWR.n2022 VPWR.n675 9.02345
R7008 VPWR.n42 VPWR.n40 8.99224
R7009 VPWR.n870 VPWR.n869 8.9761
R7010 VPWR.n1970 VPWR.n731 8.88645
R7011 VPWR.n1434 VPWR.n1359 8.77764
R7012 VPWR.n1310 VPWR.n1309 8.60378
R7013 VPWR.n2016 VPWR.n2015 8.60378
R7014 VPWR.n614 VPWR.n613 8.44958
R7015 VPWR.n2307 VPWR.n32 8.44958
R7016 VPWR.n2192 VPWR.n155 8.44958
R7017 VPWR.n2130 VPWR.n2129 8.44958
R7018 VPWR.n1241 VPWR.n1103 8.44958
R7019 VPWR.n508 VPWR.n505 8.44958
R7020 VPWR.t811 VPWR.t762 8.39273
R7021 VPWR.n2021 VPWR.n2020 8.28902
R7022 VPWR.n92 VPWR.n91 8.28285
R7023 VPWR.n1560 VPWR.n1559 8.28285
R7024 VPWR.n1446 VPWR.n1445 8.04621
R7025 VPWR.n2013 VPWR.n684 8.04017
R7026 VPWR.n604 VPWR.n603 7.98741
R7027 VPWR.n1559 VPWR.n1558 7.90638
R7028 VPWR.n1652 VPWR.n1045 7.90638
R7029 VPWR.n2209 VPWR.n155 7.75995
R7030 VPWR.n1303 VPWR.n1096 7.75995
R7031 VPWR.n1291 VPWR.n1254 7.75995
R7032 VPWR.n2010 VPWR.n2009 7.75995
R7033 VPWR.n797 VPWR.n796 7.75995
R7034 VPWR.n1791 VPWR.n1790 7.75995
R7035 VPWR.n484 VPWR.n483 7.75995
R7036 VPWR.n1088 VPWR.n1087 7.65952
R7037 VPWR.n1968 VPWR.n1967 7.51124
R7038 VPWR.n1813 VPWR.n1812 7.49704
R7039 VPWR.n1235 VPWR.n1207 7.28326
R7040 VPWR.n1233 VPWR.n1232 7.23528
R7041 VPWR.n2184 VPWR.n2183 7.21067
R7042 VPWR.n2174 VPWR.n2173 7.21067
R7043 VPWR.n1181 VPWR.n1179 7.21067
R7044 VPWR.n1214 VPWR.n1211 7.17134
R7045 VPWR.n497 VPWR.n398 7.12524
R7046 VPWR.n1319 VPWR.n1318 7.03001
R7047 VPWR.n91 VPWR.n90 6.77697
R7048 VPWR.n2217 VPWR.n152 6.77697
R7049 VPWR.n1647 VPWR.n1646 6.77697
R7050 VPWR.n912 VPWR.n911 6.73838
R7051 VPWR.t62 VPWR.t733 6.71428
R7052 VPWR.t807 VPWR.t774 6.71428
R7053 VPWR.t177 VPWR.t729 6.71428
R7054 VPWR.t105 VPWR.t101 6.71428
R7055 VPWR.t309 VPWR.t349 6.71428
R7056 VPWR.n608 VPWR.n540 6.66496
R7057 VPWR.n2307 VPWR.n2306 6.66496
R7058 VPWR.n2301 VPWR.n38 6.66496
R7059 VPWR.n2130 VPWR.n186 6.66496
R7060 VPWR.n1236 VPWR.n1104 6.66496
R7061 VPWR.n1785 VPWR.n1766 6.66496
R7062 VPWR.n505 VPWR.n337 6.66496
R7063 VPWR.n638 VPWR.n637 6.52104
R7064 VPWR.n1174 VPWR.n1173 6.52104
R7065 VPWR.n319 VPWR.n263 6.52104
R7066 VPWR.n2150 VPWR.n182 6.52104
R7067 VPWR.n2097 VPWR.n204 6.52104
R7068 VPWR.n1221 VPWR.n1220 6.50542
R7069 VPWR.n1278 VPWR.n1277 6.50542
R7070 VPWR.n609 VPWR.n607 6.48583
R7071 VPWR.n1782 VPWR.n1781 6.48583
R7072 VPWR.n1778 VPWR.n1777 6.46951
R7073 VPWR.n1516 VPWR.n1515 6.4005
R7074 VPWR VPWR.n979 6.4005
R7075 VPWR.n1777 VPWR.n1776 6.4005
R7076 VPWR.n1420 VPWR.n1417 6.3005
R7077 VPWR.n1388 VPWR.n1387 5.97436
R7078 VPWR.n606 VPWR.n605 5.8885
R7079 VPWR.n1780 VPWR.n1779 5.8885
R7080 VPWR.n1451 VPWR.n1446 5.85193
R7081 VPWR.n1321 VPWR.n1081 5.66607
R7082 VPWR.n1270 VPWR.n1269 5.66607
R7083 VPWR.n634 VPWR.n633 5.66204
R7084 VPWR.n626 VPWR.n625 5.66204
R7085 VPWR.n625 VPWR.n247 5.66204
R7086 VPWR.n536 VPWR.n528 5.66204
R7087 VPWR.n537 VPWR.n536 5.66204
R7088 VPWR.n596 VPWR.n595 5.66204
R7089 VPWR.n558 VPWR.n552 5.66204
R7090 VPWR.n559 VPWR.n558 5.66204
R7091 VPWR.n584 VPWR.n559 5.66204
R7092 VPWR.n584 VPWR.n583 5.66204
R7093 VPWR.n571 VPWR.n570 5.66204
R7094 VPWR.n567 VPWR.n566 5.66204
R7095 VPWR.n566 VPWR.n25 5.66204
R7096 VPWR.n2315 VPWR.n25 5.66204
R7097 VPWR.n2315 VPWR.n2314 5.66204
R7098 VPWR.n2186 VPWR.n166 5.66204
R7099 VPWR.n2190 VPWR.n166 5.66204
R7100 VPWR.n2197 VPWR.n2196 5.66204
R7101 VPWR.n2178 VPWR.n2177 5.66204
R7102 VPWR.n2180 VPWR.n2178 5.66204
R7103 VPWR.n2152 VPWR.n173 5.66204
R7104 VPWR.n2167 VPWR.n173 5.66204
R7105 VPWR.n2170 VPWR.n2169 5.66204
R7106 VPWR.n2107 VPWR.n200 5.66204
R7107 VPWR.n2111 VPWR.n200 5.66204
R7108 VPWR.n2115 VPWR.n2113 5.66204
R7109 VPWR.n2115 VPWR.n2114 5.66204
R7110 VPWR.n2100 VPWR.n2099 5.66204
R7111 VPWR.n1185 VPWR.n1184 5.66204
R7112 VPWR.n1186 VPWR.n1185 5.66204
R7113 VPWR.n1190 VPWR.n1189 5.66204
R7114 VPWR.n1193 VPWR.n1190 5.66204
R7115 VPWR.n1193 VPWR.n1192 5.66204
R7116 VPWR.n2340 VPWR.n2339 5.66204
R7117 VPWR.n2339 VPWR.n5 5.66204
R7118 VPWR.n2335 VPWR.n2334 5.66204
R7119 VPWR.n2334 VPWR.n2333 5.66204
R7120 VPWR.n2333 VPWR.n8 5.66204
R7121 VPWR.n359 VPWR.n8 5.66204
R7122 VPWR.n360 VPWR.n359 5.66204
R7123 VPWR.n361 VPWR.n360 5.66204
R7124 VPWR.n368 VPWR.n367 5.66204
R7125 VPWR.n369 VPWR.n368 5.66204
R7126 VPWR.n373 VPWR.n372 5.66204
R7127 VPWR.n374 VPWR.n373 5.66204
R7128 VPWR.n374 VPWR.n345 5.66204
R7129 VPWR.n383 VPWR.n345 5.66204
R7130 VPWR.n384 VPWR.n383 5.66204
R7131 VPWR.n386 VPWR.n384 5.66204
R7132 VPWR.n322 VPWR.n321 5.66204
R7133 VPWR.n329 VPWR.n259 5.66204
R7134 VPWR.n333 VPWR.n259 5.66204
R7135 VPWR.n336 VPWR.n335 5.66204
R7136 VPWR.n510 VPWR.n336 5.66204
R7137 VPWR.n469 VPWR.n468 5.66204
R7138 VPWR.n468 VPWR.n418 5.66204
R7139 VPWR.n464 VPWR.n463 5.66204
R7140 VPWR.n463 VPWR.n462 5.66204
R7141 VPWR.n462 VPWR.n421 5.66204
R7142 VPWR.n458 VPWR.n421 5.66204
R7143 VPWR.n458 VPWR.n457 5.66204
R7144 VPWR.n457 VPWR.n456 5.66204
R7145 VPWR.n581 VPWR.n560 5.48759
R7146 VPWR.n602 VPWR.n601 5.42606
R7147 VPWR.n577 VPWR.n576 5.42606
R7148 VPWR.n37 VPWR.n36 5.3712
R7149 VPWR.n634 VPWR.n243 5.29281
R7150 VPWR.n633 VPWR.n632 5.29281
R7151 VPWR.n627 VPWR.n626 5.29281
R7152 VPWR.n538 VPWR.n537 5.29281
R7153 VPWR.n598 VPWR.n542 5.29281
R7154 VPWR.n583 VPWR.n582 5.29281
R7155 VPWR.n573 VPWR.n561 5.29281
R7156 VPWR.n2314 VPWR.n26 5.29281
R7157 VPWR.n2186 VPWR.n2185 5.29281
R7158 VPWR.n2196 VPWR.n2193 5.29281
R7159 VPWR.n2177 VPWR.n170 5.29281
R7160 VPWR.n2152 VPWR.n2151 5.29281
R7161 VPWR.n2170 VPWR.n171 5.29281
R7162 VPWR.n2107 VPWR.n2106 5.29281
R7163 VPWR.n2114 VPWR.n189 5.29281
R7164 VPWR.n2099 VPWR.n2098 5.29281
R7165 VPWR.n2100 VPWR.n202 5.29281
R7166 VPWR.n1176 VPWR.n1175 5.29281
R7167 VPWR.n1176 VPWR.n1119 5.29281
R7168 VPWR.n1192 VPWR.n1191 5.29281
R7169 VPWR.n2341 VPWR.n2340 5.29281
R7170 VPWR.n361 VPWR.n350 5.29281
R7171 VPWR.n367 VPWR.n349 5.29281
R7172 VPWR.n386 VPWR.n385 5.29281
R7173 VPWR.n321 VPWR.n320 5.29281
R7174 VPWR.n322 VPWR.n261 5.29281
R7175 VPWR.n329 VPWR.n328 5.29281
R7176 VPWR.n510 VPWR.n509 5.29281
R7177 VPWR.n470 VPWR.n469 5.29281
R7178 VPWR.n456 VPWR.n423 5.29281
R7179 VPWR.n1509 VPWR.n1499 5.27109
R7180 VPWR.n1829 VPWR.n1743 5.27109
R7181 VPWR.n1134 VPWR.n1133 5.25888
R7182 VPWR.n1216 VPWR.n1079 5.2464
R7183 VPWR.n1267 VPWR.n1265 5.2464
R7184 VPWR.n2301 VPWR.n2300 5.18397
R7185 VPWR.n73 VPWR.n72 5.18397
R7186 VPWR.n1307 VPWR.n1094 5.18397
R7187 VPWR.n1967 VPWR.n732 5.18397
R7188 VPWR.n1959 VPWR.n735 5.18397
R7189 VPWR.n1219 VPWR.n1217 5.14148
R7190 VPWR.n1436 VPWR.n1435 5.1205
R7191 VPWR.n1282 VPWR.n1260 5.103
R7192 VPWR.n682 VPWR.n680 5.03657
R7193 VPWR.t390 VPWR.t776 5.03584
R7194 VPWR.t61 VPWR.t741 5.03584
R7195 VPWR.t71 VPWR.t519 5.03584
R7196 VPWR.t817 VPWR.t85 5.03584
R7197 VPWR.t821 VPWR.t140 5.03584
R7198 VPWR.n907 VPWR.n871 4.98336
R7199 VPWR.n1503 VPWR.n1500 4.9005
R7200 VPWR.n1147 VPWR.n1146 4.69218
R7201 VPWR.n2261 VPWR.n2259 4.67352
R7202 VPWR.n1983 VPWR.n1982 4.67352
R7203 VPWR.n1410 VPWR.n1409 4.67352
R7204 VPWR.n1611 VPWR.n1608 4.67352
R7205 VPWR.n1921 VPWR.n1920 4.67352
R7206 VPWR.n1920 VPWR.n829 4.67352
R7207 VPWR.n1728 VPWR.n950 4.67352
R7208 VPWR.n1734 VPWR.n1730 4.67352
R7209 VPWR.n1713 VPWR.n1712 4.67352
R7210 VPWR.n1819 VPWR.n1818 4.67352
R7211 VPWR.n1870 VPWR.n846 4.67352
R7212 VPWR.n1866 VPWR.n1865 4.67352
R7213 VPWR.n1865 VPWR.n1864 4.67352
R7214 VPWR.n917 VPWR.n916 4.67352
R7215 VPWR.n916 VPWR.n868 4.67352
R7216 VPWR.n912 VPWR.n868 4.67352
R7217 VPWR.n903 VPWR.n902 4.67352
R7218 VPWR.n902 VPWR.n873 4.67352
R7219 VPWR.n2249 VPWR.n2248 4.62124
R7220 VPWR.n1596 VPWR.n1595 4.62124
R7221 VPWR.n610 VPWR.n609 4.62124
R7222 VPWR.n603 VPWR.n541 4.62124
R7223 VPWR.n579 VPWR.n578 4.62124
R7224 VPWR.n1143 VPWR.n1134 4.62124
R7225 VPWR.n1783 VPWR.n1782 4.62124
R7226 VPWR.n1777 VPWR.n1767 4.62124
R7227 VPWR.n907 VPWR.n905 4.62124
R7228 VPWR.n1390 VPWR.n1386 4.5918
R7229 VPWR.n2258 VPWR.n2257 4.57193
R7230 VPWR.n1922 VPWR.n1921 4.57193
R7231 VPWR.n1964 VPWR.n732 4.54926
R7232 VPWR.n1962 VPWR.n735 4.54926
R7233 VPWR.n756 VPWR.n755 4.54926
R7234 VPWR.n798 VPWR.n756 4.54926
R7235 VPWR.n1228 VPWR.n1208 4.52113
R7236 VPWR.n1499 VPWR.n1498 4.51815
R7237 VPWR.n407 VPWR.n405 4.51401
R7238 VPWR.n474 VPWR.n473 4.51401
R7239 VPWR.n1857 VPWR.n1856 4.51401
R7240 VPWR.n919 VPWR.n858 4.51401
R7241 VPWR.n520 VPWR.n253 4.51401
R7242 VPWR.n258 VPWR.n257 4.51401
R7243 VPWR.n305 VPWR.n270 4.51401
R7244 VPWR.n310 VPWR.n309 4.51401
R7245 VPWR.n1947 VPWR.n814 4.51401
R7246 VPWR.n819 VPWR.n818 4.51401
R7247 VPWR.n11 VPWR.n9 4.51401
R7248 VPWR.n357 VPWR.n356 4.51401
R7249 VPWR.n381 VPWR.n380 4.51401
R7250 VPWR.n394 VPWR.n393 4.51401
R7251 VPWR.n2290 VPWR.n2289 4.51401
R7252 VPWR.n81 VPWR.n69 4.51401
R7253 VPWR.n593 VPWR.n592 4.51401
R7254 VPWR.n587 VPWR.n586 4.51401
R7255 VPWR.n622 VPWR.n621 4.51401
R7256 VPWR.n617 VPWR.n616 4.51401
R7257 VPWR.n658 VPWR.n213 4.51401
R7258 VPWR.n649 VPWR.n645 4.51401
R7259 VPWR.n107 VPWR.n106 4.51401
R7260 VPWR.n118 VPWR.n52 4.51401
R7261 VPWR.n2319 VPWR.n22 4.51401
R7262 VPWR.n2310 VPWR.n2309 4.51401
R7263 VPWR.n2230 VPWR.n2228 4.51401
R7264 VPWR.n2244 VPWR.n2243 4.51401
R7265 VPWR.n2160 VPWR.n180 4.51401
R7266 VPWR.n2165 VPWR.n2164 4.51401
R7267 VPWR.n2122 VPWR.n196 4.51401
R7268 VPWR.n2127 VPWR.n2126 4.51401
R7269 VPWR.n2083 VPWR.n2048 4.51401
R7270 VPWR.n2088 VPWR.n2087 4.51401
R7271 VPWR.n2265 VPWR.n2264 4.51401
R7272 VPWR.n2276 VPWR.n127 4.51401
R7273 VPWR.n2201 VPWR.n161 4.51401
R7274 VPWR.n2206 VPWR.n2205 4.51401
R7275 VPWR.n2038 VPWR.n669 4.51401
R7276 VPWR.n676 VPWR.n673 4.51401
R7277 VPWR.n1335 VPWR.n1074 4.51401
R7278 VPWR.n1328 VPWR.n1327 4.51401
R7279 VPWR.n1200 VPWR.n1112 4.51401
R7280 VPWR.n1205 VPWR.n1204 4.51401
R7281 VPWR.n1152 VPWR.n1151 4.51401
R7282 VPWR.n1166 VPWR.n1165 4.51401
R7283 VPWR.n697 VPWR.n695 4.51401
R7284 VPWR.n707 VPWR.n706 4.51401
R7285 VPWR.n1300 VPWR.n1299 4.51401
R7286 VPWR.n1294 VPWR.n1293 4.51401
R7287 VPWR.n740 VPWR.n738 4.51401
R7288 VPWR.n809 VPWR.n808 4.51401
R7289 VPWR.n1537 VPWR.n1341 4.51401
R7290 VPWR.n1530 VPWR.n1529 4.51401
R7291 VPWR.n1442 VPWR.n1441 4.51401
R7292 VPWR.n1459 VPWR.n1458 4.51401
R7293 VPWR.n1397 VPWR.n1396 4.51401
R7294 VPWR.n1407 VPWR.n1406 4.51401
R7295 VPWR.n788 VPWR.n787 4.51401
R7296 VPWR.n778 VPWR.n777 4.51401
R7297 VPWR.n1987 VPWR.n714 4.51401
R7298 VPWR.n1978 VPWR.n1977 4.51401
R7299 VPWR.n1602 VPWR.n1601 4.51401
R7300 VPWR.n1619 VPWR.n1618 4.51401
R7301 VPWR.n1808 VPWR.n935 4.51401
R7302 VPWR.n1799 VPWR.n936 4.51401
R7303 VPWR.n1577 VPWR.n1542 4.51401
R7304 VPWR.n1582 VPWR.n1581 4.51401
R7305 VPWR.n1035 VPWR.n1034 4.51401
R7306 VPWR.n1656 VPWR.n1655 4.51401
R7307 VPWR.n1917 VPWR.n1916 4.51401
R7308 VPWR.n1907 VPWR.n1906 4.51401
R7309 VPWR.n1697 VPWR.n994 4.51401
R7310 VPWR.n1687 VPWR.n1683 4.51401
R7311 VPWR.n1736 VPWR.n943 4.51401
R7312 VPWR.n945 VPWR.n942 4.51401
R7313 VPWR.n990 VPWR.n964 4.51401
R7314 VPWR.n1705 VPWR.n960 4.51401
R7315 VPWR.n899 VPWR.n898 4.51401
R7316 VPWR.n890 VPWR.n876 4.51401
R7317 VPWR.n1771 VPWR.n838 4.51401
R7318 VPWR.n841 VPWR.n836 4.51401
R7319 VPWR.n454 VPWR.n453 4.51401
R7320 VPWR.n443 VPWR.n427 4.51401
R7321 VPWR.n1217 VPWR.n1216 4.51198
R7322 VPWR.n2016 VPWR.n682 4.51198
R7323 VPWR.n110 VPWR.n109 4.5005
R7324 VPWR.n111 VPWR.n54 4.5005
R7325 VPWR.n120 VPWR.n119 4.5005
R7326 VPWR.n657 VPWR.n656 4.5005
R7327 VPWR.n646 VPWR.n215 4.5005
R7328 VPWR.n651 VPWR.n650 4.5005
R7329 VPWR.n529 VPWR.n249 4.5005
R7330 VPWR.n533 VPWR.n532 4.5005
R7331 VPWR.n534 VPWR.n525 4.5005
R7332 VPWR.n553 VPWR.n546 4.5005
R7333 VPWR.n556 VPWR.n555 4.5005
R7334 VPWR.n554 VPWR.n549 4.5005
R7335 VPWR.n76 VPWR.n45 4.5005
R7336 VPWR.n78 VPWR.n77 4.5005
R7337 VPWR.n83 VPWR.n82 4.5005
R7338 VPWR.n2318 VPWR.n2317 4.5005
R7339 VPWR.n28 VPWR.n24 4.5005
R7340 VPWR.n2312 VPWR.n2311 4.5005
R7341 VPWR.n2268 VPWR.n2267 4.5005
R7342 VPWR.n2269 VPWR.n129 4.5005
R7343 VPWR.n2278 VPWR.n2277 4.5005
R7344 VPWR.n2082 VPWR.n2081 4.5005
R7345 VPWR.n2052 VPWR.n2051 4.5005
R7346 VPWR.n208 VPWR.n207 4.5005
R7347 VPWR.n2121 VPWR.n2120 4.5005
R7348 VPWR.n2119 VPWR.n2118 4.5005
R7349 VPWR.n199 VPWR.n191 4.5005
R7350 VPWR.n2159 VPWR.n2158 4.5005
R7351 VPWR.n2156 VPWR.n2155 4.5005
R7352 VPWR.n175 VPWR.n174 4.5005
R7353 VPWR.n2232 VPWR.n2231 4.5005
R7354 VPWR.n2239 VPWR.n2238 4.5005
R7355 VPWR.n145 VPWR.n144 4.5005
R7356 VPWR.n2200 VPWR.n2199 4.5005
R7357 VPWR.n165 VPWR.n164 4.5005
R7358 VPWR.n2194 VPWR.n157 4.5005
R7359 VPWR.n2001 VPWR.n2000 4.5005
R7360 VPWR.n702 VPWR.n698 4.5005
R7361 VPWR.n704 VPWR.n701 4.5005
R7362 VPWR.n1149 VPWR.n1128 4.5005
R7363 VPWR.n1161 VPWR.n1160 4.5005
R7364 VPWR.n1125 VPWR.n1124 4.5005
R7365 VPWR.n1199 VPWR.n1198 4.5005
R7366 VPWR.n1197 VPWR.n1196 4.5005
R7367 VPWR.n1115 VPWR.n1106 4.5005
R7368 VPWR.n1334 VPWR.n1333 4.5005
R7369 VPWR.n1323 VPWR.n1077 4.5005
R7370 VPWR.n1326 VPWR.n1082 4.5005
R7371 VPWR.n2037 VPWR.n2036 4.5005
R7372 VPWR.n2035 VPWR.n2034 4.5005
R7373 VPWR.n2031 VPWR.n2030 4.5005
R7374 VPWR.n1098 VPWR.n1097 4.5005
R7375 VPWR.n1249 VPWR.n1248 4.5005
R7376 VPWR.n1250 VPWR.n1101 4.5005
R7377 VPWR.n764 VPWR.n761 4.5005
R7378 VPWR.n783 VPWR.n782 4.5005
R7379 VPWR.n775 VPWR.n766 4.5005
R7380 VPWR.n1394 VPWR.n1393 4.5005
R7381 VPWR.n1402 VPWR.n1401 4.5005
R7382 VPWR.n1372 VPWR.n1368 4.5005
R7383 VPWR.n1439 VPWR.n1355 4.5005
R7384 VPWR.n1454 VPWR.n1453 4.5005
R7385 VPWR.n1356 VPWR.n1352 4.5005
R7386 VPWR.n1536 VPWR.n1535 4.5005
R7387 VPWR.n1525 VPWR.n1344 4.5005
R7388 VPWR.n1528 VPWR.n1489 4.5005
R7389 VPWR.n1955 VPWR.n1954 4.5005
R7390 VPWR.n741 VPWR.n739 4.5005
R7391 VPWR.n748 VPWR.n744 4.5005
R7392 VPWR.n1986 VPWR.n1985 4.5005
R7393 VPWR.n721 VPWR.n716 4.5005
R7394 VPWR.n1980 VPWR.n1979 4.5005
R7395 VPWR.n1893 VPWR.n831 4.5005
R7396 VPWR.n1912 VPWR.n1911 4.5005
R7397 VPWR.n1904 VPWR.n1895 4.5005
R7398 VPWR.n1663 VPWR.n1662 4.5005
R7399 VPWR.n1041 VPWR.n1036 4.5005
R7400 VPWR.n1043 VPWR.n1040 4.5005
R7401 VPWR.n1576 VPWR.n1575 4.5005
R7402 VPWR.n1573 VPWR.n1572 4.5005
R7403 VPWR.n1070 VPWR.n1069 4.5005
R7404 VPWR.n1599 VPWR.n1598 4.5005
R7405 VPWR.n1614 VPWR.n1613 4.5005
R7406 VPWR.n1052 VPWR.n1048 4.5005
R7407 VPWR.n1946 VPWR.n1945 4.5005
R7408 VPWR.n1944 VPWR.n1943 4.5005
R7409 VPWR.n1940 VPWR.n1939 4.5005
R7410 VPWR.n1696 VPWR.n1695 4.5005
R7411 VPWR.n1684 VPWR.n996 4.5005
R7412 VPWR.n1689 VPWR.n1688 4.5005
R7413 VPWR.n878 VPWR.n875 4.5005
R7414 VPWR.n895 VPWR.n894 4.5005
R7415 VPWR.n881 VPWR.n880 4.5005
R7416 VPWR.n989 VPWR.n988 4.5005
R7417 VPWR.n962 VPWR.n959 4.5005
R7418 VPWR.n1707 VPWR.n1706 4.5005
R7419 VPWR.n1739 VPWR.n1738 4.5005
R7420 VPWR.n1740 VPWR.n944 4.5005
R7421 VPWR.n1832 VPWR.n1831 4.5005
R7422 VPWR.n1806 VPWR.n1805 4.5005
R7423 VPWR.n1756 VPWR.n1755 4.5005
R7424 VPWR.n1761 VPWR.n1760 4.5005
R7425 VPWR.n859 VPWR.n855 4.5005
R7426 VPWR.n927 VPWR.n926 4.5005
R7427 VPWR.n864 VPWR.n863 4.5005
R7428 VPWR.n1773 VPWR.n1772 4.5005
R7429 VPWR.n1774 VPWR.n839 4.5005
R7430 VPWR.n1881 VPWR.n1880 4.5005
R7431 VPWR.n435 VPWR.n425 4.5005
R7432 VPWR.n436 VPWR.n429 4.5005
R7433 VPWR.n445 VPWR.n444 4.5005
R7434 VPWR.n304 VPWR.n303 4.5005
R7435 VPWR.n274 VPWR.n273 4.5005
R7436 VPWR.n267 VPWR.n266 4.5005
R7437 VPWR.n519 VPWR.n518 4.5005
R7438 VPWR.n517 VPWR.n516 4.5005
R7439 VPWR.n513 VPWR.n512 4.5005
R7440 VPWR.n2331 VPWR.n2330 4.5005
R7441 VPWR.n352 VPWR.n12 4.5005
R7442 VPWR.n355 VPWR.n353 4.5005
R7443 VPWR.n378 VPWR.n377 4.5005
R7444 VPWR.n389 VPWR.n388 4.5005
R7445 VPWR.n344 VPWR.n340 4.5005
R7446 VPWR.n481 VPWR.n480 4.5005
R7447 VPWR.n408 VPWR.n406 4.5005
R7448 VPWR.n415 VPWR.n411 4.5005
R7449 VPWR.n2134 VPWR.n185 4.49637
R7450 VPWR.n1331 VPWR.n1079 4.40706
R7451 VPWR.n1272 VPWR.n1267 4.40706
R7452 VPWR.n2261 VPWR.n2260 4.36875
R7453 VPWR.n1228 VPWR.n1227 4.36875
R7454 VPWR.n1411 VPWR.n1410 4.36875
R7455 VPWR.n1923 VPWR.n826 4.36875
R7456 VPWR.n1896 VPWR.n829 4.36875
R7457 VPWR.n1723 VPWR.n950 4.36875
R7458 VPWR.n1730 VPWR.n1729 4.36875
R7459 VPWR.n1713 VPWR.n956 4.36875
R7460 VPWR.n1823 VPWR.n1822 4.36875
R7461 VPWR.n1819 VPWR.n1746 4.36875
R7462 VPWR.n1816 VPWR.n1749 4.36875
R7463 VPWR.n1873 VPWR.n845 4.36875
R7464 VPWR.n917 VPWR.n862 4.36875
R7465 VPWR.n882 VPWR.n873 4.36875
R7466 VPWR.n2300 VPWR.n2299 4.33769
R7467 VPWR.n1132 VPWR.n1131 4.29023
R7468 VPWR.n724 VPWR.n719 4.26717
R7469 VPWR.n2248 VPWR.n138 4.14168
R7470 VPWR.n224 VPWR.n220 4.02033
R7471 VPWR.n224 VPWR.n223 4.02033
R7472 VPWR.n233 VPWR.n227 4.02033
R7473 VPWR.n233 VPWR.n232 4.02033
R7474 VPWR.n116 VPWR.n65 4.02033
R7475 VPWR.n116 VPWR.n115 4.02033
R7476 VPWR.n2134 VPWR.n2133 4.02033
R7477 VPWR.n2073 VPWR.n2058 4.02033
R7478 VPWR.n2073 VPWR.n2064 4.02033
R7479 VPWR.n2072 VPWR.n2067 4.02033
R7480 VPWR.n2072 VPWR.n2071 4.02033
R7481 VPWR.n2274 VPWR.n134 4.02033
R7482 VPWR.n2274 VPWR.n2273 4.02033
R7483 VPWR.n1141 VPWR.n1137 4.02033
R7484 VPWR.n1141 VPWR.n1140 4.02033
R7485 VPWR.n694 VPWR.n690 4.02033
R7486 VPWR.n694 VPWR.n693 4.02033
R7487 VPWR.n1382 VPWR.n1378 4.02033
R7488 VPWR.n1382 VPWR.n1381 4.02033
R7489 VPWR.n780 VPWR.n771 4.02033
R7490 VPWR.n780 VPWR.n774 4.02033
R7491 VPWR.n1010 VPWR.n1006 4.02033
R7492 VPWR.n1010 VPWR.n1009 4.02033
R7493 VPWR.n1033 VPWR.n1031 4.02033
R7494 VPWR.n1648 VPWR.n1625 4.02033
R7495 VPWR.n1909 VPWR.n1900 4.02033
R7496 VPWR.n1909 VPWR.n1903 4.02033
R7497 VPWR.n978 VPWR.n973 4.02033
R7498 VPWR.n978 VPWR.n977 4.02033
R7499 VPWR.n892 VPWR.n886 4.02033
R7500 VPWR.n892 VPWR.n889 4.02033
R7501 VPWR.n3 VPWR.n2 4.02033
R7502 VPWR.n283 VPWR.n279 4.02033
R7503 VPWR.n283 VPWR.n282 4.02033
R7504 VPWR.n292 VPWR.n286 4.02033
R7505 VPWR.n292 VPWR.n291 4.02033
R7506 VPWR.n441 VPWR.n434 4.02033
R7507 VPWR.n441 VPWR.n440 4.02033
R7508 VPWR.n1330 VPWR.n1081 3.98739
R7509 VPWR.n1271 VPWR.n1270 3.98739
R7510 VPWR.n72 VPWR.n70 3.91455
R7511 VPWR.n1817 VPWR.n1816 3.86082
R7512 VPWR.n603 VPWR.n602 3.78037
R7513 VPWR.n578 VPWR.n577 3.78037
R7514 VPWR.n609 VPWR.n608 3.75517
R7515 VPWR.n35 VPWR.n34 3.75222
R7516 VPWR.n578 VPWR.n560 3.69446
R7517 VPWR.n1782 VPWR.n1766 3.66983
R7518 VPWR.n1733 VPWR.n1732 3.55606
R7519 VPWR.n1131 VPWR.n1130 3.53179
R7520 VPWR.n1533 VPWR.n1487 3.4812
R7521 VPWR.n654 VPWR.n653 3.47425
R7522 VPWR.n643 VPWR.n642 3.47425
R7523 VPWR.n642 VPWR.n641 3.47425
R7524 VPWR.n2213 VPWR.n2212 3.47425
R7525 VPWR.n2143 VPWR.n2142 3.47425
R7526 VPWR.n2146 VPWR.n2143 3.47425
R7527 VPWR.n2079 VPWR.n2078 3.47425
R7528 VPWR.n2091 VPWR.n2090 3.47425
R7529 VPWR.n2093 VPWR.n2091 3.47425
R7530 VPWR.n1168 VPWR.n1123 3.47425
R7531 VPWR.n1169 VPWR.n1168 3.47425
R7532 VPWR.n1170 VPWR.n1169 3.47425
R7533 VPWR.n1252 VPWR.n1246 3.47425
R7534 VPWR.n2006 VPWR.n2005 3.47425
R7535 VPWR.n793 VPWR.n792 3.47425
R7536 VPWR.n792 VPWR.n791 3.47425
R7537 VPWR.n791 VPWR.n759 3.47425
R7538 VPWR.n1797 VPWR.n1796 3.47425
R7539 VPWR.n301 VPWR.n300 3.47425
R7540 VPWR.n313 VPWR.n312 3.47425
R7541 VPWR.n315 VPWR.n313 3.47425
R7542 VPWR.n490 VPWR.n489 3.47425
R7543 VPWR.n489 VPWR.n488 3.47425
R7544 VPWR.n488 VPWR.n401 3.47425
R7545 VPWR.n475 VPWR.n474 3.43925
R7546 VPWR.n477 VPWR.n407 3.43925
R7547 VPWR.n257 VPWR.n251 3.43925
R7548 VPWR.n521 VPWR.n520 3.43925
R7549 VPWR.n309 VPWR.n308 3.43925
R7550 VPWR.n306 VPWR.n305 3.43925
R7551 VPWR.n818 VPWR.n811 3.43925
R7552 VPWR.n1948 VPWR.n1947 3.43925
R7553 VPWR.n356 VPWR.n14 3.43925
R7554 VPWR.n2327 VPWR.n11 3.43925
R7555 VPWR.n393 VPWR.n392 3.43925
R7556 VPWR.n380 VPWR.n379 3.43925
R7557 VPWR.n81 VPWR.n48 3.43925
R7558 VPWR.n2289 VPWR.n2288 3.43925
R7559 VPWR.n588 VPWR.n587 3.43925
R7560 VPWR.n592 VPWR.n591 3.43925
R7561 VPWR.n618 VPWR.n617 3.43925
R7562 VPWR.n621 VPWR.n620 3.43925
R7563 VPWR.n649 VPWR.n211 3.43925
R7564 VPWR.n659 VPWR.n658 3.43925
R7565 VPWR.n123 VPWR.n52 3.43925
R7566 VPWR.n107 VPWR.n51 3.43925
R7567 VPWR.n2310 VPWR.n19 3.43925
R7568 VPWR.n2320 VPWR.n2319 3.43925
R7569 VPWR.n2243 VPWR.n2242 3.43925
R7570 VPWR.n2230 VPWR.n2229 3.43925
R7571 VPWR.n2164 VPWR.n2163 3.43925
R7572 VPWR.n2161 VPWR.n2160 3.43925
R7573 VPWR.n2126 VPWR.n2125 3.43925
R7574 VPWR.n2123 VPWR.n2122 3.43925
R7575 VPWR.n2087 VPWR.n2086 3.43925
R7576 VPWR.n2084 VPWR.n2083 3.43925
R7577 VPWR.n2281 VPWR.n127 3.43925
R7578 VPWR.n2265 VPWR.n125 3.43925
R7579 VPWR.n2205 VPWR.n2204 3.43925
R7580 VPWR.n2202 VPWR.n2201 3.43925
R7581 VPWR.n673 VPWR.n666 3.43925
R7582 VPWR.n2039 VPWR.n2038 3.43925
R7583 VPWR.n1327 VPWR.n1072 3.43925
R7584 VPWR.n1336 VPWR.n1335 3.43925
R7585 VPWR.n1204 VPWR.n1203 3.43925
R7586 VPWR.n1201 VPWR.n1200 3.43925
R7587 VPWR.n1165 VPWR.n1164 3.43925
R7588 VPWR.n1151 VPWR.n1150 3.43925
R7589 VPWR.n1996 VPWR.n707 3.43925
R7590 VPWR.n699 VPWR.n697 3.43925
R7591 VPWR.n1295 VPWR.n1294 3.43925
R7592 VPWR.n1299 VPWR.n1298 3.43925
R7593 VPWR.n810 VPWR.n809 3.43925
R7594 VPWR.n1951 VPWR.n740 3.43925
R7595 VPWR.n1529 VPWR.n1339 3.43925
R7596 VPWR.n1538 VPWR.n1537 3.43925
R7597 VPWR.n1458 VPWR.n1457 3.43925
R7598 VPWR.n1441 VPWR.n1440 3.43925
R7599 VPWR.n1406 VPWR.n1405 3.43925
R7600 VPWR.n1396 VPWR.n1395 3.43925
R7601 VPWR.n777 VPWR.n776 3.43925
R7602 VPWR.n787 VPWR.n786 3.43925
R7603 VPWR.n1978 VPWR.n711 3.43925
R7604 VPWR.n1988 VPWR.n1987 3.43925
R7605 VPWR.n1618 VPWR.n1617 3.43925
R7606 VPWR.n1601 VPWR.n1600 3.43925
R7607 VPWR.n1657 VPWR.n1656 3.43925
R7608 VPWR.n1659 VPWR.n1035 3.43925
R7609 VPWR.n1906 VPWR.n1905 3.43925
R7610 VPWR.n1916 VPWR.n1915 3.43925
R7611 VPWR.n1687 VPWR.n992 3.43925
R7612 VPWR.n1698 VPWR.n1697 3.43925
R7613 VPWR.n453 VPWR.n452 3.43925
R7614 VPWR.n448 VPWR.n427 3.43925
R7615 VPWR.n1797 VPWR.n1759 3.43649
R7616 VPWR.n479 VPWR.n478 3.4105
R7617 VPWR.n410 VPWR.n409 3.4105
R7618 VPWR.n254 VPWR.n252 3.4105
R7619 VPWR.n515 VPWR.n514 3.4105
R7620 VPWR.n271 VPWR.n269 3.4105
R7621 VPWR.n272 VPWR.n268 3.4105
R7622 VPWR.n815 VPWR.n813 3.4105
R7623 VPWR.n1942 VPWR.n1941 3.4105
R7624 VPWR.n2329 VPWR.n2328 3.4105
R7625 VPWR.n354 VPWR.n13 3.4105
R7626 VPWR.n342 VPWR.n341 3.4105
R7627 VPWR.n391 VPWR.n390 3.4105
R7628 VPWR.n75 VPWR.n46 3.4105
R7629 VPWR.n80 VPWR.n79 3.4105
R7630 VPWR.n590 VPWR.n547 3.4105
R7631 VPWR.n589 VPWR.n548 3.4105
R7632 VPWR.n530 VPWR.n250 3.4105
R7633 VPWR.n531 VPWR.n524 3.4105
R7634 VPWR.n214 VPWR.n212 3.4105
R7635 VPWR.n648 VPWR.n647 3.4105
R7636 VPWR.n108 VPWR.n53 3.4105
R7637 VPWR.n122 VPWR.n121 3.4105
R7638 VPWR.n23 VPWR.n21 3.4105
R7639 VPWR.n30 VPWR.n29 3.4105
R7640 VPWR.n147 VPWR.n146 3.4105
R7641 VPWR.n2241 VPWR.n2240 3.4105
R7642 VPWR.n181 VPWR.n179 3.4105
R7643 VPWR.n2154 VPWR.n176 3.4105
R7644 VPWR.n197 VPWR.n195 3.4105
R7645 VPWR.n2117 VPWR.n192 3.4105
R7646 VPWR.n2049 VPWR.n2047 3.4105
R7647 VPWR.n2050 VPWR.n209 3.4105
R7648 VPWR.n2266 VPWR.n128 3.4105
R7649 VPWR.n2280 VPWR.n2279 3.4105
R7650 VPWR.n162 VPWR.n160 3.4105
R7651 VPWR.n163 VPWR.n158 3.4105
R7652 VPWR.n670 VPWR.n668 3.4105
R7653 VPWR.n2033 VPWR.n2032 3.4105
R7654 VPWR.n1075 VPWR.n1073 3.4105
R7655 VPWR.n1325 VPWR.n1324 3.4105
R7656 VPWR.n1113 VPWR.n1111 3.4105
R7657 VPWR.n1195 VPWR.n1107 3.4105
R7658 VPWR.n1127 VPWR.n1126 3.4105
R7659 VPWR.n1163 VPWR.n1162 3.4105
R7660 VPWR.n1999 VPWR.n1998 3.4105
R7661 VPWR.n1997 VPWR.n700 3.4105
R7662 VPWR.n1297 VPWR.n1099 3.4105
R7663 VPWR.n1296 VPWR.n1100 3.4105
R7664 VPWR.n1953 VPWR.n1952 3.4105
R7665 VPWR.n743 VPWR.n742 3.4105
R7666 VPWR.n1342 VPWR.n1340 3.4105
R7667 VPWR.n1527 VPWR.n1526 3.4105
R7668 VPWR.n1354 VPWR.n1353 3.4105
R7669 VPWR.n1456 VPWR.n1455 3.4105
R7670 VPWR.n1370 VPWR.n1369 3.4105
R7671 VPWR.n1404 VPWR.n1403 3.4105
R7672 VPWR.n785 VPWR.n784 3.4105
R7673 VPWR.n763 VPWR.n762 3.4105
R7674 VPWR.n715 VPWR.n713 3.4105
R7675 VPWR.n723 VPWR.n722 3.4105
R7676 VPWR.n1050 VPWR.n1049 3.4105
R7677 VPWR.n1616 VPWR.n1615 3.4105
R7678 VPWR.n1843 VPWR.n936 3.4105
R7679 VPWR.n1843 VPWR.n935 3.4105
R7680 VPWR.n1843 VPWR.n937 3.4105
R7681 VPWR.n1843 VPWR.n934 3.4105
R7682 VPWR.n1580 VPWR.n1579 3.4105
R7683 VPWR.n1579 VPWR.n1578 3.4105
R7684 VPWR.n1581 VPWR.n1580 3.4105
R7685 VPWR.n1578 VPWR.n1577 3.4105
R7686 VPWR.n1543 VPWR.n1541 3.4105
R7687 VPWR.n1571 VPWR.n1071 3.4105
R7688 VPWR.n1661 VPWR.n1660 3.4105
R7689 VPWR.n1039 VPWR.n1037 3.4105
R7690 VPWR.n1914 VPWR.n1913 3.4105
R7691 VPWR.n1892 VPWR.n1891 3.4105
R7692 VPWR.n995 VPWR.n993 3.4105
R7693 VPWR.n1686 VPWR.n1685 3.4105
R7694 VPWR.n1834 VPWR.n942 3.4105
R7695 VPWR.n1834 VPWR.n943 3.4105
R7696 VPWR.n1834 VPWR.n941 3.4105
R7697 VPWR.n1834 VPWR.n1833 3.4105
R7698 VPWR.n1705 VPWR.n1704 3.4105
R7699 VPWR.n1704 VPWR.n990 3.4105
R7700 VPWR.n1704 VPWR.n963 3.4105
R7701 VPWR.n1704 VPWR.n961 3.4105
R7702 VPWR.n897 VPWR.n896 3.4105
R7703 VPWR.n897 VPWR.n877 3.4105
R7704 VPWR.n897 VPWR.n876 3.4105
R7705 VPWR.n898 VPWR.n897 3.4105
R7706 VPWR.n1883 VPWR.n836 3.4105
R7707 VPWR.n1883 VPWR.n838 3.4105
R7708 VPWR.n1883 VPWR.n835 3.4105
R7709 VPWR.n1883 VPWR.n1882 3.4105
R7710 VPWR.n1855 VPWR.n858 3.4105
R7711 VPWR.n1856 VPWR.n1855 3.4105
R7712 VPWR.n1855 VPWR.n928 3.4105
R7713 VPWR.n1855 VPWR.n856 3.4105
R7714 VPWR.n428 VPWR.n426 3.4105
R7715 VPWR.n447 VPWR.n446 3.4105
R7716 VPWR.t188 VPWR.t798 3.35739
R7717 VPWR.t18 VPWR.t743 3.35739
R7718 VPWR.t341 VPWR.t217 3.35739
R7719 VPWR.t273 VPWR.t656 3.35739
R7720 VPWR.n238 VPWR.n217 3.2477
R7721 VPWR.n641 VPWR.n242 3.2477
R7722 VPWR.n2213 VPWR.n153 3.2477
R7723 VPWR.n2142 VPWR.n184 3.2477
R7724 VPWR.n2054 VPWR.n2053 3.2477
R7725 VPWR.n2093 VPWR.n2092 3.2477
R7726 VPWR.n1154 VPWR.n1129 3.2477
R7727 VPWR.n1170 VPWR.n1121 3.2477
R7728 VPWR.n1253 VPWR.n1252 3.2477
R7729 VPWR.n2005 VPWR.n2004 3.2477
R7730 VPWR.n793 VPWR.n757 3.2477
R7731 VPWR.n767 VPWR.n759 3.2477
R7732 VPWR.n1802 VPWR.n1801 3.2477
R7733 VPWR.n1794 VPWR.n1763 3.2477
R7734 VPWR.n297 VPWR.n276 3.2477
R7735 VPWR.n315 VPWR.n314 3.2477
R7736 VPWR.n496 VPWR.n495 3.2477
R7737 VPWR.n402 VPWR.n401 3.2477
R7738 VPWR.n1409 VPWR.n1367 3.2005
R7739 VPWR.n605 VPWR.n604 3.151
R7740 VPWR.n1220 VPWR.n1219 3.14804
R7741 VPWR.n1277 VPWR.n1276 3.14804
R7742 VPWR.n868 VPWR.n867 3.12116
R7743 VPWR.n228 VPWR.n224 3.05586
R7744 VPWR.n2072 VPWR.n2068 3.05586
R7745 VPWR.n1142 VPWR.n1141 3.05586
R7746 VPWR.n1383 VPWR.n1382 3.05586
R7747 VPWR.n1011 VPWR.n1010 3.05586
R7748 VPWR.n978 VPWR.n974 3.05586
R7749 VPWR.n287 VPWR.n283 3.05586
R7750 VPWR.n233 VPWR.n229 3.04861
R7751 VPWR.n104 VPWR.n62 3.04861
R7752 VPWR.n2073 VPWR.n2061 3.04861
R7753 VPWR.n1648 VPWR.n1622 3.04861
R7754 VPWR.n292 VPWR.n288 3.04861
R7755 VPWR.n2303 VPWR.n37 3.04861
R7756 VPWR.n2133 VPWR.n2132 3.04861
R7757 VPWR.n2254 VPWR.n2251 3.04861
R7758 VPWR.n1399 VPWR.n1398 3.04861
R7759 VPWR.n2344 VPWR.n3 3.04861
R7760 VPWR.n527 VPWR.n247 3.01588
R7761 VPWR.n598 VPWR.n597 3.01588
R7762 VPWR.n595 VPWR.n544 3.01588
R7763 VPWR.n573 VPWR.n572 3.01588
R7764 VPWR.n570 VPWR.n563 3.01588
R7765 VPWR.n2191 VPWR.n2190 3.01588
R7766 VPWR.n2180 VPWR.n2179 3.01588
R7767 VPWR.n2168 VPWR.n2167 3.01588
R7768 VPWR.n2112 VPWR.n2111 3.01588
R7769 VPWR.n1186 VPWR.n1116 3.01588
R7770 VPWR.n7 VPWR.n5 3.01588
R7771 VPWR.n369 VPWR.n347 3.01588
R7772 VPWR.n334 VPWR.n333 3.01588
R7773 VPWR.n420 VPWR.n418 3.01588
R7774 VPWR.n95 VPWR.n66 3.01226
R7775 VPWR.n1514 VPWR.n1513 3.01226
R7776 VPWR.n1554 VPWR.n1553 3.01226
R7777 VPWR.n1693 VPWR.n1692 3.01226
R7778 VPWR.n1628 VPWR.n1626 3.01226
R7779 VPWR.n1640 VPWR.n1631 3.01226
R7780 VPWR.n2257 VPWR.n137 2.99733
R7781 VPWR.n903 VPWR.n871 2.99733
R7782 VPWR.n62 VPWR.n58 2.91308
R7783 VPWR.n62 VPWR.n61 2.91308
R7784 VPWR.n1003 VPWR.n999 2.91308
R7785 VPWR.n1003 VPWR.n1002 2.91308
R7786 VPWR.n2254 VPWR.n2253 2.87861
R7787 VPWR.n1095 VPWR.n1094 2.8567
R7788 VPWR.n607 VPWR.n605 2.8165
R7789 VPWR.n1781 VPWR.n1779 2.8165
R7790 VPWR.n239 VPWR.n216 2.6965
R7791 VPWR.n2076 VPWR.n2075 2.6965
R7792 VPWR.n298 VPWR.n275 2.6965
R7793 VPWR.n1611 VPWR.n1610 2.69256
R7794 VPWR.n528 VPWR.n527 2.64665
R7795 VPWR.n597 VPWR.n596 2.64665
R7796 VPWR.n552 VPWR.n544 2.64665
R7797 VPWR.n572 VPWR.n571 2.64665
R7798 VPWR.n567 VPWR.n563 2.64665
R7799 VPWR.n2197 VPWR.n2191 2.64665
R7800 VPWR.n2169 VPWR.n2168 2.64665
R7801 VPWR.n2113 VPWR.n2112 2.64665
R7802 VPWR.n1180 VPWR.n1118 2.64665
R7803 VPWR.n1184 VPWR.n1118 2.64665
R7804 VPWR.n1189 VPWR.n1116 2.64665
R7805 VPWR.n2335 VPWR.n7 2.64665
R7806 VPWR.n372 VPWR.n347 2.64665
R7807 VPWR.n335 VPWR.n334 2.64665
R7808 VPWR.n464 VPWR.n420 2.64665
R7809 VPWR.n2223 VPWR.n2222 2.63579
R7810 VPWR.n220 VPWR.n218 2.63539
R7811 VPWR.n223 VPWR.n221 2.63539
R7812 VPWR.n227 VPWR.n225 2.63539
R7813 VPWR.n232 VPWR.n230 2.63539
R7814 VPWR.n65 VPWR.n63 2.63539
R7815 VPWR.n115 VPWR.n113 2.63539
R7816 VPWR.n2058 VPWR.n2056 2.63539
R7817 VPWR.n2064 VPWR.n2062 2.63539
R7818 VPWR.n2067 VPWR.n2065 2.63539
R7819 VPWR.n2071 VPWR.n2069 2.63539
R7820 VPWR.n134 VPWR.n132 2.63539
R7821 VPWR.n2273 VPWR.n2271 2.63539
R7822 VPWR.n1137 VPWR.n1135 2.63539
R7823 VPWR.n1140 VPWR.n1138 2.63539
R7824 VPWR.n690 VPWR.n688 2.63539
R7825 VPWR.n693 VPWR.n691 2.63539
R7826 VPWR.n1378 VPWR.n1376 2.63539
R7827 VPWR.n1381 VPWR.n1379 2.63539
R7828 VPWR.n771 VPWR.n769 2.63539
R7829 VPWR.n774 VPWR.n772 2.63539
R7830 VPWR.n1006 VPWR.n1004 2.63539
R7831 VPWR.n1009 VPWR.n1007 2.63539
R7832 VPWR.n1031 VPWR.n1029 2.63539
R7833 VPWR.n1625 VPWR.n1623 2.63539
R7834 VPWR.n1900 VPWR.n1898 2.63539
R7835 VPWR.n1903 VPWR.n1901 2.63539
R7836 VPWR.n867 VPWR.n865 2.63539
R7837 VPWR.n973 VPWR.n971 2.63539
R7838 VPWR.n977 VPWR.n975 2.63539
R7839 VPWR.n886 VPWR.n884 2.63539
R7840 VPWR.n889 VPWR.n887 2.63539
R7841 VPWR.n2 VPWR.n0 2.63539
R7842 VPWR.n279 VPWR.n277 2.63539
R7843 VPWR.n282 VPWR.n280 2.63539
R7844 VPWR.n286 VPWR.n284 2.63539
R7845 VPWR.n291 VPWR.n289 2.63539
R7846 VPWR.n434 VPWR.n432 2.63539
R7847 VPWR.n440 VPWR.n438 2.63539
R7848 VPWR.n1320 VPWR.n1319 2.62345
R7849 VPWR.n2252 VPWR.n137 2.61352
R7850 VPWR.n1263 VPWR.n1260 2.56175
R7851 VPWR.n849 VPWR.n846 2.54018
R7852 VPWR.n1864 VPWR.n850 2.3878
R7853 VPWR.n871 VPWR.n870 2.37764
R7854 VPWR.n222 VPWR.n221 2.37495
R7855 VPWR.n219 VPWR.n218 2.37495
R7856 VPWR.n231 VPWR.n230 2.37495
R7857 VPWR.n226 VPWR.n225 2.37495
R7858 VPWR.n114 VPWR.n113 2.37495
R7859 VPWR.n64 VPWR.n63 2.37495
R7860 VPWR.n2063 VPWR.n2062 2.37495
R7861 VPWR.n2057 VPWR.n2056 2.37495
R7862 VPWR.n2070 VPWR.n2069 2.37495
R7863 VPWR.n2066 VPWR.n2065 2.37495
R7864 VPWR.n2272 VPWR.n2271 2.37495
R7865 VPWR.n133 VPWR.n132 2.37495
R7866 VPWR.n1139 VPWR.n1138 2.37495
R7867 VPWR.n1136 VPWR.n1135 2.37495
R7868 VPWR.n692 VPWR.n691 2.37495
R7869 VPWR.n689 VPWR.n688 2.37495
R7870 VPWR.n1380 VPWR.n1379 2.37495
R7871 VPWR.n1377 VPWR.n1376 2.37495
R7872 VPWR.n773 VPWR.n772 2.37495
R7873 VPWR.n770 VPWR.n769 2.37495
R7874 VPWR.n1008 VPWR.n1007 2.37495
R7875 VPWR.n1005 VPWR.n1004 2.37495
R7876 VPWR.n1030 VPWR.n1029 2.37495
R7877 VPWR.n1624 VPWR.n1623 2.37495
R7878 VPWR.n1902 VPWR.n1901 2.37495
R7879 VPWR.n1899 VPWR.n1898 2.37495
R7880 VPWR.n866 VPWR.n865 2.37495
R7881 VPWR.n976 VPWR.n975 2.37495
R7882 VPWR.n972 VPWR.n971 2.37495
R7883 VPWR.n888 VPWR.n887 2.37495
R7884 VPWR.n885 VPWR.n884 2.37495
R7885 VPWR.n1 VPWR.n0 2.37495
R7886 VPWR.n281 VPWR.n280 2.37495
R7887 VPWR.n278 VPWR.n277 2.37495
R7888 VPWR.n290 VPWR.n289 2.37495
R7889 VPWR.n285 VPWR.n284 2.37495
R7890 VPWR.n439 VPWR.n438 2.37495
R7891 VPWR.n433 VPWR.n432 2.37495
R7892 VPWR.n1232 VPWR.n1207 2.33701
R7893 VPWR.n1983 VPWR.n717 2.33701
R7894 VPWR.n1608 VPWR.n1607 2.33701
R7895 VPWR.n1712 VPWR.n1711 2.33701
R7896 VPWR.n2133 VPWR.n186 2.32777
R7897 VPWR.n337 VPWR.n3 2.32777
R7898 VPWR.n38 VPWR.n37 2.28432
R7899 VPWR.n1399 VPWR.n1373 2.28407
R7900 VPWR.n1399 VPWR.n1375 2.28407
R7901 VPWR.n1133 VPWR.n1131 2.28374
R7902 VPWR.n2179 VPWR.n168 2.27742
R7903 VPWR.n2246 VPWR.n143 2.25932
R7904 VPWR.n2224 VPWR.n2223 2.25932
R7905 VPWR.n1012 VPWR.n1003 2.25293
R7906 VPWR.n1871 VPWR.n1870 2.23542
R7907 VPWR.n1969 VPWR.n1968 2.22199
R7908 VPWR.n1866 VPWR.n849 2.13383
R7909 VPWR.n2028 VPWR.n2027 2.0932
R7910 VPWR.n1387 VPWR.n1386 2.07374
R7911 VPWR.n1374 VPWR.n1367 2.07374
R7912 VPWR.n1504 VPWR.n717 2.03225
R7913 VPWR.n1711 VPWR.n1710 2.03225
R7914 VPWR.n58 VPWR.n56 2.01703
R7915 VPWR.n61 VPWR.n59 2.01703
R7916 VPWR.n999 VPWR.n997 2.01703
R7917 VPWR.n1002 VPWR.n1000 2.01703
R7918 VPWR.n1873 VPWR.n1872 1.98145
R7919 VPWR.n851 VPWR.n850 1.98145
R7920 VPWR.n1222 VPWR.n1214 1.88902
R7921 VPWR.n1279 VPWR.n1263 1.88902
R7922 VPWR.n60 VPWR.n59 1.88416
R7923 VPWR.n57 VPWR.n56 1.88416
R7924 VPWR.n1001 VPWR.n1000 1.88416
R7925 VPWR.n998 VPWR.n997 1.88416
R7926 VPWR.n2104 VPWR.n2103 1.88325
R7927 VPWR.n631 VPWR.n245 1.88295
R7928 VPWR.n326 VPWR.n325 1.88295
R7929 VPWR.n1522 VPWR.n1492 1.88285
R7930 VPWR.n239 VPWR.n238 1.85065
R7931 VPWR.n653 VPWR.n240 1.85065
R7932 VPWR.n2146 VPWR.n2145 1.85065
R7933 VPWR.n2076 VPWR.n2053 1.85065
R7934 VPWR.n2078 VPWR.n206 1.85065
R7935 VPWR.n1157 VPWR.n1156 1.85065
R7936 VPWR.n1796 VPWR.n1795 1.85065
R7937 VPWR.n298 VPWR.n297 1.85065
R7938 VPWR.n300 VPWR.n265 1.85065
R7939 VPWR.n493 VPWR.n399 1.85065
R7940 VPWR.n1448 VPWR.n1350 1.82907
R7941 VPWR.n1606 VPWR.n1605 1.82907
R7942 VPWR.n1155 VPWR.n1154 1.81289
R7943 VPWR.n495 VPWR.n494 1.81289
R7944 VPWR.n2212 VPWR.n2211 1.73737
R7945 VPWR.n1246 VPWR.n1245 1.73737
R7946 VPWR.n2006 VPWR.n687 1.73737
R7947 VPWR.n1304 VPWR.n1095 1.69306
R7948 VPWR.n2010 VPWR.n684 1.69306
R7949 VPWR.n1617 VPWR.n712 1.69188
R7950 VPWR.n1600 VPWR.n712 1.69188
R7951 VPWR.n1989 VPWR.n711 1.69188
R7952 VPWR.n1989 VPWR.n1988 1.69188
R7953 VPWR.n1295 VPWR.n710 1.69188
R7954 VPWR.n1298 VPWR.n710 1.69188
R7955 VPWR.n2204 VPWR.n2203 1.69188
R7956 VPWR.n2203 VPWR.n2202 1.69188
R7957 VPWR.n2321 VPWR.n19 1.69188
R7958 VPWR.n2321 VPWR.n2320 1.69188
R7959 VPWR.n392 VPWR.n18 1.69188
R7960 VPWR.n379 VPWR.n18 1.69188
R7961 VPWR.n1539 VPWR.n1339 1.69188
R7962 VPWR.n1539 VPWR.n1538 1.69188
R7963 VPWR.n1337 VPWR.n1072 1.69188
R7964 VPWR.n1337 VPWR.n1336 1.69188
R7965 VPWR.n2163 VPWR.n2162 1.69188
R7966 VPWR.n2162 VPWR.n2161 1.69188
R7967 VPWR.n588 VPWR.n15 1.69188
R7968 VPWR.n591 VPWR.n15 1.69188
R7969 VPWR.n2326 VPWR.n14 1.69188
R7970 VPWR.n2327 VPWR.n2326 1.69188
R7971 VPWR.n1579 VPWR.n1540 1.69188
R7972 VPWR.n1699 VPWR.n992 1.69188
R7973 VPWR.n1699 VPWR.n1698 1.69188
R7974 VPWR.n1405 VPWR.n991 1.69188
R7975 VPWR.n1395 VPWR.n991 1.69188
R7976 VPWR.n1164 VPWR.n664 1.69188
R7977 VPWR.n1150 VPWR.n664 1.69188
R7978 VPWR.n2086 VPWR.n2085 1.69188
R7979 VPWR.n2085 VPWR.n2084 1.69188
R7980 VPWR.n660 VPWR.n211 1.69188
R7981 VPWR.n660 VPWR.n659 1.69188
R7982 VPWR.n308 VPWR.n307 1.69188
R7983 VPWR.n307 VPWR.n306 1.69188
R7984 VPWR.n1658 VPWR.n1657 1.69188
R7985 VPWR.n1659 VPWR.n1658 1.69188
R7986 VPWR.n1457 VPWR.n1038 1.69188
R7987 VPWR.n1440 VPWR.n1038 1.69188
R7988 VPWR.n1203 VPWR.n1202 1.69188
R7989 VPWR.n1202 VPWR.n1201 1.69188
R7990 VPWR.n2125 VPWR.n2124 1.69188
R7991 VPWR.n2124 VPWR.n2123 1.69188
R7992 VPWR.n619 VPWR.n618 1.69188
R7993 VPWR.n620 VPWR.n619 1.69188
R7994 VPWR.n522 VPWR.n251 1.69188
R7995 VPWR.n522 VPWR.n521 1.69188
R7996 VPWR.n1949 VPWR.n811 1.69188
R7997 VPWR.n1949 VPWR.n1948 1.69188
R7998 VPWR.n1950 VPWR.n810 1.69188
R7999 VPWR.n1951 VPWR.n1950 1.69188
R8000 VPWR.n2040 VPWR.n666 1.69188
R8001 VPWR.n2040 VPWR.n2039 1.69188
R8002 VPWR.n2242 VPWR.n49 1.69188
R8003 VPWR.n2229 VPWR.n49 1.69188
R8004 VPWR.n2287 VPWR.n48 1.69188
R8005 VPWR.n2288 VPWR.n2287 1.69188
R8006 VPWR.n476 VPWR.n475 1.69188
R8007 VPWR.n477 VPWR.n476 1.69188
R8008 VPWR.n1915 VPWR.n1890 1.69188
R8009 VPWR.n1905 VPWR.n1890 1.69188
R8010 VPWR.n786 VPWR.n708 1.69188
R8011 VPWR.n776 VPWR.n708 1.69188
R8012 VPWR.n1995 VPWR.n699 1.69188
R8013 VPWR.n1996 VPWR.n1995 1.69188
R8014 VPWR.n2282 VPWR.n125 1.69188
R8015 VPWR.n2282 VPWR.n2281 1.69188
R8016 VPWR.n124 VPWR.n51 1.69188
R8017 VPWR.n124 VPWR.n123 1.69188
R8018 VPWR.n451 VPWR.n448 1.69188
R8019 VPWR.n452 VPWR.n451 1.69188
R8020 VPWR.t107 VPWR 1.67895
R8021 VPWR.t235 VPWR 1.67895
R8022 VPWR.n1610 VPWR.n1609 1.67669
R8023 VPWR.n1157 VPWR.n1155 1.66186
R8024 VPWR.n494 VPWR.n493 1.66186
R8025 VPWR.n1759 VPWR.n1758 1.64857
R8026 VPWR.n654 VPWR.n239 1.6241
R8027 VPWR.n643 VPWR.n240 1.6241
R8028 VPWR.n2079 VPWR.n2076 1.6241
R8029 VPWR.n2090 VPWR.n206 1.6241
R8030 VPWR.n1156 VPWR.n1123 1.6241
R8031 VPWR.n1795 VPWR.n1794 1.6241
R8032 VPWR.n301 VPWR.n298 1.6241
R8033 VPWR.n312 VPWR.n265 1.6241
R8034 VPWR.n490 VPWR.n399 1.6241
R8035 VPWR.n628 VPWR.n245 1.62167
R8036 VPWR.n327 VPWR.n326 1.62167
R8037 VPWR.n2105 VPWR.n2104 1.62136
R8038 VPWR.n2211 VPWR.n2210 1.51082
R8039 VPWR.n1245 VPWR.n1244 1.51082
R8040 VPWR.n687 VPWR.n685 1.51082
R8041 VPWR.n1508 VPWR.n1500 1.4005
R8042 VPWR.n1417 VPWR.n1416 1.4005
R8043 VPWR.n2145 VPWR.n2144 1.39755
R8044 VPWR.n1087 VPWR.n1085 1.36443
R8045 VPWR.n2022 VPWR.n2021 1.36443
R8046 VPWR.n1505 VPWR.n1503 1.3232
R8047 VPWR.n2253 VPWR.n137 1.2502
R8048 VPWR.n1779 VPWR.n1778 1.11173
R8049 VPWR.n1709 VPWR.n958 1.08324
R8050 VPWR.n235 VPWR.n234 1.05773
R8051 VPWR.n2074 VPWR.n2055 1.05773
R8052 VPWR.n1803 VPWR.n1757 1.05773
R8053 VPWR.n294 VPWR.n293 1.05773
R8054 VPWR.n1309 VPWR.n1308 1.04968
R8055 VPWR.n2015 VPWR.n2014 1.04968
R8056 VPWR.n1386 VPWR.n1373 0.992049
R8057 VPWR.n1375 VPWR.n1367 0.992049
R8058 VPWR.n2135 VPWR.n185 0.899674
R8059 VPWR.n1232 VPWR.n1231 0.863992
R8060 VPWR.n1843 VPWR.n1842 0.853
R8061 VPWR.n1835 VPWR.n1834 0.853
R8062 VPWR.n1704 VPWR.n1703 0.853
R8063 VPWR.n1884 VPWR.n1883 0.853
R8064 VPWR.n1855 VPWR.n1854 0.853
R8065 VPWR.n897 VPWR.n832 0.853
R8066 VPWR.n1734 VPWR.n1733 0.813198
R8067 VPWR.n1818 VPWR.n1817 0.813198
R8068 VPWR.n97 VPWR.n96 0.753441
R8069 VPWR.n2294 VPWR.n42 0.740996
R8070 VPWR.n751 VPWR.n750 0.706789
R8071 VPWR.n923 VPWR.n921 0.65125
R8072 VPWR.n85 VPWR.n70 0.635211
R8073 VPWR.n1225 VPWR.n1211 0.635211
R8074 VPWR.n1290 VPWR.n1289 0.635211
R8075 VPWR.n1284 VPWR.n1283 0.635211
R8076 VPWR.n730 VPWR.n727 0.635211
R8077 VPWR.n750 VPWR.n746 0.635211
R8078 VPWR.n806 VPWR.n805 0.635211
R8079 VPWR.n755 VPWR.n753 0.635211
R8080 VPWR.n398 VPWR.n396 0.635211
R8081 VPWR.n417 VPWR.n413 0.635211
R8082 VPWR.n1314 VPWR.n1088 0.630008
R8083 VPWR.n2028 VPWR.n674 0.630008
R8084 VPWR.n2025 VPWR.n675 0.630008
R8085 VPWR.n1092 VPWR.n1090 0.52509
R8086 VPWR.n1109 VPWR.n1108 0.500125
R8087 VPWR.n210 VPWR.n16 0.500125
R8088 VPWR.n663 VPWR.n662 0.500125
R8089 VPWR.n2046 VPWR.n2045 0.500125
R8090 VPWR.n1701 VPWR.n1700 0.500125
R8091 VPWR.n1839 VPWR.n939 0.500125
R8092 VPWR.n1872 VPWR.n1871 0.457643
R8093 VPWR.n2043 VPWR.n159 0.3805
R8094 VPWR.n50 VPWR.n20 0.3805
R8095 VPWR.n2323 VPWR.n2322 0.3805
R8096 VPWR.n1991 VPWR.n1990 0.3805
R8097 VPWR.n1886 VPWR.n1885 0.3805
R8098 VPWR.n938 VPWR.n833 0.3805
R8099 VPWR.n2044 VPWR.n178 0.3805
R8100 VPWR.n661 VPWR.n177 0.3805
R8101 VPWR.n2325 VPWR.n2324 0.3805
R8102 VPWR.n1338 VPWR.n709 0.3805
R8103 VPWR.n1841 VPWR.n1840 0.3805
R8104 VPWR.n931 VPWR.n929 0.3805
R8105 VPWR.n1839 VPWR.n1838 0.3805
R8106 VPWR.n1700 VPWR.n940 0.3805
R8107 VPWR.n2045 VPWR.n194 0.3805
R8108 VPWR.n662 VPWR.n193 0.3805
R8109 VPWR.n523 VPWR.n16 0.3805
R8110 VPWR.n1110 VPWR.n1109 0.3805
R8111 VPWR.n1887 VPWR.n812 0.3805
R8112 VPWR.n2042 VPWR.n2041 0.3805
R8113 VPWR.n2286 VPWR.n2285 0.3805
R8114 VPWR.n47 VPWR.n17 0.3805
R8115 VPWR.n1992 VPWR.n667 0.3805
R8116 VPWR.n1852 VPWR.n1851 0.3805
R8117 VPWR.n1850 VPWR.n1849 0.3805
R8118 VPWR.n665 VPWR.n126 0.3805
R8119 VPWR.n2284 VPWR.n2283 0.3805
R8120 VPWR.n450 VPWR.n449 0.3805
R8121 VPWR.n1994 VPWR.n1993 0.3805
R8122 VPWR.n1889 VPWR.n1888 0.3805
R8123 VPWR.n637 VPWR.n243 0.369731
R8124 VPWR.n632 VPWR.n631 0.369731
R8125 VPWR.n628 VPWR.n627 0.369731
R8126 VPWR.n614 VPWR.n538 0.369731
R8127 VPWR.n601 VPWR.n542 0.369731
R8128 VPWR.n582 VPWR.n581 0.369731
R8129 VPWR.n576 VPWR.n561 0.369731
R8130 VPWR.n32 VPWR.n26 0.369731
R8131 VPWR.n2185 VPWR.n2184 0.369731
R8132 VPWR.n2193 VPWR.n2192 0.369731
R8133 VPWR.n2174 VPWR.n170 0.369731
R8134 VPWR.n2183 VPWR.n168 0.369731
R8135 VPWR.n2151 VPWR.n2150 0.369731
R8136 VPWR.n2173 VPWR.n171 0.369731
R8137 VPWR.n2106 VPWR.n2105 0.369731
R8138 VPWR.n2129 VPWR.n189 0.369731
R8139 VPWR.n2098 VPWR.n2097 0.369731
R8140 VPWR.n2103 VPWR.n202 0.369731
R8141 VPWR.n1175 VPWR.n1174 0.369731
R8142 VPWR.n1179 VPWR.n1119 0.369731
R8143 VPWR.n1181 VPWR.n1180 0.369731
R8144 VPWR.n1191 VPWR.n1103 0.369731
R8145 VPWR.n2342 VPWR.n2341 0.369731
R8146 VPWR.n363 VPWR.n350 0.369731
R8147 VPWR.n364 VPWR.n349 0.369731
R8148 VPWR.n385 VPWR.n338 0.369731
R8149 VPWR.n320 VPWR.n319 0.369731
R8150 VPWR.n325 VPWR.n261 0.369731
R8151 VPWR.n328 VPWR.n327 0.369731
R8152 VPWR.n509 VPWR.n508 0.369731
R8153 VPWR.n471 VPWR.n470 0.369731
R8154 VPWR.n431 VPWR.n423 0.369731
R8155 VPWR.n1257 VPWR.n1255 0.317855
R8156 VPWR.n1258 VPWR.n1257 0.317855
R8157 VPWR.n2260 VPWR.n131 0.305262
R8158 VPWR.n1227 VPWR.n1226 0.305262
R8159 VPWR.n1505 VPWR.n1504 0.305262
R8160 VPWR.n725 VPWR.n724 0.305262
R8161 VPWR.n1412 VPWR.n1411 0.305262
R8162 VPWR.n1605 VPWR.n1604 0.305262
R8163 VPWR.n1609 VPWR.n1046 0.305262
R8164 VPWR.n1926 VPWR.n826 0.305262
R8165 VPWR.n1897 VPWR.n1896 0.305262
R8166 VPWR.n1724 VPWR.n1723 0.305262
R8167 VPWR.n1729 VPWR.n1728 0.305262
R8168 VPWR.n1732 VPWR.n948 0.305262
R8169 VPWR.n1710 VPWR.n1709 0.305262
R8170 VPWR.n1716 VPWR.n956 0.305262
R8171 VPWR.n1824 VPWR.n1823 0.305262
R8172 VPWR.n1822 VPWR.n1746 0.305262
R8173 VPWR.n1813 VPWR.n1749 0.305262
R8174 VPWR.n1876 VPWR.n845 0.305262
R8175 VPWR.n1861 VPWR.n851 0.305262
R8176 VPWR.n921 VPWR.n862 0.305262
R8177 VPWR.n883 VPWR.n882 0.305262
R8178 VPWR.n1704 VPWR.n933 0.297373
R8179 VPWR.n897 VPWR.n857 0.294101
R8180 VPWR.n1422 VPWR.n1420 0.25148
R8181 VPWR.n1466 VPWR.n1348 0.246654
R8182 VPWR.n1012 VPWR 0.237784
R8183 VPWR.n106 VPWR.n104 0.231913
R8184 VPWR.n235 VPWR.n217 0.227049
R8185 VPWR.n638 VPWR.n242 0.227049
R8186 VPWR.n2210 VPWR.n2209 0.227049
R8187 VPWR.n2216 VPWR.n153 0.227049
R8188 VPWR.n2144 VPWR.n182 0.227049
R8189 VPWR.n2055 VPWR.n2054 0.227049
R8190 VPWR.n2092 VPWR.n204 0.227049
R8191 VPWR.n1147 VPWR.n1129 0.227049
R8192 VPWR.n1173 VPWR.n1121 0.227049
R8193 VPWR.n1244 VPWR.n1096 0.227049
R8194 VPWR.n1254 VPWR.n1253 0.227049
R8195 VPWR.n2009 VPWR.n685 0.227049
R8196 VPWR.n2004 VPWR.n2003 0.227049
R8197 VPWR.n796 VPWR.n757 0.227049
R8198 VPWR.n768 VPWR.n767 0.227049
R8199 VPWR.n1803 VPWR.n1802 0.227049
R8200 VPWR.n1791 VPWR.n1763 0.227049
R8201 VPWR.n294 VPWR.n276 0.227049
R8202 VPWR.n314 VPWR.n263 0.227049
R8203 VPWR.n497 VPWR.n496 0.227049
R8204 VPWR.n484 VPWR.n402 0.227049
R8205 VPWR VPWR.n2303 0.217591
R8206 VPWR.n2299 VPWR.n2298 0.21207
R8207 VPWR.n731 VPWR.n730 0.21207
R8208 VPWR.n804 VPWR.n803 0.21207
R8209 VPWR.n1837 VPWR 0.209323
R8210 VPWR VPWR.n1848 0.206051
R8211 VPWR.n1607 VPWR.n1606 0.203675
R8212 VPWR VPWR.n1012 0.200023
R8213 VPWR.n857 VPWR.n837 0.196829
R8214 VPWR.n1848 VPWR.n1847 0.196829
R8215 VPWR.n1844 VPWR.n933 0.195044
R8216 VPWR.n1837 VPWR.n932 0.195044
R8217 VPWR.n1426 VPWR.n1362 0.194439
R8218 VPWR.n2249 VPWR.n140 0.180304
R8219 VPWR.n1596 VPWR.n1055 0.180304
R8220 VPWR.n2132 VPWR 0.17983
R8221 VPWR.n2251 VPWR 0.17983
R8222 VPWR.n1398 VPWR 0.17983
R8223 VPWR VPWR.n2344 0.17983
R8224 VPWR.n229 VPWR 0.179485
R8225 VPWR.n104 VPWR 0.179485
R8226 VPWR VPWR.n2061 0.179485
R8227 VPWR.n2251 VPWR 0.179485
R8228 VPWR.n1622 VPWR 0.179485
R8229 VPWR.n288 VPWR 0.179485
R8230 VPWR VPWR.n228 0.172576
R8231 VPWR.n2068 VPWR 0.172576
R8232 VPWR VPWR.n1142 0.172576
R8233 VPWR VPWR.n1383 0.172576
R8234 VPWR VPWR.n1011 0.172576
R8235 VPWR.n974 VPWR 0.172576
R8236 VPWR VPWR.n287 0.172576
R8237 VPWR.n1989 VPWR.n712 0.1603
R8238 VPWR.n1579 VPWR.n1539 0.1603
R8239 VPWR.n1699 VPWR.n991 0.1603
R8240 VPWR.n1658 VPWR.n1038 0.1603
R8241 VPWR.n1950 VPWR.n1949 0.1603
R8242 VPWR.n1890 VPWR.n708 0.1603
R8243 VPWR.n541 VPWR 0.158169
R8244 VPWR VPWR.n579 0.158169
R8245 VPWR.n1767 VPWR 0.158169
R8246 VPWR.n905 VPWR 0.158169
R8247 VPWR.n1231 VPWR.n1208 0.152881
R8248 VPWR.n1885 VPWR.n1884 0.14385
R8249 VPWR.n1842 VPWR.n938 0.14385
R8250 VPWR.n1703 VPWR.n1701 0.14385
R8251 VPWR.n1835 VPWR.n940 0.14385
R8252 VPWR.n1854 VPWR.n812 0.14385
R8253 VPWR.n1889 VPWR.n832 0.14385
R8254 VPWR.n1398 VPWR.n1397 0.143027
R8255 VPWR.n1990 VPWR.n710 0.142675
R8256 VPWR.n1338 VPWR.n1337 0.142675
R8257 VPWR.n1108 VPWR.n664 0.142675
R8258 VPWR.n1202 VPWR.n1110 0.142675
R8259 VPWR.n2040 VPWR.n667 0.142675
R8260 VPWR.n1995 VPWR.n1994 0.142675
R8261 VPWR.n229 VPWR 0.14207
R8262 VPWR.n2061 VPWR 0.14207
R8263 VPWR VPWR.n1622 0.14207
R8264 VPWR.n288 VPWR 0.14207
R8265 VPWR.n2303 VPWR 0.141725
R8266 VPWR.n2132 VPWR 0.141725
R8267 VPWR.n2344 VPWR 0.141725
R8268 VPWR VPWR.n610 0.120408
R8269 VPWR.n1143 VPWR 0.120408
R8270 VPWR VPWR.n1783 0.120408
R8271 VPWR.n905 VPWR 0.120408
R8272 VPWR.n2322 VPWR.n2321 0.12035
R8273 VPWR.n2325 VPWR.n15 0.12035
R8274 VPWR.n660 VPWR.n210 0.12035
R8275 VPWR.n619 VPWR.n523 0.12035
R8276 VPWR.n2287 VPWR.n47 0.12035
R8277 VPWR.n450 VPWR.n124 0.12035
R8278 VPWR.n237 VPWR.n236 0.120292
R8279 VPWR.n644 VPWR.n241 0.120292
R8280 VPWR.n640 VPWR.n241 0.120292
R8281 VPWR.n640 VPWR.n639 0.120292
R8282 VPWR.n636 VPWR.n635 0.120292
R8283 VPWR.n635 VPWR.n244 0.120292
R8284 VPWR.n630 VPWR.n244 0.120292
R8285 VPWR.n629 VPWR.n246 0.120292
R8286 VPWR.n624 VPWR.n246 0.120292
R8287 VPWR.n624 VPWR.n623 0.120292
R8288 VPWR.n600 VPWR.n599 0.120292
R8289 VPWR.n599 VPWR.n543 0.120292
R8290 VPWR.n594 VPWR.n543 0.120292
R8291 VPWR.n585 VPWR.n551 0.120292
R8292 VPWR.n580 VPWR.n551 0.120292
R8293 VPWR.n575 VPWR.n574 0.120292
R8294 VPWR.n574 VPWR.n562 0.120292
R8295 VPWR.n569 VPWR.n562 0.120292
R8296 VPWR.n569 VPWR.n568 0.120292
R8297 VPWR.n568 VPWR.n565 0.120292
R8298 VPWR.n565 VPWR.n564 0.120292
R8299 VPWR.n2297 VPWR.n2296 0.120292
R8300 VPWR.n2296 VPWR.n2295 0.120292
R8301 VPWR.n2295 VPWR.n41 0.120292
R8302 VPWR.n2291 VPWR.n41 0.120292
R8303 VPWR.n88 VPWR.n87 0.120292
R8304 VPWR.n89 VPWR.n88 0.120292
R8305 VPWR.n89 VPWR.n67 0.120292
R8306 VPWR.n98 VPWR.n67 0.120292
R8307 VPWR.n99 VPWR.n98 0.120292
R8308 VPWR.n100 VPWR.n99 0.120292
R8309 VPWR.n2060 VPWR.n2059 0.120292
R8310 VPWR.n2089 VPWR.n205 0.120292
R8311 VPWR.n2094 VPWR.n205 0.120292
R8312 VPWR.n2095 VPWR.n2094 0.120292
R8313 VPWR.n2096 VPWR.n203 0.120292
R8314 VPWR.n2101 VPWR.n203 0.120292
R8315 VPWR.n2102 VPWR.n2101 0.120292
R8316 VPWR.n2108 VPWR.n201 0.120292
R8317 VPWR.n2109 VPWR.n2108 0.120292
R8318 VPWR.n2110 VPWR.n2109 0.120292
R8319 VPWR.n2141 VPWR.n2140 0.120292
R8320 VPWR.n2141 VPWR.n183 0.120292
R8321 VPWR.n2147 VPWR.n183 0.120292
R8322 VPWR.n2148 VPWR.n2147 0.120292
R8323 VPWR.n2171 VPWR.n172 0.120292
R8324 VPWR.n2172 VPWR.n2171 0.120292
R8325 VPWR.n2176 VPWR.n2175 0.120292
R8326 VPWR.n2176 VPWR.n169 0.120292
R8327 VPWR.n2181 VPWR.n169 0.120292
R8328 VPWR.n2182 VPWR.n2181 0.120292
R8329 VPWR.n2187 VPWR.n167 0.120292
R8330 VPWR.n2188 VPWR.n2187 0.120292
R8331 VPWR.n2189 VPWR.n2188 0.120292
R8332 VPWR.n2208 VPWR.n154 0.120292
R8333 VPWR.n2214 VPWR.n154 0.120292
R8334 VPWR.n2215 VPWR.n2214 0.120292
R8335 VPWR.n2220 VPWR.n2219 0.120292
R8336 VPWR.n2226 VPWR.n150 0.120292
R8337 VPWR.n2227 VPWR.n2226 0.120292
R8338 VPWR.n2256 VPWR.n135 0.120292
R8339 VPWR.n2262 VPWR.n135 0.120292
R8340 VPWR.n1153 VPWR.n1148 0.120292
R8341 VPWR.n1167 VPWR.n1122 0.120292
R8342 VPWR.n1171 VPWR.n1122 0.120292
R8343 VPWR.n1172 VPWR.n1171 0.120292
R8344 VPWR.n1177 VPWR.n1120 0.120292
R8345 VPWR.n1178 VPWR.n1177 0.120292
R8346 VPWR.n1183 VPWR.n1182 0.120292
R8347 VPWR.n1183 VPWR.n1117 0.120292
R8348 VPWR.n1187 VPWR.n1117 0.120292
R8349 VPWR.n1188 VPWR.n1187 0.120292
R8350 VPWR.n1229 VPWR.n1209 0.120292
R8351 VPWR.n1224 VPWR.n1223 0.120292
R8352 VPWR.n1223 VPWR.n1212 0.120292
R8353 VPWR.n1218 VPWR.n1212 0.120292
R8354 VPWR.n1322 VPWR.n1083 0.120292
R8355 VPWR.n1317 VPWR.n1083 0.120292
R8356 VPWR.n1317 VPWR.n1316 0.120292
R8357 VPWR.n1316 VPWR.n1315 0.120292
R8358 VPWR.n1312 VPWR.n1311 0.120292
R8359 VPWR.n1311 VPWR.n1091 0.120292
R8360 VPWR.n1306 VPWR.n1091 0.120292
R8361 VPWR.n1306 VPWR.n1305 0.120292
R8362 VPWR.n1286 VPWR.n1256 0.120292
R8363 VPWR.n1281 VPWR.n1256 0.120292
R8364 VPWR.n1281 VPWR.n1280 0.120292
R8365 VPWR.n1280 VPWR.n1261 0.120292
R8366 VPWR.n1275 VPWR.n1261 0.120292
R8367 VPWR.n1275 VPWR.n1274 0.120292
R8368 VPWR.n1274 VPWR.n1273 0.120292
R8369 VPWR.n2024 VPWR.n2023 0.120292
R8370 VPWR.n2023 VPWR.n677 0.120292
R8371 VPWR.n2018 VPWR.n677 0.120292
R8372 VPWR.n2018 VPWR.n2017 0.120292
R8373 VPWR.n2017 VPWR.n681 0.120292
R8374 VPWR.n2012 VPWR.n681 0.120292
R8375 VPWR.n2012 VPWR.n2011 0.120292
R8376 VPWR.n2008 VPWR.n2007 0.120292
R8377 VPWR.n2007 VPWR.n686 0.120292
R8378 VPWR.n1413 VPWR.n1365 0.120292
R8379 VPWR.n1415 VPWR.n1414 0.120292
R8380 VPWR.n1415 VPWR.n1363 0.120292
R8381 VPWR.n1424 VPWR.n1363 0.120292
R8382 VPWR.n1427 VPWR.n1424 0.120292
R8383 VPWR.n1428 VPWR.n1427 0.120292
R8384 VPWR.n1437 VPWR.n1360 0.120292
R8385 VPWR.n1438 VPWR.n1437 0.120292
R8386 VPWR.n1469 VPWR.n1468 0.120292
R8387 VPWR.n1476 VPWR.n1475 0.120292
R8388 VPWR.n1483 VPWR.n1482 0.120292
R8389 VPWR.n1524 VPWR.n1523 0.120292
R8390 VPWR.n1519 VPWR.n1518 0.120292
R8391 VPWR.n1518 VPWR.n1495 0.120292
R8392 VPWR.n1496 VPWR.n1495 0.120292
R8393 VPWR.n1512 VPWR.n1496 0.120292
R8394 VPWR.n1512 VPWR.n1511 0.120292
R8395 VPWR.n1972 VPWR.n1971 0.120292
R8396 VPWR.n1971 VPWR.n728 0.120292
R8397 VPWR.n1966 VPWR.n728 0.120292
R8398 VPWR.n1966 VPWR.n1965 0.120292
R8399 VPWR.n1965 VPWR.n733 0.120292
R8400 VPWR.n1961 VPWR.n733 0.120292
R8401 VPWR.n1961 VPWR.n1960 0.120292
R8402 VPWR.n1960 VPWR.n736 0.120292
R8403 VPWR.n807 VPWR.n745 0.120292
R8404 VPWR.n801 VPWR.n745 0.120292
R8405 VPWR.n800 VPWR.n799 0.120292
R8406 VPWR.n799 VPWR.n754 0.120292
R8407 VPWR.n795 VPWR.n794 0.120292
R8408 VPWR.n794 VPWR.n758 0.120292
R8409 VPWR.n790 VPWR.n758 0.120292
R8410 VPWR.n790 VPWR.n789 0.120292
R8411 VPWR.n1682 VPWR.n1681 0.120292
R8412 VPWR.n1681 VPWR.n1018 0.120292
R8413 VPWR.n1677 VPWR.n1018 0.120292
R8414 VPWR.n1677 VPWR.n1676 0.120292
R8415 VPWR.n1676 VPWR.n1675 0.120292
R8416 VPWR.n1675 VPWR.n1020 0.120292
R8417 VPWR.n1671 VPWR.n1020 0.120292
R8418 VPWR.n1671 VPWR.n1670 0.120292
R8419 VPWR.n1670 VPWR.n1669 0.120292
R8420 VPWR.n1669 VPWR.n1025 0.120292
R8421 VPWR.n1027 VPWR.n1025 0.120292
R8422 VPWR.n1555 VPWR.n1550 0.120292
R8423 VPWR.n1556 VPWR.n1555 0.120292
R8424 VPWR.n1557 VPWR.n1556 0.120292
R8425 VPWR.n1557 VPWR.n1547 0.120292
R8426 VPWR.n1563 VPWR.n1547 0.120292
R8427 VPWR.n1564 VPWR.n1563 0.120292
R8428 VPWR.n1565 VPWR.n1564 0.120292
R8429 VPWR.n1565 VPWR.n1544 0.120292
R8430 VPWR.n1064 VPWR.n1061 0.120292
R8431 VPWR.n1588 VPWR.n1061 0.120292
R8432 VPWR.n1590 VPWR.n1058 0.120292
R8433 VPWR.n1058 VPWR.n1055 0.120292
R8434 VPWR.n1645 VPWR.n1644 0.120292
R8435 VPWR.n1644 VPWR.n1643 0.120292
R8436 VPWR.n1639 VPWR.n1629 0.120292
R8437 VPWR.n1639 VPWR.n1638 0.120292
R8438 VPWR.n1638 VPWR.n1632 0.120292
R8439 VPWR.n1935 VPWR.n1934 0.120292
R8440 VPWR.n1934 VPWR.n823 0.120292
R8441 VPWR.n1930 VPWR.n823 0.120292
R8442 VPWR.n1930 VPWR.n1929 0.120292
R8443 VPWR.n1929 VPWR.n1928 0.120292
R8444 VPWR.n1925 VPWR.n1924 0.120292
R8445 VPWR.n1924 VPWR.n827 0.120292
R8446 VPWR.n981 VPWR.n969 0.120292
R8447 VPWR.n983 VPWR.n966 0.120292
R8448 VPWR.n1714 VPWR.n957 0.120292
R8449 VPWR.n1720 VPWR.n1719 0.120292
R8450 VPWR.n1726 VPWR.n1725 0.120292
R8451 VPWR.n1735 VPWR.n949 0.120292
R8452 VPWR.n1820 VPWR.n1747 0.120292
R8453 VPWR.n1815 VPWR.n1747 0.120292
R8454 VPWR.n1815 VPWR.n1814 0.120292
R8455 VPWR.n1798 VPWR.n1762 0.120292
R8456 VPWR.n1793 VPWR.n1762 0.120292
R8457 VPWR.n1793 VPWR.n1792 0.120292
R8458 VPWR.n1788 VPWR.n1787 0.120292
R8459 VPWR.n1869 VPWR.n1868 0.120292
R8460 VPWR.n1868 VPWR.n1867 0.120292
R8461 VPWR.n1867 VPWR.n847 0.120292
R8462 VPWR.n1863 VPWR.n1862 0.120292
R8463 VPWR.n915 VPWR.n914 0.120292
R8464 VPWR.n914 VPWR.n913 0.120292
R8465 VPWR.n296 VPWR.n295 0.120292
R8466 VPWR.n311 VPWR.n264 0.120292
R8467 VPWR.n316 VPWR.n264 0.120292
R8468 VPWR.n317 VPWR.n316 0.120292
R8469 VPWR.n318 VPWR.n262 0.120292
R8470 VPWR.n323 VPWR.n262 0.120292
R8471 VPWR.n324 VPWR.n323 0.120292
R8472 VPWR.n330 VPWR.n260 0.120292
R8473 VPWR.n331 VPWR.n330 0.120292
R8474 VPWR.n332 VPWR.n331 0.120292
R8475 VPWR.n2343 VPWR.n4 0.120292
R8476 VPWR.n2338 VPWR.n4 0.120292
R8477 VPWR.n2338 VPWR.n2337 0.120292
R8478 VPWR.n2337 VPWR.n2336 0.120292
R8479 VPWR.n2336 VPWR.n6 0.120292
R8480 VPWR.n362 VPWR.n351 0.120292
R8481 VPWR VPWR.n362 0.120292
R8482 VPWR.n366 VPWR.n365 0.120292
R8483 VPWR.n366 VPWR.n348 0.120292
R8484 VPWR.n370 VPWR.n348 0.120292
R8485 VPWR.n371 VPWR.n370 0.120292
R8486 VPWR.n371 VPWR.n346 0.120292
R8487 VPWR.n375 VPWR.n346 0.120292
R8488 VPWR.n376 VPWR.n375 0.120292
R8489 VPWR.n382 VPWR.n376 0.120292
R8490 VPWR.n498 VPWR.n397 0.120292
R8491 VPWR.n492 VPWR.n397 0.120292
R8492 VPWR.n492 VPWR.n491 0.120292
R8493 VPWR.n491 VPWR.n400 0.120292
R8494 VPWR.n487 VPWR.n400 0.120292
R8495 VPWR.n487 VPWR.n486 0.120292
R8496 VPWR.n486 VPWR.n485 0.120292
R8497 VPWR.n472 VPWR.n412 0.120292
R8498 VPWR.n467 VPWR.n412 0.120292
R8499 VPWR.n467 VPWR.n466 0.120292
R8500 VPWR.n466 VPWR.n465 0.120292
R8501 VPWR.n465 VPWR.n419 0.120292
R8502 VPWR.n461 VPWR.n419 0.120292
R8503 VPWR.n461 VPWR.n460 0.120292
R8504 VPWR.n460 VPWR.n459 0.120292
R8505 VPWR.n459 VPWR.n422 0.120292
R8506 VPWR.n455 VPWR.n422 0.120292
R8507 VPWR.n1109 VPWR.n709 0.120125
R8508 VPWR.n1991 VPWR.n709 0.120125
R8509 VPWR.n1992 VPWR.n1991 0.120125
R8510 VPWR.n1993 VPWR.n1992 0.120125
R8511 VPWR.n2324 VPWR.n16 0.120125
R8512 VPWR.n2324 VPWR.n2323 0.120125
R8513 VPWR.n2323 VPWR.n17 0.120125
R8514 VPWR.n449 VPWR.n17 0.120125
R8515 VPWR.n662 VPWR.n661 0.120125
R8516 VPWR.n661 VPWR.n50 0.120125
R8517 VPWR.n2285 VPWR.n50 0.120125
R8518 VPWR.n2285 VPWR.n2284 0.120125
R8519 VPWR.n2045 VPWR.n2044 0.120125
R8520 VPWR.n2044 VPWR.n2043 0.120125
R8521 VPWR.n2043 VPWR.n2042 0.120125
R8522 VPWR.n2042 VPWR.n665 0.120125
R8523 VPWR.n1700 VPWR.n833 0.120125
R8524 VPWR.n1886 VPWR.n833 0.120125
R8525 VPWR.n1887 VPWR.n1886 0.120125
R8526 VPWR.n1888 VPWR.n1887 0.120125
R8527 VPWR.n1840 VPWR.n1839 0.120125
R8528 VPWR.n1840 VPWR.n929 0.120125
R8529 VPWR.n1851 VPWR.n929 0.120125
R8530 VPWR.n1851 VPWR.n1850 0.120125
R8531 VPWR.n2139 VPWR.n2138 0.113774
R8532 VPWR.n2138 VPWR.n184 0.113774
R8533 VPWR.n695 VPWR.n686 0.112479
R8534 VPWR.n789 VPWR.n788 0.112479
R8535 VPWR.n1918 VPWR.n1917 0.112479
R8536 VPWR.n900 VPWR.n899 0.112479
R8537 VPWR.n455 VPWR.n454 0.112479
R8538 VPWR.n2203 VPWR.n159 0.1086
R8539 VPWR.n2162 VPWR.n178 0.1086
R8540 VPWR.n2085 VPWR.n2046 0.1086
R8541 VPWR.n2124 VPWR.n194 0.1086
R8542 VPWR.n2041 VPWR.n49 0.1086
R8543 VPWR.n2282 VPWR.n126 0.1086
R8544 VPWR.n594 VPWR.n593 0.107271
R8545 VPWR.n2149 VPWR.n180 0.107271
R8546 VPWR.n1218 VPWR.n1074 0.107271
R8547 VPWR.n1483 VPWR.n1341 0.107271
R8548 VPWR.n1544 VPWR.n1542 0.107271
R8549 VPWR.n9 VPWR.n6 0.107271
R8550 VPWR.n1845 VPWR.n1844 0.10625
R8551 VPWR.n1846 VPWR.n932 0.10625
R8552 VPWR.n1313 VPWR.n1090 0.105418
R8553 VPWR.n2019 VPWR.n680 0.105418
R8554 VPWR.n228 VPWR 0.105238
R8555 VPWR.n2068 VPWR 0.105238
R8556 VPWR.n1142 VPWR 0.105238
R8557 VPWR.n1383 VPWR 0.105238
R8558 VPWR.n1011 VPWR 0.105238
R8559 VPWR.n974 VPWR 0.105238
R8560 VPWR.n287 VPWR 0.105238
R8561 VPWR.n2259 VPWR.n2258 0.102087
R8562 VPWR.n1982 VPWR.n719 0.102087
R8563 VPWR.n1923 VPWR.n1922 0.102087
R8564 VPWR VPWR.n629 0.0981562
R8565 VPWR.n612 VPWR 0.0981562
R8566 VPWR.n575 VPWR 0.0981562
R8567 VPWR VPWR.n2308 0.0981562
R8568 VPWR.n2297 VPWR 0.0981562
R8569 VPWR VPWR.n201 0.0981562
R8570 VPWR.n2131 VPWR 0.0981562
R8571 VPWR.n2140 VPWR 0.0981562
R8572 VPWR.n2175 VPWR 0.0981562
R8573 VPWR VPWR.n167 0.0981562
R8574 VPWR.n2207 VPWR 0.0981562
R8575 VPWR.n2219 VPWR 0.0981562
R8576 VPWR.n2256 VPWR 0.0981562
R8577 VPWR.n1182 VPWR 0.0981562
R8578 VPWR.n1240 VPWR 0.0981562
R8579 VPWR.n1230 VPWR 0.0981562
R8580 VPWR VPWR.n1229 0.0981562
R8581 VPWR.n1312 VPWR 0.0981562
R8582 VPWR VPWR.n1286 0.0981562
R8583 VPWR VPWR.n1365 0.0981562
R8584 VPWR.n1475 VPWR 0.0981562
R8585 VPWR VPWR.n1519 0.0981562
R8586 VPWR VPWR.n1064 0.0981562
R8587 VPWR.n1719 VPWR 0.0981562
R8588 VPWR VPWR.n949 0.0981562
R8589 VPWR VPWR.n1820 0.0981562
R8590 VPWR.n1752 VPWR 0.0981562
R8591 VPWR VPWR.n1788 0.0981562
R8592 VPWR.n1869 VPWR 0.0981562
R8593 VPWR VPWR.n1858 0.0981562
R8594 VPWR VPWR.n900 0.0981562
R8595 VPWR VPWR.n260 0.0981562
R8596 VPWR VPWR.n506 0.0981562
R8597 VPWR.n365 VPWR 0.0981562
R8598 VPWR.n395 VPWR 0.0981562
R8599 VPWR.n1844 VPWR.n1843 0.0977722
R8600 VPWR.n1834 VPWR.n933 0.0977722
R8601 VPWR.n1883 VPWR.n837 0.0977722
R8602 VPWR.n1855 VPWR.n857 0.0977722
R8603 VPWR.n1482 VPWR 0.0968542
R8604 VPWR VPWR.n1918 0.0968542
R8605 VPWR.n480 VPWR.n407 0.0950946
R8606 VPWR.n474 VPWR.n411 0.0950946
R8607 VPWR.n1856 VPWR.n855 0.0950946
R8608 VPWR.n863 VPWR.n858 0.0950946
R8609 VPWR.n520 VPWR.n519 0.0950946
R8610 VPWR.n513 VPWR.n257 0.0950946
R8611 VPWR.n305 VPWR.n304 0.0950946
R8612 VPWR.n309 VPWR.n267 0.0950946
R8613 VPWR.n1947 VPWR.n1946 0.0950946
R8614 VPWR.n1940 VPWR.n818 0.0950946
R8615 VPWR.n2330 VPWR.n11 0.0950946
R8616 VPWR.n356 VPWR.n355 0.0950946
R8617 VPWR.n380 VPWR.n378 0.0950946
R8618 VPWR.n393 VPWR.n340 0.0950946
R8619 VPWR.n2289 VPWR.n45 0.0950946
R8620 VPWR.n82 VPWR.n81 0.0950946
R8621 VPWR.n592 VPWR.n546 0.0950946
R8622 VPWR.n587 VPWR.n549 0.0950946
R8623 VPWR.n621 VPWR.n249 0.0950946
R8624 VPWR.n617 VPWR.n525 0.0950946
R8625 VPWR.n658 VPWR.n657 0.0950946
R8626 VPWR.n650 VPWR.n649 0.0950946
R8627 VPWR.n109 VPWR.n107 0.0950946
R8628 VPWR.n120 VPWR.n52 0.0950946
R8629 VPWR.n2319 VPWR.n2318 0.0950946
R8630 VPWR.n2311 VPWR.n2310 0.0950946
R8631 VPWR.n2231 VPWR.n2230 0.0950946
R8632 VPWR.n2243 VPWR.n145 0.0950946
R8633 VPWR.n2160 VPWR.n2159 0.0950946
R8634 VPWR.n2164 VPWR.n175 0.0950946
R8635 VPWR.n2122 VPWR.n2121 0.0950946
R8636 VPWR.n2126 VPWR.n191 0.0950946
R8637 VPWR.n2083 VPWR.n2082 0.0950946
R8638 VPWR.n2087 VPWR.n208 0.0950946
R8639 VPWR.n2267 VPWR.n2265 0.0950946
R8640 VPWR.n2278 VPWR.n127 0.0950946
R8641 VPWR.n2201 VPWR.n2200 0.0950946
R8642 VPWR.n2205 VPWR.n157 0.0950946
R8643 VPWR.n2038 VPWR.n2037 0.0950946
R8644 VPWR.n2031 VPWR.n673 0.0950946
R8645 VPWR.n1335 VPWR.n1334 0.0950946
R8646 VPWR.n1327 VPWR.n1326 0.0950946
R8647 VPWR.n1200 VPWR.n1199 0.0950946
R8648 VPWR.n1204 VPWR.n1106 0.0950946
R8649 VPWR.n1151 VPWR.n1149 0.0950946
R8650 VPWR.n1165 VPWR.n1125 0.0950946
R8651 VPWR.n2000 VPWR.n697 0.0950946
R8652 VPWR.n707 VPWR.n701 0.0950946
R8653 VPWR.n1299 VPWR.n1098 0.0950946
R8654 VPWR.n1294 VPWR.n1101 0.0950946
R8655 VPWR.n1954 VPWR.n740 0.0950946
R8656 VPWR.n809 VPWR.n744 0.0950946
R8657 VPWR.n1537 VPWR.n1536 0.0950946
R8658 VPWR.n1529 VPWR.n1528 0.0950946
R8659 VPWR.n1441 VPWR.n1439 0.0950946
R8660 VPWR.n1458 VPWR.n1352 0.0950946
R8661 VPWR.n1396 VPWR.n1394 0.0950946
R8662 VPWR.n1406 VPWR.n1368 0.0950946
R8663 VPWR.n787 VPWR.n761 0.0950946
R8664 VPWR.n777 VPWR.n775 0.0950946
R8665 VPWR.n1987 VPWR.n1986 0.0950946
R8666 VPWR.n1979 VPWR.n1978 0.0950946
R8667 VPWR.n1601 VPWR.n1599 0.0950946
R8668 VPWR.n1618 VPWR.n1048 0.0950946
R8669 VPWR.n1805 VPWR.n935 0.0950946
R8670 VPWR.n1760 VPWR.n936 0.0950946
R8671 VPWR.n1577 VPWR.n1576 0.0950946
R8672 VPWR.n1581 VPWR.n1070 0.0950946
R8673 VPWR.n1662 VPWR.n1035 0.0950946
R8674 VPWR.n1656 VPWR.n1040 0.0950946
R8675 VPWR.n1916 VPWR.n831 0.0950946
R8676 VPWR.n1906 VPWR.n1904 0.0950946
R8677 VPWR.n1697 VPWR.n1696 0.0950946
R8678 VPWR.n1688 VPWR.n1687 0.0950946
R8679 VPWR.n1738 VPWR.n943 0.0950946
R8680 VPWR.n1832 VPWR.n942 0.0950946
R8681 VPWR.n990 VPWR.n989 0.0950946
R8682 VPWR.n1706 VPWR.n1705 0.0950946
R8683 VPWR.n898 VPWR.n875 0.0950946
R8684 VPWR.n880 VPWR.n876 0.0950946
R8685 VPWR.n1772 VPWR.n838 0.0950946
R8686 VPWR.n1881 VPWR.n836 0.0950946
R8687 VPWR.n453 VPWR.n425 0.0950946
R8688 VPWR.n445 VPWR.n427 0.0950946
R8689 VPWR VPWR.n1143 0.0930646
R8690 VPWR.n1845 VPWR.n837 0.0913766
R8691 VPWR.n1847 VPWR.n1846 0.0913766
R8692 VPWR.n2203 VPWR.n20 0.086275
R8693 VPWR.n2162 VPWR.n177 0.086275
R8694 VPWR.n2085 VPWR.n663 0.086275
R8695 VPWR.n2124 VPWR.n193 0.086275
R8696 VPWR.n2286 VPWR.n49 0.086275
R8697 VPWR.n2283 VPWR.n2282 0.086275
R8698 VPWR.n656 VPWR.n213 0.0838333
R8699 VPWR.n651 VPWR.n645 0.0838333
R8700 VPWR.n533 VPWR.n529 0.0838333
R8701 VPWR.n556 VPWR.n554 0.0838333
R8702 VPWR.n2317 VPWR.n22 0.0838333
R8703 VPWR.n77 VPWR.n76 0.0838333
R8704 VPWR.n119 VPWR.n118 0.0838333
R8705 VPWR.n2081 VPWR.n2048 0.0838333
R8706 VPWR.n2088 VPWR.n207 0.0838333
R8707 VPWR.n2120 VPWR.n2119 0.0838333
R8708 VPWR.n2156 VPWR.n174 0.0838333
R8709 VPWR.n2199 VPWR.n161 0.0838333
R8710 VPWR.n2277 VPWR.n2276 0.0838333
R8711 VPWR.n1152 VPWR.n1128 0.0838333
R8712 VPWR.n1166 VPWR.n1124 0.0838333
R8713 VPWR.n1198 VPWR.n1197 0.0838333
R8714 VPWR.n1082 VPWR.n1077 0.0838333
R8715 VPWR.n1300 VPWR.n1097 0.0838333
R8716 VPWR.n2036 VPWR.n2035 0.0838333
R8717 VPWR.n706 VPWR.n704 0.0838333
R8718 VPWR.n1397 VPWR.n1393 0.0838333
R8719 VPWR.n1453 VPWR.n1355 0.0838333
R8720 VPWR.n1489 VPWR.n1344 0.0838333
R8721 VPWR.n1985 VPWR.n714 0.0838333
R8722 VPWR.n1955 VPWR.n739 0.0838333
R8723 VPWR.n778 VPWR.n766 0.0838333
R8724 VPWR.n1695 VPWR.n994 0.0838333
R8725 VPWR.n1689 VPWR.n1683 0.0838333
R8726 VPWR.n1573 VPWR.n1069 0.0838333
R8727 VPWR.n1602 VPWR.n1598 0.0838333
R8728 VPWR.n1945 VPWR.n1944 0.0838333
R8729 VPWR.n1907 VPWR.n1895 0.0838333
R8730 VPWR.n988 VPWR.n964 0.0838333
R8731 VPWR.n1707 VPWR.n960 0.0838333
R8732 VPWR.n1761 VPWR.n1756 0.0838333
R8733 VPWR.n890 VPWR.n881 0.0838333
R8734 VPWR.n303 VPWR.n270 0.0838333
R8735 VPWR.n310 VPWR.n266 0.0838333
R8736 VPWR.n518 VPWR.n517 0.0838333
R8737 VPWR.n353 VPWR.n352 0.0838333
R8738 VPWR.n381 VPWR.n377 0.0838333
R8739 VPWR.n481 VPWR.n406 0.0838333
R8740 VPWR.n444 VPWR.n443 0.0838333
R8741 VPWR.n834 VPWR 0.08275
R8742 VPWR.n1702 VPWR 0.08275
R8743 VPWR.n1836 VPWR 0.08275
R8744 VPWR.n1853 VPWR 0.08275
R8745 VPWR.n930 VPWR 0.08275
R8746 VPWR VPWR.n2249 0.082648
R8747 VPWR VPWR.n1596 0.082648
R8748 VPWR.n610 VPWR 0.082648
R8749 VPWR VPWR.n541 0.082648
R8750 VPWR.n579 VPWR 0.082648
R8751 VPWR.n1783 VPWR 0.082648
R8752 VPWR VPWR.n1767 0.082648
R8753 VPWR.n616 VPWR.n615 0.0812292
R8754 VPWR.n586 VPWR.n550 0.0812292
R8755 VPWR.n2312 VPWR.n27 0.0812292
R8756 VPWR.n83 VPWR.n74 0.0812292
R8757 VPWR.n111 VPWR.n55 0.0812292
R8758 VPWR.n2128 VPWR.n2127 0.0812292
R8759 VPWR.n2166 VPWR.n2165 0.0812292
R8760 VPWR.n2194 VPWR.n156 0.0812292
R8761 VPWR.n2237 VPWR.n144 0.0812292
R8762 VPWR.n2269 VPWR.n130 0.0812292
R8763 VPWR.n1206 VPWR.n1205 0.0812292
R8764 VPWR.n1329 VPWR.n1328 0.0812292
R8765 VPWR.n1250 VPWR.n1102 0.0812292
R8766 VPWR.n2030 VPWR.n672 0.0812292
R8767 VPWR.n703 VPWR.n702 0.0812292
R8768 VPWR.n1460 VPWR.n1459 0.0812292
R8769 VPWR.n1531 VPWR.n1530 0.0812292
R8770 VPWR.n1980 VPWR.n720 0.0812292
R8771 VPWR.n748 VPWR.n747 0.0812292
R8772 VPWR.n782 VPWR.n781 0.0812292
R8773 VPWR.n1655 VPWR.n1654 0.0812292
R8774 VPWR.n1052 VPWR.n1047 0.0812292
R8775 VPWR.n1939 VPWR.n817 0.0812292
R8776 VPWR.n1911 VPWR.n1910 0.0812292
R8777 VPWR.n1827 VPWR.n945 0.0812292
R8778 VPWR.n1800 VPWR.n1799 0.0812292
R8779 VPWR.n1880 VPWR.n1879 0.0812292
R8780 VPWR.n894 VPWR.n893 0.0812292
R8781 VPWR.n507 VPWR.n258 0.0812292
R8782 VPWR.n358 VPWR.n357 0.0812292
R8783 VPWR.n344 VPWR.n339 0.0812292
R8784 VPWR.n415 VPWR.n414 0.0812292
R8785 VPWR.n436 VPWR.n430 0.0812292
R8786 VPWR.n535 VPWR.n534 0.0760208
R8787 VPWR.n2316 VPWR.n24 0.0760208
R8788 VPWR.n87 VPWR.n69 0.0760208
R8789 VPWR.n2116 VPWR.n199 0.0760208
R8790 VPWR.n2198 VPWR.n165 0.0760208
R8791 VPWR.n2244 VPWR.n140 0.0760208
R8792 VPWR.n1194 VPWR.n1115 0.0760208
R8793 VPWR.n1249 VPWR.n1247 0.0760208
R8794 VPWR.n2024 VPWR.n676 0.0760208
R8795 VPWR.n1452 VPWR.n1356 0.0760208
R8796 VPWR.n1984 VPWR.n716 0.0760208
R8797 VPWR.n808 VPWR.n807 0.0760208
R8798 VPWR.n1043 VPWR.n1042 0.0760208
R8799 VPWR.n1613 VPWR.n1051 0.0760208
R8800 VPWR.n1935 VPWR.n819 0.0760208
R8801 VPWR.n919 VPWR.n918 0.0760208
R8802 VPWR.n512 VPWR.n256 0.0760208
R8803 VPWR.n388 VPWR.n343 0.0760208
R8804 VPWR.n2321 VPWR.n20 0.074525
R8805 VPWR.n177 VPWR.n15 0.074525
R8806 VPWR.n663 VPWR.n660 0.074525
R8807 VPWR.n619 VPWR.n193 0.074525
R8808 VPWR.n2287 VPWR.n2286 0.074525
R8809 VPWR.n2283 VPWR.n124 0.074525
R8810 VPWR.n655 VPWR.n215 0.0708125
R8811 VPWR.n553 VPWR.n545 0.0708125
R8812 VPWR.n2291 VPWR.n2290 0.0708125
R8813 VPWR.n2080 VPWR.n2052 0.0708125
R8814 VPWR.n2158 VPWR.n2153 0.0708125
R8815 VPWR.n2228 VPWR.n2227 0.0708125
R8816 VPWR.n1160 VPWR.n1158 0.0708125
R8817 VPWR.n1333 VPWR.n1076 0.0708125
R8818 VPWR.n1273 VPWR.n669 0.0708125
R8819 VPWR.n1401 VPWR.n1371 0.0708125
R8820 VPWR.n1535 VPWR.n1343 0.0708125
R8821 VPWR.n738 VPWR.n736 0.0708125
R8822 VPWR.n1694 VPWR.n996 0.0708125
R8823 VPWR.n1575 VPWR.n1570 0.0708125
R8824 VPWR.n1632 VPWR.n814 0.0708125
R8825 VPWR.n1858 VPWR.n1857 0.0708125
R8826 VPWR.n302 VPWR.n274 0.0708125
R8827 VPWR.n2332 VPWR.n2331 0.0708125
R8828 VPWR.n479 VPWR.n408 0.0680676
R8829 VPWR.n410 VPWR.n408 0.0680676
R8830 VPWR.n928 VPWR.n927 0.0680676
R8831 VPWR.n927 VPWR.n856 0.0680676
R8832 VPWR.n516 VPWR.n254 0.0680676
R8833 VPWR.n516 VPWR.n515 0.0680676
R8834 VPWR.n273 VPWR.n271 0.0680676
R8835 VPWR.n273 VPWR.n272 0.0680676
R8836 VPWR.n1943 VPWR.n815 0.0680676
R8837 VPWR.n1943 VPWR.n1942 0.0680676
R8838 VPWR.n2329 VPWR.n12 0.0680676
R8839 VPWR.n354 VPWR.n12 0.0680676
R8840 VPWR.n389 VPWR.n342 0.0680676
R8841 VPWR.n390 VPWR.n389 0.0680676
R8842 VPWR.n78 VPWR.n75 0.0680676
R8843 VPWR.n80 VPWR.n78 0.0680676
R8844 VPWR.n555 VPWR.n547 0.0680676
R8845 VPWR.n555 VPWR.n548 0.0680676
R8846 VPWR.n532 VPWR.n530 0.0680676
R8847 VPWR.n532 VPWR.n531 0.0680676
R8848 VPWR.n646 VPWR.n214 0.0680676
R8849 VPWR.n648 VPWR.n646 0.0680676
R8850 VPWR.n108 VPWR.n54 0.0680676
R8851 VPWR.n121 VPWR.n54 0.0680676
R8852 VPWR.n28 VPWR.n23 0.0680676
R8853 VPWR.n30 VPWR.n28 0.0680676
R8854 VPWR.n2239 VPWR.n147 0.0680676
R8855 VPWR.n2240 VPWR.n2239 0.0680676
R8856 VPWR.n2155 VPWR.n181 0.0680676
R8857 VPWR.n2155 VPWR.n2154 0.0680676
R8858 VPWR.n2118 VPWR.n197 0.0680676
R8859 VPWR.n2118 VPWR.n2117 0.0680676
R8860 VPWR.n2051 VPWR.n2049 0.0680676
R8861 VPWR.n2051 VPWR.n2050 0.0680676
R8862 VPWR.n2266 VPWR.n129 0.0680676
R8863 VPWR.n2279 VPWR.n129 0.0680676
R8864 VPWR.n164 VPWR.n162 0.0680676
R8865 VPWR.n164 VPWR.n163 0.0680676
R8866 VPWR.n2034 VPWR.n670 0.0680676
R8867 VPWR.n2034 VPWR.n2033 0.0680676
R8868 VPWR.n1323 VPWR.n1075 0.0680676
R8869 VPWR.n1325 VPWR.n1323 0.0680676
R8870 VPWR.n1196 VPWR.n1113 0.0680676
R8871 VPWR.n1196 VPWR.n1195 0.0680676
R8872 VPWR.n1161 VPWR.n1127 0.0680676
R8873 VPWR.n1162 VPWR.n1161 0.0680676
R8874 VPWR.n1999 VPWR.n698 0.0680676
R8875 VPWR.n700 VPWR.n698 0.0680676
R8876 VPWR.n1248 VPWR.n1099 0.0680676
R8877 VPWR.n1248 VPWR.n1100 0.0680676
R8878 VPWR.n1953 VPWR.n741 0.0680676
R8879 VPWR.n743 VPWR.n741 0.0680676
R8880 VPWR.n1525 VPWR.n1342 0.0680676
R8881 VPWR.n1527 VPWR.n1525 0.0680676
R8882 VPWR.n1454 VPWR.n1354 0.0680676
R8883 VPWR.n1455 VPWR.n1454 0.0680676
R8884 VPWR.n1402 VPWR.n1370 0.0680676
R8885 VPWR.n1403 VPWR.n1402 0.0680676
R8886 VPWR.n784 VPWR.n783 0.0680676
R8887 VPWR.n783 VPWR.n763 0.0680676
R8888 VPWR.n721 VPWR.n715 0.0680676
R8889 VPWR.n723 VPWR.n721 0.0680676
R8890 VPWR.n1614 VPWR.n1050 0.0680676
R8891 VPWR.n1615 VPWR.n1614 0.0680676
R8892 VPWR.n1755 VPWR.n937 0.0680676
R8893 VPWR.n1755 VPWR.n934 0.0680676
R8894 VPWR.n1572 VPWR.n1543 0.0680676
R8895 VPWR.n1572 VPWR.n1571 0.0680676
R8896 VPWR.n1661 VPWR.n1036 0.0680676
R8897 VPWR.n1039 VPWR.n1036 0.0680676
R8898 VPWR.n1913 VPWR.n1912 0.0680676
R8899 VPWR.n1912 VPWR.n1892 0.0680676
R8900 VPWR.n1684 VPWR.n995 0.0680676
R8901 VPWR.n1686 VPWR.n1684 0.0680676
R8902 VPWR.n944 VPWR.n941 0.0680676
R8903 VPWR.n1833 VPWR.n944 0.0680676
R8904 VPWR.n963 VPWR.n962 0.0680676
R8905 VPWR.n962 VPWR.n961 0.0680676
R8906 VPWR.n896 VPWR.n895 0.0680676
R8907 VPWR.n895 VPWR.n877 0.0680676
R8908 VPWR.n839 VPWR.n835 0.0680676
R8909 VPWR.n1882 VPWR.n839 0.0680676
R8910 VPWR.n429 VPWR.n428 0.0680676
R8911 VPWR.n446 VPWR.n429 0.0680676
R8912 VPWR.n623 VPWR.n622 0.0656042
R8913 VPWR.n2110 VPWR.n196 0.0656042
R8914 VPWR.n1188 VPWR.n1112 0.0656042
R8915 VPWR.n1442 VPWR.n1438 0.0656042
R8916 VPWR.n1034 VPWR.n1027 0.0656042
R8917 VPWR.n1736 VPWR.n1735 0.0656042
R8918 VPWR.n332 VPWR.n253 0.0656042
R8919 VPWR.n236 VPWR 0.0603958
R8920 VPWR.n636 VPWR 0.0603958
R8921 VPWR VPWR.n611 0.0603958
R8922 VPWR.n600 VPWR 0.0603958
R8923 VPWR.n2304 VPWR 0.0603958
R8924 VPWR VPWR.n2302 0.0603958
R8925 VPWR.n103 VPWR 0.0603958
R8926 VPWR VPWR.n2060 0.0603958
R8927 VPWR.n2096 VPWR 0.0603958
R8928 VPWR.n2149 VPWR 0.0603958
R8929 VPWR.n2208 VPWR 0.0603958
R8930 VPWR.n2218 VPWR 0.0603958
R8931 VPWR VPWR.n150 0.0603958
R8932 VPWR.n2250 VPWR 0.0603958
R8933 VPWR.n2255 VPWR 0.0603958
R8934 VPWR VPWR.n2262 0.0603958
R8935 VPWR.n1144 VPWR 0.0603958
R8936 VPWR.n1148 VPWR 0.0603958
R8937 VPWR VPWR.n1120 0.0603958
R8938 VPWR VPWR.n1239 0.0603958
R8939 VPWR VPWR.n1238 0.0603958
R8940 VPWR.n1224 VPWR 0.0603958
R8941 VPWR.n1305 VPWR 0.0603958
R8942 VPWR.n1302 VPWR 0.0603958
R8943 VPWR VPWR.n1301 0.0603958
R8944 VPWR VPWR.n1292 0.0603958
R8945 VPWR.n1288 VPWR 0.0603958
R8946 VPWR VPWR.n1287 0.0603958
R8947 VPWR.n2011 VPWR 0.0603958
R8948 VPWR.n2008 VPWR 0.0603958
R8949 VPWR.n1384 VPWR 0.0603958
R8950 VPWR.n1392 VPWR 0.0603958
R8951 VPWR.n1414 VPWR 0.0603958
R8952 VPWR VPWR.n1360 0.0603958
R8953 VPWR.n1461 VPWR 0.0603958
R8954 VPWR.n1468 VPWR 0.0603958
R8955 VPWR.n1470 VPWR 0.0603958
R8956 VPWR VPWR.n1476 0.0603958
R8957 VPWR.n1477 VPWR 0.0603958
R8958 VPWR.n1481 VPWR 0.0603958
R8959 VPWR.n1523 VPWR 0.0603958
R8960 VPWR.n1520 VPWR 0.0603958
R8961 VPWR.n1511 VPWR 0.0603958
R8962 VPWR VPWR.n1510 0.0603958
R8963 VPWR.n1510 VPWR 0.0603958
R8964 VPWR.n1507 VPWR 0.0603958
R8965 VPWR VPWR.n1506 0.0603958
R8966 VPWR VPWR.n1976 0.0603958
R8967 VPWR.n1973 VPWR 0.0603958
R8968 VPWR VPWR.n1972 0.0603958
R8969 VPWR VPWR.n800 0.0603958
R8970 VPWR.n795 VPWR 0.0603958
R8971 VPWR.n1013 VPWR 0.0603958
R8972 VPWR VPWR.n1653 0.0603958
R8973 VPWR.n1550 VPWR 0.0603958
R8974 VPWR.n1589 VPWR 0.0603958
R8975 VPWR VPWR.n1589 0.0603958
R8976 VPWR.n1590 VPWR 0.0603958
R8977 VPWR.n1597 VPWR 0.0603958
R8978 VPWR.n1603 VPWR 0.0603958
R8979 VPWR.n1620 VPWR 0.0603958
R8980 VPWR.n1645 VPWR 0.0603958
R8981 VPWR.n1643 VPWR 0.0603958
R8982 VPWR.n1629 VPWR 0.0603958
R8983 VPWR.n1925 VPWR 0.0603958
R8984 VPWR.n1919 VPWR 0.0603958
R8985 VPWR VPWR.n969 0.0603958
R8986 VPWR.n982 VPWR 0.0603958
R8987 VPWR.n983 VPWR 0.0603958
R8988 VPWR VPWR.n1714 0.0603958
R8989 VPWR.n1715 VPWR 0.0603958
R8990 VPWR VPWR.n955 0.0603958
R8991 VPWR VPWR.n1720 0.0603958
R8992 VPWR.n1721 VPWR 0.0603958
R8993 VPWR.n1725 VPWR 0.0603958
R8994 VPWR VPWR.n1726 0.0603958
R8995 VPWR.n1727 VPWR 0.0603958
R8996 VPWR.n1827 VPWR 0.0603958
R8997 VPWR VPWR.n1826 0.0603958
R8998 VPWR VPWR.n1825 0.0603958
R8999 VPWR.n1821 VPWR 0.0603958
R9000 VPWR.n1751 VPWR 0.0603958
R9001 VPWR VPWR.n1752 0.0603958
R9002 VPWR.n1809 VPWR 0.0603958
R9003 VPWR.n1809 VPWR 0.0603958
R9004 VPWR.n1789 VPWR 0.0603958
R9005 VPWR.n1787 VPWR 0.0603958
R9006 VPWR.n1784 VPWR 0.0603958
R9007 VPWR.n843 VPWR 0.0603958
R9008 VPWR.n1875 VPWR 0.0603958
R9009 VPWR VPWR.n1874 0.0603958
R9010 VPWR VPWR.n847 0.0603958
R9011 VPWR.n1863 VPWR 0.0603958
R9012 VPWR.n1859 VPWR 0.0603958
R9013 VPWR.n915 VPWR 0.0603958
R9014 VPWR.n909 VPWR 0.0603958
R9015 VPWR VPWR.n908 0.0603958
R9016 VPWR VPWR.n904 0.0603958
R9017 VPWR.n901 VPWR 0.0603958
R9018 VPWR.n295 VPWR 0.0603958
R9019 VPWR.n318 VPWR 0.0603958
R9020 VPWR VPWR.n2343 0.0603958
R9021 VPWR.n500 VPWR 0.0603958
R9022 VPWR VPWR.n499 0.0603958
R9023 VPWR VPWR.n498 0.0603958
R9024 VPWR VPWR.n472 0.0603958
R9025 VPWR.n2238 VPWR 0.0577917
R9026 VPWR.n1407 VPWR 0.0577917
R9027 VPWR.n926 VPWR 0.0577917
R9028 VPWR.n478 VPWR.n409 0.0574697
R9029 VPWR.n514 VPWR.n252 0.0574697
R9030 VPWR.n269 VPWR.n268 0.0574697
R9031 VPWR.n1941 VPWR.n813 0.0574697
R9032 VPWR.n2328 VPWR.n13 0.0574697
R9033 VPWR.n391 VPWR.n341 0.0574697
R9034 VPWR.n79 VPWR.n46 0.0574697
R9035 VPWR.n590 VPWR.n589 0.0574697
R9036 VPWR.n524 VPWR.n250 0.0574697
R9037 VPWR.n647 VPWR.n212 0.0574697
R9038 VPWR.n122 VPWR.n53 0.0574697
R9039 VPWR.n29 VPWR.n21 0.0574697
R9040 VPWR.n2241 VPWR.n146 0.0574697
R9041 VPWR.n179 VPWR.n176 0.0574697
R9042 VPWR.n195 VPWR.n192 0.0574697
R9043 VPWR.n2047 VPWR.n209 0.0574697
R9044 VPWR.n2280 VPWR.n128 0.0574697
R9045 VPWR.n160 VPWR.n158 0.0574697
R9046 VPWR.n2032 VPWR.n668 0.0574697
R9047 VPWR.n1324 VPWR.n1073 0.0574697
R9048 VPWR.n1111 VPWR.n1107 0.0574697
R9049 VPWR.n1163 VPWR.n1126 0.0574697
R9050 VPWR.n1998 VPWR.n1997 0.0574697
R9051 VPWR.n1297 VPWR.n1296 0.0574697
R9052 VPWR.n1952 VPWR.n742 0.0574697
R9053 VPWR.n1526 VPWR.n1340 0.0574697
R9054 VPWR.n1456 VPWR.n1353 0.0574697
R9055 VPWR.n1404 VPWR.n1369 0.0574697
R9056 VPWR.n785 VPWR.n762 0.0574697
R9057 VPWR.n722 VPWR.n713 0.0574697
R9058 VPWR.n1616 VPWR.n1049 0.0574697
R9059 VPWR.n1578 VPWR.n1541 0.0574697
R9060 VPWR.n1580 VPWR.n1071 0.0574697
R9061 VPWR.n1660 VPWR.n1037 0.0574697
R9062 VPWR.n1914 VPWR.n1891 0.0574697
R9063 VPWR.n1685 VPWR.n993 0.0574697
R9064 VPWR.n447 VPWR.n426 0.0574697
R9065 VPWR.n622 VPWR.n248 0.0551875
R9066 VPWR.n198 VPWR.n196 0.0551875
R9067 VPWR.n1114 VPWR.n1112 0.0551875
R9068 VPWR.n1443 VPWR.n1442 0.0551875
R9069 VPWR.n1664 VPWR.n1034 0.0551875
R9070 VPWR.n1737 VPWR.n1736 0.0551875
R9071 VPWR.n255 VPWR.n253 0.0551875
R9072 VPWR.n1831 VPWR 0.0538854
R9073 VPWR VPWR.n1774 0.0538854
R9074 VPWR.n435 VPWR 0.0538854
R9075 VPWR.n2264 VPWR 0.0525833
R9076 VPWR.n1041 VPWR 0.0525833
R9077 VPWR.n1740 VPWR 0.0525833
R9078 VPWR.n1773 VPWR 0.0525833
R9079 VPWR.n710 VPWR.n159 0.0522
R9080 VPWR.n1337 VPWR.n178 0.0522
R9081 VPWR.n2046 VPWR.n664 0.0522
R9082 VPWR.n1202 VPWR.n194 0.0522
R9083 VPWR.n2041 VPWR.n2040 0.0522
R9084 VPWR.n1995 VPWR.n126 0.0522
R9085 VPWR.n1842 VPWR.n1841 0.051025
R9086 VPWR.n652 VPWR.n215 0.0499792
R9087 VPWR.n557 VPWR.n553 0.0499792
R9088 VPWR.n2290 VPWR.n44 0.0499792
R9089 VPWR.n2077 VPWR.n2052 0.0499792
R9090 VPWR.n2158 VPWR.n2157 0.0499792
R9091 VPWR VPWR.n2228 0.0499792
R9092 VPWR.n1160 VPWR.n1159 0.0499792
R9093 VPWR.n1333 VPWR.n1332 0.0499792
R9094 VPWR.n671 VPWR.n669 0.0499792
R9095 VPWR.n1401 VPWR.n1400 0.0499792
R9096 VPWR.n1535 VPWR.n1534 0.0499792
R9097 VPWR.n1956 VPWR.n738 0.0499792
R9098 VPWR.n1690 VPWR.n996 0.0499792
R9099 VPWR.n1575 VPWR.n1574 0.0499792
R9100 VPWR.n816 VPWR.n814 0.0499792
R9101 VPWR.n1708 VPWR.n959 0.0499792
R9102 VPWR.n1806 VPWR.n1804 0.0499792
R9103 VPWR.n1857 VPWR.n854 0.0499792
R9104 VPWR.n299 VPWR.n274 0.0499792
R9105 VPWR.n2331 VPWR.n10 0.0499792
R9106 VPWR.n482 VPWR.n405 0.0499792
R9107 VPWR VPWR.n1808 0.047375
R9108 VPWR.n931 VPWR.n834 0.0460404
R9109 VPWR.n1853 VPWR.n1852 0.0460404
R9110 VPWR.n1849 VPWR.n930 0.0460404
R9111 VPWR.n1702 VPWR.n939 0.0454816
R9112 VPWR.n534 VPWR.n526 0.0447708
R9113 VPWR.n2313 VPWR.n24 0.0447708
R9114 VPWR.n112 VPWR.n110 0.0447708
R9115 VPWR.n199 VPWR.n190 0.0447708
R9116 VPWR.n2195 VPWR.n165 0.0447708
R9117 VPWR.n2245 VPWR.n2244 0.0447708
R9118 VPWR.n2270 VPWR.n2268 0.0447708
R9119 VPWR.n1115 VPWR.n1105 0.0447708
R9120 VPWR.n1251 VPWR.n1249 0.0447708
R9121 VPWR.n2001 VPWR.n696 0.0447708
R9122 VPWR.n1356 VPWR.n1351 0.0447708
R9123 VPWR.n1981 VPWR.n716 0.0447708
R9124 VPWR.n765 VPWR.n764 0.0447708
R9125 VPWR.n1044 VPWR.n1043 0.0447708
R9126 VPWR.n1613 VPWR.n1612 0.0447708
R9127 VPWR.n1938 VPWR.n819 0.0447708
R9128 VPWR.n1894 VPWR.n1893 0.0447708
R9129 VPWR.n1831 VPWR.n1830 0.0447708
R9130 VPWR.n1774 VPWR.n840 0.0447708
R9131 VPWR.n920 VPWR.n919 0.0447708
R9132 VPWR.n879 VPWR.n878 0.0447708
R9133 VPWR.n512 VPWR.n511 0.0447708
R9134 VPWR.n388 VPWR.n387 0.0447708
R9135 VPWR.n437 VPWR.n435 0.0447708
R9136 VPWR.n1838 VPWR.n1836 0.0446687
R9137 VPWR.n480 VPWR.n479 0.0410405
R9138 VPWR.n411 VPWR.n410 0.0410405
R9139 VPWR.n928 VPWR.n855 0.0410405
R9140 VPWR.n863 VPWR.n856 0.0410405
R9141 VPWR.n519 VPWR.n254 0.0410405
R9142 VPWR.n515 VPWR.n513 0.0410405
R9143 VPWR.n304 VPWR.n271 0.0410405
R9144 VPWR.n272 VPWR.n267 0.0410405
R9145 VPWR.n1946 VPWR.n815 0.0410405
R9146 VPWR.n1942 VPWR.n1940 0.0410405
R9147 VPWR.n2330 VPWR.n2329 0.0410405
R9148 VPWR.n355 VPWR.n354 0.0410405
R9149 VPWR.n378 VPWR.n342 0.0410405
R9150 VPWR.n390 VPWR.n340 0.0410405
R9151 VPWR.n75 VPWR.n45 0.0410405
R9152 VPWR.n82 VPWR.n80 0.0410405
R9153 VPWR.n547 VPWR.n546 0.0410405
R9154 VPWR.n549 VPWR.n548 0.0410405
R9155 VPWR.n530 VPWR.n249 0.0410405
R9156 VPWR.n531 VPWR.n525 0.0410405
R9157 VPWR.n657 VPWR.n214 0.0410405
R9158 VPWR.n650 VPWR.n648 0.0410405
R9159 VPWR.n109 VPWR.n108 0.0410405
R9160 VPWR.n121 VPWR.n120 0.0410405
R9161 VPWR.n2318 VPWR.n23 0.0410405
R9162 VPWR.n2311 VPWR.n30 0.0410405
R9163 VPWR.n2231 VPWR.n147 0.0410405
R9164 VPWR.n2240 VPWR.n145 0.0410405
R9165 VPWR.n2159 VPWR.n181 0.0410405
R9166 VPWR.n2154 VPWR.n175 0.0410405
R9167 VPWR.n2121 VPWR.n197 0.0410405
R9168 VPWR.n2117 VPWR.n191 0.0410405
R9169 VPWR.n2082 VPWR.n2049 0.0410405
R9170 VPWR.n2050 VPWR.n208 0.0410405
R9171 VPWR.n2267 VPWR.n2266 0.0410405
R9172 VPWR.n2279 VPWR.n2278 0.0410405
R9173 VPWR.n2200 VPWR.n162 0.0410405
R9174 VPWR.n163 VPWR.n157 0.0410405
R9175 VPWR.n2037 VPWR.n670 0.0410405
R9176 VPWR.n2033 VPWR.n2031 0.0410405
R9177 VPWR.n1334 VPWR.n1075 0.0410405
R9178 VPWR.n1326 VPWR.n1325 0.0410405
R9179 VPWR.n1199 VPWR.n1113 0.0410405
R9180 VPWR.n1195 VPWR.n1106 0.0410405
R9181 VPWR.n1149 VPWR.n1127 0.0410405
R9182 VPWR.n1162 VPWR.n1125 0.0410405
R9183 VPWR.n2000 VPWR.n1999 0.0410405
R9184 VPWR.n701 VPWR.n700 0.0410405
R9185 VPWR.n1099 VPWR.n1098 0.0410405
R9186 VPWR.n1101 VPWR.n1100 0.0410405
R9187 VPWR.n1954 VPWR.n1953 0.0410405
R9188 VPWR.n744 VPWR.n743 0.0410405
R9189 VPWR.n1536 VPWR.n1342 0.0410405
R9190 VPWR.n1528 VPWR.n1527 0.0410405
R9191 VPWR.n1439 VPWR.n1354 0.0410405
R9192 VPWR.n1455 VPWR.n1352 0.0410405
R9193 VPWR.n1394 VPWR.n1370 0.0410405
R9194 VPWR.n1403 VPWR.n1368 0.0410405
R9195 VPWR.n784 VPWR.n761 0.0410405
R9196 VPWR.n775 VPWR.n763 0.0410405
R9197 VPWR.n1986 VPWR.n715 0.0410405
R9198 VPWR.n1979 VPWR.n723 0.0410405
R9199 VPWR.n1599 VPWR.n1050 0.0410405
R9200 VPWR.n1615 VPWR.n1048 0.0410405
R9201 VPWR.n1805 VPWR.n937 0.0410405
R9202 VPWR.n1760 VPWR.n934 0.0410405
R9203 VPWR.n1576 VPWR.n1543 0.0410405
R9204 VPWR.n1571 VPWR.n1070 0.0410405
R9205 VPWR.n1662 VPWR.n1661 0.0410405
R9206 VPWR.n1040 VPWR.n1039 0.0410405
R9207 VPWR.n1913 VPWR.n831 0.0410405
R9208 VPWR.n1904 VPWR.n1892 0.0410405
R9209 VPWR.n1696 VPWR.n995 0.0410405
R9210 VPWR.n1688 VPWR.n1686 0.0410405
R9211 VPWR.n1738 VPWR.n941 0.0410405
R9212 VPWR.n1833 VPWR.n1832 0.0410405
R9213 VPWR.n989 VPWR.n963 0.0410405
R9214 VPWR.n1706 VPWR.n961 0.0410405
R9215 VPWR.n896 VPWR.n875 0.0410405
R9216 VPWR.n880 VPWR.n877 0.0410405
R9217 VPWR.n1772 VPWR.n835 0.0410405
R9218 VPWR.n1882 VPWR.n1881 0.0410405
R9219 VPWR.n428 VPWR.n425 0.0410405
R9220 VPWR.n446 VPWR.n445 0.0410405
R9221 VPWR.n2322 VPWR.n18 0.04045
R9222 VPWR.n2326 VPWR.n2325 0.04045
R9223 VPWR.n307 VPWR.n210 0.04045
R9224 VPWR.n523 VPWR.n522 0.04045
R9225 VPWR.n476 VPWR.n47 0.04045
R9226 VPWR.n451 VPWR.n450 0.04045
R9227 VPWR.n616 VPWR.n526 0.0395625
R9228 VPWR.n586 VPWR.n585 0.0395625
R9229 VPWR.n2313 VPWR.n2312 0.0395625
R9230 VPWR.n84 VPWR.n83 0.0395625
R9231 VPWR.n112 VPWR.n111 0.0395625
R9232 VPWR.n2127 VPWR.n190 0.0395625
R9233 VPWR.n2165 VPWR.n172 0.0395625
R9234 VPWR.n2195 VPWR.n2194 0.0395625
R9235 VPWR.n2245 VPWR.n144 0.0395625
R9236 VPWR.n2270 VPWR.n2269 0.0395625
R9237 VPWR.n1205 VPWR.n1105 0.0395625
R9238 VPWR.n1328 VPWR.n1322 0.0395625
R9239 VPWR.n1251 VPWR.n1250 0.0395625
R9240 VPWR.n2030 VPWR.n2029 0.0395625
R9241 VPWR.n702 VPWR.n696 0.0395625
R9242 VPWR.n1459 VPWR.n1351 0.0395625
R9243 VPWR.n1530 VPWR.n1524 0.0395625
R9244 VPWR.n1981 VPWR.n1980 0.0395625
R9245 VPWR.n749 VPWR.n748 0.0395625
R9246 VPWR.n782 VPWR.n765 0.0395625
R9247 VPWR.n1655 VPWR.n1044 0.0395625
R9248 VPWR.n1582 VPWR.n1065 0.0395625
R9249 VPWR.n1612 VPWR.n1052 0.0395625
R9250 VPWR.n1939 VPWR.n1938 0.0395625
R9251 VPWR.n1911 VPWR.n1894 0.0395625
R9252 VPWR.n1830 VPWR.n945 0.0395625
R9253 VPWR.n1799 VPWR.n1798 0.0395625
R9254 VPWR.n1880 VPWR.n840 0.0395625
R9255 VPWR.n920 VPWR.n864 0.0395625
R9256 VPWR.n894 VPWR.n879 0.0395625
R9257 VPWR.n511 VPWR.n258 0.0395625
R9258 VPWR.n357 VPWR.n351 0.0395625
R9259 VPWR.n387 VPWR.n344 0.0395625
R9260 VPWR.n416 VPWR.n415 0.0395625
R9261 VPWR.n437 VPWR.n436 0.0395625
R9262 VPWR.n1801 VPWR.n1759 0.0382581
R9263 VPWR.n1841 VPWR 0.036925
R9264 VPWR VPWR.n931 0.0366988
R9265 VPWR.n1852 VPWR 0.0366988
R9266 VPWR.n1849 VPWR 0.0366988
R9267 VPWR VPWR.n939 0.0362546
R9268 VPWR.n1838 VPWR 0.0356084
R9269 VPWR.n652 VPWR.n651 0.0343542
R9270 VPWR.n557 VPWR.n556 0.0343542
R9271 VPWR.n76 VPWR.n44 0.0343542
R9272 VPWR.n118 VPWR.n117 0.0343542
R9273 VPWR.n2077 VPWR.n207 0.0343542
R9274 VPWR.n2157 VPWR.n2156 0.0343542
R9275 VPWR.n2276 VPWR.n2275 0.0343542
R9276 VPWR.n1159 VPWR.n1124 0.0343542
R9277 VPWR.n1332 VPWR.n1077 0.0343542
R9278 VPWR.n2036 VPWR.n671 0.0343542
R9279 VPWR.n706 VPWR.n705 0.0343542
R9280 VPWR.n1534 VPWR.n1344 0.0343542
R9281 VPWR.n1956 VPWR.n1955 0.0343542
R9282 VPWR.n779 VPWR.n778 0.0343542
R9283 VPWR.n1690 VPWR.n1689 0.0343542
R9284 VPWR.n1574 VPWR.n1573 0.0343542
R9285 VPWR.n1945 VPWR.n816 0.0343542
R9286 VPWR.n1908 VPWR.n1907 0.0343542
R9287 VPWR.n1708 VPWR.n1707 0.0343542
R9288 VPWR.n1804 VPWR.n1756 0.0343542
R9289 VPWR.n859 VPWR.n854 0.0343542
R9290 VPWR.n891 VPWR.n890 0.0343542
R9291 VPWR.n299 VPWR.n266 0.0343542
R9292 VPWR.n352 VPWR.n10 0.0343542
R9293 VPWR.n443 VPWR.n442 0.0343542
R9294 VPWR VPWR.n1392 0.0330521
R9295 VPWR VPWR.n1469 0.0330521
R9296 VPWR.n1973 VPWR 0.0330521
R9297 VPWR VPWR.n981 0.0330521
R9298 VPWR.n1875 VPWR 0.0330521
R9299 VPWR.n499 VPWR 0.0330521
R9300 VPWR.n612 VPWR 0.03175
R9301 VPWR.n611 VPWR 0.03175
R9302 VPWR.n2308 VPWR 0.03175
R9303 VPWR VPWR.n103 0.03175
R9304 VPWR VPWR.n2131 0.03175
R9305 VPWR VPWR.n2207 0.03175
R9306 VPWR VPWR.n2250 0.03175
R9307 VPWR.n1240 VPWR 0.03175
R9308 VPWR.n1239 VPWR 0.03175
R9309 VPWR.n1302 VPWR 0.03175
R9310 VPWR.n1292 VPWR 0.03175
R9311 VPWR.n1384 VPWR 0.03175
R9312 VPWR.n1461 VPWR 0.03175
R9313 VPWR.n1507 VPWR 0.03175
R9314 VPWR.n1976 VPWR 0.03175
R9315 VPWR.n1663 VPWR 0.03175
R9316 VPWR.n1653 VPWR 0.03175
R9317 VPWR.n1721 VPWR 0.03175
R9318 VPWR VPWR.n1739 0.03175
R9319 VPWR.n1826 VPWR 0.03175
R9320 VPWR.n1825 VPWR 0.03175
R9321 VPWR.n1807 VPWR 0.03175
R9322 VPWR.n1784 VPWR 0.03175
R9323 VPWR VPWR.n1771 0.03175
R9324 VPWR VPWR.n843 0.03175
R9325 VPWR.n925 VPWR 0.03175
R9326 VPWR.n904 VPWR 0.03175
R9327 VPWR.n506 VPWR 0.03175
R9328 VPWR VPWR.n395 0.03175
R9329 VPWR.n500 VPWR 0.03175
R9330 VPWR.n53 VPWR.n51 0.0292489
R9331 VPWR.n123 VPWR.n122 0.0292489
R9332 VPWR.n128 VPWR.n125 0.0292489
R9333 VPWR.n2281 VPWR.n2280 0.0292489
R9334 VPWR.n1998 VPWR.n699 0.0292489
R9335 VPWR.n1997 VPWR.n1996 0.0292489
R9336 VPWR.n786 VPWR.n785 0.0292489
R9337 VPWR.n776 VPWR.n762 0.0292489
R9338 VPWR.n1600 VPWR.n1049 0.0292489
R9339 VPWR.n1617 VPWR.n1616 0.0292489
R9340 VPWR.n1988 VPWR.n713 0.0292489
R9341 VPWR.n722 VPWR.n711 0.0292489
R9342 VPWR.n1298 VPWR.n1297 0.0292489
R9343 VPWR.n1296 VPWR.n1295 0.0292489
R9344 VPWR.n2202 VPWR.n160 0.0292489
R9345 VPWR.n2204 VPWR.n158 0.0292489
R9346 VPWR.n2320 VPWR.n21 0.0292489
R9347 VPWR.n29 VPWR.n19 0.0292489
R9348 VPWR.n379 VPWR.n341 0.0292489
R9349 VPWR.n392 VPWR.n391 0.0292489
R9350 VPWR.n1538 VPWR.n1340 0.0292489
R9351 VPWR.n1526 VPWR.n1339 0.0292489
R9352 VPWR.n1336 VPWR.n1073 0.0292489
R9353 VPWR.n1324 VPWR.n1072 0.0292489
R9354 VPWR.n2161 VPWR.n179 0.0292489
R9355 VPWR.n2163 VPWR.n176 0.0292489
R9356 VPWR.n591 VPWR.n590 0.0292489
R9357 VPWR.n589 VPWR.n588 0.0292489
R9358 VPWR.n2328 VPWR.n2327 0.0292489
R9359 VPWR.n14 VPWR.n13 0.0292489
R9360 VPWR.n1540 VPWR.n1071 0.0292489
R9361 VPWR.n1541 VPWR.n1540 0.0292489
R9362 VPWR.n1915 VPWR.n1914 0.0292489
R9363 VPWR.n1905 VPWR.n1891 0.0292489
R9364 VPWR.n1698 VPWR.n993 0.0292489
R9365 VPWR.n1685 VPWR.n992 0.0292489
R9366 VPWR.n1395 VPWR.n1369 0.0292489
R9367 VPWR.n1405 VPWR.n1404 0.0292489
R9368 VPWR.n1150 VPWR.n1126 0.0292489
R9369 VPWR.n1164 VPWR.n1163 0.0292489
R9370 VPWR.n2084 VPWR.n2047 0.0292489
R9371 VPWR.n2086 VPWR.n209 0.0292489
R9372 VPWR.n659 VPWR.n212 0.0292489
R9373 VPWR.n647 VPWR.n211 0.0292489
R9374 VPWR.n306 VPWR.n269 0.0292489
R9375 VPWR.n308 VPWR.n268 0.0292489
R9376 VPWR.n1660 VPWR.n1659 0.0292489
R9377 VPWR.n1657 VPWR.n1037 0.0292489
R9378 VPWR.n1440 VPWR.n1353 0.0292489
R9379 VPWR.n1457 VPWR.n1456 0.0292489
R9380 VPWR.n1201 VPWR.n1111 0.0292489
R9381 VPWR.n1203 VPWR.n1107 0.0292489
R9382 VPWR.n2123 VPWR.n195 0.0292489
R9383 VPWR.n2125 VPWR.n192 0.0292489
R9384 VPWR.n620 VPWR.n250 0.0292489
R9385 VPWR.n618 VPWR.n524 0.0292489
R9386 VPWR.n521 VPWR.n252 0.0292489
R9387 VPWR.n514 VPWR.n251 0.0292489
R9388 VPWR.n1948 VPWR.n813 0.0292489
R9389 VPWR.n1941 VPWR.n811 0.0292489
R9390 VPWR.n1952 VPWR.n1951 0.0292489
R9391 VPWR.n810 VPWR.n742 0.0292489
R9392 VPWR.n2039 VPWR.n668 0.0292489
R9393 VPWR.n2032 VPWR.n666 0.0292489
R9394 VPWR.n2229 VPWR.n146 0.0292489
R9395 VPWR.n2242 VPWR.n2241 0.0292489
R9396 VPWR.n2288 VPWR.n46 0.0292489
R9397 VPWR.n79 VPWR.n48 0.0292489
R9398 VPWR.n478 VPWR.n477 0.0292489
R9399 VPWR.n475 VPWR.n409 0.0292489
R9400 VPWR.n452 VPWR.n426 0.0292489
R9401 VPWR.n448 VPWR.n447 0.0292489
R9402 VPWR.n529 VPWR.n248 0.0291458
R9403 VPWR.n564 VPWR.n22 0.0291458
R9404 VPWR.n2120 VPWR.n198 0.0291458
R9405 VPWR.n2189 VPWR.n161 0.0291458
R9406 VPWR.n1198 VPWR.n1114 0.0291458
R9407 VPWR.n1301 VPWR.n1300 0.0291458
R9408 VPWR.n1443 VPWR.n1355 0.0291458
R9409 VPWR.n1506 VPWR.n714 0.0291458
R9410 VPWR.n1603 VPWR.n1602 0.0291458
R9411 VPWR.n518 VPWR.n255 0.0291458
R9412 VPWR.n382 VPWR.n381 0.0291458
R9413 VPWR.n2232 VPWR 0.0265417
R9414 VPWR.n1372 VPWR 0.0265417
R9415 VPWR VPWR.n859 0.0265417
R9416 VPWR.n237 VPWR.n213 0.0239375
R9417 VPWR.n2059 VPWR.n2048 0.0239375
R9418 VPWR.n1153 VPWR.n1152 0.0239375
R9419 VPWR VPWR.n1481 0.0239375
R9420 VPWR.n1013 VPWR.n994 0.0239375
R9421 VPWR.n1919 VPWR 0.0239375
R9422 VPWR.n966 VPWR.n964 0.0239375
R9423 VPWR.n296 VPWR.n270 0.0239375
R9424 VPWR.n1993 VPWR 0.022975
R9425 VPWR.n449 VPWR 0.022975
R9426 VPWR.n2284 VPWR 0.022975
R9427 VPWR.n665 VPWR 0.022975
R9428 VPWR.n1888 VPWR 0.022975
R9429 VPWR.n1850 VPWR 0.022975
R9430 VPWR.n639 VPWR 0.0226354
R9431 VPWR.n630 VPWR 0.0226354
R9432 VPWR.n615 VPWR 0.0226354
R9433 VPWR.n580 VPWR 0.0226354
R9434 VPWR.n2304 VPWR 0.0226354
R9435 VPWR.n2302 VPWR 0.0226354
R9436 VPWR.n84 VPWR 0.0226354
R9437 VPWR VPWR.n69 0.0226354
R9438 VPWR.n100 VPWR 0.0226354
R9439 VPWR.n105 VPWR 0.0226354
R9440 VPWR.n117 VPWR 0.0226354
R9441 VPWR VPWR.n2095 0.0226354
R9442 VPWR.n2102 VPWR 0.0226354
R9443 VPWR.n2128 VPWR 0.0226354
R9444 VPWR VPWR.n2148 0.0226354
R9445 VPWR.n2172 VPWR 0.0226354
R9446 VPWR.n2182 VPWR 0.0226354
R9447 VPWR.n2215 VPWR 0.0226354
R9448 VPWR VPWR.n2218 0.0226354
R9449 VPWR VPWR.n2255 0.0226354
R9450 VPWR.n2263 VPWR 0.0226354
R9451 VPWR.n2275 VPWR 0.0226354
R9452 VPWR.n1144 VPWR 0.0226354
R9453 VPWR.n1172 VPWR 0.0226354
R9454 VPWR.n1178 VPWR 0.0226354
R9455 VPWR VPWR.n1206 0.0226354
R9456 VPWR.n1238 VPWR 0.0226354
R9457 VPWR.n1230 VPWR 0.0226354
R9458 VPWR VPWR.n1209 0.0226354
R9459 VPWR.n1315 VPWR 0.0226354
R9460 VPWR.n1288 VPWR 0.0226354
R9461 VPWR.n1287 VPWR 0.0226354
R9462 VPWR.n2029 VPWR 0.0226354
R9463 VPWR.n676 VPWR 0.0226354
R9464 VPWR.n2002 VPWR 0.0226354
R9465 VPWR.n705 VPWR 0.0226354
R9466 VPWR.n1400 VPWR 0.0226354
R9467 VPWR.n1408 VPWR 0.0226354
R9468 VPWR VPWR.n1413 0.0226354
R9469 VPWR.n1428 VPWR 0.0226354
R9470 VPWR VPWR.n1460 0.0226354
R9471 VPWR.n1470 VPWR 0.0226354
R9472 VPWR.n1477 VPWR 0.0226354
R9473 VPWR.n1520 VPWR 0.0226354
R9474 VPWR.n749 VPWR 0.0226354
R9475 VPWR.n808 VPWR 0.0226354
R9476 VPWR.n801 VPWR 0.0226354
R9477 VPWR VPWR.n760 0.0226354
R9478 VPWR.n779 VPWR 0.0226354
R9479 VPWR.n1664 VPWR 0.0226354
R9480 VPWR.n1654 VPWR 0.0226354
R9481 VPWR.n1583 VPWR 0.0226354
R9482 VPWR.n1065 VPWR 0.0226354
R9483 VPWR VPWR.n1588 0.0226354
R9484 VPWR VPWR.n1620 0.0226354
R9485 VPWR.n1928 VPWR 0.0226354
R9486 VPWR VPWR.n827 0.0226354
R9487 VPWR VPWR.n830 0.0226354
R9488 VPWR.n1908 VPWR 0.0226354
R9489 VPWR VPWR.n982 0.0226354
R9490 VPWR.n987 VPWR 0.0226354
R9491 VPWR.n1715 VPWR 0.0226354
R9492 VPWR.n955 VPWR 0.0226354
R9493 VPWR.n1727 VPWR 0.0226354
R9494 VPWR VPWR.n1737 0.0226354
R9495 VPWR.n1741 VPWR 0.0226354
R9496 VPWR.n1821 VPWR 0.0226354
R9497 VPWR.n1814 VPWR 0.0226354
R9498 VPWR VPWR.n1751 0.0226354
R9499 VPWR.n1792 VPWR 0.0226354
R9500 VPWR.n1789 VPWR 0.0226354
R9501 VPWR.n1775 VPWR 0.0226354
R9502 VPWR.n1874 VPWR 0.0226354
R9503 VPWR.n1862 VPWR 0.0226354
R9504 VPWR.n1859 VPWR 0.0226354
R9505 VPWR.n918 VPWR 0.0226354
R9506 VPWR.n913 VPWR 0.0226354
R9507 VPWR.n909 VPWR 0.0226354
R9508 VPWR.n908 VPWR 0.0226354
R9509 VPWR.n901 VPWR 0.0226354
R9510 VPWR VPWR.n874 0.0226354
R9511 VPWR.n891 VPWR 0.0226354
R9512 VPWR VPWR.n317 0.0226354
R9513 VPWR.n324 VPWR 0.0226354
R9514 VPWR.n507 VPWR 0.0226354
R9515 VPWR.n485 VPWR 0.0226354
R9516 VPWR.n482 VPWR 0.0226354
R9517 VPWR.n416 VPWR 0.0226354
R9518 VPWR.n473 VPWR 0.0226354
R9519 VPWR VPWR.n424 0.0226354
R9520 VPWR.n442 VPWR 0.0226354
R9521 VPWR.n1846 VPWR.n1845 0.0218125
R9522 VPWR.n2220 VPWR 0.0213333
R9523 VPWR VPWR.n754 0.0213333
R9524 VPWR VPWR.n1582 0.0213333
R9525 VPWR VPWR.n1597 0.0213333
R9526 VPWR.n864 VPWR 0.0213333
R9527 VPWR.n2309 VPWR 0.0200312
R9528 VPWR VPWR.n2206 0.0200312
R9529 VPWR.n1293 VPWR 0.0200312
R9530 VPWR.n1977 VPWR 0.0200312
R9531 VPWR VPWR.n1619 0.0200312
R9532 VPWR VPWR.n841 0.0200312
R9533 VPWR VPWR.n394 0.0200312
R9534 VPWR.n1990 VPWR.n1989 0.018125
R9535 VPWR.n1539 VPWR.n1338 0.018125
R9536 VPWR.n1108 VPWR.n991 0.018125
R9537 VPWR.n1110 VPWR.n1038 0.018125
R9538 VPWR.n1950 VPWR.n667 0.018125
R9539 VPWR.n1994 VPWR.n708 0.018125
R9540 VPWR.n1885 VPWR.n712 0.01695
R9541 VPWR.n1579 VPWR.n938 0.01695
R9542 VPWR.n1701 VPWR.n1699 0.01695
R9543 VPWR.n1658 VPWR.n940 0.01695
R9544 VPWR.n1949 VPWR.n812 0.01695
R9545 VPWR.n1890 VPWR.n1889 0.01695
R9546 VPWR.n110 VPWR 0.016125
R9547 VPWR.n2268 VPWR 0.016125
R9548 VPWR VPWR.n2001 0.016125
R9549 VPWR.n764 VPWR 0.016125
R9550 VPWR.n1893 VPWR 0.016125
R9551 VPWR.n878 VPWR 0.016125
R9552 VPWR.n473 VPWR 0.016125
R9553 VPWR.n656 VPWR.n655 0.0135208
R9554 VPWR.n593 VPWR.n545 0.0135208
R9555 VPWR.n2081 VPWR.n2080 0.0135208
R9556 VPWR.n2153 VPWR.n180 0.0135208
R9557 VPWR.n1158 VPWR.n1128 0.0135208
R9558 VPWR.n1076 VPWR.n1074 0.0135208
R9559 VPWR.n1393 VPWR.n1371 0.0135208
R9560 VPWR.n1343 VPWR.n1341 0.0135208
R9561 VPWR.n1695 VPWR.n1694 0.0135208
R9562 VPWR.n1570 VPWR.n1542 0.0135208
R9563 VPWR.n988 VPWR.n987 0.0135208
R9564 VPWR.n1808 VPWR.n1807 0.0135208
R9565 VPWR.n303 VPWR.n302 0.0135208
R9566 VPWR.n2332 VPWR.n9 0.0135208
R9567 VPWR VPWR.n2232 0.0122188
R9568 VPWR VPWR.n1372 0.0122188
R9569 VPWR VPWR.n481 0.0122188
R9570 VPWR VPWR.n959 0.0109167
R9571 VPWR VPWR.n1806 0.0109167
R9572 VPWR.n405 VPWR 0.0109167
R9573 VPWR.n1847 VPWR 0.00972152
R9574 VPWR VPWR.n932 0.00972152
R9575 VPWR VPWR.n1837 0.00972152
R9576 VPWR.n1848 VPWR 0.00972152
R9577 VPWR.n535 VPWR.n533 0.0083125
R9578 VPWR.n2317 VPWR.n2316 0.0083125
R9579 VPWR.n106 VPWR.n105 0.0083125
R9580 VPWR.n2119 VPWR.n2116 0.0083125
R9581 VPWR.n2199 VPWR.n2198 0.0083125
R9582 VPWR.n2264 VPWR.n2263 0.0083125
R9583 VPWR.n1197 VPWR.n1194 0.0083125
R9584 VPWR.n1247 VPWR.n1097 0.0083125
R9585 VPWR.n2002 VPWR.n695 0.0083125
R9586 VPWR.n1453 VPWR.n1452 0.0083125
R9587 VPWR.n1985 VPWR.n1984 0.0083125
R9588 VPWR.n788 VPWR.n760 0.0083125
R9589 VPWR.n1042 VPWR.n1041 0.0083125
R9590 VPWR.n1598 VPWR.n1051 0.0083125
R9591 VPWR.n1917 VPWR.n830 0.0083125
R9592 VPWR.n1741 VPWR.n1740 0.0083125
R9593 VPWR.n1775 VPWR.n1773 0.0083125
R9594 VPWR.n899 VPWR.n874 0.0083125
R9595 VPWR.n517 VPWR.n256 0.0083125
R9596 VPWR.n377 VPWR.n343 0.0083125
R9597 VPWR.n454 VPWR.n424 0.0083125
R9598 VPWR VPWR.n1663 0.00701042
R9599 VPWR.n1739 VPWR 0.00701042
R9600 VPWR.n1771 VPWR 0.00701042
R9601 VPWR.n1884 VPWR.n834 0.0052
R9602 VPWR.n1703 VPWR.n1702 0.0052
R9603 VPWR.n1836 VPWR.n1835 0.0052
R9604 VPWR.n1854 VPWR.n1853 0.0052
R9605 VPWR.n930 VPWR.n832 0.0052
R9606 VPWR.n645 VPWR.n644 0.00310417
R9607 VPWR.n554 VPWR.n550 0.00310417
R9608 VPWR.n2309 VPWR.n27 0.00310417
R9609 VPWR.n77 VPWR.n74 0.00310417
R9610 VPWR.n119 VPWR.n55 0.00310417
R9611 VPWR.n2089 VPWR.n2088 0.00310417
R9612 VPWR.n2166 VPWR.n174 0.00310417
R9613 VPWR.n2206 VPWR.n156 0.00310417
R9614 VPWR.n2238 VPWR.n2237 0.00310417
R9615 VPWR.n2277 VPWR.n130 0.00310417
R9616 VPWR.n1167 VPWR.n1166 0.00310417
R9617 VPWR.n1329 VPWR.n1082 0.00310417
R9618 VPWR.n1293 VPWR.n1102 0.00310417
R9619 VPWR.n2035 VPWR.n672 0.00310417
R9620 VPWR.n704 VPWR.n703 0.00310417
R9621 VPWR.n1408 VPWR.n1407 0.00310417
R9622 VPWR.n1531 VPWR.n1489 0.00310417
R9623 VPWR.n1977 VPWR.n720 0.00310417
R9624 VPWR.n747 VPWR.n739 0.00310417
R9625 VPWR.n781 VPWR.n766 0.00310417
R9626 VPWR.n1683 VPWR.n1682 0.00310417
R9627 VPWR.n1583 VPWR.n1069 0.00310417
R9628 VPWR.n1619 VPWR.n1047 0.00310417
R9629 VPWR.n1944 VPWR.n817 0.00310417
R9630 VPWR.n1910 VPWR.n1895 0.00310417
R9631 VPWR.n960 VPWR.n957 0.00310417
R9632 VPWR.n1800 VPWR.n1761 0.00310417
R9633 VPWR.n1879 VPWR.n841 0.00310417
R9634 VPWR.n926 VPWR.n925 0.00310417
R9635 VPWR.n893 VPWR.n881 0.00310417
R9636 VPWR.n311 VPWR.n310 0.00310417
R9637 VPWR.n358 VPWR.n353 0.00310417
R9638 VPWR.n394 VPWR.n339 0.00310417
R9639 VPWR.n414 VPWR.n406 0.00310417
R9640 VPWR.n444 VPWR.n430 0.00310417
R9641 clknet_1_1__leaf_clk.n30 clknet_1_1__leaf_clk.n28 333.392
R9642 clknet_1_1__leaf_clk.n39 clknet_1_1__leaf_clk.n27 301.392
R9643 clknet_1_1__leaf_clk.n30 clknet_1_1__leaf_clk.n29 301.392
R9644 clknet_1_1__leaf_clk.n32 clknet_1_1__leaf_clk.n31 301.392
R9645 clknet_1_1__leaf_clk.n34 clknet_1_1__leaf_clk.n33 301.392
R9646 clknet_1_1__leaf_clk.n36 clknet_1_1__leaf_clk.n35 301.392
R9647 clknet_1_1__leaf_clk.n38 clknet_1_1__leaf_clk.n37 301.392
R9648 clknet_1_1__leaf_clk.n40 clknet_1_1__leaf_clk.n26 297.863
R9649 clknet_1_1__leaf_clk.n18 clknet_1_1__leaf_clk.t32 294.557
R9650 clknet_1_1__leaf_clk.n15 clknet_1_1__leaf_clk.t40 294.557
R9651 clknet_1_1__leaf_clk.n13 clknet_1_1__leaf_clk.t35 294.557
R9652 clknet_1_1__leaf_clk.n11 clknet_1_1__leaf_clk.t39 294.557
R9653 clknet_1_1__leaf_clk.n10 clknet_1_1__leaf_clk.t41 294.557
R9654 clknet_1_1__leaf_clk.n2 clknet_1_1__leaf_clk.n0 248.638
R9655 clknet_1_1__leaf_clk.n18 clknet_1_1__leaf_clk.t36 211.01
R9656 clknet_1_1__leaf_clk.n15 clknet_1_1__leaf_clk.t37 211.01
R9657 clknet_1_1__leaf_clk.n13 clknet_1_1__leaf_clk.t38 211.01
R9658 clknet_1_1__leaf_clk.n11 clknet_1_1__leaf_clk.t34 211.01
R9659 clknet_1_1__leaf_clk.n10 clknet_1_1__leaf_clk.t33 211.01
R9660 clknet_1_1__leaf_clk.n2 clknet_1_1__leaf_clk.n1 203.463
R9661 clknet_1_1__leaf_clk.n4 clknet_1_1__leaf_clk.n3 203.463
R9662 clknet_1_1__leaf_clk.n8 clknet_1_1__leaf_clk.n7 203.463
R9663 clknet_1_1__leaf_clk.n25 clknet_1_1__leaf_clk.n24 203.463
R9664 clknet_1_1__leaf_clk.n6 clknet_1_1__leaf_clk.n5 202.456
R9665 clknet_1_1__leaf_clk clknet_1_1__leaf_clk.n42 199.607
R9666 clknet_1_1__leaf_clk.n22 clknet_1_1__leaf_clk.n9 188.201
R9667 clknet_1_1__leaf_clk clknet_1_1__leaf_clk.n13 156.207
R9668 clknet_1_1__leaf_clk clknet_1_1__leaf_clk.n10 156.207
R9669 clknet_1_1__leaf_clk.n19 clknet_1_1__leaf_clk.n18 153.097
R9670 clknet_1_1__leaf_clk.n16 clknet_1_1__leaf_clk.n15 152.296
R9671 clknet_1_1__leaf_clk.n12 clknet_1_1__leaf_clk.n11 152.296
R9672 clknet_1_1__leaf_clk.n4 clknet_1_1__leaf_clk.n2 45.177
R9673 clknet_1_1__leaf_clk.n23 clknet_1_1__leaf_clk.n8 45.177
R9674 clknet_1_1__leaf_clk.n25 clknet_1_1__leaf_clk.n23 45.177
R9675 clknet_1_1__leaf_clk.n6 clknet_1_1__leaf_clk.n4 44.0476
R9676 clknet_1_1__leaf_clk.n8 clknet_1_1__leaf_clk.n6 44.0476
R9677 clknet_1_1__leaf_clk.n0 clknet_1_1__leaf_clk.t29 40.0005
R9678 clknet_1_1__leaf_clk.n0 clknet_1_1__leaf_clk.t30 40.0005
R9679 clknet_1_1__leaf_clk.n1 clknet_1_1__leaf_clk.t25 40.0005
R9680 clknet_1_1__leaf_clk.n1 clknet_1_1__leaf_clk.t27 40.0005
R9681 clknet_1_1__leaf_clk.n3 clknet_1_1__leaf_clk.t28 40.0005
R9682 clknet_1_1__leaf_clk.n3 clknet_1_1__leaf_clk.t23 40.0005
R9683 clknet_1_1__leaf_clk.n5 clknet_1_1__leaf_clk.t24 40.0005
R9684 clknet_1_1__leaf_clk.n5 clknet_1_1__leaf_clk.t26 40.0005
R9685 clknet_1_1__leaf_clk.n7 clknet_1_1__leaf_clk.t21 40.0005
R9686 clknet_1_1__leaf_clk.n7 clknet_1_1__leaf_clk.t22 40.0005
R9687 clknet_1_1__leaf_clk.n9 clknet_1_1__leaf_clk.t31 40.0005
R9688 clknet_1_1__leaf_clk.n9 clknet_1_1__leaf_clk.t20 40.0005
R9689 clknet_1_1__leaf_clk.n24 clknet_1_1__leaf_clk.t17 40.0005
R9690 clknet_1_1__leaf_clk.n24 clknet_1_1__leaf_clk.t18 40.0005
R9691 clknet_1_1__leaf_clk.n42 clknet_1_1__leaf_clk.t19 40.0005
R9692 clknet_1_1__leaf_clk.n42 clknet_1_1__leaf_clk.t16 40.0005
R9693 clknet_1_1__leaf_clk.n21 clknet_1_1__leaf_clk 34.5053
R9694 clknet_1_1__leaf_clk.n14 clknet_1_1__leaf_clk 33.8485
R9695 clknet_1_1__leaf_clk.n32 clknet_1_1__leaf_clk.n30 32.0005
R9696 clknet_1_1__leaf_clk.n34 clknet_1_1__leaf_clk.n32 32.0005
R9697 clknet_1_1__leaf_clk.n38 clknet_1_1__leaf_clk.n36 32.0005
R9698 clknet_1_1__leaf_clk.n39 clknet_1_1__leaf_clk.n38 32.0005
R9699 clknet_1_1__leaf_clk.n36 clknet_1_1__leaf_clk.n34 31.2005
R9700 clknet_1_1__leaf_clk.n27 clknet_1_1__leaf_clk.t12 27.5805
R9701 clknet_1_1__leaf_clk.n27 clknet_1_1__leaf_clk.t13 27.5805
R9702 clknet_1_1__leaf_clk.n26 clknet_1_1__leaf_clk.t14 27.5805
R9703 clknet_1_1__leaf_clk.n26 clknet_1_1__leaf_clk.t11 27.5805
R9704 clknet_1_1__leaf_clk.n28 clknet_1_1__leaf_clk.t8 27.5805
R9705 clknet_1_1__leaf_clk.n28 clknet_1_1__leaf_clk.t9 27.5805
R9706 clknet_1_1__leaf_clk.n29 clknet_1_1__leaf_clk.t4 27.5805
R9707 clknet_1_1__leaf_clk.n29 clknet_1_1__leaf_clk.t6 27.5805
R9708 clknet_1_1__leaf_clk.n31 clknet_1_1__leaf_clk.t7 27.5805
R9709 clknet_1_1__leaf_clk.n31 clknet_1_1__leaf_clk.t2 27.5805
R9710 clknet_1_1__leaf_clk.n33 clknet_1_1__leaf_clk.t3 27.5805
R9711 clknet_1_1__leaf_clk.n33 clknet_1_1__leaf_clk.t5 27.5805
R9712 clknet_1_1__leaf_clk.n35 clknet_1_1__leaf_clk.t0 27.5805
R9713 clknet_1_1__leaf_clk.n35 clknet_1_1__leaf_clk.t1 27.5805
R9714 clknet_1_1__leaf_clk.n37 clknet_1_1__leaf_clk.t10 27.5805
R9715 clknet_1_1__leaf_clk.n37 clknet_1_1__leaf_clk.t15 27.5805
R9716 clknet_1_1__leaf_clk.n23 clknet_1_1__leaf_clk.n22 15.262
R9717 clknet_1_1__leaf_clk.n20 clknet_1_1__leaf_clk.n19 13.8005
R9718 clknet_1_1__leaf_clk.n41 clknet_1_1__leaf_clk.n25 13.177
R9719 clknet_1_1__leaf_clk.n14 clknet_1_1__leaf_clk.n12 11.6482
R9720 clknet_1_1__leaf_clk.n22 clknet_1_1__leaf_clk.n21 10.8268
R9721 clknet_1_1__leaf_clk.n40 clknet_1_1__leaf_clk.n39 10.4484
R9722 clknet_1_1__leaf_clk.n17 clknet_1_1__leaf_clk.n16 9.3005
R9723 clknet_1_1__leaf_clk.n20 clknet_1_1__leaf_clk.n17 8.37704
R9724 clknet_1_1__leaf_clk.n21 clknet_1_1__leaf_clk 5.19349
R9725 clknet_1_1__leaf_clk.n17 clknet_1_1__leaf_clk.n14 3.99105
R9726 clknet_1_1__leaf_clk.n41 clknet_1_1__leaf_clk 3.13183
R9727 clknet_1_1__leaf_clk.n19 clknet_1_1__leaf_clk 3.10907
R9728 clknet_1_1__leaf_clk clknet_1_1__leaf_clk.n40 1.75844
R9729 clknet_1_1__leaf_clk.n16 clknet_1_1__leaf_clk 1.67435
R9730 clknet_1_1__leaf_clk.n12 clknet_1_1__leaf_clk 1.67435
R9731 clknet_1_1__leaf_clk clknet_1_1__leaf_clk.n20 0.693495
R9732 clknet_1_1__leaf_clk clknet_1_1__leaf_clk.n41 0.604792
R9733 counter[6].n0 counter[6].t0 368.521
R9734 counter[6].n1 counter[6].t1 216.155
R9735 counter[6].n1 counter[6] 78.8791
R9736 counter[6].n2 counter[6] 18.0287
R9737 counter[6] counter[6].n0 10.5563
R9738 counter[6].n0 counter[6] 5.48477
R9739 counter[6] counter[6].n2 4.18512
R9740 counter[6].n2 counter[6].n1 0.985115
R9741 counter[3].n0 counter[3].t0 368.521
R9742 counter[3].n1 counter[3].t1 216.155
R9743 counter[3].n1 counter[3] 78.8791
R9744 counter[3].n2 counter[3] 18.8501
R9745 counter[3] counter[3].n0 10.5563
R9746 counter[3].n0 counter[3] 5.48477
R9747 counter[3] counter[3].n2 4.18512
R9748 counter[3].n2 counter[3].n1 0.985115
R9749 clknet_1_0__leaf_clk.n6 clknet_1_0__leaf_clk.n4 333.392
R9750 clknet_1_0__leaf_clk.n6 clknet_1_0__leaf_clk.n5 301.392
R9751 clknet_1_0__leaf_clk.n8 clknet_1_0__leaf_clk.n7 301.392
R9752 clknet_1_0__leaf_clk.n10 clknet_1_0__leaf_clk.n9 301.392
R9753 clknet_1_0__leaf_clk.n12 clknet_1_0__leaf_clk.n11 301.392
R9754 clknet_1_0__leaf_clk.n31 clknet_1_0__leaf_clk.n13 301.392
R9755 clknet_1_0__leaf_clk.n30 clknet_1_0__leaf_clk.n14 297.863
R9756 clknet_1_0__leaf_clk.n2 clknet_1_0__leaf_clk.t33 294.557
R9757 clknet_1_0__leaf_clk.n0 clknet_1_0__leaf_clk.t37 294.557
R9758 clknet_1_0__leaf_clk.n41 clknet_1_0__leaf_clk.t36 294.557
R9759 clknet_1_0__leaf_clk.n38 clknet_1_0__leaf_clk.t34 294.557
R9760 clknet_1_0__leaf_clk.n36 clknet_1_0__leaf_clk.t32 294.557
R9761 clknet_1_0__leaf_clk.n34 clknet_1_0__leaf_clk.n33 287.303
R9762 clknet_1_0__leaf_clk.n17 clknet_1_0__leaf_clk.n15 248.638
R9763 clknet_1_0__leaf_clk.n2 clknet_1_0__leaf_clk.t38 211.01
R9764 clknet_1_0__leaf_clk.n0 clknet_1_0__leaf_clk.t41 211.01
R9765 clknet_1_0__leaf_clk.n41 clknet_1_0__leaf_clk.t40 211.01
R9766 clknet_1_0__leaf_clk.n38 clknet_1_0__leaf_clk.t39 211.01
R9767 clknet_1_0__leaf_clk.n36 clknet_1_0__leaf_clk.t35 211.01
R9768 clknet_1_0__leaf_clk.n17 clknet_1_0__leaf_clk.n16 203.463
R9769 clknet_1_0__leaf_clk.n19 clknet_1_0__leaf_clk.n18 203.463
R9770 clknet_1_0__leaf_clk.n23 clknet_1_0__leaf_clk.n22 203.463
R9771 clknet_1_0__leaf_clk.n25 clknet_1_0__leaf_clk.n24 203.463
R9772 clknet_1_0__leaf_clk.n27 clknet_1_0__leaf_clk.n26 203.463
R9773 clknet_1_0__leaf_clk.n21 clknet_1_0__leaf_clk.n20 202.456
R9774 clknet_1_0__leaf_clk clknet_1_0__leaf_clk.n28 199.607
R9775 clknet_1_0__leaf_clk clknet_1_0__leaf_clk.n2 156.207
R9776 clknet_1_0__leaf_clk.n37 clknet_1_0__leaf_clk.n36 153.097
R9777 clknet_1_0__leaf_clk.n39 clknet_1_0__leaf_clk.n38 152.296
R9778 clknet_1_0__leaf_clk.n1 clknet_1_0__leaf_clk.n0 152
R9779 clknet_1_0__leaf_clk.n42 clknet_1_0__leaf_clk.n41 152
R9780 clknet_1_0__leaf_clk.n19 clknet_1_0__leaf_clk.n17 45.177
R9781 clknet_1_0__leaf_clk.n25 clknet_1_0__leaf_clk.n23 45.177
R9782 clknet_1_0__leaf_clk.n27 clknet_1_0__leaf_clk.n25 45.177
R9783 clknet_1_0__leaf_clk.n21 clknet_1_0__leaf_clk.n19 44.0476
R9784 clknet_1_0__leaf_clk.n23 clknet_1_0__leaf_clk.n21 44.0476
R9785 clknet_1_0__leaf_clk.n15 clknet_1_0__leaf_clk.t26 40.0005
R9786 clknet_1_0__leaf_clk.n15 clknet_1_0__leaf_clk.t28 40.0005
R9787 clknet_1_0__leaf_clk.n16 clknet_1_0__leaf_clk.t30 40.0005
R9788 clknet_1_0__leaf_clk.n16 clknet_1_0__leaf_clk.t31 40.0005
R9789 clknet_1_0__leaf_clk.n18 clknet_1_0__leaf_clk.t29 40.0005
R9790 clknet_1_0__leaf_clk.n18 clknet_1_0__leaf_clk.t17 40.0005
R9791 clknet_1_0__leaf_clk.n20 clknet_1_0__leaf_clk.t19 40.0005
R9792 clknet_1_0__leaf_clk.n20 clknet_1_0__leaf_clk.t16 40.0005
R9793 clknet_1_0__leaf_clk.n22 clknet_1_0__leaf_clk.t22 40.0005
R9794 clknet_1_0__leaf_clk.n22 clknet_1_0__leaf_clk.t18 40.0005
R9795 clknet_1_0__leaf_clk.n24 clknet_1_0__leaf_clk.t20 40.0005
R9796 clknet_1_0__leaf_clk.n24 clknet_1_0__leaf_clk.t21 40.0005
R9797 clknet_1_0__leaf_clk.n26 clknet_1_0__leaf_clk.t23 40.0005
R9798 clknet_1_0__leaf_clk.n26 clknet_1_0__leaf_clk.t24 40.0005
R9799 clknet_1_0__leaf_clk.n28 clknet_1_0__leaf_clk.t25 40.0005
R9800 clknet_1_0__leaf_clk.n28 clknet_1_0__leaf_clk.t27 40.0005
R9801 clknet_1_0__leaf_clk.n8 clknet_1_0__leaf_clk.n6 32.0005
R9802 clknet_1_0__leaf_clk.n10 clknet_1_0__leaf_clk.n8 32.0005
R9803 clknet_1_0__leaf_clk.n32 clknet_1_0__leaf_clk.n12 32.0005
R9804 clknet_1_0__leaf_clk.n32 clknet_1_0__leaf_clk.n31 32.0005
R9805 clknet_1_0__leaf_clk.n12 clknet_1_0__leaf_clk.n10 31.2005
R9806 clknet_1_0__leaf_clk.n35 clknet_1_0__leaf_clk.n34 28.6283
R9807 clknet_1_0__leaf_clk.n3 clknet_1_0__leaf_clk 28.0697
R9808 clknet_1_0__leaf_clk.n14 clknet_1_0__leaf_clk.t1 27.5805
R9809 clknet_1_0__leaf_clk.n14 clknet_1_0__leaf_clk.t3 27.5805
R9810 clknet_1_0__leaf_clk.n4 clknet_1_0__leaf_clk.t2 27.5805
R9811 clknet_1_0__leaf_clk.n4 clknet_1_0__leaf_clk.t4 27.5805
R9812 clknet_1_0__leaf_clk.n5 clknet_1_0__leaf_clk.t6 27.5805
R9813 clknet_1_0__leaf_clk.n5 clknet_1_0__leaf_clk.t7 27.5805
R9814 clknet_1_0__leaf_clk.n7 clknet_1_0__leaf_clk.t5 27.5805
R9815 clknet_1_0__leaf_clk.n7 clknet_1_0__leaf_clk.t9 27.5805
R9816 clknet_1_0__leaf_clk.n9 clknet_1_0__leaf_clk.t11 27.5805
R9817 clknet_1_0__leaf_clk.n9 clknet_1_0__leaf_clk.t8 27.5805
R9818 clknet_1_0__leaf_clk.n11 clknet_1_0__leaf_clk.t14 27.5805
R9819 clknet_1_0__leaf_clk.n11 clknet_1_0__leaf_clk.t10 27.5805
R9820 clknet_1_0__leaf_clk.n33 clknet_1_0__leaf_clk.t12 27.5805
R9821 clknet_1_0__leaf_clk.n33 clknet_1_0__leaf_clk.t13 27.5805
R9822 clknet_1_0__leaf_clk.n13 clknet_1_0__leaf_clk.t15 27.5805
R9823 clknet_1_0__leaf_clk.n13 clknet_1_0__leaf_clk.t0 27.5805
R9824 clknet_1_0__leaf_clk.n43 clknet_1_0__leaf_clk.n42 27.3319
R9825 clknet_1_0__leaf_clk.n40 clknet_1_0__leaf_clk.n39 21.4985
R9826 clknet_1_0__leaf_clk.n3 clknet_1_0__leaf_clk.n1 21.401
R9827 clknet_1_0__leaf_clk.n34 clknet_1_0__leaf_clk.n32 14.0898
R9828 clknet_1_0__leaf_clk.n29 clknet_1_0__leaf_clk.n27 13.177
R9829 clknet_1_0__leaf_clk.n40 clknet_1_0__leaf_clk.n37 11.0654
R9830 clknet_1_0__leaf_clk.n31 clknet_1_0__leaf_clk.n30 10.4484
R9831 clknet_1_0__leaf_clk.n43 clknet_1_0__leaf_clk.n40 7.18319
R9832 clknet_1_0__leaf_clk.n35 clknet_1_0__leaf_clk.n3 5.63649
R9833 clknet_1_0__leaf_clk clknet_1_0__leaf_clk.n29 3.13183
R9834 clknet_1_0__leaf_clk.n37 clknet_1_0__leaf_clk 3.10907
R9835 clknet_1_0__leaf_clk clknet_1_0__leaf_clk.n43 2.66671
R9836 clknet_1_0__leaf_clk clknet_1_0__leaf_clk.n35 2.66671
R9837 clknet_1_0__leaf_clk.n42 clknet_1_0__leaf_clk 2.01193
R9838 clknet_1_0__leaf_clk.n30 clknet_1_0__leaf_clk 1.75844
R9839 clknet_1_0__leaf_clk.n39 clknet_1_0__leaf_clk 1.67435
R9840 clknet_1_0__leaf_clk.n1 clknet_1_0__leaf_clk 1.37896
R9841 clknet_1_0__leaf_clk.n29 clknet_1_0__leaf_clk 0.604792
R9842 _11_ _11_.n0 623.909
R9843 _11_.n24 _11_.t18 334.723
R9844 _11_.n5 _11_.t4 334.723
R9845 _11_.n18 _11_.t19 261.887
R9846 _11_.n14 _11_.t10 256.07
R9847 _11_.n8 _11_.t7 241.536
R9848 _11_.n3 _11_.t13 241.536
R9849 _11_.n1 _11_.t17 231.835
R9850 _11_.n21 _11_.t5 230.363
R9851 _11_ _11_.n30 216.464
R9852 _11_.n24 _11_.t9 206.19
R9853 _11_.n5 _11_.t14 206.19
R9854 _11_.n11 _11_.t8 183.505
R9855 _11_.n8 _11_.t20 169.237
R9856 _11_.n3 _11_.t6 169.237
R9857 _11_.n21 _11_.t16 158.064
R9858 _11_ _11_.n3 157.555
R9859 _11_ _11_.n8 157.166
R9860 _11_.n1 _11_.t11 157.07
R9861 _11_.n18 _11_.t15 155.847
R9862 _11_.n22 _11_.n21 154.048
R9863 _11_.n12 _11_.n11 153.863
R9864 _11_.n19 _11_.n18 153.13
R9865 _11_.n25 _11_.n24 152
R9866 _11_.n15 _11_.n14 152
R9867 _11_.n6 _11_.n5 152
R9868 _11_.n2 _11_.n1 152
R9869 _11_.n14 _11_.t21 150.03
R9870 _11_.n11 _11_.t12 114.532
R9871 _11_.n27 _11_.n26 41.0809
R9872 _11_.n30 _11_.t3 38.5719
R9873 _11_.n30 _11_.t2 38.5719
R9874 _11_.n0 _11_.t0 26.5955
R9875 _11_.n0 _11_.t1 26.5955
R9876 _11_.n17 _11_.n16 25.2401
R9877 _11_.n20 _11_.n19 22.3199
R9878 _11_.n10 _11_.n9 21.8442
R9879 _11_.n10 _11_.n7 20.8523
R9880 _11_.n28 _11_.n27 13.7699
R9881 _11_.n28 _11_.n2 12.7179
R9882 _11_.n4 _11_ 12.3175
R9883 _11_.n9 _11_ 11.4531
R9884 _11_.n7 _11_.n4 11.4418
R9885 _11_.n23 _11_.n20 10.8618
R9886 _11_.n7 _11_.n6 10.3976
R9887 _11_.n25 _11_ 9.6005
R9888 _11_.n29 _11_ 9.6005
R9889 _11_ _11_.n22 9.39918
R9890 _11_.n13 _11_.n12 9.3005
R9891 _11_.n29 _11_.n28 9.3005
R9892 _11_.n23 _11_ 8.80957
R9893 _11_.n6 _11_ 8.22907
R9894 _11_.n15 _11_ 7.6805
R9895 _11_.n16 _11_.n15 4.6085
R9896 _11_.n16 _11_ 4.58918
R9897 _11_.n22 _11_ 4.3525
R9898 _11_.n4 _11_ 4.10616
R9899 _11_.n9 _11_ 3.81804
R9900 _11_.n26 _11_ 3.62717
R9901 _11_.n19 _11_ 3.2005
R9902 _11_ _11_.n29 3.2005
R9903 _11_.n17 _11_.n13 2.49494
R9904 _11_.n2 _11_ 2.3045
R9905 _11_.n12 _11_ 1.97868
R9906 _11_.n13 _11_.n10 1.71582
R9907 _11_.n27 _11_.n23 1.38649
R9908 _11_.n26 _11_.n25 1.2805
R9909 _11_.n20 _11_.n17 1.24753
R9910 counter[2].n0 counter[2].t0 368.521
R9911 counter[2].n1 counter[2].t1 216.155
R9912 counter[2].n1 counter[2] 78.8791
R9913 counter[2].n2 counter[2] 18.0287
R9914 counter[2] counter[2].n0 10.5563
R9915 counter[2].n0 counter[2] 5.48477
R9916 counter[2] counter[2].n2 4.18512
R9917 counter[2].n2 counter[2].n1 0.985115
R9918 counter[0].n0 counter[0].t0 368.521
R9919 counter[0].n1 counter[0].t1 216.155
R9920 counter[0].n1 counter[0] 78.8791
R9921 counter[0].n2 counter[0] 20.493
R9922 counter[0] counter[0].n0 10.5563
R9923 counter[0].n0 counter[0] 5.48477
R9924 counter[0] counter[0].n2 4.18512
R9925 counter[0].n2 counter[0].n1 0.985115
R9926 net2.n14 net2.t0 315.034
R9927 net2.t1 net2.n14 265.769
R9928 net2 net2.t1 262.318
R9929 net2.n4 net2.t7 260.322
R9930 net2.n9 net2.t4 241.536
R9931 net2.n0 net2.t5 212.081
R9932 net2.n1 net2.t10 212.081
R9933 net2.n6 net2.t9 183.505
R9934 net2.n4 net2.t8 175.169
R9935 net2.n9 net2.t11 169.237
R9936 net2.n10 net2.n9 159.952
R9937 net2.n7 net2.n6 153.863
R9938 net2.n3 net2.n2 152.698
R9939 net2.n5 net2.n4 152
R9940 net2.n0 net2.t2 139.78
R9941 net2.n1 net2.t6 139.78
R9942 net2.n6 net2.t3 114.532
R9943 net2.n2 net2.n0 37.246
R9944 net2.n8 net2.n5 34.4715
R9945 net2.n2 net2.n1 24.1005
R9946 net2.n12 net2.n3 18.9449
R9947 net2.n13 net2.n12 14.916
R9948 net2.n11 net2.n10 13.8005
R9949 net2 net2.n7 10.8927
R9950 net2.n14 net2.n13 8.72777
R9951 net2.n8 net2 6.07742
R9952 net2.n10 net2 3.33963
R9953 net2.n10 net2 3.29747
R9954 net2 net2.n13 3.29747
R9955 net2.n11 net2.n8 3.19006
R9956 net2.n3 net2 1.97868
R9957 net2.n7 net2 1.97868
R9958 net2.n5 net2 1.55726
R9959 net2.n12 net2.n11 1.38649
R9960 net3.t5 net3.t6 395.01
R9961 net3 net3.t5 320.745
R9962 net3.n3 net3.t2 260.322
R9963 net3.n0 net3.t4 229.369
R9964 net3.n7 net3.t0 222.68
R9965 net3.n3 net3.t3 175.169
R9966 net3.n0 net3.t7 157.07
R9967 net3.n4 net3.n3 152
R9968 net3.n1 net3.n0 152
R9969 net3.n8 net3.t1 132.322
R9970 net3.n8 net3.n7 95.0273
R9971 net3.n5 net3 25.2581
R9972 net3.n5 net3 20.1696
R9973 net3.n7 net3.n6 12.7813
R9974 net3.n1 net3 12.0005
R9975 net3 net3.n4 11.2497
R9976 net3.n6 net3.n2 9.79203
R9977 net3.n6 net3.n5 5.9277
R9978 net3.n2 net3 4.53383
R9979 net3 net3.n8 2.70465
R9980 net3.n2 net3.n1 1.6005
R9981 net3.n4 net3 1.55726
R9982 clk.n3 clk.t2 184.768
R9983 clk.n2 clk.t1 184.768
R9984 clk.n1 clk.t3 184.768
R9985 clk.n0 clk.t0 184.768
R9986 clk.n4 clk.n3 171.375
R9987 clk.n3 clk.t6 146.208
R9988 clk.n2 clk.t5 146.208
R9989 clk.n1 clk.t7 146.208
R9990 clk.n0 clk.t4 146.208
R9991 clk.n3 clk.n2 40.6397
R9992 clk.n2 clk.n1 40.6397
R9993 clk.n1 clk.n0 40.6397
R9994 clk clk.n4 12.3171
R9995 clk.n4 clk 2.23542
R9996 _16_.n12 _16_.t0 339.418
R9997 _16_ _16_.t1 269.426
R9998 _16_.n1 _16_.t7 264.029
R9999 _16_ _16_.n5 241.976
R10000 _16_.n3 _16_.t3 241.536
R10001 _16_.n5 _16_.t8 241.536
R10002 _16_.n1 _16_.t2 206.19
R10003 _16_.n4 _16_.n3 171.332
R10004 _16_.n3 _16_.t9 169.237
R10005 _16_.n5 _16_.t6 169.237
R10006 _16_.n2 _16_.n1 160.96
R10007 _16_.n9 _16_.n8 153.165
R10008 _16_.n8 _16_.t5 144.548
R10009 _16_.n8 _16_.t4 128.482
R10010 _16_.n7 _16_.n2 21.45
R10011 _16_.n7 _16_.n6 16.7975
R10012 _16_.n10 _16_ 15.8161
R10013 _16_.n11 _16_.n10 14.0946
R10014 _16_ _16_.n0 11.2645
R10015 _16_ _16_.n9 9.55788
R10016 _16_.n6 _16_ 6.4005
R10017 _16_.n0 _16_ 6.1445
R10018 _16_.n2 _16_ 5.4405
R10019 _16_.n0 _16_ 4.63498
R10020 _16_.n4 _16_ 4.44132
R10021 _16_.n11 _16_ 4.3525
R10022 _16_.n13 _16_.n12 4.0914
R10023 _16_ _16_.n13 3.61789
R10024 _16_.n9 _16_ 3.29747
R10025 _16_.n13 _16_.n11 2.3045
R10026 _16_.n12 _16_ 1.74382
R10027 _16_.n6 _16_.n4 1.50638
R10028 _16_.n10 _16_.n7 1.38649
R10029 net6.n3 net6.t3 323.342
R10030 net6.n0 net6.t2 323.342
R10031 net6.n1 net6.t10 260.322
R10032 net6.n8 net6.t12 241.536
R10033 net6.n17 net6.t0 222.679
R10034 net6.n12 net6.t14 212.081
R10035 net6.n13 net6.t4 212.081
R10036 net6.n3 net6.t9 194.809
R10037 net6.n0 net6.t5 194.809
R10038 net6.n5 net6.t8 183.505
R10039 net6.n1 net6.t11 175.169
R10040 net6.n8 net6.t6 169.237
R10041 net6 net6.n3 158.133
R10042 net6 net6.n0 158.133
R10043 net6 net6.n8 157.555
R10044 net6.n15 net6.n14 155.52
R10045 net6.n6 net6.n5 153.863
R10046 net6.n2 net6.n1 152
R10047 net6.n12 net6.t7 139.78
R10048 net6.n13 net6.t15 139.78
R10049 net6.n18 net6.t1 129.078
R10050 net6.n5 net6.t13 114.532
R10051 net6.n18 net6.n17 96.7191
R10052 net6.n11 net6 55.2785
R10053 net6.n14 net6.n13 37.246
R10054 net6.n14 net6.n12 24.1005
R10055 net6.n10 net6.n9 21.4124
R10056 net6.n16 net6.n15 21.1949
R10057 net6.n4 net6.n2 20.043
R10058 net6.n7 net6.n6 15.2615
R10059 net6.n17 net6.n16 12.4213
R10060 net6.n9 net6 12.3175
R10061 net6.n16 net6.n11 8.09819
R10062 net6.n11 net6.n10 7.53948
R10063 net6.n4 net6 7.39885
R10064 net6 net6.n18 5.84085
R10065 net6.n15 net6 5.4405
R10066 net6.n9 net6 4.10616
R10067 net6.n7 net6.n4 2.60421
R10068 net6.n10 net6.n7 2.43577
R10069 net6.n6 net6 1.97868
R10070 net6.n2 net6 1.55726
R10071 counter[8].n0 counter[8].t0 368.521
R10072 counter[8].n1 counter[8].t1 216.155
R10073 counter[8].n1 counter[8] 78.8791
R10074 counter[8].n2 counter[8] 18.0834
R10075 counter[8] counter[8].n0 10.5563
R10076 counter[8].n0 counter[8] 5.48477
R10077 counter[8] counter[8].n2 4.18512
R10078 counter[8].n2 counter[8].n1 0.985115
R10079 counter[4].n0 counter[4].t0 368.521
R10080 counter[4].n1 counter[4].t1 216.155
R10081 counter[4].n1 counter[4] 78.8791
R10082 counter[4].n2 counter[4] 18.7251
R10083 counter[4] counter[4].n0 10.5563
R10084 counter[4].n0 counter[4] 5.48477
R10085 counter[4] counter[4].n2 4.18512
R10086 counter[4].n2 counter[4].n1 0.985115
R10087 counter[5].n0 counter[5].t0 368.521
R10088 counter[5].n1 counter[5].t1 216.155
R10089 counter[5].n1 counter[5] 78.8791
R10090 counter[5].n2 counter[5] 18.0287
R10091 counter[5] counter[5].n0 10.5563
R10092 counter[5].n0 counter[5] 5.48477
R10093 counter[5] counter[5].n2 4.18512
R10094 counter[5].n2 counter[5].n1 0.985115
R10095 counter[1].n0 counter[1].t0 368.521
R10096 counter[1].n1 counter[1].t1 216.155
R10097 counter[1].n1 counter[1] 78.8791
R10098 counter[1].n2 counter[1] 18.0287
R10099 counter[1] counter[1].n0 10.5563
R10100 counter[1].n0 counter[1] 5.48477
R10101 counter[1] counter[1].n2 4.18512
R10102 counter[1].n2 counter[1].n1 0.985115
R10103 counter[7].n0 counter[7].t0 368.521
R10104 counter[7].n1 counter[7].t1 216.155
R10105 counter[7].n1 counter[7] 78.8791
R10106 counter[7].n2 counter[7] 19.5465
R10107 counter[7] counter[7].n0 10.5563
R10108 counter[7].n0 counter[7] 5.48477
R10109 counter[7] counter[7].n2 4.18512
R10110 counter[7].n2 counter[7].n1 0.985115
R10111 enable.n0 enable.t0 260.322
R10112 enable.n0 enable.t1 175.169
R10113 enable.n1 enable.n0 153.13
R10114 enable.n1 enable 9.86591
R10115 enable enable.n1 3.2005
R10116 counter[9].n0 counter[9].t0 368.521
R10117 counter[9].n2 counter[9].t1 216.155
R10118 counter[9] counter[9].n2 78.8791
R10119 counter[9].n1 counter[9] 22.9394
R10120 counter[9].n1 counter[9].n0 6.52665
R10121 counter[9].n0 counter[9] 5.48477
R10122 counter[9].n2 counter[9] 5.16973
R10123 counter[9] counter[9].n1 4.03013
C0 clknet_1_0__leaf_clk a_2401_4399# 0.020113f
C1 a_3979_4943# a_4779_5161# 2.3e-20
C2 _11_ a_4811_3861# 1.58e-19
C3 a_4399_5175# a_4495_5175# 0.310858f
C4 a_5814_4399# a_7005_3311# 1.26e-19
C5 _18_ _16_ 0.283975f
C6 _11_ a_7216_3311# 4.03e-21
C7 net8 a_3831_3105# 9.57e-20
C8 net9 a_4995_4399# 0.063508f
C9 a_4520_4373# a_4220_3829# 8.74e-19
C10 _21_ _06_ 0.224771f
C11 net2 a_2302_7937# 4.89e-19
C12 a_4259_3311# a_4341_3311# 0.005167f
C13 _11_ a_5077_4721# 4.38e-19
C14 _16_ a_3601_3855# 0.010038f
C15 _17_ a_5162_4943# 0.002153f
C16 net5 a_3849_2388# 0.233889f
C17 _12_ _11_ 0.214271f
C18 a_2849_7497# a_2678_7119# 0.001229f
C19 a_3831_3339# VPWR 0.254188f
C20 clknet_0_clk a_4714_5309# 1.49e-19
C21 a_1683_3861# a_2471_2741# 3.4e-19
C22 net6 a_1849_3861# 1.26e-19
C23 net3 _13_ 0.031667f
C24 _17_ a_4811_3861# 1.12e-20
C25 a_4329_5461# a_4977_3861# 4.98e-20
C26 a_2849_7663# VPWR 0.080219f
C27 net9 a_7641_3311# 6.87e-19
C28 a_1845_5461# a_1849_3861# 1.82e-21
C29 a_3215_3829# net5 0.001034f
C30 a_7723_2741# VPWR 0.230416f
C31 _11_ _14_ 0.007676f
C32 _17_ a_5077_4721# 4.44e-20
C33 a_4329_5461# _22_ 7.51e-19
C34 a_1915_7815# a_1915_7351# 0.025128f
C35 net7 a_4520_4373# 0.003377f
C36 a_4454_4649# a_4995_4399# 4.72e-19
C37 _15_ a_5376_4233# 0.002542f
C38 a_6817_3311# a_7171_2767# 1.65e-19
C39 _24_ a_7185_3677# 7.21e-19
C40 _19_ _23_ 2.58e-20
C41 net7 clk 6.87e-19
C42 a_2295_7637# a_2695_6575# 4.52e-21
C43 a_6817_3311# a_7258_3423# 0.118966f
C44 _11_ a_2614_2883# 1e-19
C45 VPWR enable 0.196543f
C46 net2 a_2295_7337# 3.07e-19
C47 _16_ a_5179_3311# 1.25e-20
C48 net3 counter[2] 7.38e-19
C49 net8 a_4287_4399# 0.057781f
C50 a_1875_8207# a_2125_8207# 0.025037f
C51 _23_ a_7619_5162# 6.47e-19
C52 a_6375_5309# _25_ 1.87e-19
C53 net7 a_5891_3133# 0.006602f
C54 _11_ _20_ 0.174111f
C55 a_3099_4765# a_3183_4765# 0.008508f
C56 a_2566_3423# a_2313_3311# 3.39e-19
C57 a_2991_3579# a_4259_3311# 3.71e-21
C58 a_1683_3861# a_1505_3855# 5.87e-19
C59 a_2674_4765# a_1959_3311# 5.5e-20
C60 a_2235_4399# a_2398_3677# 8.98e-19
C61 _23_ a_6651_3311# 0.029061f
C62 net10 a_8109_2767# 0.003077f
C63 clknet_1_0__leaf_clk a_2991_3579# 1.1e-19
C64 clknet_1_1__leaf_clk a_7258_3423# 2.7e-19
C65 a_2217_3855# VPWR 0.003619f
C66 a_2991_3579# a_2840_3087# 0.001062f
C67 _16_ a_2715_3829# 7.03e-19
C68 a_2678_8029# a_2849_7663# 0.001229f
C69 a_7345_2388# counter[8] 6.92e-19
C70 a_2253_8029# clknet_1_0__leaf_clk 7.44e-19
C71 net6 a_3099_4765# 0.021756f
C72 _17_ _20_ 1.89e-19
C73 a_5814_4399# _09_ 3.55e-20
C74 net10 a_7683_3579# 0.008159f
C75 _15_ a_7171_2767# 0.038186f
C76 a_7077_2767# a_7723_2741# 0.016298f
C77 a_2561_9514# a_2502_7637# 2.02e-20
C78 net1 a_2295_7637# 0.003904f
C79 _23_ a_7683_3829# 1.75e-20
C80 a_3831_3105# a_3917_3105# 0.006584f
C81 counter[4] counter[5] 0.068962f
C82 _21_ VPWR 0.492491f
C83 a_4779_5161# a_5165_3855# 6.17e-21
C84 clknet_0_clk a_3267_4667# 3.43e-19
C85 _12_ a_2849_7497# 0.023132f
C86 a_2295_7337# _11_ 9.54e-19
C87 _15_ a_7258_3423# 0.002208f
C88 _03_ VPWR 0.393273f
C89 a_2302_7241# a_2695_6575# 0.011211f
C90 _05_ a_6375_5309# 1.27e-19
C91 _11_ a_2673_4233# 6.78e-19
C92 net4 a_2566_3423# 0.007782f
C93 _11_ a_6375_5309# 0.087773f
C94 a_6817_3861# a_7599_3855# 6.32e-19
C95 a_5179_3311# a_5533_3311# 0.062224f
C96 a_4399_5175# _21_ 0.001295f
C97 net3 a_2471_2741# 0.002183f
C98 a_5786_3423# a_6211_3579# 1.28e-19
C99 _05_ a_5814_4399# 0.003024f
C100 a_5345_3311# a_6043_3677# 0.193199f
C101 net4 a_3831_3105# 0.083888f
C102 _11_ a_5814_4399# 0.049204f
C103 a_7753_2767# VPWR 0.283149f
C104 net9 a_5997_3133# 6.77e-19
C105 a_4786_5065# net6 0.001918f
C106 _17_ a_6375_5309# 0.139841f
C107 a_2302_7937# a_2849_7497# 4.5e-20
C108 _00_ a_2695_6575# 5.19e-20
C109 clknet_1_0__leaf_clk _01_ 0.05158f
C110 a_4977_3861# a_5345_3311# 1.17e-19
C111 a_5135_5309# VPWR 0.002269f
C112 a_4811_3861# a_5786_3423# 3.92e-19
C113 a_5418_3829# a_5179_3311# 1.62e-19
C114 a_6211_3579# a_6169_3311# 7.84e-20
C115 clknet_0_clk a_4779_5161# 0.043419f
C116 VPWR counter[6] 0.462317f
C117 net1 a_2302_7241# 0.00338f
C118 _22_ a_5345_3311# 0.02378f
C119 a_1849_3861# VPWR 0.341027f
C120 a_7090_3677# VPWR 0.248502f
C121 _07_ a_4767_3463# 1.81e-19
C122 _11_ a_3145_6825# 0.002858f
C123 _17_ a_5814_4399# 0.002308f
C124 a_1959_3311# a_3831_3339# 7.98e-21
C125 a_6817_3861# a_6817_3311# 0.027195f
C126 a_6651_3861# a_7258_3423# 1.99e-20
C127 a_4495_5175# a_4714_5309# 0.006169f
C128 _03_ a_2823_3677# 0.001345f
C129 net8 net10 1.02e-19
C130 clknet_1_0__leaf_clk a_2800_4399# 3.26e-19
C131 _11_ a_6719_3133# 0.006396f
C132 net2 _16_ 5.41e-20
C133 net7 a_5618_3677# 0.005696f
C134 net3 a_2011_7351# 0.006429f
C135 net2 _10_ 0.006086f
C136 a_4786_5065# _06_ 1.63e-21
C137 net6 a_4767_3463# 0.173962f
C138 net4 a_4349_4175# 7.88e-20
C139 net6 a_2235_4399# 0.006287f
C140 net7 a_7289_5309# 1.83e-19
C141 net1 _00_ 0.056053f
C142 a_1845_5461# a_2235_4399# 5.49e-20
C143 clknet_1_0__leaf_clk clknet_0_clk 0.004956f
C144 net7 a_7599_3677# 3.05e-20
C145 a_2842_4511# a_3099_4765# 0.036838f
C146 a_2431_7497# a_2230_7485# 4.67e-20
C147 a_2401_4399# net8 0.001542f
C148 _18_ a_4349_4175# 9.76e-19
C149 a_2302_7241# a_2651_7485# 2.36e-19
C150 clknet_1_1__leaf_clk a_6817_3861# 0.026802f
C151 a_2295_7337# a_2849_7497# 0.057611f
C152 net7 a_4220_3829# 0.142058f
C153 a_2011_7351# a_2253_7119# 0.008508f
C154 a_2125_3311# a_2745_2388# 7.04e-21
C155 a_4779_5161# clknet_1_1__leaf_clk 0.228247f
C156 net1 a_2317_6575# 0.00162f
C157 _14_ a_3215_3829# 1.74e-20
C158 _05_ _16_ 0.001611f
C159 net7 a_5213_4664# 1.85e-20
C160 a_5213_4664# a_5436_4399# 3.74e-19
C161 _18_ a_4287_4399# 0.002103f
C162 a_7683_3829# a_7641_4233# 7.84e-20
C163 a_7090_3855# net10 3.33e-19
C164 VPWR counter[1] 0.340796f
C165 a_5077_4721# a_4995_4399# 2.78e-19
C166 _11_ _16_ 0.223435f
C167 _20_ a_5786_3423# 6.25e-20
C168 a_2122_3855# a_2398_3677# 4.47e-19
C169 a_2715_3829# a_2566_3423# 0.001344f
C170 a_2547_3855# a_2125_3311# 0.003824f
C171 net8 a_4341_3311# 4.38e-20
C172 _06_ a_4767_3463# 2.49e-19
C173 _10_ _11_ 0.033565f
C174 a_7090_3677# a_7077_2767# 2.47e-19
C175 _15_ a_6817_3861# 0.058771f
C176 _19_ a_5250_3855# 6.46e-21
C177 a_3099_4765# VPWR 0.169689f
C178 a_4779_5161# _15_ 3.85e-20
C179 a_1915_7815# _12_ 6.08e-20
C180 net8 a_5843_3829# 0.084103f
C181 _17_ _16_ 0.048058f
C182 net9 a_6211_3579# 0.115737f
C183 clknet_1_1__leaf_clk a_4259_3311# 2.42e-19
C184 a_6127_3677# VPWR 0.004788f
C185 net6 a_3245_3855# 0.007899f
C186 net2 counter[0] 0.010591f
C187 a_1959_3311# _03_ 0.095111f
C188 net9 a_4811_3861# 5.55e-19
C189 net9 a_7216_3311# 0.002793f
C190 _15_ a_4259_3311# 0.080244f
C191 a_7258_3829# VPWR 0.182123f
C192 net9 a_5077_4721# 0.004319f
C193 a_2125_8207# a_2295_7637# 5.23e-20
C194 a_1915_7815# a_2302_7937# 0.034054f
C195 _11_ a_5533_3311# 0.016192f
C196 _24_ a_7005_3855# 4.8e-19
C197 a_5814_4399# a_5786_3423# 2.72e-20
C198 a_6375_5309# a_6651_5309# 0.00119f
C199 a_4786_5065# VPWR 0.321592f
C200 a_5149_4721# a_5618_3677# 5.18e-21
C201 a_6651_3861# a_6817_3861# 0.970499f
C202 _15_ a_2840_3087# 8.81e-20
C203 a_3099_4765# a_2823_3677# 2.6e-20
C204 _23_ a_7185_3677# 8.32e-19
C205 a_2235_4399# a_2842_4511# 0.136461f
C206 a_1915_7351# _12_ 0.027335f
C207 _04_ a_2401_4399# 0.215918f
C208 net3 a_2235_6575# 0.079675f
C209 _05_ a_5418_3829# 8.7e-19
C210 _14_ _02_ 0.166596f
C211 a_4399_5175# a_4786_5065# 0.034054f
C212 clknet_1_0__leaf_clk a_2674_4765# 0.002436f
C213 a_4495_5175# a_4779_5161# 0.030894f
C214 _11_ a_5418_3829# 7.26e-20
C215 net8 a_6427_2741# 0.004343f
C216 a_2674_4765# a_2840_3087# 4.44e-21
C217 a_4454_4649# a_4811_3861# 4.26e-19
C218 net2 a_2502_7637# 1.88e-19
C219 a_1849_3861# a_1959_3311# 0.010101f
C220 a_1683_3861# a_2125_3311# 2.24e-19
C221 a_5149_4721# a_5213_4664# 0.266837f
C222 net6 a_4737_4943# 1.73e-19
C223 a_4767_3463# VPWR 0.226919f
C224 net6 a_2122_3855# 6.57e-20
C225 a_2235_4399# VPWR 0.6434f
C226 clknet_0_clk a_5333_5321# 0.004448f
C227 net4 a_2401_4399# 0.34974f
C228 a_4329_5461# a_5250_3855# 5.07e-19
C229 _17_ a_5418_3829# 1.03e-20
C230 net7 a_5149_4721# 6.37e-20
C231 a_2011_7637# a_2011_7351# 0.015931f
C232 a_1845_5461# a_2122_3855# 7.35e-19
C233 a_3389_3105# VPWR 3.83e-21
C234 net10 counter[8] 0.009948f
C235 a_5149_4721# a_5436_4399# 3.14e-19
C236 net9 _20_ 1.35e-20
C237 a_7090_3677# a_7171_2767# 7.6e-20
C238 _18_ a_2401_4399# 8.49e-20
C239 _24_ a_7599_3677# 8.56e-19
C240 _11_ a_2566_3423# 0.004479f
C241 _22_ a_5891_3133# 0.002353f
C242 a_6817_3311# a_7683_3579# 0.034054f
C243 a_7258_3423# a_7090_3677# 0.239923f
C244 _11_ a_3831_3105# 0.002917f
C245 net8 a_5165_3855# 0.005878f
C246 net2 a_2502_7396# 3.35e-21
C247 _16_ a_5786_3423# 8.82e-22
C248 _14_ net5 0.258421f
C249 a_1875_8207# a_2011_7637# 7.31e-19
C250 a_3799_4943# VPWR 0.252612f
C251 _00_ a_2125_8207# 0.07841f
C252 a_4454_4649# _20_ 4.3e-20
C253 net7 a_6623_3133# 6.49e-19
C254 net7 _24_ 2.68e-19
C255 a_3267_4667# _21_ 1.76e-19
C256 a_2398_3677# a_2493_3677# 0.007724f
C257 _16_ a_3849_2388# 3.59e-21
C258 a_3831_3339# a_4259_3311# 0.00155f
C259 a_2566_3423# a_2907_3677# 9.73e-19
C260 a_2125_3311# a_2524_3311# 0.001351f
C261 clknet_1_1__leaf_clk a_5333_5321# 3.41e-20
C262 _19_ net6 0.04173f
C263 _04_ a_2991_3579# 7.11e-19
C264 net8 a_7599_3855# 2.29e-20
C265 a_2235_4399# a_2823_3677# 0.001131f
C266 a_2230_7485# VPWR 3.44e-19
C267 a_1915_7351# a_2295_7337# 0.048748f
C268 clknet_1_1__leaf_clk a_7683_3579# 1.1e-19
C269 a_3245_3855# VPWR 0.261491f
C270 clknet_0_clk a_5871_5162# 0.012442f
C271 _08_ a_7005_3855# 0.134213f
C272 net5 a_2614_2883# 3.95e-20
C273 _16_ a_3215_3829# 0.243866f
C274 _18_ a_3979_4943# 0.190808f
C275 a_8265_2388# counter[8] 0.111116f
C276 a_6425_2388# counter[7] 8.38e-19
C277 a_2849_7663# clknet_1_0__leaf_clk 0.012004f
C278 a_2589_4399# a_1683_3861# 3.23e-19
C279 a_5418_3829# a_5801_4233# 4.67e-20
C280 net5 _20_ 8.42e-21
C281 clknet_0_clk net8 8.45e-19
C282 a_5814_4399# net9 0.111158f
C283 net1 a_2431_7663# 0.002441f
C284 net6 a_7619_5162# 1.17e-21
C285 net11 counter[7] 1.31e-19
C286 net4 a_2991_3579# 0.020834f
C287 net3 a_2125_3311# 0.00115f
C288 _22_ counter[7] 1.31e-20
C289 clknet_0_clk a_7199_4943# 1.5e-20
C290 net6 a_6651_3311# 5.6e-22
C291 _16_ a_4995_4399# 0.036674f
C292 _19_ _06_ 7.42e-21
C293 a_2431_7663# a_2230_7663# 4.67e-20
C294 a_2502_7637# a_2651_7663# 0.005525f
C295 a_2401_4399# a_2715_3829# 0.003783f
C296 a_1875_8207# a_2011_7351# 6.59e-20
C297 _11_ a_4287_4399# 3.73e-19
C298 a_5786_3423# a_5533_3311# 3.39e-19
C299 a_4779_5161# _21_ 8.19e-20
C300 net8 a_6817_3311# 1.04e-19
C301 _11_ a_2769_4765# 0.00121f
C302 a_3917_3339# VPWR 0.00273f
C303 a_7199_4943# a_6817_3311# 3.03e-21
C304 a_4915_5321# net6 0.001158f
C305 clknet_1_1__leaf_clk a_5871_5162# 0.035969f
C306 a_1457_2388# VPWR 0.25802f
C307 a_4341_3311# counter[4] 4.37e-20
C308 a_5250_3855# a_5345_3311# 8.92e-19
C309 a_5843_3829# a_5179_3311# 0.002274f
C310 a_4737_4943# VPWR 0.004852f
C311 a_4977_3861# a_5618_3677# 7.62e-19
C312 clknet_1_0__leaf_clk a_2217_3855# 0.001355f
C313 clknet_0_clk a_4986_5220# 0.004436f
C314 _17_ a_4287_4399# 0.060488f
C315 _22_ a_5618_3677# 0.002895f
C316 clknet_1_1__leaf_clk net8 0.073766f
C317 a_7515_3677# VPWR 0.215619f
C318 net1 a_2431_7497# 0.001727f
C319 a_2122_3855# VPWR 0.259474f
C320 a_4811_3861# a_5505_2388# 1.7e-21
C321 _11_ a_2389_6575# 2.12e-19
C322 _08_ a_7599_3677# 1.22e-19
C323 _21_ a_4259_3311# 0.087922f
C324 a_7090_3855# a_6817_3311# 1.54e-19
C325 a_6817_3861# a_7090_3677# 1.54e-19
C326 _04_ a_2800_4399# 2.91e-19
C327 a_7258_3829# a_7258_3423# 0.012451f
C328 clknet_1_1__leaf_clk a_7199_4943# 3.65e-19
C329 a_2235_4399# a_1959_3311# 2.82e-20
C330 a_5213_4664# a_4977_3861# 0.003413f
C331 net7 a_6043_3677# 0.040127f
C332 net3 a_2302_7241# 0.005586f
C333 a_4329_5461# net6 8.49e-19
C334 clknet_1_1__leaf_clk a_5744_3311# 4.82e-19
C335 clknet_1_0__leaf_clk _03_ 0.00668f
C336 _16_ _02_ 3.22e-20
C337 a_7019_4943# a_5814_4399# 0.010673f
C338 _03_ a_2840_3087# 9.33e-19
C339 a_5213_4664# _22_ 0.155189f
C340 a_4915_5321# _06_ 4.29e-19
C341 net9 _16_ 0.243936f
C342 _15_ net8 0.048599f
C343 net7 a_6425_2388# 4.41e-19
C344 net7 _08_ 1.97e-19
C345 net10 _09_ 0.081678f
C346 _15_ a_7199_4943# 0.001357f
C347 net7 net11 2.47e-20
C348 net7 a_4977_3861# 0.456298f
C349 clknet_1_1__leaf_clk a_7090_3855# 0.001015f
C350 a_2502_7396# a_2849_7497# 0.037333f
C351 a_3267_4667# a_3099_4765# 0.310858f
C352 a_2295_7337# a_2678_7119# 0.001632f
C353 a_2431_7497# a_2651_7485# 4.62e-19
C354 a_2302_7241# a_2253_7119# 4.04e-19
C355 a_2674_4765# net8 4.11e-20
C356 net1 a_1845_5461# 0.001584f
C357 a_5345_3311# a_5599_2741# 0.002313f
C358 a_4986_5220# clknet_1_1__leaf_clk 4.65e-20
C359 net7 _22_ 0.179589f
C360 a_7723_2741# a_8109_2767# 0.006406f
C361 a_2547_3855# a_2398_3677# 0.001152f
C362 _22_ a_5436_4399# 0.006962f
C363 a_2715_3829# a_2991_3579# 0.007214f
C364 a_4443_4175# a_4349_3855# 1.26e-19
C365 _19_ VPWR 0.197759f
C366 a_7515_3855# net10 0.00375f
C367 net8 a_4929_3311# 0.002158f
C368 _20_ a_6211_3579# 3.47e-20
C369 a_4329_5461# _06_ 1.96e-20
C370 _23_ a_7005_3855# 0.014354f
C371 a_4454_4649# _16_ 0.029136f
C372 clknet_1_0__leaf_clk a_1849_3861# 0.158653f
C373 a_7683_3579# a_7723_2741# 0.005283f
C374 _15_ a_7090_3855# 0.001174f
C375 a_7515_3677# a_7077_2767# 2.58e-19
C376 _23_ counter[7] 0.004833f
C377 net3 a_2317_6575# 1.25e-19
C378 a_4986_5220# _15_ 1.61e-21
C379 _11_ net10 0.36244f
C380 a_4399_5175# _19_ 0.065395f
C381 a_1875_8207# a_2235_6575# 2.44e-21
C382 a_2302_7937# _12_ 0.003541f
C383 a_7619_5162# VPWR 0.28996f
C384 clknet_0_clk _18_ 0.002702f
C385 net8 a_6651_3861# 0.001229f
C386 a_6651_3311# VPWR 0.667506f
C387 net9 a_5533_3311# 1.61e-19
C388 _16_ net5 0.096932f
C389 clknet_1_1__leaf_clk _04_ 1.67e-21
C390 a_4495_5175# net8 1.55e-19
C391 net6 a_4349_3855# 0.044713f
C392 a_7199_4943# a_6651_3861# 6.06e-21
C393 net9 a_7345_2388# 0.202772f
C394 _11_ a_2401_4399# 0.082924f
C395 _13_ a_2589_4399# 5.97e-20
C396 _14_ a_2614_2883# 0.089653f
C397 net9 a_5418_3829# 2.05e-20
C398 _07_ a_5345_3311# 0.195848f
C399 a_7683_3829# VPWR 0.48745f
C400 a_2125_3311# a_2471_2741# 0.010515f
C401 _15_ _04_ 3.75e-19
C402 a_2011_7637# a_2295_7637# 0.032244f
C403 a_4915_5321# VPWR 0.191062f
C404 _11_ a_4341_3311# 0.002312f
C405 a_5814_4399# a_6211_3579# 0.001883f
C406 _15_ a_3917_3105# 0.001523f
C407 a_6651_3861# a_7090_3855# 0.273138f
C408 a_2695_6575# VPWR 0.292813f
C409 a_6817_3861# a_7258_3829# 0.118966f
C410 a_1849_3861# a_2631_3855# 6.32e-19
C411 _17_ a_2401_4399# 9.29e-21
C412 _06_ a_4349_3855# 2.02e-19
C413 a_2235_4399# a_3267_4667# 0.048608f
C414 _04_ a_2674_4765# 0.01404f
C415 a_2295_7337# _12_ 0.062549f
C416 a_4399_5175# a_4915_5321# 1.28e-19
C417 a_3979_4943# _05_ 4.91e-20
C418 net6 a_5345_3311# 0.045685f
C419 _18_ clknet_1_1__leaf_clk 3.06e-19
C420 clknet_1_0__leaf_clk a_3099_4765# 6.75e-21
C421 a_4779_5161# a_4786_5065# 0.961627f
C422 a_5149_4721# a_4977_3861# 1.08e-19
C423 _11_ a_5843_3829# 1.18e-19
C424 clknet_0_clk a_5179_3311# 1.17e-21
C425 a_4767_3463# a_5001_3311# 0.005167f
C426 _11_ a_3979_4943# 0.001495f
C427 a_2122_3855# a_1959_3311# 4.57e-19
C428 a_1683_3861# a_2398_3677# 0.001041f
C429 a_5149_4721# _22_ 0.019192f
C430 a_2290_3829# _03_ 0.009555f
C431 _15_ net4 0.003757f
C432 a_4329_5461# VPWR 1.29479f
C433 clknet_1_1__leaf_clk a_3601_3855# 8.24e-20
C434 a_6651_3311# a_7077_2767# 9.12e-19
C435 net7 _23_ 0.074369f
C436 a_2493_3677# VPWR 0.005794f
C437 _09_ a_6427_2741# 1.89e-19
C438 clknet_0_clk a_6457_5309# 5.18e-20
C439 net6 a_2547_3855# 5.09e-19
C440 net4 a_2674_4765# 0.034877f
C441 _17_ a_5843_3829# 4.35e-22
C442 _18_ _15_ 0.045245f
C443 a_5179_3311# a_6817_3311# 8.05e-21
C444 a_2295_7637# a_2011_7351# 9.64e-20
C445 a_2302_7937# a_2295_7337# 3.36e-19
C446 a_2011_7637# a_2302_7241# 1.53e-19
C447 a_2936_2767# VPWR 0.012117f
C448 _17_ a_3979_4943# 0.043588f
C449 _24_ _08_ 0.423487f
C450 net1 VPWR 1.47718f
C451 a_4329_5461# a_4399_5175# 0.022122f
C452 a_4779_5161# a_4767_3463# 8.37e-20
C453 a_7683_3579# a_7753_2767# 1.25e-19
C454 _24_ net11 0.002712f
C455 _18_ a_2674_4765# 5.13e-20
C456 _12_ a_3145_6825# 0.001754f
C457 _11_ a_2991_3579# 0.065594f
C458 _22_ a_6623_3133# 0.001961f
C459 a_6817_3311# a_7005_3311# 0.097994f
C460 a_7258_3423# a_7515_3677# 0.036838f
C461 a_1849_3861# a_2290_3829# 0.127288f
C462 _24_ _22_ 0.01067f
C463 _11_ a_6427_2741# 0.19543f
C464 a_2230_7663# VPWR 4.59e-19
C465 clknet_1_1__leaf_clk a_5179_3311# 0.319108f
C466 net2 _01_ 9.85e-20
C467 a_1875_8207# a_2295_7637# 0.001828f
C468 _00_ a_2011_7637# 0.001635f
C469 net7 a_6825_3133# 6.33e-20
C470 net8 _21_ 0.333812f
C471 a_4259_3311# a_4767_3463# 0.017774f
C472 a_2566_3423# net5 0.001073f
C473 a_2398_3677# a_2524_3311# 0.005525f
C474 a_2651_7485# VPWR 0.002269f
C475 clknet_1_1__leaf_clk a_7005_3311# 6.27e-19
C476 a_2041_4649# a_2235_4399# 5.05e-19
C477 a_4349_3855# VPWR 0.206364f
C478 a_2011_7351# a_2302_7241# 0.192341f
C479 clknet_1_0__leaf_clk a_2235_4399# 0.245743f
C480 _15_ a_5179_3311# 4.49e-20
C481 net5 a_3831_3105# 0.201023f
C482 _16_ a_4811_3861# 1.57e-19
C483 _18_ a_4495_5175# 2.33e-19
C484 a_3799_4943# a_4779_5161# 6.46e-21
C485 a_7939_2223# counter[7] 3.7e-19
C486 a_2235_4399# a_2840_3087# 4.07e-21
C487 a_5505_2388# counter[5] 0.1107f
C488 a_5599_2741# a_5891_3133# 0.001675f
C489 a_2745_2388# counter[3] 4.98e-19
C490 a_5843_3829# a_5801_4233# 7.84e-20
C491 net1 a_2678_8029# 4.16e-19
C492 a_7599_3855# _09_ 1.2e-19
C493 a_4399_5175# a_4349_3855# 2.76e-21
C494 _19_ a_4714_5309# 1.38e-19
C495 _15_ counter[4] 9.07e-20
C496 _15_ a_7005_3311# 0.005742f
C497 _12_ _10_ 0.002721f
C498 _01_ _11_ 0.20957f
C499 _15_ a_2715_3829# 1.37e-19
C500 net4 a_3831_3339# 4.87e-19
C501 net3 a_2398_3677# 3.32e-20
C502 net6 a_1683_3861# 1.88e-19
C503 net8 counter[6] 0.079257f
C504 a_7515_3855# a_7599_3855# 0.008508f
C505 a_5618_3677# a_5713_3677# 0.007724f
C506 a_6375_5309# a_5814_4399# 0.010774f
C507 _16_ _14_ 0.202586f
C508 a_4986_5220# _21_ 0.0043f
C509 a_2674_4765# a_2715_3829# 0.004197f
C510 a_2842_4511# a_2547_3855# 0.004484f
C511 _18_ a_3831_3339# 1.7e-19
C512 a_4454_4649# a_4287_4399# 0.046138f
C513 _11_ a_2800_4399# 0.003523f
C514 a_5533_3311# a_5505_2388# 7.39e-20
C515 _09_ a_7941_3087# 0.002954f
C516 a_5345_3311# VPWR 0.323392f
C517 net6 a_2037_3855# 1.35e-20
C518 a_6043_3677# a_6425_2388# 3.85e-20
C519 a_2561_9514# enable 0.231636f
C520 a_2745_2388# VPWR 0.317416f
C521 _16_ a_2614_2883# 0.146025f
C522 _09_ a_6817_3311# 0.413296f
C523 a_6545_5309# VPWR 0.002069f
C524 a_5843_3829# a_5786_3423# 6.84e-19
C525 clknet_1_0__leaf_clk a_2230_7485# 0.001172f
C526 a_5675_3855# a_5345_3311# 1.5e-19
C527 a_6651_3311# a_7258_3423# 0.141453f
C528 clknet_0_clk _05_ 0.067252f
C529 a_2547_3855# VPWR 0.228175f
C530 a_7185_3677# VPWR 0.002923f
C531 net6 a_4520_4373# 0.016498f
C532 _16_ _20_ 0.011071f
C533 _22_ a_6043_3677# 6.29e-19
C534 _08_ a_4977_3861# 8.29e-20
C535 _11_ clknet_0_clk 0.042991f
C536 _22_ a_6425_2388# 2.78e-19
C537 a_7723_2741# counter[8] 0.001844f
C538 _23_ _24_ 0.206353f
C539 a_1875_8207# _00_ 0.167554f
C540 a_1959_3311# a_2493_3677# 0.002698f
C541 a_4811_3861# a_5418_3829# 0.136009f
C542 a_7090_3855# a_7090_3677# 0.013839f
C543 a_4786_5065# a_5333_5321# 0.095025f
C544 _08_ _22_ 1.19e-20
C545 a_6817_3861# a_7515_3677# 1.3e-19
C546 a_4915_5321# a_4714_5309# 4.67e-20
C547 a_4986_5220# a_5135_5309# 0.005525f
C548 a_7515_3855# a_6817_3311# 1.3e-19
C549 _03_ a_2313_3311# 0.13856f
C550 net6 clk 2.01e-20
C551 _11_ a_4069_5309# 1.46e-19
C552 _22_ a_4977_3861# 0.015364f
C553 net3 a_2431_7497# 2.06e-19
C554 clknet_1_1__leaf_clk _09_ 0.003413f
C555 net7 a_5713_3677# 5.23e-19
C556 a_5213_4664# a_5250_3855# 1.41e-19
C557 _22_ net11 1.96e-19
C558 _03_ a_3917_3105# 5.07e-20
C559 _11_ a_6817_3311# 7.13e-19
C560 clknet_0_clk _17_ 0.029087f
C561 _15_ _25_ 0.003323f
C562 a_4520_4373# _06_ 0.004838f
C563 clknet_1_1__leaf_clk a_7515_3855# 1.84e-19
C564 net7 a_5250_3855# 0.034093f
C565 net9 net10 0.022804f
C566 a_2302_7241# a_2235_6575# 1.58e-19
C567 a_2502_7396# a_2678_7119# 0.007724f
C568 _17_ a_4069_5309# 7.93e-19
C569 a_2431_7497# a_2253_7119# 9.73e-19
C570 _01_ a_2849_7497# 0.121379f
C571 a_2295_7337# _10_ 0.011255f
C572 _15_ _09_ 0.030214f
C573 a_3099_4765# net8 3.5e-19
C574 net4 _03_ 0.031989f
C575 a_5618_3677# a_5599_2741# 1.83e-19
C576 _05_ clknet_1_1__leaf_clk 0.143201f
C577 a_2125_8207# VPWR 0.262851f
C578 _11_ clknet_1_1__leaf_clk 0.367667f
C579 a_2547_3855# a_2823_3677# 5.06e-19
C580 a_3215_3829# a_2991_3579# 0.002391f
C581 a_2398_3677# counter[2] 1.99e-20
C582 _20_ a_5533_3311# 5.09e-20
C583 _18_ _21_ 0.005609f
C584 _04_ a_1849_3861# 0.011144f
C585 clknet_1_0__leaf_clk a_2122_3855# 0.032164f
C586 a_2235_4399# a_2290_3829# 0.002941f
C587 a_5814_4399# _16_ 0.001016f
C588 _15_ a_7515_3855# 2.78e-19
C589 _05_ _15_ 9.02e-20
C590 net3 a_1845_5461# 0.011213f
C591 a_4779_5161# _19_ 0.074331f
C592 _11_ _15_ 1.40124f
C593 _17_ clknet_1_1__leaf_clk 0.044595f
C594 a_2502_7637# _12_ 5.69e-20
C595 a_7005_3855# a_7185_3855# 0.001229f
C596 net8 a_7258_3829# 8.61e-20
C597 a_1683_3861# VPWR 0.684183f
C598 a_7199_4943# a_7258_3829# 2.48e-20
C599 a_4786_5065# net8 4.93e-19
C600 a_2235_6575# a_2317_6575# 0.005167f
C601 _25_ a_6651_3861# 1.01e-19
C602 _14_ a_2566_3423# 1.1e-19
C603 net4 a_1849_3861# 0.002039f
C604 net6 a_7005_3855# 3.93e-20
C605 net7 a_5599_2741# 0.212284f
C606 _14_ a_3831_3105# 9.06e-21
C607 a_6817_3861# a_6651_3311# 2.64e-19
C608 _11_ a_2674_4765# 0.054008f
C609 a_2401_4399# a_4454_4649# 1.23e-20
C610 a_6651_3861# _09_ 1.11e-19
C611 _23_ a_6043_3677# 0.001187f
C612 net9 a_5843_3829# 0.007609f
C613 _17_ _15_ 0.083602f
C614 a_2398_3677# a_2471_2741# 3.53e-19
C615 _23_ a_6425_2388# 2.99e-20
C616 _07_ a_5618_3677# 0.008539f
C617 a_2566_3423# a_2614_2883# 5.83e-19
C618 a_2037_3855# VPWR 0.075425f
C619 a_2011_7637# a_2431_7663# 0.036838f
C620 a_2302_7937# a_2502_7637# 0.074815f
C621 _23_ _08_ 0.030554f
C622 _11_ a_4929_3311# 0.001677f
C623 _21_ a_5179_3311# 5.62e-21
C624 _15_ a_5795_3133# 2.85e-21
C625 net6 _13_ 2.81e-21
C626 a_4220_3829# a_4443_4175# 0.011458f
C627 counter[7] counter[9] 2.14e-19
C628 _23_ net11 0.257634f
C629 a_7258_3829# a_7090_3855# 0.239923f
C630 a_6817_3861# a_7683_3829# 0.034054f
C631 a_6651_3861# a_7515_3855# 0.032244f
C632 a_4520_4373# VPWR 0.084816f
C633 net8 a_4767_3463# 0.236033f
C634 a_2401_4399# net5 3.57e-21
C635 a_2235_4399# net8 9.67e-20
C636 _04_ a_3099_4765# 0.006456f
C637 a_2502_7396# _12_ 0.032034f
C638 a_1959_3311# a_2745_2388# 8.97e-21
C639 a_4786_5065# a_4986_5220# 0.074815f
C640 a_4495_5175# _05_ 9.72e-20
C641 _23_ _22_ 0.511385f
C642 a_4779_5161# a_4915_5321# 0.136009f
C643 net6 a_5618_3677# 6.05e-21
C644 a_5149_4721# a_5250_3855# 0.001605f
C645 _11_ a_6651_3861# 3.54e-20
C646 a_5213_4664# _07_ 0.001092f
C647 clknet_0_clk a_5786_3423# 8.09e-19
C648 _11_ a_4495_5175# 1.82e-19
C649 VPWR clk 1.81336f
C650 net4 counter[1] 3.68e-19
C651 net2 a_2849_7663# 1.04e-19
C652 net6 a_4585_2388# 0.195979f
C653 a_4399_5175# a_4520_4373# 0.002561f
C654 a_2547_3855# a_1959_3311# 0.002525f
C655 a_2524_3311# VPWR 0.003212f
C656 a_5675_3855# clk 2.32e-21
C657 _09_ a_7723_2741# 0.17213f
C658 clknet_0_clk a_6651_5309# 6.75e-20
C659 net6 a_4220_3829# 0.050235f
C660 net4 a_3099_4765# 0.002624f
C661 net7 _07_ 0.047771f
C662 net9 a_6427_2741# 9.8e-19
C663 clknet_0_clk a_3215_3829# 4.87e-21
C664 net6 a_5213_4664# 0.027058f
C665 a_2302_7937# a_2502_7396# 1.26e-19
C666 a_2295_7637# a_2302_7241# 3.36e-19
C667 a_2502_7637# a_2295_7337# 6.88e-20
C668 _17_ a_4495_5175# 0.036473f
C669 a_4329_5461# a_4779_5161# 0.022305f
C670 _15_ a_5801_4233# 0.00162f
C671 a_7515_3855# a_7723_2741# 9.49e-21
C672 _18_ a_3099_4765# 3.43e-19
C673 _11_ a_3831_3339# 0.163973f
C674 net6 net7 0.905861f
C675 _22_ a_6825_3133# 2.76e-20
C676 a_7090_3677# a_7005_3311# 0.037333f
C677 a_7683_3579# a_7515_3677# 0.310858f
C678 _11_ a_7723_2741# 2.01e-20
C679 net3 VPWR 2.1402f
C680 clknet_1_0__leaf_clk a_2695_6575# 0.00537f
C681 a_2849_7663# _11_ 2.48e-19
C682 a_2290_3829# a_2122_3855# 0.239923f
C683 net6 a_5436_4399# 0.001357f
C684 a_1849_3861# a_2715_3829# 0.034054f
C685 _06_ a_4220_3829# 0.002127f
C686 clknet_1_1__leaf_clk a_5786_3423# 0.046669f
C687 _16_ a_5533_3311# 1.98e-21
C688 a_4287_4399# _20_ 6.22e-20
C689 _06_ a_5213_4664# 9.69e-19
C690 _17_ a_3831_3339# 6.88e-22
C691 _00_ a_2295_7637# 0.118744f
C692 a_2991_3579# net5 0.13266f
C693 a_2253_7119# VPWR 0.004522f
C694 clknet_1_1__leaf_clk a_3215_3829# 1.5e-19
C695 a_2235_4399# _04_ 0.09532f
C696 a_7005_3855# VPWR 0.078044f
C697 a_2011_7351# a_2431_7497# 0.036838f
C698 a_1915_7351# _01_ 1.56e-19
C699 net9 a_5165_3855# 1.41e-19
C700 a_2295_7337# a_2502_7396# 0.260055f
C701 clknet_1_0__leaf_clk a_2493_3677# 5.04e-19
C702 _16_ a_5418_3829# 0.001117f
C703 net7 _06_ 0.141876f
C704 _08_ a_7641_4233# 7.43e-19
C705 _15_ a_5786_3423# 4.59e-21
C706 _18_ a_4786_5065# 1.59e-19
C707 VPWR counter[7] 0.49968f
C708 net2 _03_ 5.34e-20
C709 a_5250_3855# a_5345_3855# 0.007724f
C710 a_2840_3087# a_2936_2767# 0.002032f
C711 a_5418_3829# a_5759_3855# 9.73e-19
C712 _06_ a_5436_4399# 6.53e-20
C713 a_1825_2388# counter[1] 0.1107f
C714 a_1683_3861# a_1959_3311# 0.001876f
C715 _15_ a_6651_5309# 0.001194f
C716 net1 clknet_1_0__leaf_clk 0.561165f
C717 _19_ a_5333_5321# 0.014678f
C718 net9 a_7599_3855# 1.06e-19
C719 _15_ a_3215_3829# 8.84e-19
C720 a_5418_3829# counter[5] 2.7e-21
C721 counter[2] counter[3] 0.070133f
C722 net3 a_2823_3677# 1.53e-21
C723 _13_ VPWR 0.524973f
C724 _11_ a_2217_3855# 3.45e-19
C725 net4 a_2235_4399# 0.071607f
C726 clknet_1_1__leaf_clk a_4995_4399# 3.57e-20
C727 a_2037_3855# a_1959_3311# 2.5e-19
C728 clknet_1_0__leaf_clk a_2230_7663# 0.001704f
C729 _00_ a_2302_7241# 4.06e-19
C730 clknet_0_clk net9 0.132797f
C731 a_5149_4721# _07_ 0.096566f
C732 _18_ a_2235_4399# 7.56e-20
C733 a_5618_3677# VPWR 0.256044f
C734 _09_ a_7753_2767# 0.07143f
C735 _11_ _21_ 0.059807f
C736 _16_ a_2566_3423# 0.005579f
C737 _11_ _03_ 0.00174f
C738 a_4585_2388# VPWR 0.287214f
C739 _16_ a_3831_3105# 0.039613f
C740 a_4349_3855# a_4259_3311# 8.68e-19
C741 _09_ a_7090_3677# 0.0221f
C742 a_7289_5309# VPWR 6.35e-19
C743 a_6651_3311# a_7683_3579# 0.048748f
C744 a_5675_3855# a_5618_3677# 7.26e-19
C745 clknet_1_0__leaf_clk a_2651_7485# 4.64e-19
C746 _04_ a_3245_3855# 0.072162f
C747 net9 a_6817_3311# 0.047741f
C748 a_7599_3677# VPWR 0.005629f
C749 VPWR counter[2] 0.494839f
C750 a_4779_5161# a_5345_3311# 4.79e-20
C751 a_4220_3829# VPWR 0.17068f
C752 net6 a_5149_4721# 0.09145f
C753 net11 a_7939_2223# 0.250513f
C754 _08_ a_5250_3855# 1.22e-20
C755 _23_ a_6825_3133# 1.08e-20
C756 _17_ _21_ 0.019243f
C757 a_5213_4664# VPWR 0.129866f
C758 a_7077_2767# counter[7] 1.91e-19
C759 clknet_0_clk a_4454_4649# 2.03e-19
C760 a_2401_4399# _14_ 3.24e-22
C761 a_4977_3861# a_5250_3855# 0.074815f
C762 a_4915_5321# a_5333_5321# 3.39e-19
C763 a_7683_3829# a_7683_3579# 0.026048f
C764 a_4811_3861# a_5843_3829# 0.048748f
C765 a_1582_7439# VPWR 4.93e-19
C766 a_5871_5162# _19_ 0.214472f
C767 _22_ a_5250_3855# 0.006172f
C768 a_4399_5175# a_4220_3829# 8.51e-20
C769 _11_ counter[6] 0.002692f
C770 net4 a_3245_3855# 0.005199f
C771 _11_ a_1849_3861# 0.008371f
C772 clknet_1_1__leaf_clk net9 0.461828f
C773 _24_ a_7185_3855# 7.21e-19
C774 _11_ a_7090_3677# 5.04e-19
C775 a_3799_4943# _18_ 0.09549f
C776 net7 VPWR 1.83862f
C777 a_5436_4399# VPWR 1.76e-19
C778 _19_ net8 2.14e-19
C779 a_4767_3463# a_5179_3311# 0.020429f
C780 a_5149_4721# _06_ 0.003245f
C781 net7 a_5675_3855# 0.054488f
C782 net2 counter[1] 0.015257f
C783 net6 _24_ 0.002355f
C784 _18_ a_3245_3855# 4.57e-20
C785 _16_ a_4349_4175# 0.001343f
C786 _01_ a_2678_7119# 5.75e-19
C787 a_2502_7396# _10_ 2.11e-19
C788 a_4329_5461# a_5333_5321# 8.9e-19
C789 a_6211_3579# a_6427_2741# 0.001105f
C790 a_4399_5175# net7 0.114197f
C791 clknet_0_clk a_7019_4943# 2.96e-20
C792 net3 a_1959_3311# 0.005671f
C793 a_2011_7637# VPWR 0.19379f
C794 _15_ net9 0.08758f
C795 a_2471_2741# VPWR 0.377321f
C796 _16_ a_4287_4399# 0.061172f
C797 clknet_1_1__leaf_clk a_4454_4649# 0.007927f
C798 _24_ a_7363_3087# 0.002926f
C799 net8 a_6651_3311# 3.27e-19
C800 a_2235_4399# a_2715_3829# 4.12e-19
C801 a_7199_4943# a_7619_5162# 0.017591f
C802 _04_ a_2122_3855# 3.3e-20
C803 clknet_1_0__leaf_clk a_2547_3855# 0.004501f
C804 a_2949_3311# VPWR 4.65e-19
C805 a_2547_3855# a_2840_3087# 3.78e-21
C806 a_7199_4943# a_6651_3311# 3.35e-21
C807 a_5814_4399# net10 3.58e-19
C808 _22_ a_5599_2741# 0.106132f
C809 a_4986_5220# _19_ 0.034076f
C810 _15_ a_4454_4649# 5.11e-20
C811 net8 a_7683_3829# 4.93e-20
C812 net9 a_4929_3311# 8.5e-21
C813 net4 a_2122_3855# 4.27e-19
C814 a_2235_6575# a_1845_5461# 5.68e-19
C815 _10_ a_2389_6575# 5.49e-20
C816 _14_ a_2991_3579# 1.14e-20
C817 net6 a_5345_3855# 0.001259f
C818 a_4915_5321# net8 0.00192f
C819 a_7090_3855# a_6651_3311# 1.73e-19
C820 a_2125_3311# a_2398_3677# 0.081834f
C821 clknet_1_1__leaf_clk a_7019_4943# 7.87e-19
C822 _11_ a_3099_4765# 0.043928f
C823 a_3267_4667# a_4520_4373# 2.22e-20
C824 a_2011_7351# VPWR 0.181976f
C825 net9 a_6651_3861# 8.34e-19
C826 _13_ a_1959_3311# 6.65e-20
C827 _15_ net5 0.016962f
C828 a_1505_3855# VPWR 0.006911f
C829 _23_ a_7939_2223# 9.55e-20
C830 a_4329_5461# a_5871_5162# 1.59e-19
C831 _07_ a_6043_3677# 5.62e-20
C832 a_2295_7637# a_2431_7663# 0.141453f
C833 a_2302_7937# a_2253_8029# 6.32e-19
C834 a_2125_8207# clknet_1_0__leaf_clk 2.59e-19
C835 _15_ a_5997_3133# 5.62e-21
C836 a_2823_3677# a_2949_3311# 0.006169f
C837 a_4811_3861# a_5165_3855# 0.057611f
C838 _15_ a_7019_4943# 0.001697f
C839 a_4329_5461# net8 0.001938f
C840 a_7258_3829# a_7515_3855# 0.036838f
C841 a_2547_3855# a_2631_3855# 0.008508f
C842 _17_ a_3099_4765# 1.03e-20
C843 a_2715_3829# a_3245_3855# 2.84e-19
C844 a_2674_4765# net5 1.47e-19
C845 a_5149_4721# VPWR 0.2552f
C846 _08_ _07_ 9.41e-21
C847 a_7258_3423# counter[7] 1.4e-19
C848 _01_ _12_ 0.353697f
C849 net6 a_6043_3677# 4.38e-19
C850 _07_ a_4977_3861# 0.029939f
C851 a_4786_5065# _05_ 0.181338f
C852 a_4986_5220# a_4915_5321# 0.239923f
C853 a_1875_8207# VPWR 0.260172f
C854 a_5814_4399# a_5843_3829# 0.009572f
C855 _22_ _07_ 0.503878f
C856 net2 a_2235_4399# 2.26e-20
C857 _11_ a_4786_5065# 3.7e-19
C858 a_4495_5175# a_4454_4649# 0.001715f
C859 net7 a_5376_4233# 2.79e-19
C860 net6 _08_ 5.42e-20
C861 clknet_1_0__leaf_clk a_1683_3861# 0.318658f
C862 clknet_0_clk a_5162_4943# 4.01e-19
C863 net6 a_4977_3861# 0.048602f
C864 net9 a_7723_2741# 0.001158f
C865 a_6623_3133# VPWR 0.001618f
C866 a_4779_5161# clk 4.16e-19
C867 a_1457_2388# a_1825_2388# 2.48e-19
C868 a_2302_7937# _01_ 8.68e-20
C869 a_2295_7637# a_2431_7497# 5.28e-20
C870 _18_ _19_ 0.036736f
C871 _24_ VPWR 0.6956f
C872 a_6211_3579# a_6817_3311# 8.52e-19
C873 clknet_0_clk a_4811_3861# 0.009291f
C874 net6 _22_ 0.641715f
C875 a_2502_7637# a_2502_7396# 0.013851f
C876 _17_ a_4786_5065# 0.050404f
C877 a_6425_2388# counter[9] 2.37e-20
C878 a_4329_5461# a_4986_5220# 0.007109f
C879 clknet_1_0__leaf_clk a_2037_3855# 0.03291f
C880 clknet_0_clk a_5077_4721# 2.68e-20
C881 _21_ a_4995_4399# 0.053333f
C882 _15_ a_7216_4233# 4.15e-19
C883 _23_ a_5599_2741# 2.79e-19
C884 _11_ a_4767_3463# 0.046716f
C885 net11 counter[9] 0.066386f
C886 a_2401_4399# _16_ 1.01e-19
C887 a_4520_4373# a_4259_3311# 7.94e-19
C888 _22_ a_7363_3087# 3.67e-19
C889 a_7258_3423# a_7599_3677# 9.73e-19
C890 _11_ a_2235_4399# 0.205946f
C891 net8 a_4349_3855# 2.79e-20
C892 a_2290_3829# a_2547_3855# 0.036838f
C893 _11_ a_3389_3105# 8.14e-19
C894 clknet_1_1__leaf_clk a_6211_3579# 0.084941f
C895 _06_ a_4977_3861# 0.183131f
C896 a_5814_4399# a_6427_2741# 4.57e-20
C897 _16_ a_4341_3311# 0.00109f
C898 a_1959_3311# a_2471_2741# 2.64e-19
C899 _00_ a_2431_7663# 0.005564f
C900 _06_ _22_ 0.004416f
C901 clknet_1_1__leaf_clk a_5505_2388# 4.13e-21
C902 _17_ a_4767_3463# 1.09e-21
C903 a_3831_3339# net5 4.5e-19
C904 a_2313_3311# a_2493_3677# 0.001229f
C905 net7 a_4714_5309# 0.001683f
C906 _17_ a_2235_4399# 1.5e-21
C907 net6 a_3215_2999# 5.34e-20
C908 a_2235_6575# VPWR 0.266078f
C909 net10 a_7345_2388# 2.65e-20
C910 net7 a_7258_3423# 1.23e-19
C911 a_2295_7337# _01_ 0.092611f
C912 a_5345_3855# VPWR 0.004219f
C913 clknet_1_1__leaf_clk a_4811_3861# 0.670964f
C914 a_2302_7241# a_2431_7497# 0.124967f
C915 _15_ a_6211_3579# 7.77e-19
C916 _18_ a_4915_5321# 7.52e-20
C917 a_3979_4943# _16_ 1.86e-20
C918 a_3799_4943# _05_ 4.45e-20
C919 a_6427_2741# a_6719_3133# 0.001675f
C920 _11_ a_3799_4943# 0.001422f
C921 a_6817_3861# a_7005_3855# 0.097994f
C922 _21_ net9 0.170283f
C923 _24_ a_7077_2767# 0.085832f
C924 net8 a_5345_3311# 0.003497f
C925 _15_ a_4811_3861# 0.034785f
C926 a_2561_9514# net1 0.10983f
C927 _11_ a_3245_3855# 2.49e-20
C928 net3 a_2041_4649# 0.001185f
C929 a_5179_3311# a_6651_3311# 0.003146f
C930 clknet_1_0__leaf_clk net3 0.373279f
C931 a_5786_3423# a_6127_3677# 9.73e-19
C932 net4 a_2936_2767# 0.003167f
C933 net3 a_2840_3087# 9.94e-20
C934 a_3099_4765# a_3215_3829# 0.001534f
C935 _17_ a_3799_4943# 0.250762f
C936 net2 a_1457_2388# 0.223155f
C937 _23_ a_7185_3855# 8.32e-19
C938 net6 a_3433_4175# 0.001315f
C939 a_4454_4649# _21_ 0.128337f
C940 _16_ a_2991_3579# 1.37e-19
C941 a_6043_3677# VPWR 0.1878f
C942 _01_ a_3145_6825# 0.012244f
C943 net9 a_7753_2767# 0.005829f
C944 net6 _23_ 0.023006f
C945 a_6425_2388# VPWR 0.309637f
C946 _15_ _14_ 1.65e-19
C947 net6 a_3225_4399# 5.88e-19
C948 a_5675_3855# a_6043_3677# 3.78e-19
C949 _09_ a_7515_3677# 0.024482f
C950 a_6651_3311# a_7005_3311# 0.062224f
C951 _08_ VPWR 0.467036f
C952 clknet_0_clk a_6375_5309# 1.5e-19
C953 _02_ a_1849_3861# 0.275992f
C954 a_1683_3861# a_2290_3829# 0.141453f
C955 clknet_1_0__leaf_clk a_2253_7119# 0.002574f
C956 net9 counter[6] 3.69e-19
C957 net9 a_7090_3677# 0.023502f
C958 net6 a_2589_4399# 5.63e-21
C959 net1 a_1499_7119# 0.060735f
C960 a_4977_3861# VPWR 0.300379f
C961 a_4779_5161# a_5618_3677# 7.91e-22
C962 net11 VPWR 0.794015f
C963 clknet_1_1__leaf_clk _20_ 0.0051f
C964 _23_ a_7363_3087# 2.44e-19
C965 _08_ a_5675_3855# 7.33e-20
C966 clknet_0_clk a_5814_4399# 0.316676f
C967 _22_ VPWR 0.56354f
C968 a_2674_4765# _14_ 5.19e-22
C969 _11_ a_3917_3339# 0.003027f
C970 _21_ net5 2.83e-22
C971 _23_ counter[9] 7.62e-19
C972 _15_ a_2614_2883# 4.86e-20
C973 a_4811_3861# a_6651_3861# 0.002059f
C974 a_4977_3861# a_5675_3855# 0.192206f
C975 _03_ net5 3.86e-19
C976 a_1849_3861# a_2248_4233# 8.12e-19
C977 a_7515_3855# a_7515_3677# 0.01464f
C978 a_2290_3829# a_2037_3855# 3.39e-19
C979 a_3215_2999# counter[3] 6.79e-20
C980 a_5418_3829# a_5843_3829# 1.28e-19
C981 _22_ a_5675_3855# 1.1e-21
C982 a_4495_5175# a_4811_3861# 1.16e-21
C983 _15_ _20_ 0.093509f
C984 _13_ a_2041_4649# 0.01129f
C985 clknet_1_0__leaf_clk _13_ 0.02176f
C986 a_4779_5161# a_5213_4664# 0.00484f
C987 _11_ a_7515_3677# 3.81e-21
C988 _11_ a_2122_3855# 0.003174f
C989 a_5814_4399# a_6817_3311# 2.14e-19
C990 _18_ a_4349_3855# 3.94e-20
C991 net7 a_6817_3861# 2.99e-20
C992 _19_ _25_ 9.05e-21
C993 _01_ _10_ 0.002197f
C994 clknet_1_1__leaf_clk a_6375_5309# 0.001522f
C995 a_2125_3311# VPWR 0.342267f
C996 _17_ a_4737_4943# 0.002375f
C997 a_4779_5161# net7 0.035144f
C998 a_2295_7637# VPWR 0.721856f
C999 a_3215_2999# VPWR 0.201367f
C1000 a_4220_3829# a_4259_3311# 2.2e-19
C1001 clknet_1_1__leaf_clk a_5814_4399# 1.80017f
C1002 a_7619_5162# _25_ 0.227897f
C1003 _04_ a_2547_3855# 0.001211f
C1004 a_2235_4399# a_3215_3829# 0.002539f
C1005 a_2800_4399# _16_ 2.63e-21
C1006 _15_ a_6375_5309# 0.142876f
C1007 net11 a_7077_2767# 2.78e-19
C1008 _24_ a_7258_3423# 0.014122f
C1009 _05_ _19_ 0.284135f
C1010 _22_ a_7077_2767# 0.140356f
C1011 a_6651_3311# _09_ 0.098799f
C1012 net4 a_2745_2388# 0.202764f
C1013 _15_ a_5814_4399# 0.047247f
C1014 net7 a_4259_3311# 0.003261f
C1015 _11_ _19_ 0.032711f
C1016 net9 a_6127_3677# 8.89e-19
C1017 clknet_0_clk _16_ 0.019509f
C1018 a_4495_5175# _20_ 1.76e-19
C1019 net4 a_2547_3855# 0.006897f
C1020 a_2842_4511# a_3225_4399# 4.67e-20
C1021 clknet_1_1__leaf_clk a_6719_3133# 3.29e-19
C1022 a_7683_3829# _09_ 5.87e-19
C1023 a_2842_4511# a_2589_4399# 3.39e-19
C1024 net8 a_4520_4373# 0.028641f
C1025 a_2566_3423# a_2991_3579# 1.28e-19
C1026 a_7515_3855# a_6651_3311# 1.29e-19
C1027 a_2125_3311# a_2823_3677# 0.195152f
C1028 a_5871_5162# clk 0.012863f
C1029 a_2302_7241# VPWR 0.309635f
C1030 net9 a_7258_3829# 2.66e-21
C1031 _17_ _19_ 0.214371f
C1032 net2 a_2695_6575# 3.45e-20
C1033 a_2823_3677# a_3215_2999# 0.001309f
C1034 _07_ a_5713_3677# 2.91e-19
C1035 _23_ VPWR 1.70159f
C1036 a_3433_4175# VPWR 0.001324f
C1037 net10 a_7267_3087# 8.38e-19
C1038 _11_ a_6651_3311# 0.012822f
C1039 a_2011_7637# clknet_1_0__leaf_clk 0.038899f
C1040 a_2302_7937# a_2849_7663# 0.095025f
C1041 a_4786_5065# net9 1.52e-20
C1042 a_2295_7637# a_2678_8029# 0.002698f
C1043 _15_ a_6719_3133# 0.00403f
C1044 a_4349_3855# counter[4] 4.47e-20
C1045 net1 a_1957_8207# 0.010028f
C1046 a_3215_3829# a_3245_3855# 0.025037f
C1047 a_3831_3339# _20_ 3.41e-19
C1048 a_2715_3829# a_4349_3855# 2.67e-21
C1049 a_7683_3829# a_7515_3855# 0.310858f
C1050 a_5418_3829# a_5165_3855# 3.39e-19
C1051 a_2471_2741# a_2840_3087# 0.046138f
C1052 a_3099_4765# net5 4.89e-20
C1053 a_2589_4399# VPWR 0.093135f
C1054 _07_ a_5250_3855# 0.002926f
C1055 a_4915_5321# _05_ 0.001005f
C1056 _00_ VPWR 0.655201f
C1057 a_5814_4399# a_6651_3861# 0.016172f
C1058 net8 a_5891_3133# 0.001229f
C1059 clknet_1_1__leaf_clk _16_ 0.001692f
C1060 _21_ a_4811_3861# 0.016583f
C1061 _11_ a_4915_5321# 5.19e-20
C1062 a_4779_5161# a_5149_4721# 0.007926f
C1063 a_4786_5065# a_4454_4649# 0.002652f
C1064 a_5179_3311# a_5345_3311# 0.966391f
C1065 net9 a_4767_3463# 3.24e-20
C1066 a_2695_6575# _11_ 0.201886f
C1067 _04_ a_1683_3861# 0.001469f
C1068 a_2317_6575# VPWR 2.01e-19
C1069 clknet_1_1__leaf_clk a_5759_3855# 0.001538f
C1070 a_2302_7937# enable 4.56e-21
C1071 net1 net2 0.722672f
C1072 net6 a_5250_3855# 0.019975f
C1073 _15_ _16_ 0.656968f
C1074 a_6825_3133# VPWR 1.16e-19
C1075 a_6211_3579# counter[6] 4.54e-21
C1076 a_1825_2388# a_2745_2388# 1.37e-20
C1077 clknet_0_clk a_5418_3829# 3.18e-19
C1078 a_2431_7663# a_2431_7497# 0.013661f
C1079 clknet_1_0__leaf_clk a_2011_7351# 0.044938f
C1080 _17_ a_4915_5321# 0.016441f
C1081 a_4329_5461# _05_ 0.005813f
C1082 a_5505_2388# counter[6] 4.98e-19
C1083 _04_ a_2037_3855# 3.27e-21
C1084 a_7939_2223# counter[9] 0.109832f
C1085 _11_ a_4329_5461# 4.59e-19
C1086 net2 a_2230_7663# 2.28e-19
C1087 clknet_1_0__leaf_clk a_1505_3855# 1.21e-20
C1088 _24_ a_6817_3861# 0.035946f
C1089 _14_ _03_ 0.071143f
C1090 a_2674_4765# _16_ 1.81e-20
C1091 _11_ a_2493_3677# 6.67e-19
C1092 _23_ a_7077_2767# 0.04546f
C1093 net4 a_1683_3861# 0.007432f
C1094 a_4454_4649# a_4767_3463# 2.49e-20
C1095 a_7090_3677# a_7216_3311# 0.005525f
C1096 a_7005_3311# a_7185_3677# 0.001229f
C1097 a_2235_4399# a_4454_4649# 1.89e-21
C1098 _22_ a_7171_2767# 0.063386f
C1099 _04_ a_4520_4373# 8.65e-21
C1100 a_2715_3829# a_2547_3855# 0.310858f
C1101 a_1959_3311# a_2125_3311# 0.970278f
C1102 _07_ a_5599_2741# 9.24e-19
C1103 net8 a_7005_3855# 1.28e-19
C1104 _18_ a_1683_3861# 3.08e-21
C1105 _22_ a_7258_3423# 8.71e-19
C1106 _06_ a_5250_3855# 3.32e-19
C1107 clknet_1_1__leaf_clk a_5533_3311# 0.011819f
C1108 net1 _11_ 0.002334f
C1109 _03_ a_2614_2883# 0.005187f
C1110 _16_ a_4929_3311# 7.06e-20
C1111 net8 counter[7] 5.9e-19
C1112 net4 a_2037_3855# 1.97e-19
C1113 a_1875_8207# clknet_1_0__leaf_clk 3.24e-19
C1114 a_4329_5461# _17_ 7.15e-19
C1115 _00_ a_2678_8029# 8.32e-19
C1116 _21_ _20_ 0.296715f
C1117 net7 a_5333_5321# 0.019182f
C1118 a_1683_3861# a_3601_3855# 4.04e-20
C1119 net6 a_5599_2741# 0.211407f
C1120 a_2235_4399# net5 1.51e-20
C1121 net7 a_7683_3579# 8.32e-20
C1122 a_2502_7396# _01_ 0.004715f
C1123 a_7641_4233# VPWR 7.83e-19
C1124 clknet_1_1__leaf_clk a_5418_3829# 0.01748f
C1125 a_1915_7351# a_2230_7485# 7.84e-20
C1126 _15_ a_5533_3311# 7.24e-21
C1127 net10 a_8265_2388# 0.219068f
C1128 _14_ a_1849_3861# 4.89e-20
C1129 net5 a_3389_3105# 0.002311f
C1130 a_4495_5175# _16_ 1.29e-20
C1131 a_7258_3829# a_7216_4233# 4.62e-19
C1132 a_7090_3855# a_7005_3855# 0.037333f
C1133 _15_ a_7345_2388# 0.006207f
C1134 _18_ a_4520_4373# 7.58e-19
C1135 a_2849_7497# a_2695_6575# 6.31e-19
C1136 net8 a_5618_3677# 0.001808f
C1137 a_7515_3677# a_7641_3311# 0.006169f
C1138 _15_ a_5418_3829# 0.03519f
C1139 _11_ a_4349_3855# 0.07562f
C1140 net3 a_2313_3311# 7.76e-19
C1141 net4 a_2524_3311# 6.57e-19
C1142 net3 _04_ 5.28e-22
C1143 a_5618_3677# a_5744_3311# 0.005525f
C1144 a_7199_4943# a_7289_5309# 0.004764f
C1145 net8 a_4220_3829# 2.76e-19
C1146 _16_ a_3831_3339# 0.113241f
C1147 a_5713_3677# VPWR 0.003234f
C1148 a_5814_4399# _21_ 3.33e-20
C1149 net8 a_5213_4664# 0.003744f
C1150 a_2431_7497# a_1845_5461# 1.29e-20
C1151 _17_ a_4349_3855# 9.12e-21
C1152 a_5871_5162# net7 0.030401f
C1153 a_7939_2223# VPWR 0.293517f
C1154 a_1683_3861# a_2715_3829# 0.048748f
C1155 _14_ counter[1] 1.03e-21
C1156 net6 _07_ 0.066033f
C1157 clknet_1_0__leaf_clk a_2235_6575# 0.024338f
C1158 _02_ a_2122_3855# 8.22e-19
C1159 net3 net4 0.0313f
C1160 net9 a_7515_3677# 0.020729f
C1161 a_5250_3855# VPWR 0.255475f
C1162 net10 a_6427_2741# 0.158335f
C1163 net7 net8 1.22349f
C1164 net1 a_2849_7497# 6.38e-20
C1165 _23_ a_7171_2767# 0.038842f
C1166 _08_ a_6817_3861# 0.415957f
C1167 _11_ a_5345_3311# 0.042209f
C1168 net8 a_5436_4399# 1.76e-19
C1169 a_2122_3855# a_2248_4233# 0.005525f
C1170 net7 a_7199_4943# 5.4e-19
C1171 _15_ a_3831_3105# 0.110742f
C1172 a_4977_3861# a_6817_3861# 0.001861f
C1173 a_2401_4399# a_2991_3579# 8.13e-20
C1174 _11_ a_2745_2388# 3.83e-19
C1175 _23_ a_7258_3423# 0.005759f
C1176 _06_ a_4443_4175# 6.56e-20
C1177 _13_ _04_ 1.41e-19
C1178 _11_ a_6545_5309# 0.001703f
C1179 a_4779_5161# a_4977_3861# 3.93e-19
C1180 net3 a_1499_7119# 0.042192f
C1181 a_4786_5065# a_4811_3861# 1.6e-20
C1182 _22_ a_6817_3861# 4.96e-21
C1183 a_5814_4399# a_7090_3677# 6.58e-20
C1184 a_4779_5161# _22_ 1.01e-19
C1185 a_4986_5220# a_5213_4664# 3.7e-19
C1186 _11_ a_2547_3855# 0.017838f
C1187 _17_ a_5345_3311# 6.74e-21
C1188 _06_ _07_ 5.11e-20
C1189 net5 a_3917_3339# 2.72e-19
C1190 net2 a_2125_8207# 0.008042f
C1191 a_2398_3677# VPWR 0.286549f
C1192 a_4986_5220# net7 0.026259f
C1193 a_2431_7663# VPWR 0.211499f
C1194 a_4915_5321# a_4995_4399# 1.71e-20
C1195 net4 _13_ 0.050083f
C1196 net6 _06_ 0.037389f
C1197 a_5599_2741# VPWR 0.405792f
C1198 _19_ net9 4.58e-20
C1199 a_4811_3861# a_4767_3463# 1.28e-19
C1200 _21_ _16_ 0.249175f
C1201 _15_ a_4349_4175# 0.005043f
C1202 counter[7] counter[8] 0.067503f
C1203 _16_ _03_ 0.005745f
C1204 a_5675_3855# a_5599_2741# 3.32e-21
C1205 _24_ a_7683_3579# 0.009415f
C1206 net10 a_7599_3855# 3.67e-19
C1207 net2 a_1683_3861# 3.28e-19
C1208 _15_ a_4287_4399# 9.44e-19
C1209 net3 a_1825_2388# 0.233128f
C1210 a_4329_5461# a_4995_4399# 2.81e-20
C1211 net9 a_6651_3311# 0.11266f
C1212 net4 a_4220_3829# 1.34e-19
C1213 net4 counter[2] 0.006188f
C1214 a_3267_4667# a_3225_4399# 7.84e-20
C1215 net6 counter[3] 1.1e-21
C1216 a_2674_4765# a_2769_4765# 0.007724f
C1217 _14_ a_3389_3105# 5.76e-19
C1218 net8 a_5149_4721# 0.003186f
C1219 a_2842_4511# a_3183_4765# 9.73e-19
C1220 a_2431_7497# VPWR 0.211083f
C1221 _18_ a_4220_3829# 0.079699f
C1222 net10 a_7941_3087# 0.002502f
C1223 a_4443_4175# VPWR 2.25e-21
C1224 clknet_1_0__leaf_clk a_2125_3311# 0.021572f
C1225 a_3831_3339# a_3831_3105# 0.012876f
C1226 _16_ a_1849_3861# 8.97e-20
C1227 a_2125_3311# a_2840_3087# 4.63e-19
C1228 a_2295_7637# clknet_1_0__leaf_clk 0.308902f
C1229 _11_ a_1683_3861# 0.00462f
C1230 a_4915_5321# net9 0.004659f
C1231 a_2502_7637# a_2849_7663# 0.037333f
C1232 _07_ VPWR 0.322336f
C1233 net10 a_6817_3311# 0.003321f
C1234 _15_ a_7267_3087# 0.004129f
C1235 net6 a_2842_4511# 3.85e-19
C1236 a_5250_3855# a_5376_4233# 0.005525f
C1237 _23_ a_6817_3861# 0.031087f
C1238 a_3215_2999# a_2840_3087# 4e-20
C1239 a_4767_3463# _20_ 0.113204f
C1240 net1 a_1915_7815# 0.045364f
C1241 a_7005_3311# counter[7] 2.77e-20
C1242 a_5871_5162# _24_ 1.86e-20
C1243 a_3183_4765# VPWR 0.004177f
C1244 counter[5] counter[6] 0.070133f
C1245 _12_ a_2230_7485# 0.001666f
C1246 a_7185_3855# VPWR 0.002923f
C1247 a_1582_7439# a_1499_7119# 2.42e-19
C1248 _18_ net7 0.004371f
C1249 _07_ a_5675_3855# 0.009837f
C1250 _11_ a_2037_3855# 2.52e-19
C1251 a_5814_4399# a_7258_3829# 0.006157f
C1252 a_4495_5175# a_4287_4399# 9.42e-20
C1253 _24_ net8 1.23e-20
C1254 a_1915_7815# a_2230_7663# 7.84e-20
C1255 net6 VPWR 3.11824f
C1256 a_5179_3311# a_5618_3677# 0.273138f
C1257 a_4329_5461# net9 1.97e-19
C1258 a_5345_3311# a_5786_3423# 0.110715f
C1259 net4 a_2471_2741# 0.021386f
C1260 a_1845_5461# VPWR 1.52032f
C1261 clknet_1_1__leaf_clk net10 6.99e-20
C1262 _24_ a_7199_4943# 0.197975f
C1263 _11_ a_4520_4373# 0.002559f
C1264 a_2502_7637# enable 1.46e-21
C1265 net4 a_2949_3311# 0.00133f
C1266 net6 a_5675_3855# 8.63e-19
C1267 a_4399_5175# net6 1.76e-19
C1268 a_7363_3087# VPWR 4.51e-19
C1269 _05_ clk 0.0016f
C1270 a_2745_2388# a_3849_2388# 9e-21
C1271 clknet_1_0__leaf_clk a_2302_7241# 0.083453f
C1272 clknet_0_clk a_5843_3829# 0.01296f
C1273 _11_ clk 1.2e-19
C1274 clknet_0_clk a_3979_4943# 8e-19
C1275 VPWR counter[9] 0.449609f
C1276 net2 net3 1.28152f
C1277 a_1825_2388# counter[2] 4.98e-19
C1278 _15_ net10 0.289356f
C1279 net11 a_8109_2767# 0.004987f
C1280 clknet_1_0__leaf_clk a_3433_4175# 1.8e-20
C1281 net1 a_1915_7351# 0.081622f
C1282 a_4585_2388# counter[4] 0.110403f
C1283 a_7090_3677# a_7345_2388# 6.36e-19
C1284 a_4329_5461# a_4454_4649# 1.01e-19
C1285 _17_ a_4520_4373# 0.062168f
C1286 a_3099_4765# _16_ 0.003542f
C1287 a_5333_5321# a_4977_3861# 1.11e-20
C1288 _24_ a_7090_3855# 0.010979f
C1289 _06_ VPWR 0.276236f
C1290 a_7683_3579# net11 0.092457f
C1291 a_1959_3311# a_2398_3677# 0.273138f
C1292 _03_ a_2566_3423# 0.006259f
C1293 a_5333_5321# _22_ 0.001069f
C1294 a_3979_4943# a_4069_5309# 0.004764f
C1295 a_2715_3829# a_4220_3829# 1e-20
C1296 net8 a_5345_3855# 4.84e-19
C1297 clknet_1_0__leaf_clk a_2589_4399# 0.003123f
C1298 _17_ clk 1.68e-19
C1299 net7 a_5179_3311# 0.003956f
C1300 _06_ a_5675_3855# 9.38e-20
C1301 _03_ a_3831_3105# 2.93e-20
C1302 _00_ clknet_1_0__leaf_clk 0.144154f
C1303 net7 a_6457_5309# 0.003849f
C1304 net6 a_7077_2767# 5.59e-20
C1305 _14_ a_1457_2388# 0.001394f
C1306 _09_ counter[7] 5.27e-21
C1307 net7 a_7005_3311# 2.26e-19
C1308 a_2401_4399# a_2674_4765# 0.074434f
C1309 clknet_1_1__leaf_clk a_5843_3829# 0.005058f
C1310 net3 _11_ 0.005186f
C1311 clknet_1_0__leaf_clk a_2317_6575# 2.61e-19
C1312 _15_ a_4341_3311# 1.25e-19
C1313 a_3979_4943# clknet_1_1__leaf_clk 1.19e-21
C1314 a_4786_5065# _16_ 6.29e-20
C1315 VPWR counter[3] 0.49419f
C1316 a_6651_3861# net10 4.73e-19
C1317 net2 _13_ 0.197255f
C1318 a_7077_2767# a_7363_3087# 0.010132f
C1319 a_1849_3861# a_2566_3423# 0.001879f
C1320 a_2290_3829# a_2125_3311# 3.46e-19
C1321 net8 a_6043_3677# 0.007067f
C1322 _15_ a_5843_3829# 0.031321f
C1323 a_2715_3829# a_2471_2741# 2.52e-20
C1324 counter[0] counter[1] 0.079742f
C1325 net8 a_6425_2388# 0.2272f
C1326 a_2842_4511# VPWR 0.177502f
C1327 _19_ a_4811_3861# 9.86e-21
C1328 _21_ a_4349_4175# 2.03e-19
C1329 a_3979_4943# _15_ 2e-21
C1330 _08_ net8 2.38e-19
C1331 a_6211_3579# a_6651_3311# 0.001745f
C1332 _11_ counter[7] 2.36e-19
C1333 net8 a_4977_3861# 0.031957f
C1334 _25_ a_7289_5309# 8.17e-20
C1335 a_7199_4943# _08_ 0.001905f
C1336 _21_ a_4287_4399# 0.002821f
C1337 net9 a_5345_3311# 0.017191f
C1338 a_4413_3311# VPWR 3.08e-19
C1339 _16_ a_4767_3463# 1.3e-19
C1340 net8 _22_ 0.137056f
C1341 net6 a_5376_4233# 0.001426f
C1342 clknet_1_1__leaf_clk a_6427_2741# 3.39e-19
C1343 a_2235_4399# _16_ 6.86e-20
C1344 _11_ _13_ 0.217373f
C1345 _09_ a_7599_3677# 6.12e-19
C1346 a_1683_3861# a_3215_3829# 1.05e-19
C1347 _02_ a_2547_3855# 3.18e-19
C1348 _15_ a_2991_3579# 2.99e-20
C1349 net2 a_1582_7439# 0.010623f
C1350 a_5675_3855# VPWR 0.182006f
C1351 _22_ a_5744_3311# 6.82e-19
C1352 net10 a_7723_2741# 0.104575f
C1353 net6 a_4382_4649# 0.002624f
C1354 _08_ a_7090_3855# 0.030723f
C1355 _11_ a_5618_3677# 0.026293f
C1356 _23_ a_8109_2767# 0.009249f
C1357 a_5149_4721# a_5179_3311# 5.07e-21
C1358 a_2125_8207# a_1915_7815# 3.08e-19
C1359 a_4399_5175# VPWR 0.376761f
C1360 net7 _25_ 3.01e-19
C1361 a_5843_3829# a_6651_3861# 4.62e-19
C1362 _15_ a_6427_2741# 0.086673f
C1363 a_2674_4765# a_2991_3579# 2.18e-19
C1364 _23_ a_7683_3579# 2.3e-19
C1365 a_4779_5161# a_5250_3855# 8.34e-21
C1366 net7 _09_ 2.46e-19
C1367 a_4986_5220# a_4977_3861# 8.21e-21
C1368 a_4915_5321# a_4811_3861# 5.48e-20
C1369 net3 a_2849_7497# 4.27e-20
C1370 _11_ a_4220_3829# 0.058411f
C1371 _05_ a_5213_4664# 2.43e-19
C1372 _11_ a_5213_4664# 0.004209f
C1373 net6 a_7171_2767# 7.2e-20
C1374 net2 a_2011_7637# 0.019416f
C1375 net6 a_4714_5309# 1.91e-20
C1376 clknet_1_1__leaf_clk a_5165_3855# 0.017223f
C1377 a_2823_3677# VPWR 0.183311f
C1378 _16_ a_3245_3855# 0.059496f
C1379 _12_ a_2695_6575# 0.026119f
C1380 clknet_0_clk a_4069_5309# 9.48e-20
C1381 _05_ net7 0.232588f
C1382 a_4329_5461# a_4811_3861# 3.84e-19
C1383 _17_ a_4220_3829# 1.33e-19
C1384 a_2678_8029# VPWR 0.005789f
C1385 a_7077_2767# VPWR 0.152186f
C1386 a_7363_3087# a_7171_2767# 6.96e-20
C1387 _11_ net7 0.966176f
C1388 _17_ a_5213_4664# 2.72e-19
C1389 _15_ a_5165_3855# 0.019231f
C1390 _24_ a_7005_3311# 3.3e-19
C1391 a_5871_5162# _23_ 1.03e-19
C1392 _17_ net7 0.072785f
C1393 a_2302_7937# a_2695_6575# 6.42e-21
C1394 a_1683_3861# _02_ 0.184941f
C1395 _11_ a_2471_2741# 7.66e-19
C1396 clknet_0_clk clknet_1_1__leaf_clk 0.335671f
C1397 _23_ net8 0.011201f
C1398 _19_ a_5814_4399# 6.04e-19
C1399 _16_ a_3917_3339# 5.76e-19
C1400 net2 a_2011_7351# 0.00144f
C1401 net1 _12_ 0.312817f
C1402 _11_ a_2949_3311# 5.7e-19
C1403 net2 a_1505_3855# 0.002977f
C1404 a_1875_8207# a_1957_8207# 0.006406f
C1405 _23_ a_7199_4943# 0.007723f
C1406 a_2401_4399# _21_ 2.75e-21
C1407 a_2674_4765# a_2800_4399# 0.005525f
C1408 a_2991_3579# a_3831_3339# 7.43e-20
C1409 _14_ a_2936_2767# 0.003598f
C1410 a_2125_3311# a_2313_3311# 0.097994f
C1411 _02_ a_2037_3855# 0.114994f
C1412 a_2401_4399# _03_ 3.92e-19
C1413 clknet_1_0__leaf_clk a_2398_3677# 0.003461f
C1414 a_5376_4233# VPWR 0.001185f
C1415 clknet_0_clk _15_ 4.05e-19
C1416 clknet_1_1__leaf_clk a_6817_3311# 0.031849f
C1417 net10 a_7753_2767# 0.001384f
C1418 _16_ a_2122_3855# 1.68e-20
C1419 a_2431_7663# clknet_1_0__leaf_clk 0.050329f
C1420 _04_ a_3215_2999# 1.25e-20
C1421 net6 a_3267_4667# 0.129987f
C1422 a_5814_4399# a_6651_3311# 6.92e-20
C1423 net10 a_7090_3677# 5.45e-19
C1424 _23_ a_7090_3855# 0.012578f
C1425 a_2561_9514# a_2295_7637# 6.9e-23
C1426 net1 a_2302_7937# 0.006588f
C1427 a_4811_3861# a_4349_3855# 1.44e-19
C1428 net2 a_1875_8207# 0.107098f
C1429 net11 counter[8] 0.024563f
C1430 a_4382_4649# VPWR 0.011634f
C1431 a_2295_7337# a_2695_6575# 4.04e-19
C1432 a_1959_3311# VPWR 0.741952f
C1433 _15_ a_6817_3311# 0.036316f
C1434 _12_ a_2651_7485# 0.002771f
C1435 net4 a_2125_3311# 0.019846f
C1436 net6 a_5001_3311# 7.29e-19
C1437 net9 clk 4.05e-20
C1438 a_4779_5161# _07_ 5.99e-19
C1439 a_1915_7815# net3 9.98e-20
C1440 a_5345_3311# a_6211_3579# 0.034054f
C1441 _05_ a_5149_4721# 3.16e-19
C1442 a_5179_3311# a_6043_3677# 0.032244f
C1443 net4 a_3215_2999# 0.130038f
C1444 a_5786_3423# a_5618_3677# 0.239923f
C1445 _24_ _25_ 0.095329f
C1446 net7 a_5801_4233# 1.38e-19
C1447 a_2401_4399# a_1849_3861# 5.5e-20
C1448 a_3267_4667# _06_ 1.81e-20
C1449 _11_ a_5149_4721# 0.042839f
C1450 a_5345_3311# a_5505_2388# 1.2e-20
C1451 a_4520_4373# a_4454_4649# 0.221119f
C1452 net6 a_6817_3861# 1.27e-19
C1453 clknet_1_1__leaf_clk _15_ 0.471647f
C1454 _24_ _09_ 0.151845f
C1455 a_3849_2388# a_4585_2388# 2.31e-20
C1456 a_7171_2767# VPWR 0.191262f
C1457 a_4779_5161# net6 0.001597f
C1458 net9 a_5891_3133# 6.97e-19
C1459 a_4714_5309# VPWR 7.65e-20
C1460 a_4811_3861# a_5345_3311# 0.003047f
C1461 _19_ _16_ 0.001191f
C1462 clknet_1_0__leaf_clk a_2431_7497# 0.024273f
C1463 a_4977_3861# a_5179_3311# 0.003672f
C1464 clknet_0_clk a_4495_5175# 0.00222f
C1465 _04_ a_3433_4175# 0.002919f
C1466 a_7683_3579# a_7939_2223# 3.35e-20
C1467 a_7258_3423# VPWR 0.186041f
C1468 _22_ a_5179_3311# 0.019806f
C1469 net1 a_2295_7337# 0.002755f
C1470 _07_ a_4259_3311# 1.81e-20
C1471 _24_ a_7515_3855# 0.013075f
C1472 _17_ a_5149_4721# 7.49e-19
C1473 a_1457_2388# counter[0] 0.109791f
C1474 net3 _02_ 0.031079f
C1475 a_2235_4399# a_4287_4399# 9.88e-21
C1476 _21_ a_2991_3579# 1.79e-21
C1477 _04_ a_3225_4399# 6.79e-19
C1478 _03_ a_2991_3579# 3.08e-19
C1479 _04_ a_2589_4399# 0.126198f
C1480 a_4399_5175# a_4714_5309# 7.84e-20
C1481 a_4349_3855# _20_ 1.05e-19
C1482 a_2235_4399# a_2769_4765# 0.002698f
C1483 a_1959_3311# a_2823_3677# 0.032244f
C1484 a_6651_3861# a_6817_3311# 2.64e-19
C1485 _05_ _24_ 2.08e-20
C1486 _11_ a_6623_3133# 7.08e-19
C1487 net7 a_5786_3423# 0.005145f
C1488 _11_ _24_ 4.57e-19
C1489 net3 a_1915_7351# 0.115857f
C1490 net2 a_2235_6575# 0.165774f
C1491 net4 a_3433_4175# 5.3e-19
C1492 net6 a_4259_3311# 0.005791f
C1493 a_4779_5161# _06_ 0.002324f
C1494 net7 a_6651_5309# 5.71e-19
C1495 net6 a_2041_4649# 4.71e-21
C1496 net1 a_2125_8527# 0.003019f
C1497 a_2524_3311# net5 3e-19
C1498 a_2561_9514# _00_ 4.57e-22
C1499 _14_ a_2745_2388# 4.42e-19
C1500 clknet_1_0__leaf_clk net6 6.56e-20
C1501 a_2842_4511# a_3267_4667# 1.28e-19
C1502 net4 a_2589_4399# 0.011292f
C1503 a_2401_4399# a_3099_4765# 0.194203f
C1504 clknet_1_0__leaf_clk a_1845_5461# 1.67275f
C1505 _17_ _24_ 0.004444f
C1506 clknet_1_1__leaf_clk a_6651_3861# 0.285659f
C1507 _14_ a_2547_3855# 2.97e-21
C1508 net9 counter[7] 0.006102f
C1509 a_4495_5175# clknet_1_1__leaf_clk 1.54e-20
C1510 a_4915_5321# _16_ 2.16e-20
C1511 a_7077_2767# a_7171_2767# 0.062574f
C1512 a_2614_2883# a_2745_2388# 0.002548f
C1513 a_7258_3829# net10 2.56e-19
C1514 a_7723_2741# a_7941_3087# 0.007234f
C1515 a_5213_4664# a_4995_4399# 0.004465f
C1516 a_2715_3829# a_2125_3311# 0.00183f
C1517 _20_ a_5345_3311# 0.003428f
C1518 _13_ _02_ 0.053355f
C1519 _10_ a_2695_6575# 0.423817f
C1520 a_2235_6575# _11_ 0.005192f
C1521 _23_ counter[8] 9.18e-19
C1522 _15_ a_6651_3861# 0.069151f
C1523 a_7258_3423# a_7077_2767# 3.15e-19
C1524 a_3267_4667# VPWR 0.386139f
C1525 net3 net5 9.15e-21
C1526 a_4495_5175# _15_ 1.09e-20
C1527 net7 a_4995_4399# 2.13e-20
C1528 a_6043_3677# _09_ 1.4e-19
C1529 a_4329_5461# _16_ 4.51e-19
C1530 net8 a_5250_3855# 0.003635f
C1531 _25_ _08_ 0.208467f
C1532 clknet_1_1__leaf_clk a_3831_3339# 2.67e-20
C1533 net9 a_5618_3677# 0.003585f
C1534 a_5001_3311# VPWR 9.47e-20
C1535 a_6651_3311# a_7345_2388# 4.75e-20
C1536 _08_ _09_ 0.013938f
C1537 _09_ net11 0.071633f
C1538 _16_ a_2936_2767# 0.00427f
C1539 _23_ a_5179_3311# 3.56e-21
C1540 net9 a_7599_3677# 1.5e-19
C1541 _15_ a_3831_3339# 0.22097f
C1542 _22_ _09_ 0.009594f
C1543 net1 _10_ 0.033245f
C1544 a_6817_3861# VPWR 0.31297f
C1545 net9 a_5213_4664# 0.122363f
C1546 _08_ a_7515_3855# 0.013878f
C1547 _11_ a_6043_3677# 0.045045f
C1548 a_6375_5309# a_6545_5309# 0.001675f
C1549 a_1915_7815# a_2011_7637# 0.310858f
C1550 a_4779_5161# VPWR 0.438492f
C1551 a_2125_8207# a_2302_7937# 0.001655f
C1552 a_5814_4399# a_5345_3311# 1.98e-20
C1553 clknet_0_clk _21_ 4.86e-19
C1554 a_5675_3855# a_6817_3861# 8.68e-20
C1555 a_2547_3855# a_2673_4233# 0.006169f
C1556 _11_ a_6425_2388# 2.18e-19
C1557 _23_ a_7005_3311# 0.012973f
C1558 a_2235_4399# a_2401_4399# 0.966818f
C1559 _11_ _08_ 1.44e-20
C1560 _05_ a_4977_3861# 2.65e-21
C1561 _14_ a_1683_3861# 0.001276f
C1562 clknet_1_0__leaf_clk a_2842_4511# 5.16e-19
C1563 net7 net9 0.742565f
C1564 _11_ a_4977_3861# 8.46e-20
C1565 net2 a_2125_3311# 3.95e-20
C1566 net8 a_5599_2741# 0.1454f
C1567 _05_ _22_ 0.001519f
C1568 a_4399_5175# a_4779_5161# 0.048635f
C1569 _11_ net11 2.31e-19
C1570 net2 a_2295_7637# 4.59e-19
C1571 _11_ _22_ 0.420712f
C1572 a_4259_3311# a_4413_3311# 0.004009f
C1573 net6 a_5333_5321# 9.51e-20
C1574 net5 a_4585_2388# 0.001724f
C1575 _16_ a_4349_3855# 0.008193f
C1576 a_4259_3311# VPWR 0.211123f
C1577 a_2041_4649# VPWR 0.006535f
C1578 net6 a_2290_3829# 6.4e-20
C1579 clknet_0_clk a_5135_5309# 4.62e-19
C1580 a_4329_5461# a_5418_3829# 8.05e-21
C1581 _17_ a_4977_3861# 1.22e-20
C1582 clknet_1_0__leaf_clk VPWR 3.74806f
C1583 a_2840_3087# VPWR 0.007674f
C1584 a_1915_7815# a_2011_7351# 6.79e-19
C1585 a_2011_7637# a_1915_7351# 6.79e-19
C1586 a_1845_5461# a_2290_3829# 3.17e-20
C1587 _17_ _22_ 1.76e-19
C1588 net7 a_4454_4649# 3.79e-19
C1589 clknet_1_1__leaf_clk _21_ 0.038033f
C1590 a_5149_4721# a_4995_4399# 0.049785f
C1591 a_7258_3423# a_7171_2767# 5.71e-20
C1592 _11_ a_2125_3311# 0.03376f
C1593 _22_ a_5795_3133# 0.002279f
C1594 a_6817_3311# a_7090_3677# 0.078545f
C1595 a_2295_7637# _11_ 8.58e-21
C1596 _11_ a_3215_2999# 0.159397f
C1597 _15_ _21_ 0.054317f
C1598 _16_ a_5345_3311# 4.88e-21
C1599 net2 a_2302_7241# 8.79e-19
C1600 a_1875_8207# a_1915_7815# 1.32e-19
C1601 _00_ a_1957_8207# 6.18e-19
C1602 net8 _07_ 0.001136f
C1603 _23_ _25_ 0.0063f
C1604 net7 a_5997_3133# 0.001525f
C1605 a_2398_3677# a_2313_3311# 0.037333f
C1606 _16_ a_2745_2388# 4.24e-19
C1607 a_2125_3311# a_2907_3677# 3.14e-19
C1608 _02_ a_1505_3855# 0.01416f
C1609 net7 a_7019_4943# 6.19e-19
C1610 a_2235_4399# a_2991_3579# 3.85e-19
C1611 _04_ a_2398_3677# 3.52e-21
C1612 a_5871_5162# net6 0.019537f
C1613 net8 a_7185_3855# 7.49e-20
C1614 _23_ _09_ 0.130147f
C1615 a_1915_7351# a_2011_7351# 0.310858f
C1616 net3 _12_ 0.271994f
C1617 a_2631_3855# VPWR 0.007439f
C1618 clknet_1_0__leaf_clk a_2823_3677# 6.12e-19
C1619 clknet_1_1__leaf_clk a_7090_3677# 3.02e-19
C1620 net5 a_2471_2741# 0.006016f
C1621 _16_ a_2547_3855# 1.35e-19
C1622 a_7939_2223# counter[8] 0.006251f
C1623 a_3799_4943# a_3979_4943# 0.185422f
C1624 net10 a_7515_3677# 0.003817f
C1625 net6 net8 0.806426f
C1626 net2 _00_ 0.002662f
C1627 net5 a_2949_3311# 6.03e-19
C1628 a_4811_3861# a_7005_3855# 2.33e-21
C1629 a_5149_4721# net9 0.170073f
C1630 net1 a_2502_7637# 0.002893f
C1631 net6 a_7199_4943# 7.38e-20
C1632 net3 _14_ 0.471315f
C1633 _05_ _23_ 9.36e-20
C1634 a_2502_7396# a_2695_6575# 2.48e-20
C1635 _12_ a_2253_7119# 1.13e-19
C1636 a_2302_7241# _11_ 4.06e-19
C1637 _15_ a_7090_3677# 0.001788f
C1638 net4 a_2398_3677# 0.004091f
C1639 net2 a_2317_6575# 6.45e-19
C1640 _11_ _23_ 0.090724f
C1641 a_7090_3855# a_7185_3855# 0.007724f
C1642 a_7258_3829# a_7599_3855# 9.73e-19
C1643 net8 counter[9] 1.68e-20
C1644 a_5786_3423# a_6043_3677# 0.036838f
C1645 a_4495_5175# _21_ 9.57e-19
C1646 a_5345_3311# a_5533_3311# 0.095025f
C1647 _11_ a_3225_4399# 8.02e-19
C1648 a_5179_3311# a_5713_3677# 0.002698f
C1649 net3 a_2614_2883# 8.22e-19
C1650 a_2401_4399# a_2122_3855# 0.001124f
C1651 _11_ a_2589_4399# 0.020189f
C1652 net8 _06_ 0.209874f
C1653 a_4454_4649# a_5149_4721# 5.89e-19
C1654 a_6375_5309# clk 1.34e-19
C1655 a_8109_2767# VPWR 0.009314f
C1656 _17_ _23_ 0.082072f
C1657 a_4585_2388# a_5505_2388# 1.37e-20
C1658 a_4986_5220# net6 6.81e-19
C1659 a_3245_3855# a_2991_3579# 0.001352f
C1660 _00_ _11_ 0.003231f
C1661 a_5418_3829# a_5345_3311# 0.001607f
C1662 _24_ net9 0.165357f
C1663 a_4811_3861# a_5618_3677# 4.58e-19
C1664 a_4977_3861# a_5786_3423# 6.74e-19
C1665 a_5250_3855# a_5179_3311# 2.14e-19
C1666 a_5333_5321# VPWR 0.085296f
C1667 a_6043_3677# a_6169_3311# 0.006169f
C1668 clknet_0_clk a_4786_5065# 0.025079f
C1669 a_2290_3829# VPWR 0.200136f
C1670 a_7683_3579# VPWR 0.462064f
C1671 _22_ a_5786_3423# 0.001181f
C1672 a_5814_4399# clk 1.27e-19
C1673 net1 a_2502_7396# 1.33e-19
C1674 a_4329_5461# a_4287_4399# 1.78e-20
C1675 _11_ a_2317_6575# 1.17e-19
C1676 _13_ _14_ 0.074354f
C1677 a_7258_3829# a_6817_3311# 2.96e-21
C1678 a_6817_3861# a_7258_3423# 2.96e-21
C1679 _03_ a_3831_3339# 2.2e-20
C1680 a_1959_3311# a_4259_3311# 1.62e-21
C1681 a_6651_3861# a_7090_3677# 1.73e-19
C1682 _11_ a_6825_3133# 0.001561f
C1683 a_4220_3829# a_4811_3861# 0.044245f
C1684 _22_ a_6169_3311# 7.63e-20
C1685 net3 a_2295_7337# 0.008811f
C1686 clknet_1_1__leaf_clk a_6127_3677# 1.62e-19
C1687 net7 a_6211_3579# 0.064911f
C1688 clknet_1_0__leaf_clk a_1959_3311# 0.293401f
C1689 _16_ a_1683_3861# 0.001516f
C1690 a_1959_3311# a_2840_3087# 3.11e-19
C1691 a_5213_4664# a_4811_3861# 0.004179f
C1692 net7 a_5505_2388# 0.201574f
C1693 a_4986_5220# _06_ 2.41e-19
C1694 net6 _04_ 0.050232f
C1695 net10 a_6651_3311# 0.001924f
C1696 a_7641_4233# _09_ 1.66e-19
C1697 a_1845_5461# _04_ 0.00168f
C1698 _18_ a_4443_4175# 6.01e-19
C1699 a_1915_7351# a_2235_6575# 3.66e-19
C1700 a_2302_7241# a_2849_7497# 0.099725f
C1701 a_1582_7439# _12_ 0.001776f
C1702 _16_ a_2037_3855# 4.26e-21
C1703 a_2502_7396# a_2651_7485# 0.005525f
C1704 clknet_1_1__leaf_clk a_7258_3829# 5.16e-19
C1705 net7 a_4811_3861# 0.088061f
C1706 a_2842_4511# net8 1.22e-20
C1707 a_5179_3311# a_5599_2741# 0.009169f
C1708 net1 a_2389_6575# 0.002601f
C1709 a_4786_5065# clknet_1_1__leaf_clk 0.013843f
C1710 _22_ a_4995_4399# 9.75e-19
C1711 a_7515_3855# a_7641_4233# 0.006169f
C1712 a_7683_3829# net10 0.084593f
C1713 a_4349_4175# a_4349_3855# 6.96e-20
C1714 a_7723_2741# a_7753_2767# 0.025037f
C1715 net6 net4 0.008308f
C1716 _20_ a_5618_3677# 9.2e-20
C1717 _18_ a_3183_4765# 1.72e-19
C1718 a_2547_3855# a_2566_3423# 3.73e-19
C1719 a_5871_5162# VPWR 0.209324f
C1720 a_2715_3829# a_2398_3677# 0.005602f
C1721 a_4520_4373# _16_ 0.035189f
C1722 a_7019_4943# _24_ 0.095435f
C1723 net8 a_4413_3311# 8.5e-20
C1724 a_1845_5461# net4 4.87e-19
C1725 net11 a_7641_3311# 3e-19
C1726 _15_ a_7258_3829# 4.57e-19
C1727 a_3215_3829# a_3215_2999# 8.07e-19
C1728 a_2614_2883# counter[2] 6.46e-19
C1729 a_4786_5065# _15_ 1.53e-20
C1730 net8 VPWR 1.78891f
C1731 a_5814_4399# a_7005_3855# 9.53e-19
C1732 _18_ net6 0.081404f
C1733 a_3979_4943# _19_ 0.082191f
C1734 a_4220_3829# _20_ 3.36e-20
C1735 a_2011_7637# _12_ 1.23e-19
C1736 a_7199_4943# VPWR 0.178246f
C1737 _00_ a_2849_7497# 0.001531f
C1738 clknet_1_1__leaf_clk a_4767_3463# 0.050301f
C1739 clknet_0_clk a_3799_4943# 2.32e-20
C1740 net8 a_5675_3855# 0.00311f
C1741 a_5744_3311# VPWR 1.42e-19
C1742 net9 a_6043_3677# 0.031858f
C1743 a_4399_5175# net8 1.16e-19
C1744 net6 a_3601_3855# 7.79e-20
C1745 net9 a_6425_2388# 7.77e-19
C1746 _08_ net9 0.003243f
C1747 _14_ a_2471_2741# 0.134293f
C1748 net9 net11 0.055197f
C1749 net9 a_4977_3861# 0.002182f
C1750 net7 _20_ 0.035834f
C1751 _15_ a_4767_3463# 2.8e-19
C1752 a_7090_3855# VPWR 0.247111f
C1753 a_1915_7815# a_2295_7637# 0.048748f
C1754 _18_ _06_ 3.12e-20
C1755 net9 _22_ 0.369389f
C1756 a_2011_7637# a_2302_7937# 0.194892f
C1757 _24_ a_7216_4233# 9.29e-19
C1758 _07_ a_5179_3311# 0.112051f
C1759 a_4986_5220# VPWR 0.266088f
C1760 net3 _16_ 6.72e-19
C1761 counter[9] counter[8] 0.299988f
C1762 a_2471_2741# a_2614_2883# 0.221119f
C1763 _15_ a_3389_3105# 1.81e-19
C1764 a_3215_3829# a_3433_4175# 0.007234f
C1765 a_6651_3861# a_7258_3829# 0.141453f
C1766 a_2235_4399# a_2674_4765# 0.269567f
C1767 _04_ a_2842_4511# 0.04931f
C1768 net3 _10_ 0.003052f
C1769 _05_ a_5250_3855# 6.05e-21
C1770 a_2011_7351# _12_ 0.036321f
C1771 net6 a_5179_3311# 0.083542f
C1772 a_4495_5175# a_4786_5065# 0.192261f
C1773 clknet_1_0__leaf_clk a_3267_4667# 1.77e-20
C1774 _11_ a_5250_3855# 2.99e-20
C1775 a_5149_4721# a_4811_3861# 0.001396f
C1776 net8 a_7077_2767# 4.33e-20
C1777 a_1683_3861# a_2566_3423# 0.001786f
C1778 net2 a_2431_7663# 3.46e-19
C1779 net4 counter[3] 6.72e-19
C1780 a_2290_3829# a_1959_3311# 0.001425f
C1781 a_4767_3463# a_4929_3311# 0.004009f
C1782 a_1849_3861# _03_ 1.23e-19
C1783 clknet_1_1__leaf_clk a_3245_3855# 7.11e-20
C1784 _14_ a_1505_3855# 6.31e-19
C1785 a_2313_3311# VPWR 0.083158f
C1786 net6 counter[4] 0.003133f
C1787 a_6651_3311# a_6427_2741# 2.81e-20
C1788 net7 a_6375_5309# 0.168744f
C1789 net6 a_2715_3829# 6.37e-19
C1790 clknet_0_clk a_4737_4943# 2.01e-19
C1791 _04_ VPWR 0.27578f
C1792 net4 a_2842_4511# 0.034264f
C1793 _17_ a_5250_3855# 9.6e-21
C1794 a_1875_8207# _12_ 1.27e-21
C1795 net7 a_5814_4399# 0.037674f
C1796 a_3917_3105# VPWR 0.002731f
C1797 a_2011_7637# a_2295_7337# 9.64e-20
C1798 a_2302_7937# a_2011_7351# 1.53e-19
C1799 a_2561_9514# VPWR 0.305606f
C1800 _22_ net5 4.26e-20
C1801 a_4495_5175# a_4767_3463# 5.98e-21
C1802 _18_ a_2842_4511# 1.41e-19
C1803 _24_ a_7216_3311# 6.57e-19
C1804 _11_ a_2398_3677# 0.00274f
C1805 _22_ a_5997_3133# 0.002069f
C1806 a_6817_3311# a_7515_3677# 0.194892f
C1807 a_7258_3423# a_7683_3579# 1.28e-19
C1808 _11_ a_5599_2741# 2.67e-19
C1809 net4 VPWR 1.18326f
C1810 net8 a_5376_4233# 4.88e-19
C1811 net2 a_2431_7497# 8.2e-21
C1812 _16_ a_5618_3677# 7.37e-22
C1813 _00_ a_1915_7815# 0.001095f
C1814 a_1875_8207# a_2302_7937# 0.00324f
C1815 net7 a_6719_3133# 5.42e-19
C1816 _18_ VPWR 0.686881f
C1817 a_2566_3423# a_2524_3311# 4.62e-19
C1818 a_3099_4765# _21_ 8.88e-21
C1819 a_2125_3311# net5 8.3e-19
C1820 net8 a_4382_4649# 0.001644f
C1821 _04_ a_2823_3677# 0.001409f
C1822 a_1499_7119# VPWR 0.229121f
C1823 a_3601_3855# VPWR 0.009139f
C1824 a_1915_7351# a_2302_7241# 0.034054f
C1825 _23_ net9 0.065132f
C1826 a_2011_7351# a_2295_7337# 0.030894f
C1827 clknet_1_1__leaf_clk a_7515_3677# 2.2e-19
C1828 _16_ counter[2] 3.86e-19
C1829 clknet_1_0__leaf_clk a_2041_4649# 0.001585f
C1830 _16_ a_4220_3829# 0.01721f
C1831 _15_ a_3917_3339# 7.85e-19
C1832 _08_ a_7216_4233# 0.001882f
C1833 net5 a_3215_2999# 0.081136f
C1834 clknet_0_clk _19_ 0.038005f
C1835 _18_ a_4399_5175# 0.006776f
C1836 VPWR counter[8] 0.228646f
C1837 a_7345_2388# counter[7] 0.110188f
C1838 a_4811_3861# a_5345_3855# 0.001632f
C1839 a_4585_2388# counter[5] 4.98e-19
C1840 a_5213_4664# _16_ 0.060109f
C1841 a_5599_2741# a_5795_3133# 0.00119f
C1842 net1 a_2253_8029# 8.57e-19
C1843 _19_ a_4069_5309# 8.17e-20
C1844 net6 _25_ 2.22e-20
C1845 counter[3] counter[4] 0.077431f
C1846 _12_ a_2235_6575# 0.001375f
C1847 _01_ a_2695_6575# 0.014882f
C1848 net8 a_7171_2767# 6.89e-20
C1849 net6 _09_ 1.5e-20
C1850 _11_ a_4443_4175# 5.64e-19
C1851 net4 a_2823_3677# 0.022715f
C1852 net3 a_2566_3423# 3.22e-20
C1853 net7 _16_ 5.07e-19
C1854 _16_ a_5436_4399# 3.12e-19
C1855 a_6211_3579# a_6043_3677# 0.310858f
C1856 a_5618_3677# a_5533_3311# 0.037333f
C1857 a_2431_7663# a_2651_7663# 4.62e-19
C1858 net7 a_5759_3855# 0.001255f
C1859 a_2842_4511# a_2715_3829# 0.002135f
C1860 a_4786_5065# _21_ 0.001538f
C1861 _11_ _07_ 0.161717f
C1862 a_2401_4399# a_2547_3855# 3.42e-19
C1863 _13_ counter[0] 3.39e-20
C1864 a_4520_4373# a_4287_4399# 0.005961f
C1865 _11_ a_3183_4765# 0.002344f
C1866 a_5179_3311# VPWR 0.727748f
C1867 a_6211_3579# a_6425_2388# 2.93e-21
C1868 net7 counter[5] 0.002945f
C1869 a_4329_5461# a_5165_3855# 2.19e-20
C1870 a_7199_4943# a_7258_3423# 1.02e-20
C1871 _17_ a_4443_4175# 3.09e-20
C1872 a_1825_2388# VPWR 0.272145f
C1873 _05_ net6 0.03493f
C1874 _16_ a_2471_2741# 0.184103f
C1875 a_4413_3311# counter[4] 4.17e-20
C1876 clknet_1_1__leaf_clk _19_ 0.060342f
C1877 a_5505_2388# a_6425_2388# 1.37e-20
C1878 a_5843_3829# a_5345_3311# 0.002689f
C1879 a_5675_3855# a_5179_3311# 0.004606f
C1880 a_6457_5309# VPWR 0.001434f
C1881 a_6651_3311# a_6817_3311# 0.970499f
C1882 _17_ _07_ 3.97e-20
C1883 _11_ net6 2.01574f
C1884 clknet_1_0__leaf_clk a_2631_3855# 3.7e-19
C1885 clknet_0_clk a_4915_5321# 0.003343f
C1886 net1 _01_ 1.96e-19
C1887 VPWR counter[4] 0.454642f
C1888 a_2715_3829# VPWR 0.421579f
C1889 a_4977_3861# a_5505_2388# 7.09e-22
C1890 _22_ a_6211_3579# 3.11e-19
C1891 a_7005_3311# VPWR 0.079695f
C1892 _11_ a_1845_5461# 0.055744f
C1893 _08_ a_4811_3861# 3.42e-20
C1894 a_6375_5309# _24_ 4.18e-19
C1895 _21_ a_4767_3463# 0.011629f
C1896 a_1875_8207# a_2125_8527# 0.007234f
C1897 _23_ a_7019_4943# 0.213625f
C1898 _22_ a_5505_2388# 8.8e-19
C1899 a_6651_3861# a_7515_3677# 1.29e-19
C1900 a_4811_3861# a_4977_3861# 0.961627f
C1901 a_7258_3829# a_7090_3677# 3.15e-19
C1902 a_4495_5175# a_4737_4943# 0.008508f
C1903 a_1959_3311# a_2313_3311# 0.062224f
C1904 a_4779_5161# a_5333_5321# 0.057611f
C1905 _19_ _15_ 6.2e-22
C1906 a_7090_3855# a_7258_3423# 3.15e-19
C1907 a_2235_4399# _03_ 4.31e-20
C1908 _04_ a_1959_3311# 2.08e-19
C1909 _22_ a_4811_3861# 0.016414f
C1910 a_5213_4664# a_5418_3829# 1.06e-19
C1911 net7 a_5533_3311# 4.68e-19
C1912 net3 a_2502_7396# 3.02e-19
C1913 clknet_1_1__leaf_clk a_6651_3311# 0.306202f
C1914 _17_ net6 0.277113f
C1915 _03_ a_3389_3105# 1.17e-19
C1916 _24_ a_5814_4399# 0.025563f
C1917 clknet_0_clk a_4329_5461# 1.74729f
C1918 a_3831_3339# a_3917_3339# 0.006584f
C1919 _15_ a_7619_5162# 8.98e-20
C1920 _11_ _06_ 0.020042f
C1921 clknet_1_1__leaf_clk a_7683_3829# 9.45e-20
C1922 net7 a_5418_3829# 0.040813f
C1923 _15_ a_6651_3311# 0.02569f
C1924 a_2295_7337# a_2235_6575# 4.35e-19
C1925 a_2431_7497# a_2849_7497# 3.39e-19
C1926 a_3267_4667# net8 5.45e-19
C1927 net4 a_1959_3311# 0.008383f
C1928 a_5786_3423# a_5599_2741# 3.07e-19
C1929 a_4915_5321# clknet_1_1__leaf_clk 1.17e-20
C1930 a_1957_8207# VPWR 0.008578f
C1931 net8 a_5001_3311# 5.79e-19
C1932 _18_ a_4382_4649# 0.00112f
C1933 _20_ a_6043_3677# 1.2e-20
C1934 _17_ _06_ 0.001225f
C1935 _23_ a_7216_4233# 9.59e-19
C1936 a_2401_4399# a_1683_3861# 9.16e-19
C1937 clknet_1_0__leaf_clk a_2290_3829# 0.01796f
C1938 a_5149_4721# _16_ 0.113309f
C1939 a_2235_4399# a_1849_3861# 1.36e-19
C1940 _07_ a_5801_4233# 5.27e-19
C1941 a_7515_3677# a_7723_2741# 0.003595f
C1942 _15_ a_7683_3829# 1.61e-19
C1943 a_4915_5321# _15_ 2.35e-21
C1944 net3 a_2389_6575# 8.45e-20
C1945 a_4495_5175# _19_ 0.046625f
C1946 a_4779_5161# a_5871_5162# 5.23e-20
C1947 _11_ counter[3] 1.03e-19
C1948 _25_ VPWR 0.22908f
C1949 a_2295_7637# _12_ 2.52e-19
C1950 a_4329_5461# clknet_1_1__leaf_clk 0.002451f
C1951 net2 VPWR 2.41286f
C1952 net8 a_6817_3861# 5.19e-19
C1953 _09_ VPWR 0.262387f
C1954 _22_ _20_ 2.69e-20
C1955 a_7619_5162# a_6651_3861# 7.7e-20
C1956 _14_ a_2125_3311# 5.98e-19
C1957 a_7199_4943# a_6817_3861# 6.98e-21
C1958 a_4779_5161# net8 0.001356f
C1959 net7 a_3831_3105# 2.04e-20
C1960 net9 a_7939_2223# 0.003439f
C1961 _11_ a_2842_4511# 0.032361f
C1962 a_2401_4399# a_4520_4373# 8.39e-21
C1963 a_6651_3861# a_6651_3311# 0.037572f
C1964 _14_ a_3215_2999# 0.112679f
C1965 _23_ a_6211_3579# 1.37e-20
C1966 net9 a_5250_3855# 6.38e-21
C1967 a_4329_5461# _15_ 2.08e-20
C1968 a_2566_3423# a_2471_2741# 1.66e-20
C1969 a_7515_3855# VPWR 0.233266f
C1970 a_2125_3311# a_2614_2883# 0.010312f
C1971 _07_ a_5786_3423# 0.004454f
C1972 a_2302_7937# a_2295_7637# 0.966391f
C1973 a_1915_7815# a_2431_7663# 1.28e-19
C1974 _11_ a_4413_3311# 0.001879f
C1975 _05_ VPWR 0.240335f
C1976 a_5814_4399# a_6043_3677# 0.001605f
C1977 _11_ VPWR 5.18499f
C1978 a_2290_3829# a_2631_3855# 9.73e-19
C1979 a_2122_3855# a_2217_3855# 0.007724f
C1980 a_6817_3861# a_7090_3855# 0.078545f
C1981 _17_ a_2842_4511# 2.52e-22
C1982 a_6651_3861# a_7683_3829# 0.048748f
C1983 a_4220_3829# a_4349_4175# 0.010132f
C1984 a_2566_3423# a_2949_3311# 4.67e-20
C1985 _23_ a_7216_3311# 6.82e-19
C1986 net8 a_4259_3311# 7.44e-19
C1987 _23_ a_4811_3861# 1.94e-21
C1988 a_2302_7241# _12_ 0.206007f
C1989 a_4737_4943# _21_ 1.26e-19
C1990 a_2235_4399# a_3099_4765# 0.030894f
C1991 _04_ a_3267_4667# 0.003723f
C1992 _08_ a_5814_4399# 0.011527f
C1993 a_4495_5175# a_4915_5321# 0.036838f
C1994 a_4399_5175# _05_ 1.85e-19
C1995 a_4779_5161# a_4986_5220# 0.260055f
C1996 net6 a_5786_3423# 6.78e-21
C1997 _11_ a_5675_3855# 7.12e-21
C1998 a_5149_4721# a_5418_3829# 1e-18
C1999 clknet_0_clk a_5345_3311# 3.43e-21
C2000 _11_ a_4399_5175# 8.65e-19
C2001 net6 a_3849_2388# 3.58e-19
C2002 a_2715_3829# a_1959_3311# 0.00142f
C2003 a_2122_3855# _03_ 0.001262f
C2004 a_5814_4399# _22_ 8.12e-19
C2005 clknet_1_1__leaf_clk a_4349_3855# 0.001857f
C2006 _17_ VPWR 2.38225f
C2007 a_2235_6575# _10_ 0.107891f
C2008 _09_ a_7077_2767# 0.001692f
C2009 a_5843_3829# clk 1.4e-22
C2010 a_2907_3677# VPWR 0.004797f
C2011 clknet_0_clk a_6545_5309# 9.17e-20
C2012 net6 a_3215_3829# 0.080758f
C2013 net4 a_3267_4667# 7.5e-19
C2014 a_7005_3855# net10 6.3e-20
C2015 net9 a_5599_2741# 0.125008f
C2016 _17_ a_5675_3855# 8.73e-21
C2017 _00_ _12_ 4.17e-19
C2018 a_2295_7637# a_2295_7337# 0.040702f
C2019 _24_ a_7345_2388# 0.00116f
C2020 a_5345_3311# a_6817_3311# 0.002814f
C2021 a_2302_7937# a_2302_7241# 0.027204f
C2022 net10 counter[7] 4.65e-20
C2023 a_4329_5461# a_4495_5175# 0.017149f
C2024 _17_ a_4399_5175# 0.0702f
C2025 _15_ a_4349_3855# 0.046541f
C2026 a_4786_5065# a_4767_3463# 2.42e-19
C2027 a_7515_3677# a_7753_2767# 3.93e-20
C2028 _18_ a_3267_4667# 0.001543f
C2029 a_7683_3829# a_7723_2741# 1.35e-20
C2030 _11_ a_2823_3677# 0.045224f
C2031 a_7258_3423# a_7005_3311# 3.39e-19
C2032 _22_ a_6719_3133# 6.12e-20
C2033 net6 a_4995_4399# 0.00514f
C2034 a_2849_7663# a_2695_6575# 9.03e-20
C2035 a_2651_7663# VPWR 0.003202f
C2036 _11_ a_7077_2767# 0.054652f
C2037 a_3099_4765# a_3245_3855# 1.65e-19
C2038 a_1849_3861# a_2122_3855# 0.078737f
C2039 clknet_1_1__leaf_clk a_5345_3311# 0.486375f
C2040 _06_ a_3215_3829# 1.6e-20
C2041 _19_ _21_ 7.87e-20
C2042 _00_ a_2302_7937# 0.208988f
C2043 a_2823_3677# a_2907_3677# 0.008508f
C2044 a_2398_3677# net5 4.4e-19
C2045 a_2849_7497# VPWR 0.074934f
C2046 a_2295_7337# a_2302_7241# 0.969092f
C2047 clknet_1_0__leaf_clk a_2313_3311# 0.003207f
C2048 _13_ a_2401_4399# 7.99e-20
C2049 a_1915_7351# a_2431_7497# 1.28e-19
C2050 _16_ a_4977_3861# 9.89e-20
C2051 clknet_1_0__leaf_clk _04_ 0.005301f
C2052 net5 a_5599_2741# 1.18e-20
C2053 _15_ a_5345_3311# 2.57e-20
C2054 net2 a_1959_3311# 5.19e-20
C2055 _18_ a_4779_5161# 6.58e-19
C2056 _22_ _16_ 0.135659f
C2057 a_1457_2388# counter[1] 0.057818f
C2058 a_5675_3855# a_5801_4233# 0.006169f
C2059 a_5599_2741# a_5997_3133# 0.005781f
C2060 a_4977_3861# a_5759_3855# 3.14e-19
C2061 net9 _07_ 0.03749f
C2062 a_3849_2388# counter[3] 0.110188f
C2063 _06_ a_4995_4399# 0.046896f
C2064 net10 a_7599_3677# 3.08e-19
C2065 net1 a_2849_7663# 5.53e-20
C2066 a_6375_5309# _23_ 0.026998f
C2067 a_4495_5175# a_4349_3855# 4.21e-21
C2068 _19_ a_5135_5309# 2.79e-19
C2069 _15_ a_2547_3855# 7.5e-20
C2070 net6 _02_ 0.001309f
C2071 _23_ a_5814_4399# 0.042503f
C2072 a_5179_3311# a_5001_3311# 1.43e-19
C2073 net6 net9 0.566537f
C2074 clknet_1_0__leaf_clk net4 0.158995f
C2075 a_4915_5321# _21_ 1.21e-19
C2076 _00_ a_2295_7337# 8.76e-20
C2077 net7 net10 6.54e-19
C2078 a_2674_4765# a_2547_3855# 0.002298f
C2079 net4 a_2840_3087# 0.01239f
C2080 _09_ a_7171_2767# 2.04e-21
C2081 a_5786_3423# VPWR 0.183641f
C2082 _11_ a_4382_4649# 0.002546f
C2083 _16_ a_2125_3311# 2.51e-21
C2084 net1 enable 0.067176f
C2085 _11_ a_1959_3311# 0.005486f
C2086 _16_ a_3215_2999# 0.01632f
C2087 a_6425_2388# a_7345_2388# 1.37e-20
C2088 a_3849_2388# VPWR 0.316408f
C2089 a_6651_3311# a_7090_3677# 0.273138f
C2090 a_5843_3829# a_5618_3677# 0.003655f
C2091 a_6651_5309# VPWR 0.002272f
C2092 net9 counter[9] 5.19e-19
C2093 _09_ a_7258_3423# 0.039926f
C2094 a_5675_3855# a_5786_3423# 0.001204f
C2095 clknet_1_0__leaf_clk a_1499_7119# 3.26e-19
C2096 a_3215_3829# VPWR 0.252112f
C2097 net11 a_7345_2388# 3.2e-20
C2098 a_6169_3311# VPWR 2.75e-19
C2099 _22_ a_5533_3311# 0.012798f
C2100 net6 a_4454_4649# 0.074355f
C2101 a_5250_3855# a_5505_2388# 3e-19
C2102 a_4779_5161# a_5179_3311# 2.6e-21
C2103 _08_ a_5418_3829# 9.82e-20
C2104 _06_ net9 0.017291f
C2105 _17_ a_4382_4649# 0.002503f
C2106 a_4329_5461# _21_ 0.001038f
C2107 _22_ a_7345_2388# 1.85e-19
C2108 a_2125_8527# _00_ 0.002065f
C2109 clknet_0_clk a_4520_4373# 7.65e-20
C2110 a_4986_5220# a_5333_5321# 0.037333f
C2111 a_4786_5065# a_4737_4943# 4.04e-19
C2112 a_4977_3861# a_5418_3829# 0.110715f
C2113 a_4915_5321# a_5135_5309# 4.62e-19
C2114 a_6817_3861# a_7005_3311# 1.41e-20
C2115 a_4811_3861# a_5250_3855# 0.260055f
C2116 _11_ a_7171_2767# 0.039972f
C2117 _22_ a_5418_3829# 0.01767f
C2118 a_3979_4943# a_4220_3829# 6.83e-19
C2119 net3 _01_ 0.006403f
C2120 clknet_0_clk clk 0.00889f
C2121 net6 net5 0.003368f
C2122 _11_ a_7258_3423# 8.51e-19
C2123 a_4995_4399# VPWR 0.011033f
C2124 a_4259_3311# a_5179_3311# 2.37e-21
C2125 a_4454_4649# _06_ 0.111795f
C2126 net6 a_7019_4943# 2.84e-19
C2127 net7 a_5843_3829# 0.08513f
C2128 a_2302_7241# _10_ 6.77e-19
C2129 a_2502_7396# a_2235_6575# 0.0033f
C2130 _15_ a_1683_3861# 8.17e-21
C2131 _16_ a_3433_4175# 3.98e-19
C2132 _01_ a_2253_7119# 2.39e-19
C2133 _23_ _16_ 3.32e-22
C2134 a_3979_4943# net7 0.002934f
C2135 a_1915_7815# VPWR 0.415615f
C2136 a_5599_2741# a_5505_2388# 3.27e-19
C2137 a_4259_3311# counter[4] 2.6e-19
C2138 a_3215_3829# a_2823_3677# 0.006202f
C2139 a_2290_3829# a_2313_3311# 6.87e-19
C2140 _16_ a_3225_4399# 4.87e-20
C2141 a_7641_3311# VPWR 4.71e-19
C2142 _24_ a_7267_3087# 9.33e-19
C2143 clknet_1_0__leaf_clk a_2715_3829# 0.002373f
C2144 a_2235_4399# a_2122_3855# 0.002054f
C2145 _04_ a_2290_3829# 8.38e-20
C2146 clknet_1_1__leaf_clk clk 0.008913f
C2147 a_4786_5065# _19_ 0.457296f
C2148 a_2431_7663# _12_ 7.61e-20
C2149 net8 a_7090_3855# 2.79e-19
C2150 _15_ a_4520_4373# 6.77e-20
C2151 _02_ VPWR 0.325572f
C2152 _25_ a_6817_3861# 1.11e-19
C2153 a_2235_6575# a_2389_6575# 0.004009f
C2154 net4 a_2290_3829# 5.24e-19
C2155 _10_ a_2317_6575# 4.63e-20
C2156 _14_ a_2398_3677# 9.43e-20
C2157 a_4986_5220# net8 5.83e-19
C2158 net7 a_6427_2741# 0.023542f
C2159 net9 VPWR 0.964697f
C2160 a_7258_3829# a_6651_3311# 1.99e-20
C2161 _13_ a_2800_4399# 2.65e-20
C2162 _18_ a_5333_5321# 2.19e-20
C2163 _15_ clk 0.005511f
C2164 a_2125_3311# a_2566_3423# 0.127288f
C2165 _11_ a_3267_4667# 0.052724f
C2166 a_1915_7351# VPWR 0.399249f
C2167 net9 a_5675_3855# 0.002503f
C2168 _07_ a_6211_3579# 3.3e-20
C2169 a_2248_4233# VPWR 4.21e-19
C2170 _23_ a_7345_2388# 7.52e-20
C2171 a_2398_3677# a_2614_2883# 0.003601f
C2172 net5 counter[3] 0.082806f
C2173 _24_ net10 0.13484f
C2174 a_2295_7637# a_2502_7637# 0.273138f
C2175 _19_ a_4767_3463# 4.85e-22
C2176 a_2302_7937# a_2431_7663# 0.110715f
C2177 a_2011_7637# a_2253_8029# 0.008508f
C2178 _11_ a_5001_3311# 0.001398f
C2179 a_8109_2767# counter[8] 1.28e-20
C2180 _15_ a_5891_3133# 3.42e-21
C2181 _07_ a_5505_2388# 7.51e-19
C2182 a_6817_3861# a_7515_3855# 0.194892f
C2183 a_3215_2999# a_3831_3105# 0.013543f
C2184 a_2991_3579# a_2949_3311# 7.84e-20
C2185 _17_ a_3267_4667# 1.35e-20
C2186 a_7005_3855# a_6817_3311# 1.41e-20
C2187 a_7258_3829# a_7683_3829# 1.28e-19
C2188 a_6817_3311# counter[7] 5.88e-20
C2189 a_4454_4649# VPWR 0.316019f
C2190 a_2842_4511# net5 1.47e-21
C2191 _04_ net8 7.52e-21
C2192 a_5213_4664# a_5165_3855# 1.39e-19
C2193 a_2431_7497# _12_ 0.039032f
C2194 _07_ a_4811_3861# 0.022853f
C2195 a_4786_5065# a_4915_5321# 0.110715f
C2196 net6 a_6211_3579# 3.96e-21
C2197 a_4779_5161# _05_ 0.196756f
C2198 _11_ a_6817_3861# 2.03e-20
C2199 _11_ a_4779_5161# 2.33e-19
C2200 net5 a_4413_3311# 1.04e-20
C2201 clknet_0_clk a_5618_3677# 4.63e-19
C2202 net6 a_5505_2388# 0.013611f
C2203 net2 clknet_1_0__leaf_clk 0.026712f
C2204 a_4399_5175# a_4454_4649# 3.4e-19
C2205 a_4495_5175# a_4520_4373# 0.006438f
C2206 net7 a_5165_3855# 0.014734f
C2207 clknet_1_1__leaf_clk a_7005_3855# 3.58e-19
C2208 net5 VPWR 0.923749f
C2209 net6 a_4811_3861# 0.0618f
C2210 net9 a_7077_2767# 0.008597f
C2211 net4 net8 0.001699f
C2212 a_7019_4943# VPWR 0.206381f
C2213 a_2295_7637# a_2502_7396# 6.88e-20
C2214 net6 a_5077_4721# 4.57e-19
C2215 a_3799_4943# _19_ 0.001413f
C2216 a_2431_7663# a_2295_7337# 5.28e-20
C2217 clknet_0_clk a_4220_3829# 8.98e-21
C2218 a_2502_7637# a_2302_7241# 1.26e-19
C2219 _17_ a_4779_5161# 0.42661f
C2220 a_4329_5461# a_4786_5065# 0.016444f
C2221 clknet_0_clk a_5213_4664# 7.62e-19
C2222 _15_ a_7005_3855# 0.007874f
C2223 _18_ net8 0.01511f
C2224 _12_ a_1845_5461# 4.42e-19
C2225 _15_ counter[7] 0.003538f
C2226 _11_ a_4259_3311# 0.222369f
C2227 _11_ a_2041_4649# 0.002118f
C2228 _22_ a_7267_3087# 1.37e-20
C2229 a_6817_3311# a_7599_3677# 6.32e-19
C2230 a_7090_3677# a_7185_3677# 0.007724f
C2231 _11_ a_2840_3087# 9.44e-19
C2232 clknet_1_0__leaf_clk _11_ 0.317456f
C2233 a_1849_3861# a_2547_3855# 0.196846f
C2234 a_2290_3829# a_2715_3829# 1.28e-19
C2235 clknet_0_clk net7 0.043959f
C2236 _06_ a_4811_3861# 0.091082f
C2237 clknet_1_1__leaf_clk a_5618_3677# 0.042872f
C2238 _07_ _20_ 1.72e-19
C2239 _17_ a_4259_3311# 1e-20
C2240 _00_ a_2502_7637# 0.00938f
C2241 a_1683_3861# a_2217_3855# 0.002698f
C2242 a_2823_3677# net5 0.019334f
C2243 net7 a_4069_5309# 5.91e-19
C2244 clknet_1_0__leaf_clk _17_ 3.38e-20
C2245 a_2678_7119# VPWR 0.004407f
C2246 a_2011_7351# _01_ 8.93e-19
C2247 net7 a_6817_3311# 0.001362f
C2248 a_2295_7337# a_2431_7497# 0.136009f
C2249 _13_ a_2674_4765# 5.02e-20
C2250 clknet_1_1__leaf_clk a_4220_3829# 0.048773f
C2251 a_2302_7241# a_2502_7396# 0.080195f
C2252 _08_ net10 0.001321f
C2253 _16_ a_5250_3855# 0.00213f
C2254 _18_ a_4986_5220# 5.4e-20
C2255 net6 _20_ 0.00624f
C2256 a_6427_2741# a_6623_3133# 0.00119f
C2257 a_2037_3855# a_2217_3855# 0.001229f
C2258 net10 net11 0.310558f
C2259 a_6651_3861# a_7005_3855# 0.062224f
C2260 a_1683_3861# _03_ 0.001727f
C2261 _02_ a_1959_3311# 3.71e-19
C2262 _19_ a_4737_4943# 1.83e-19
C2263 net8 a_5179_3311# 0.009204f
C2264 _22_ net10 0.074459f
C2265 a_7258_3423# a_7641_3311# 4.67e-20
C2266 _15_ a_4220_3829# 0.229149f
C2267 clknet_1_1__leaf_clk net7 0.397702f
C2268 _11_ a_2631_3855# 7.61e-19
C2269 net4 a_2313_3311# 4.45e-19
C2270 _15_ a_5213_4664# 1.57e-19
C2271 net4 _04_ 0.689049f
C2272 a_5345_3311# a_6127_3677# 3.14e-19
C2273 a_5533_3311# a_5713_3677# 0.001229f
C2274 clknet_1_0__leaf_clk a_2651_7663# 0.002297f
C2275 a_3267_4667# a_3215_3829# 0.004132f
C2276 a_5814_4399# _07_ 0.022424f
C2277 a_4454_4649# a_4382_4649# 0.005941f
C2278 _18_ _04_ 0.003255f
C2279 a_2589_4399# a_2769_4765# 0.001229f
C2280 a_4520_4373# _21_ 0.114705f
C2281 _16_ a_2398_3677# 2.79e-19
C2282 _09_ a_8109_2767# 2.25e-19
C2283 a_6211_3579# VPWR 0.400861f
C2284 net7 _15_ 0.590844f
C2285 a_2295_7337# a_1845_5461# 6.92e-20
C2286 net6 a_6375_5309# 0.157729f
C2287 net9 a_7171_2767# 0.003753f
C2288 a_5505_2388# VPWR 0.315151f
C2289 a_6651_3311# a_7515_3677# 0.032244f
C2290 clknet_1_0__leaf_clk a_2849_7497# 0.018091f
C2291 a_5162_4943# VPWR 0.004407f
C2292 a_5250_3855# a_5533_3311# 0.001307f
C2293 a_5843_3829# a_6043_3677# 4.17e-19
C2294 a_1683_3861# a_1849_3861# 0.968904f
C2295 _09_ a_7683_3579# 0.010518f
C2296 _04_ a_3601_3855# 2.55e-19
C2297 net9 a_7258_3423# 0.022365f
C2298 a_4811_3861# VPWR 0.421866f
C2299 net6 a_5814_4399# 0.047825f
C2300 net1 a_2230_7485# 1.42e-19
C2301 a_7216_3311# VPWR -4.73e-35
C2302 net11 a_8265_2388# 0.003661f
C2303 _08_ a_5843_3829# 9.54e-19
C2304 _23_ a_7267_3087# 4.18e-19
C2305 clknet_0_clk a_5149_4721# 0.034583f
C2306 a_5077_4721# VPWR 0.001301f
C2307 a_4915_5321# a_4737_4943# 9.73e-19
C2308 a_7683_3829# a_7515_3677# 7.04e-19
C2309 a_5418_3829# a_5250_3855# 0.239923f
C2310 _18_ net4 3.06e-19
C2311 a_7515_3855# a_7683_3579# 7.04e-19
C2312 _05_ a_5333_5321# 0.114695f
C2313 a_4811_3861# a_5675_3855# 0.030894f
C2314 a_1959_3311# net5 8.46e-19
C2315 _15_ a_2471_2741# 3.5e-20
C2316 _03_ a_2524_3311# 0.001074f
C2317 a_4977_3861# a_5843_3829# 0.034054f
C2318 a_1849_3861# a_2037_3855# 0.097818f
C2319 _12_ VPWR 0.307826f
C2320 a_4495_5175# a_4220_3829# 7.28e-21
C2321 net7 a_4929_3311# 1.98e-19
C2322 _11_ a_5333_5321# 7.39e-21
C2323 _22_ a_5843_3829# 4.4e-21
C2324 net4 a_3601_3855# 6.79e-19
C2325 _11_ a_2290_3829# 0.005658f
C2326 _11_ a_7683_3579# 5.38e-21
C2327 _24_ a_7599_3855# 8.56e-19
C2328 _14_ VPWR 0.685574f
C2329 a_4767_3463# a_5345_3311# 0.00145f
C2330 net7 a_6651_3861# 8.61e-20
C2331 a_5871_5162# _25_ 6.03e-21
C2332 _18_ a_3601_3855# 2.06e-20
C2333 _01_ a_2235_6575# 3.94e-19
C2334 _16_ a_4443_4175# 3.31e-19
C2335 a_2431_7497# _10_ 6.67e-19
C2336 _17_ a_5333_5321# 0.016586f
C2337 a_4495_5175# net7 0.037726f
C2338 net3 _03_ 0.019455f
C2339 a_6043_3677# a_6427_2741# 0.009905f
C2340 a_4779_5161# a_4995_4399# 2.84e-21
C2341 a_2302_7937# VPWR 0.335402f
C2342 a_2614_2883# VPWR 0.108977f
C2343 _16_ _07_ 0.003808f
C2344 a_6427_2741# a_6425_2388# 0.01226f
C2345 a_5165_3855# a_5345_3855# 0.001229f
C2346 _20_ a_4413_3311# 0.001506f
C2347 _23_ net10 0.188811f
C2348 clknet_1_1__leaf_clk a_5149_4721# 7.2e-19
C2349 _24_ a_7941_3087# 5.3e-19
C2350 net8 _09_ 2.1e-20
C2351 clknet_1_0__leaf_clk a_3215_3829# 1.95e-19
C2352 _04_ a_2715_3829# 0.008333f
C2353 a_7199_4943# _25_ 0.082413f
C2354 a_2235_4399# a_2547_3855# 0.001393f
C2355 net11 a_6427_2741# 1.29e-21
C2356 _20_ VPWR 0.175404f
C2357 a_7199_4943# _09_ 2.51e-21
C2358 _24_ a_6817_3311# 0.03707f
C2359 _05_ a_5871_5162# 0.121098f
C2360 a_4915_5321# _19_ 0.040707f
C2361 _22_ a_6427_2741# 0.191159f
C2362 _07_ counter[5] 1.62e-19
C2363 net6 _16_ 0.291584f
C2364 net4 a_1825_2388# 7.77e-19
C2365 _11_ a_5871_5162# 0.004334f
C2366 net8 a_7515_3855# 1.1e-19
C2367 _15_ a_5149_4721# 2.91e-20
C2368 a_4399_5175# _20_ 1.63e-20
C2369 _14_ a_2823_3677# 0.002114f
C2370 net4 a_2715_3829# 0.110738f
C2371 net3 a_1849_3861# 0.007798f
C2372 a_2401_4399# a_2589_4399# 0.095025f
C2373 a_2125_3311# a_2991_3579# 0.034054f
C2374 _05_ a_7199_4943# 4.21e-20
C2375 clknet_1_1__leaf_clk _24_ 0.041474f
C2376 a_3267_4667# a_4454_4649# 1.25e-19
C2377 _11_ net8 0.418201f
C2378 a_2566_3423# a_2398_3677# 0.239923f
C2379 net6 counter[5] 0.080069f
C2380 a_2295_7337# VPWR 0.446206f
C2381 net9 a_6817_3861# 0.001054f
C2382 _18_ a_2715_3829# 3.26e-20
C2383 _17_ a_5871_5162# 0.019971f
C2384 a_4329_5461# _19_ 5.98e-19
C2385 a_6375_5309# VPWR 0.455589f
C2386 a_2673_4233# VPWR 0.002609f
C2387 _07_ a_5533_3311# 0.128255f
C2388 a_2991_3579# a_3215_2999# 0.001036f
C2389 a_4779_5161# net9 6.06e-20
C2390 a_1915_7815# clknet_1_0__leaf_clk 0.007095f
C2391 a_2502_7637# a_2431_7663# 0.239923f
C2392 _11_ a_5744_3311# 0.002651f
C2393 _15_ a_6623_3133# 0.006963f
C2394 _06_ _16_ 0.064563f
C2395 counter[6] counter[7] 0.079796f
C2396 a_4977_3861# a_5165_3855# 0.095025f
C2397 _15_ _24_ 0.032103f
C2398 _17_ net8 0.172731f
C2399 a_5814_4399# VPWR 1.3575f
C2400 _17_ a_7199_4943# 8.24e-19
C2401 a_4986_5220# _05_ 3.36e-19
C2402 _07_ a_5418_3829# 0.011124f
C2403 _08_ a_7599_3855# 2.34e-19
C2404 net6 a_5533_3311# 0.00565f
C2405 a_5814_4399# a_5675_3855# 5.73e-19
C2406 _21_ a_4220_3829# 0.005326f
C2407 net8 a_5795_3133# 0.005557f
C2408 a_2125_8527# VPWR 5.43e-19
C2409 _11_ a_7090_3855# 6.96e-20
C2410 _11_ a_4986_5220# 3.53e-20
C2411 net2 _04_ 4.09e-22
C2412 a_4779_5161# a_4454_4649# 0.001895f
C2413 _21_ a_5213_4664# 1.69e-19
C2414 net3 counter[1] 0.103986f
C2415 a_2235_4399# a_1683_3861# 0.002682f
C2416 clknet_1_1__leaf_clk a_5345_3855# 0.002214f
C2417 _13_ a_1849_3861# 1.58e-19
C2418 clknet_1_0__leaf_clk _02_ 0.254839f
C2419 a_2011_7637# enable 2.06e-20
C2420 a_3145_6825# VPWR 0.006514f
C2421 net6 a_5418_3829# 0.012704f
C2422 a_6719_3133# VPWR 0.001259f
C2423 _16_ counter[3] 9.14e-20
C2424 a_6043_3677# a_6817_3311# 2.56e-19
C2425 clknet_1_0__leaf_clk a_1915_7351# 0.01132f
C2426 net7 _21_ 0.326643f
C2427 clknet_0_clk a_4977_3861# 5.94e-19
C2428 a_2502_7637# a_2431_7497# 1.77e-19
C2429 a_5179_3311# a_7005_3311# 4.76e-21
C2430 a_2431_7663# a_2502_7396# 1.77e-19
C2431 _17_ a_4986_5220# 0.032936f
C2432 a_2295_7637# _01_ 6.79e-20
C2433 a_4329_5461# a_4915_5321# 0.013455f
C2434 a_7345_2388# counter[9] 2.34e-19
C2435 clknet_0_clk _22_ 0.003156f
C2436 net11 a_7941_3087# 0.001149f
C2437 net2 net4 8.49e-21
C2438 clknet_1_0__leaf_clk a_2248_4233# 0.001807f
C2439 _14_ a_1959_3311# 0.008544f
C2440 _23_ a_6427_2741# 0.130093f
C2441 _08_ a_6817_3311# 0.001269f
C2442 _11_ a_2313_3311# 4.78e-19
C2443 a_2842_4511# _16_ 1.01e-19
C2444 _24_ a_6651_3861# 0.031818f
C2445 a_4454_4649# a_4259_3311# 5.65e-20
C2446 a_6817_3311# net11 2.58e-19
C2447 _22_ a_7941_3087# 3.34e-21
C2448 a_7258_3423# a_7216_3311# 4.62e-19
C2449 _11_ _04_ 0.257603f
C2450 _11_ a_3917_3105# 6.46e-19
C2451 a_2235_4399# a_4520_4373# 1.55e-21
C2452 a_5814_4399# a_7077_2767# 1.15e-20
C2453 net1 a_2695_6575# 4.64e-19
C2454 _06_ a_5418_3829# 0.001008f
C2455 clknet_1_1__leaf_clk a_6043_3677# 0.044904f
C2456 _16_ a_4413_3311# 5.12e-19
C2457 a_1959_3311# a_2614_2883# 0.00127f
C2458 net2 a_1499_7119# 0.07281f
C2459 _22_ a_6817_3311# 3.15e-20
C2460 _03_ a_2471_2741# 0.112166f
C2461 _00_ a_2253_8029# 3.7e-19
C2462 net7 a_5135_5309# 0.002551f
C2463 _16_ VPWR 2.17996f
C2464 clknet_1_1__leaf_clk _08_ 0.00277f
C2465 _17_ _04_ 6.62e-21
C2466 a_1959_3311# _20_ 1.9e-21
C2467 _03_ a_2949_3311# 9.96e-20
C2468 a_1683_3861# a_3245_3855# 2.77e-19
C2469 a_4259_3311# net5 5.06e-20
C2470 net7 counter[6] 1.8e-19
C2471 _10_ VPWR 0.249351f
C2472 _11_ net4 0.952686f
C2473 net6 a_3831_3105# 1.4e-20
C2474 clknet_1_1__leaf_clk net11 1.82e-20
C2475 a_5759_3855# VPWR 0.004428f
C2476 clknet_1_1__leaf_clk a_4977_3861# 0.079788f
C2477 clknet_1_0__leaf_clk net5 6.12e-20
C2478 net7 a_7090_3677# 4.39e-19
C2479 a_2302_7241# _01_ 0.239739f
C2480 a_2502_7396# a_2431_7497# 0.239923f
C2481 net10 a_7939_2223# 1.3e-21
C2482 _15_ a_6043_3677# 1.98e-20
C2483 net5 a_2840_3087# 0.075434f
C2484 _18_ _05_ 1.11e-19
C2485 clknet_1_1__leaf_clk _22_ 0.031888f
C2486 VPWR counter[5] 0.450193f
C2487 a_4399_5175# _16_ 3.45e-20
C2488 a_5675_3855# a_5759_3855# 0.008508f
C2489 a_6427_2741# a_6825_3133# 0.005781f
C2490 _11_ _18_ 0.035586f
C2491 a_7258_3829# a_7005_3855# 3.39e-19
C2492 _24_ a_7723_2741# 0.003347f
C2493 _15_ _08_ 0.030258f
C2494 net8 a_5786_3423# 0.00264f
C2495 _15_ net11 1.7e-19
C2496 _15_ a_4977_3861# 0.027322f
C2497 counter[1] counter[2] 0.070133f
C2498 _17_ net4 9.08e-20
C2499 a_7683_3579# a_7641_3311# 7.84e-20
C2500 net4 a_2907_3677# 8.77e-19
C2501 _11_ a_3601_3855# 0.00137f
C2502 _15_ _22_ 0.422897f
C2503 net3 a_2235_4399# 1.48e-19
C2504 a_5786_3423# a_5744_3311# 4.62e-19
C2505 a_5345_3311# a_6651_3311# 3.23e-19
C2506 _00_ _01_ 0.014628f
C2507 net2 a_1825_2388# 0.016821f
C2508 net8 a_6169_3311# 5.67e-20
C2509 _17_ _18_ 0.181987f
C2510 net1 a_2230_7663# 2.14e-19
C2511 a_5149_4721# _21_ 0.001146f
C2512 _16_ a_2823_3677# 6.21e-20
C2513 a_5533_3311# VPWR 0.079731f
C2514 a_2502_7396# a_1845_5461# 2.84e-19
C2515 net9 a_8109_2767# 3.29e-19
C2516 a_7939_2223# a_8265_2388# 0.024477f
C2517 a_7345_2388# VPWR 0.303091f
C2518 a_1683_3861# a_2122_3855# 0.273138f
C2519 net6 a_4287_4399# 4.02e-19
C2520 _02_ a_2290_3829# 4.65e-19
C2521 clknet_1_0__leaf_clk a_2678_7119# 0.002447f
C2522 _09_ a_7005_3311# 0.129132f
C2523 clknet_0_clk _23_ 2.29e-20
C2524 a_6651_3311# a_7185_3677# 0.002698f
C2525 net9 a_7683_3579# 0.001937f
C2526 a_5418_3829# VPWR 0.185172f
C2527 VPWR counter[0] 0.375177f
C2528 _23_ a_7941_3087# 3.52e-19
C2529 net8 a_4995_4399# 0.009814f
C2530 _08_ a_6651_3861# 0.097891f
C2531 _11_ a_5179_3311# 0.029022f
C2532 _15_ a_3215_2999# 1.84e-19
C2533 a_4779_5161# a_5162_4943# 0.001632f
C2534 a_2122_3855# a_2037_3855# 0.037333f
C2535 a_2290_3829# a_2248_4233# 4.62e-19
C2536 a_4977_3861# a_6651_3861# 1.33e-19
C2537 a_5418_3829# a_5675_3855# 0.036838f
C2538 a_4811_3861# a_6817_3861# 3.42e-21
C2539 _23_ a_6817_3311# 0.031117f
C2540 net7 a_6127_3677# 0.002598f
C2541 a_4779_5161# a_4811_3861# 0.001493f
C2542 _11_ a_6457_5309# 2.28e-19
C2543 _22_ a_6651_3861# 5.82e-21
C2544 _13_ a_2235_4399# 0.002226f
C2545 _11_ counter[4] 6.77e-20
C2546 _11_ a_7005_3311# 2.79e-20
C2547 a_4786_5065# a_5213_4664# 0.003687f
C2548 _11_ a_2715_3829# 0.033019f
C2549 a_5814_4399# a_7258_3423# 7.13e-20
C2550 _06_ a_4287_4399# 4.79e-19
C2551 _17_ a_5179_3311# 1.69e-21
C2552 net2 a_1957_8207# 0.00492f
C2553 clknet_1_1__leaf_clk _23_ 0.071442f
C2554 a_2566_3423# VPWR 0.219675f
C2555 a_4786_5065# net7 0.027472f
C2556 a_2502_7637# VPWR 0.286747f
C2557 a_4986_5220# a_4995_4399# 1.55e-20
C2558 a_3831_3105# VPWR 0.2419f
C2559 a_5871_5162# net9 3.61e-20
C2560 a_7077_2767# a_7345_2388# 1.23e-19
C2561 _04_ a_3215_3829# 0.171873f
C2562 _15_ a_3433_4175# 1.54e-19
C2563 _16_ a_1959_3311# 1.96e-20
C2564 net8 net9 0.748324f
C2565 _15_ _23_ 0.683594f
C2566 net11 a_7723_2741# 0.088145f
C2567 _24_ a_7090_3677# 0.010089f
C2568 net10 a_7185_3855# 8.52e-20
C2569 a_7199_4943# net9 7.48e-22
C2570 _22_ a_7723_2741# 4.31e-19
C2571 net4 a_3849_2388# 0.003224f
C2572 net3 a_1457_2388# 0.006292f
C2573 clknet_1_0__leaf_clk _12_ 0.075464f
C2574 net7 a_4767_3463# 0.084753f
C2575 net9 a_5744_3311# 3.93e-19
C2576 net6 net10 1.08e-19
C2577 net4 a_3215_3829# 0.005124f
C2578 net3 a_2122_3855# 8.21e-19
C2579 clknet_1_0__leaf_clk _14_ 0.088295f
C2580 clknet_1_1__leaf_clk a_6825_3133# 5.67e-20
C2581 _05_ _25_ 4.6e-21
C2582 a_2566_3423# a_2823_3677# 0.036838f
C2583 a_2401_4399# a_3183_4765# 4.04e-19
C2584 _14_ a_2840_3087# 0.122283f
C2585 net8 a_4454_4649# 0.063158f
C2586 a_7515_3855# _09_ 0.001217f
C2587 a_2674_4765# a_2589_4399# 0.037333f
C2588 a_2502_7396# VPWR 0.271061f
C2589 _19_ clk 0.013619f
C2590 _11_ _25_ 2.54e-20
C2591 _18_ a_3215_3829# 0.002375f
C2592 net2 _11_ 0.001125f
C2593 a_4349_4175# VPWR 5.6e-19
C2594 net10 a_7363_3087# 0.002966f
C2595 a_2502_7637# a_2678_8029# 0.007724f
C2596 net10 counter[9] 0.092658f
C2597 a_2295_7637# a_2849_7663# 0.062224f
C2598 a_4986_5220# net9 4.56e-19
C2599 a_2302_7937# clknet_1_0__leaf_clk 0.470509f
C2600 _11_ _09_ 0.004259f
C2601 a_2431_7663# a_2253_8029# 9.73e-19
C2602 net6 a_2401_4399# 0.004467f
C2603 _15_ a_6825_3133# 0.002119f
C2604 a_4287_4399# VPWR 0.004487f
C2605 a_3215_3829# a_3601_3855# 0.006406f
C2606 a_2614_2883# a_2840_3087# 0.005961f
C2607 a_5418_3829# a_5376_4233# 4.62e-19
C2608 a_5250_3855# a_5165_3855# 0.037333f
C2609 a_4259_3311# _20_ 0.237238f
C2610 _23_ a_6651_3861# 0.029216f
C2611 net1 a_2125_8207# 0.073427f
C2612 a_2769_4765# VPWR 0.003961f
C2613 net8 net5 0.002187f
C2614 a_1845_5461# a_2401_4399# 1.63e-19
C2615 a_4779_5161# a_6375_5309# 2.69e-21
C2616 _17_ _25_ 1.89e-19
C2617 _07_ a_5843_3829# 0.008579f
C2618 net8 a_5997_3133# 1.72e-20
C2619 a_3799_4943# net7 2.88e-19
C2620 a_4399_5175# a_4287_4399# 2.76e-20
C2621 a_5814_4399# a_6817_3861# 0.008007f
C2622 _21_ a_4977_3861# 0.002388f
C2623 _11_ _05_ 0.023537f
C2624 a_5179_3311# a_5786_3423# 0.141453f
C2625 a_4786_5065# a_5149_4721# 6.47e-19
C2626 _21_ _22_ 2.96e-19
C2627 _04_ _02_ 1.6e-19
C2628 a_2389_6575# VPWR 3.14e-19
C2629 a_7019_4943# a_7199_4943# 0.185422f
C2630 a_2295_7637# enable 1.25e-19
C2631 net6 a_5843_3829# 0.002597f
C2632 a_6043_3677# counter[6] 2e-19
C2633 a_3979_4943# net6 1.5e-19
C2634 a_7171_2767# a_7345_2388# 2.21e-19
C2635 _17_ _05_ 0.0576f
C2636 a_2849_7663# a_2302_7241# 4.5e-20
C2637 clknet_0_clk a_5250_3855# 4.59e-20
C2638 clknet_1_0__leaf_clk a_2295_7337# 0.683552f
C2639 a_8265_2388# counter[9] 0.039377f
C2640 a_6425_2388# counter[6] 0.1107f
C2641 a_5333_5321# a_5162_4943# 0.001229f
C2642 _15_ a_7641_4233# 6.51e-20
C2643 _11_ _17_ 0.113734f
C2644 a_7258_3423# a_7345_2388# 2.21e-20
C2645 clknet_1_0__leaf_clk a_2673_4233# 4.11e-19
C2646 net2 a_2651_7663# 1.37e-19
C2647 a_3849_2388# counter[4] 0.001146f
C2648 net11 a_7753_2767# 0.01512f
C2649 _23_ a_7723_2741# 0.220841f
C2650 a_4329_5461# a_4520_4373# 3.15e-19
C2651 a_3267_4667# _16_ 0.001048f
C2652 net4 _02_ 1.19e-19
C2653 _24_ a_7258_3829# 0.015657f
C2654 _11_ a_2907_3677# 0.002515f
C2655 _22_ a_7753_2767# 6.52e-20
C2656 _03_ a_2125_3311# 0.260627f
C2657 a_1959_3311# a_2566_3423# 0.141453f
C2658 a_7515_3677# a_7599_3677# 0.008508f
C2659 _04_ a_4454_4649# 3.15e-21
C2660 a_2715_3829# a_3215_3829# 0.016344f
C2661 a_4329_5461# clk 0.318051f
C2662 clknet_1_1__leaf_clk a_5713_3677# 0.001835f
C2663 _06_ a_5843_3829# 1.75e-19
C2664 _22_ a_7090_3677# 0.004398f
C2665 _22_ counter[6] 9.35e-22
C2666 _03_ a_3215_2999# 1.19e-19
C2667 net2 a_2849_7497# 1.01e-21
C2668 _00_ a_2849_7663# 0.139872f
C2669 net4 a_2248_4233# 1.81e-19
C2670 net7 a_4737_4943# 6.13e-20
C2671 a_2313_3311# net5 2.02e-19
C2672 net6 a_6427_2741# 0.009771f
C2673 net7 a_7515_3677# 1.49e-19
C2674 _04_ net5 0.003846f
C2675 net3 a_2695_6575# 0.001478f
C2676 a_2401_4399# a_2842_4511# 0.111047f
C2677 a_2011_7351# a_2230_7485# 0.006169f
C2678 clknet_1_1__leaf_clk a_5250_3855# 0.033626f
C2679 a_1915_7351# a_1499_7119# 5.03e-19
C2680 net5 a_3917_3105# 0.001706f
C2681 net10 VPWR 1.28398f
C2682 a_2431_7497# _01_ 0.00226f
C2683 a_6651_3311# counter[7] 2.09e-20
C2684 net9 counter[8] 2.39e-19
C2685 _14_ a_2290_3829# 8.48e-21
C2686 a_4779_5161# _16_ 1.49e-19
C2687 a_7090_3855# a_7216_4233# 0.005525f
C2688 a_7077_2767# a_7267_3087# 0.011458f
C2689 _18_ a_4454_4649# 5.77e-19
C2690 a_1849_3861# a_2125_3311# 6.25e-19
C2691 net8 a_6211_3579# 0.020836f
C2692 a_2849_7497# _11_ 0.001319f
C2693 _00_ enable 2.67e-19
C2694 _15_ a_5250_3855# 0.026278f
C2695 _19_ a_4220_3829# 8.51e-20
C2696 net8 a_5505_2388# 3.76e-19
C2697 net4 net5 0.483177f
C2698 a_2401_4399# VPWR 0.304738f
C2699 a_4520_4373# a_4349_3855# 1.06e-19
C2700 a_6043_3677# a_6127_3677# 0.008508f
C2701 net8 a_4811_3861# 0.036074f
C2702 net3 a_2936_2767# 1.66e-19
C2703 a_4382_4649# a_4287_4399# 0.002032f
C2704 net1 net3 0.313425f
C2705 a_4341_3311# VPWR 2.86e-19
C2706 net9 a_5179_3311# 0.006834f
C2707 _16_ a_4259_3311# 0.105405f
C2708 net6 a_5165_3855# 0.008614f
C2709 clknet_1_0__leaf_clk _16_ 4.14e-20
C2710 clknet_1_1__leaf_clk a_5599_2741# 1.84e-19
C2711 _01_ a_1845_5461# 3.77e-19
C2712 a_8265_2388# VPWR 0.276039f
C2713 _19_ net7 0.552257f
C2714 _16_ a_2840_3087# 3.76e-19
C2715 a_1683_3861# a_2547_3855# 0.032244f
C2716 clknet_1_0__leaf_clk _10_ 0.006812f
C2717 _02_ a_2715_3829# 1.8e-19
C2718 net9 a_7005_3311# 0.016338f
C2719 net10 a_7077_2767# 0.27342f
C2720 clknet_0_clk _07_ 0.114561f
C2721 a_5843_3829# VPWR 0.406789f
C2722 _23_ a_7753_2767# 0.113094f
C2723 _11_ a_5786_3423# 0.039242f
C2724 _08_ a_7258_3829# 0.047112f
C2725 a_3979_4943# VPWR 0.185924f
C2726 a_2290_3829# a_2673_4233# 4.67e-20
C2727 a_5843_3829# a_5675_3855# 0.310858f
C2728 a_4986_5220# a_5162_4943# 0.007724f
C2729 _15_ a_5599_2741# 1.2e-20
C2730 net7 a_7619_5162# 2.85e-19
C2731 a_2842_4511# a_2991_3579# 8.5e-21
C2732 a_2674_4765# a_2398_3677# 9.19e-21
C2733 a_2401_4399# a_2823_3677# 0.001133f
C2734 _23_ a_7090_3677# 0.011058f
C2735 _06_ a_5165_3855# 0.114717f
C2736 net7 a_6651_3311# 0.007864f
C2737 _11_ a_6651_5309# 0.005861f
C2738 a_4779_5161# a_5418_3829# 2.9e-20
C2739 a_4986_5220# a_4811_3861# 2.08e-22
C2740 _22_ a_7258_3829# 9.3e-20
C2741 a_4786_5065# a_4977_3861# 6.46e-19
C2742 clknet_0_clk net6 0.087511f
C2743 _11_ a_3215_3829# 0.001227f
C2744 _11_ a_6169_3311# 2.44e-19
C2745 a_3979_4943# a_4399_5175# 0.017007f
C2746 a_3099_4765# a_3215_2999# 3.06e-22
C2747 a_4786_5065# _22_ 8.56e-19
C2748 a_1845_5461# clknet_0_clk 0.317755f
C2749 a_2589_4399# a_1849_3861# 2.83e-19
C2750 net2 a_1915_7815# 0.092265f
C2751 net8 _20_ 0.027217f
C2752 _09_ a_7641_3311# 0.001794f
C2753 _17_ a_6651_5309# 3.01e-19
C2754 a_2991_3579# VPWR 0.391294f
C2755 a_4915_5321# net7 0.035198f
C2756 net5 counter[4] 0.001223f
C2757 clknet_1_1__leaf_clk _07_ 0.44529f
C2758 a_2253_8029# VPWR 0.005315f
C2759 a_4329_5461# a_4220_3829# 4.81e-21
C2760 a_7723_2741# a_7939_2223# 1.29e-21
C2761 a_6427_2741# VPWR 0.419035f
C2762 a_2715_3829# net5 6.71e-21
C2763 a_7267_3087# a_7171_2767# 1.26e-19
C2764 _11_ a_4995_4399# 1.22e-19
C2765 a_4329_5461# a_5213_4664# 1.03e-20
C2766 _15_ a_4443_4175# 0.004604f
C2767 clknet_0_clk _06_ 2.8e-19
C2768 _24_ a_7515_3677# 0.012283f
C2769 net2 _02_ 0.035742f
C2770 _15_ _07_ 0.022092f
C2771 clknet_1_1__leaf_clk net6 0.323735f
C2772 a_4329_5461# net7 0.002812f
C2773 net3 a_2745_2388# 0.001252f
C2774 net9 _09_ 0.571636f
C2775 _11_ a_7641_3311# 9.67e-22
C2776 _19_ a_5149_4721# 1.87e-20
C2777 net1 a_1582_7439# 0.001512f
C2778 net2 a_1915_7351# 0.004306f
C2779 a_3099_4765# a_3225_4399# 0.006169f
C2780 a_3267_4667# a_4287_4399# 3.28e-20
C2781 _04_ _14_ 4.63e-22
C2782 a_2401_4399# a_4382_4649# 1.01e-20
C2783 net8 a_5814_4399# 0.001798f
C2784 a_1683_3861# a_2037_3855# 0.062224f
C2785 a_2842_4511# a_2800_4399# 4.62e-19
C2786 net6 _15_ 0.117386f
C2787 a_2991_3579# a_2823_3677# 0.310858f
C2788 a_2235_4399# a_2125_3311# 3.23e-21
C2789 a_2401_4399# a_1959_3311# 1.21e-19
C2790 _01_ VPWR 0.468919f
C2791 clknet_1_0__leaf_clk a_2566_3423# 0.001507f
C2792 net9 a_7515_3855# 2.45e-19
C2793 net10 a_7171_2767# 0.007482f
C2794 a_5165_3855# VPWR 0.084103f
C2795 _18_ a_4811_3861# 5.99e-21
C2796 _16_ a_2290_3829# 1.76e-20
C2797 a_7199_4943# a_5814_4399# 0.006666f
C2798 _11_ _02_ 0.012298f
C2799 a_2502_7637# clknet_1_0__leaf_clk 0.040993f
C2800 clknet_1_1__leaf_clk _06_ 0.005269f
C2801 a_2431_7663# a_2849_7663# 3.39e-19
C2802 _05_ net9 1.93e-19
C2803 net10 a_7258_3423# 1.26e-19
C2804 _15_ a_7363_3087# 0.001637f
C2805 net6 a_2674_4765# 3.12e-19
C2806 a_2471_2741# a_2936_2767# 0.005941f
C2807 _11_ net9 0.233741f
C2808 a_4220_3829# a_4349_3855# 0.062574f
C2809 a_2561_9514# a_2302_7937# 4.65e-23
C2810 net4 _14_ 0.209869f
C2811 net1 a_2011_7637# 0.017118f
C2812 a_3215_2999# a_3389_3105# 0.006584f
C2813 a_6427_2741# a_7077_2767# 0.010893f
C2814 _23_ a_7258_3829# 0.006211f
C2815 a_2800_4399# VPWR 3.37e-19
C2816 _19_ _24_ 8.27e-21
C2817 a_7599_3855# VPWR 0.00533f
C2818 _12_ a_1499_7119# 0.090947f
C2819 net6 a_4929_3311# 1.78e-19
C2820 _11_ a_2248_4233# 4.01e-19
C2821 a_5814_4399# a_7090_3855# 0.01166f
C2822 _15_ _06_ 0.139237f
C2823 net2 net5 7.09e-21
C2824 a_2011_7637# a_2230_7663# 0.006169f
C2825 a_6651_3861# a_7185_3855# 0.002698f
C2826 a_4915_5321# a_5149_4721# 1.61e-19
C2827 net4 a_2614_2883# 0.007901f
C2828 _17_ net9 7.02e-19
C2829 a_5179_3311# a_6211_3579# 0.048748f
C2830 a_5345_3311# a_5618_3677# 0.074022f
C2831 _24_ a_7619_5162# 0.006166f
C2832 clknet_0_clk VPWR 2.53166f
C2833 a_7019_4943# _25_ 0.001476f
C2834 net7 a_4349_3855# 0.006434f
C2835 _11_ a_4454_4649# 0.043142f
C2836 a_2431_7663# enable 2.79e-20
C2837 a_5179_3311# a_5505_2388# 1.63e-21
C2838 _24_ a_6651_3311# 0.03301f
C2839 net6 a_6651_3861# 2.14e-19
C2840 a_4495_5175# net6 8.38e-19
C2841 net9 a_5795_3133# 0.001755f
C2842 a_7941_3087# VPWR 0.003335f
C2843 a_5786_3423# a_6169_3311# 4.67e-20
C2844 a_4811_3861# a_5179_3311# 0.012779f
C2845 clknet_1_0__leaf_clk a_2502_7396# 0.037641f
C2846 clknet_0_clk a_5675_3855# 0.013741f
C2847 a_4069_5309# VPWR 0.002157f
C2848 clknet_0_clk a_4399_5175# 0.002548f
C2849 a_3245_3855# a_3215_2999# 6.77e-20
C2850 a_2745_2388# counter[2] 0.1107f
C2851 a_6817_3311# VPWR 0.31984f
C2852 net1 a_2011_7351# 0.030538f
C2853 _07_ a_3831_3339# 2.73e-21
C2854 _11_ net5 0.388184f
C2855 _17_ a_4454_4649# 0.076419f
C2856 net8 _16_ 0.193029f
C2857 _24_ a_7683_3829# 0.009415f
C2858 a_4329_5461# a_5149_4721# 6.61e-19
C2859 _08_ a_7515_3677# 3.02e-19
C2860 net3 a_1683_3861# 0.023332f
C2861 a_2235_4399# a_2589_4399# 0.062224f
C2862 a_1959_3311# a_2991_3579# 0.048748f
C2863 _03_ a_2398_3677# 0.010537f
C2864 a_7515_3677# net11 0.003417f
C2865 _05_ a_7019_4943# 6.38e-20
C2866 clknet_1_0__leaf_clk a_2769_4765# 4.17e-19
C2867 net8 a_5759_3855# 9.28e-20
C2868 net7 a_5345_3311# 0.030766f
C2869 _06_ a_6651_3861# 4.19e-21
C2870 net6 a_3831_3339# 4.93e-21
C2871 clknet_1_1__leaf_clk VPWR 3.34801f
C2872 net4 a_2673_4233# 3.33e-19
C2873 net3 a_2037_3855# 0.003111f
C2874 net7 a_6545_5309# 0.00717f
C2875 net6 a_7723_2741# 4.97e-21
C2876 net1 a_1875_8207# 0.224922f
C2877 net9 a_5801_4233# 3.81e-19
C2878 net7 a_7185_3677# 1.13e-19
C2879 a_2401_4399# a_3267_4667# 0.034054f
C2880 clknet_1_0__leaf_clk a_2389_6575# 3.8e-19
C2881 _17_ a_7019_4943# 0.056144f
C2882 clknet_1_1__leaf_clk a_5675_3855# 0.024694f
C2883 _15_ a_4413_3311# 2.18e-19
C2884 a_2842_4511# a_2674_4765# 0.239923f
C2885 _14_ a_2715_3829# 1.02e-20
C2886 a_4399_5175# clknet_1_1__leaf_clk 1.77e-20
C2887 a_4986_5220# _16_ 1.35e-21
C2888 _15_ VPWR 1.72333f
C2889 a_2471_2741# a_2745_2388# 4.71e-19
C2890 a_7258_3829# a_7641_4233# 4.67e-20
C2891 a_6817_3861# net10 5.04e-19
C2892 a_1849_3861# a_2398_3677# 0.002f
C2893 a_2122_3855# a_2125_3311# 0.004962f
C2894 _20_ a_5179_3311# 0.004564f
C2895 a_2235_6575# a_2695_6575# 0.001479f
C2896 _13_ a_1683_3861# 3.88e-19
C2897 a_6817_3311# a_7077_2767# 0.008374f
C2898 a_2715_3829# a_2614_2883# 6.81e-19
C2899 _15_ a_5675_3855# 0.0351f
C2900 a_2674_4765# VPWR 0.255338f
C2901 _19_ a_4977_3861# 4.93e-21
C2902 net8 a_7345_2388# 7.5e-19
C2903 _21_ a_4443_4175# 4.25e-19
C2904 a_4399_5175# _15_ 1.78e-19
C2905 a_6043_3677# a_6651_3311# 3.54e-19
C2906 a_6211_3579# _09_ 0.001669f
C2907 _19_ _22_ 7e-20
C2908 a_7619_5162# _08_ 0.109717f
C2909 net8 a_5418_3829# 0.001066f
C2910 net9 a_5786_3423# 0.007121f
C2911 _21_ _07_ 4.77e-20
C2912 a_4929_3311# VPWR 4.84e-19
C2913 _08_ a_6651_3311# 1.13e-19
C2914 _04_ _16_ 0.025302f
C2915 _09_ a_7216_3311# 3.07e-19
C2916 a_6651_3311# net11 3.07e-19
C2917 _16_ a_3917_3105# 8.82e-20
C2918 _02_ a_3215_3829# 7.66e-20
C2919 net9 a_6169_3311# 0.001933f
C2920 net6 _21_ 0.083542f
C2921 net2 _12_ 0.10227f
C2922 a_6651_3861# VPWR 0.714632f
C2923 _22_ a_6651_3311# 4.68e-20
C2924 _15_ a_2823_3677# 1.6e-20
C2925 net1 a_2235_6575# 0.232539f
C2926 _08_ a_7683_3829# 0.004928f
C2927 _11_ a_6211_3579# 0.028602f
C2928 a_5814_4399# a_5179_3311# 4.21e-21
C2929 a_6375_5309# a_6457_5309# 0.005781f
C2930 a_2125_8207# a_2011_7637# 1.96e-19
C2931 a_5149_4721# a_5345_3311# 8.41e-19
C2932 a_4495_5175# VPWR 0.175351f
C2933 a_7683_3829# net11 1.16e-19
C2934 net4 _16_ 0.442589f
C2935 a_5843_3829# a_6817_3861# 2.73e-19
C2936 a_2715_3829# a_2673_4233# 7.84e-20
C2937 a_5675_3855# a_6651_3861# 1.07e-19
C2938 _15_ a_7077_2767# 0.087822f
C2939 _23_ a_7515_3677# 0.006274f
C2940 a_2674_4765# a_2823_3677# 1.06e-19
C2941 a_4786_5065# a_5250_3855# 9.47e-20
C2942 net2 _14_ 0.45134f
C2943 counter[8] VGND 0.587415f
C2944 counter[9] VGND 0.871549f
C2945 counter[7] VGND 0.919615f
C2946 counter[6] VGND 0.662885f
C2947 counter[5] VGND 0.638642f
C2948 counter[4] VGND 0.794555f
C2949 counter[3] VGND 0.823254f
C2950 counter[2] VGND 0.636768f
C2951 counter[1] VGND 0.621106f
C2952 counter[0] VGND 0.997297f
C2953 clk VGND 3.38597f
C2954 enable VGND 1.15467f
C2955 VPWR VGND 0.363098p
C2956 a_8265_2388# VGND 0.269609f
C2957 a_7939_2223# VGND 0.257101f
C2958 a_7345_2388# VGND 0.296141f
C2959 a_6425_2388# VGND 0.269288f
C2960 a_5505_2388# VGND 0.278393f
C2961 a_4585_2388# VGND 0.327843f
C2962 a_3849_2388# VGND 0.269041f
C2963 a_2745_2388# VGND 0.276333f
C2964 a_1825_2388# VGND 0.316834f
C2965 a_1457_2388# VGND 0.25238f
C2966 a_8109_2767# VGND 8.84e-19
C2967 a_7753_2767# VGND 0.004608f
C2968 a_7171_2767# VGND 0.01879f
C2969 a_7941_3087# VGND 0.005268f
C2970 a_7363_3087# VGND 0.00969f
C2971 a_7267_3087# VGND 0.006323f
C2972 a_6825_3133# VGND 0.001553f
C2973 a_6719_3133# VGND 0.003693f
C2974 a_6623_3133# VGND 0.003656f
C2975 a_5997_3133# VGND 0.003203f
C2976 a_5891_3133# VGND 0.005457f
C2977 a_5795_3133# VGND 0.005167f
C2978 a_2936_2767# VGND 0.001114f
C2979 a_3917_3105# VGND 0.004685f
C2980 a_3389_3105# VGND 0.007506f
C2981 a_2840_3087# VGND 0.183329f
C2982 a_7723_2741# VGND 0.363777f
C2983 a_7077_2767# VGND 0.343017f
C2984 a_6427_2741# VGND 0.260798f
C2985 a_5599_2741# VGND 0.294745f
C2986 a_3831_3105# VGND 0.255389f
C2987 a_3215_2999# VGND 0.284107f
C2988 a_2614_2883# VGND 0.207092f
C2989 a_2471_2741# VGND 0.20644f
C2990 a_7641_3311# VGND 0.004786f
C2991 net11 VGND 0.755509f
C2992 a_7216_3311# VGND 0.009087f
C2993 a_7599_3677# VGND 3.75e-19
C2994 a_6169_3311# VGND 0.004164f
C2995 a_7185_3677# VGND 0.002645f
C2996 a_7005_3311# VGND 0.063765f
C2997 a_7515_3677# VGND 0.268634f
C2998 a_7683_3579# VGND 0.376509f
C2999 a_7090_3677# VGND 0.227724f
C3000 a_7258_3423# VGND 0.257495f
C3001 a_6817_3311# VGND 0.334487f
C3002 _09_ VGND 0.540883f
C3003 a_6651_3311# VGND 0.496464f
C3004 a_5744_3311# VGND 0.008691f
C3005 a_6127_3677# VGND 2.5e-19
C3006 a_5001_3311# VGND 7.68e-19
C3007 a_4929_3311# VGND 0.002515f
C3008 a_4413_3311# VGND 0.002664f
C3009 a_4341_3311# VGND 7.95e-19
C3010 a_5713_3677# VGND 7.5e-19
C3011 a_5533_3311# VGND 0.062716f
C3012 a_6043_3677# VGND 0.275541f
C3013 a_6211_3579# VGND 0.356576f
C3014 a_5618_3677# VGND 0.218254f
C3015 a_5786_3423# VGND 0.278138f
C3016 a_5345_3311# VGND 0.323857f
C3017 a_5179_3311# VGND 0.485385f
C3018 a_3917_3339# VGND 0.004685f
C3019 _20_ VGND 0.296302f
C3020 a_2949_3311# VGND 0.004794f
C3021 net5 VGND 1.52242f
C3022 a_2524_3311# VGND 0.007478f
C3023 a_2907_3677# VGND 3.28e-19
C3024 a_2313_3311# VGND 0.069011f
C3025 a_4767_3463# VGND 0.233023f
C3026 a_4259_3311# VGND 0.25233f
C3027 a_3831_3339# VGND 0.250617f
C3028 a_2823_3677# VGND 0.29125f
C3029 a_2991_3579# VGND 0.405228f
C3030 a_2398_3677# VGND 0.210325f
C3031 a_2566_3423# VGND 0.255348f
C3032 a_2125_3311# VGND 0.417108f
C3033 _03_ VGND 0.578555f
C3034 a_1959_3311# VGND 0.557931f
C3035 a_7599_3855# VGND 0.001033f
C3036 a_7185_3855# VGND 0.002645f
C3037 net10 VGND 1.52118f
C3038 a_7641_4233# VGND 0.005282f
C3039 a_5759_3855# VGND 0.002002f
C3040 a_7216_4233# VGND 0.010952f
C3041 a_7005_3855# VGND 0.070151f
C3042 a_5801_4233# VGND 0.005844f
C3043 a_4349_3855# VGND 0.014804f
C3044 a_3601_3855# VGND 0.001519f
C3045 a_3245_3855# VGND 0.026188f
C3046 a_2631_3855# VGND 4.07e-19
C3047 a_2217_3855# VGND 6.93e-19
C3048 a_5376_4233# VGND 0.006941f
C3049 a_5165_3855# VGND 0.060618f
C3050 a_4443_4175# VGND 0.006538f
C3051 a_4349_4175# VGND 0.008165f
C3052 a_3433_4175# VGND 0.007253f
C3053 a_2673_4233# VGND 0.004473f
C3054 a_1505_3855# VGND 4.64e-19
C3055 a_2248_4233# VGND 0.008558f
C3056 a_2037_3855# VGND 0.080622f
C3057 a_7515_3855# VGND 0.275172f
C3058 a_7683_3829# VGND 0.371259f
C3059 a_7090_3855# VGND 0.237292f
C3060 a_7258_3829# VGND 0.266551f
C3061 a_6817_3861# VGND 0.344626f
C3062 a_6651_3861# VGND 0.532322f
C3063 a_5675_3855# VGND 0.288597f
C3064 a_5843_3829# VGND 0.391747f
C3065 a_5250_3855# VGND 0.200127f
C3066 a_5418_3829# VGND 0.247676f
C3067 a_4977_3861# VGND 0.312142f
C3068 a_4811_3861# VGND 0.480598f
C3069 a_4220_3829# VGND 0.352433f
C3070 a_3215_3829# VGND 0.430766f
C3071 a_2547_3855# VGND 0.280567f
C3072 a_2715_3829# VGND 0.367396f
C3073 a_2122_3855# VGND 0.214988f
C3074 a_2290_3829# VGND 0.263107f
C3075 a_1849_3861# VGND 0.41156f
C3076 _02_ VGND 0.385543f
C3077 a_1683_3861# VGND 0.551857f
C3078 _14_ VGND 1.2474f
C3079 a_5436_4399# VGND 0.004249f
C3080 a_4995_4399# VGND 0.154917f
C3081 _07_ VGND 0.467795f
C3082 a_4287_4399# VGND 0.204157f
C3083 a_3225_4399# VGND 0.00681f
C3084 _16_ VGND 2.102403f
C3085 _22_ VGND 1.56987f
C3086 a_5077_4721# VGND 8.25e-20
C3087 a_5213_4664# VGND 0.189132f
C3088 net9 VGND 1.97499f
C3089 _06_ VGND 0.355082f
C3090 _21_ VGND 0.491639f
C3091 a_4382_4649# VGND 9.9e-19
C3092 a_2800_4399# VGND 0.007439f
C3093 a_3183_4765# VGND 0.002478f
C3094 a_2769_4765# VGND 5.31e-19
C3095 a_2589_4399# VGND 0.062654f
C3096 a_5814_4399# VGND 2.07482f
C3097 a_5149_4721# VGND 0.166512f
C3098 a_4454_4649# VGND 0.208373f
C3099 a_4520_4373# VGND 0.228425f
C3100 net8 VGND 1.78641f
C3101 a_3099_4765# VGND 0.331871f
C3102 a_3267_4667# VGND 0.427232f
C3103 a_2674_4765# VGND 0.220057f
C3104 a_2842_4511# VGND 0.267836f
C3105 a_2401_4399# VGND 0.384412f
C3106 _04_ VGND 0.647447f
C3107 a_2235_4399# VGND 0.561386f
C3108 a_2041_4649# VGND 0.005123f
C3109 _13_ VGND 1.1383f
C3110 net4 VGND 1.31662f
C3111 _08_ VGND 0.727548f
C3112 a_7289_5309# VGND 0.00819f
C3113 a_6651_5309# VGND 0.003851f
C3114 a_6545_5309# VGND 0.003674f
C3115 a_6457_5309# VGND 0.001688f
C3116 a_4737_4943# VGND 7.93e-19
C3117 a_5333_5321# VGND 0.060853f
C3118 a_5135_5309# VGND 0.006624f
C3119 a_4714_5309# VGND 0.005539f
C3120 a_4069_5309# VGND 0.005238f
C3121 _25_ VGND 0.366822f
C3122 a_7619_5162# VGND 0.272105f
C3123 a_7199_4943# VGND 0.262291f
C3124 _24_ VGND 0.696921f
C3125 a_7019_4943# VGND 0.271218f
C3126 _23_ VGND 0.973323f
C3127 a_6375_5309# VGND 0.264312f
C3128 _15_ VGND 3.54853f
C3129 net7 VGND 2.72082f
C3130 net6 VGND 3.218744f
C3131 _19_ VGND 0.32708f
C3132 a_5871_5162# VGND 0.252712f
C3133 clknet_1_1__leaf_clk VGND 3.414301f
C3134 _05_ VGND 0.318608f
C3135 a_4915_5321# VGND 0.241882f
C3136 a_4986_5220# VGND 0.198121f
C3137 a_4786_5065# VGND 0.303545f
C3138 a_4779_5161# VGND 0.46613f
C3139 a_4495_5175# VGND 0.281525f
C3140 a_4399_5175# VGND 0.378965f
C3141 a_3979_4943# VGND 0.234926f
C3142 _18_ VGND 0.468402f
C3143 a_3799_4943# VGND 0.254342f
C3144 _17_ VGND 0.622186f
C3145 a_4329_5461# VGND 2.29287f
C3146 clknet_0_clk VGND 4.193551f
C3147 a_1845_5461# VGND 2.29289f
C3148 a_2389_6575# VGND 0.002457f
C3149 a_2317_6575# VGND 0.001303f
C3150 a_3145_6825# VGND 0.005104f
C3151 _11_ VGND 5.669386f
C3152 a_2695_6575# VGND 0.298451f
C3153 _10_ VGND 0.339714f
C3154 a_2235_6575# VGND 0.252154f
C3155 a_2253_7119# VGND 6.89e-19
C3156 a_2849_7497# VGND 0.064411f
C3157 a_2651_7485# VGND 0.006624f
C3158 a_1499_7119# VGND 0.017559f
C3159 a_2230_7485# VGND 0.004183f
C3160 _12_ VGND 1.2616f
C3161 a_1582_7439# VGND 0.004429f
C3162 _01_ VGND 0.405148f
C3163 a_2431_7497# VGND 0.238144f
C3164 a_2502_7396# VGND 0.195482f
C3165 a_2302_7241# VGND 0.31379f
C3166 a_2295_7337# VGND 0.552106f
C3167 a_2011_7351# VGND 0.279727f
C3168 a_1915_7351# VGND 0.390267f
C3169 net3 VGND 2.298238f
C3170 a_2651_7663# VGND 0.007478f
C3171 a_2230_7663# VGND 0.004654f
C3172 clknet_1_0__leaf_clk VGND 4.010709f
C3173 a_2849_7663# VGND 0.069779f
C3174 a_2253_8029# VGND 6.84e-19
C3175 a_2431_7663# VGND 0.264386f
C3176 a_2502_7637# VGND 0.210923f
C3177 a_2295_7637# VGND 0.580201f
C3178 a_2302_7937# VGND 0.340144f
C3179 a_2011_7637# VGND 0.287469f
C3180 a_1915_7815# VGND 0.412387f
C3181 a_2125_8207# VGND 0.013142f
C3182 a_1957_8207# VGND 0.006974f
C3183 _00_ VGND 0.757573f
C3184 a_2125_8527# VGND 0.006222f
C3185 a_1875_8207# VGND 0.393994f
C3186 net2 VGND 3.503971f
C3187 net1 VGND 1.81106f
C3188 a_2561_9514# VGND 0.293097f
C3189 net6.t5 VGND 0.023291f
C3190 net6.t2 VGND 0.034395f
C3191 net6.n0 VGND 0.095831f
C3192 net6.t10 VGND 0.040459f
C3193 net6.t11 VGND 0.025233f
C3194 net6.n1 VGND 0.081347f
C3195 net6.n2 VGND 0.124436f
C3196 net6.t9 VGND 0.023291f
C3197 net6.t3 VGND 0.034395f
C3198 net6.n3 VGND 0.095831f
C3199 net6.n4 VGND 0.41789f
C3200 net6.t8 VGND 0.021456f
C3201 net6.t13 VGND 0.017754f
C3202 net6.n5 VGND 0.093771f
C3203 net6.n6 VGND 0.080526f
C3204 net6.n7 VGND 0.286209f
C3205 net6.t6 VGND 0.027524f
C3206 net6.t12 VGND 0.043832f
C3207 net6.n8 VGND 0.059723f
C3208 net6.n9 VGND 0.146037f
C3209 net6.n10 VGND 0.772479f
C3210 net6.n11 VGND 0.732404f
C3211 net6.t7 VGND 0.023842f
C3212 net6.t14 VGND 0.040459f
C3213 net6.n12 VGND 0.051672f
C3214 net6.t15 VGND 0.023842f
C3215 net6.t4 VGND 0.040459f
C3216 net6.n13 VGND 0.057394f
C3217 net6.n14 VGND 0.027196f
C3218 net6.n15 VGND 0.1061f
C3219 net6.n16 VGND 0.491563f
C3220 net6.t0 VGND 0.092732f
C3221 net6.n17 VGND 0.127274f
C3222 net6.t1 VGND 0.050895f
C3223 net6.n18 VGND 0.064268f
C3224 _16_.t1 VGND 0.046376f
C3225 _16_.n0 VGND 0.026397f
C3226 _16_.t7 VGND 0.021164f
C3227 _16_.t2 VGND 0.017507f
C3228 _16_.n1 VGND 0.047954f
C3229 _16_.n2 VGND 0.154756f
C3230 _16_.t9 VGND 0.020065f
C3231 _16_.t3 VGND 0.031953f
C3232 _16_.n3 VGND 0.045672f
C3233 _16_.n4 VGND 0.0375f
C3234 _16_.t6 VGND 0.020065f
C3235 _16_.t8 VGND 0.031953f
C3236 _16_.n5 VGND 0.058943f
C3237 _16_.n6 VGND 0.063595f
C3238 _16_.n7 VGND 0.426096f
C3239 _16_.t4 VGND 0.012893f
C3240 _16_.t5 VGND 0.013824f
C3241 _16_.n8 VGND 0.03796f
C3242 _16_.n9 VGND 0.022428f
C3243 _16_.n10 VGND 0.327394f
C3244 _16_.n11 VGND 0.020414f
C3245 _16_.t0 VGND 0.119992f
C3246 _16_.n12 VGND 0.021583f
C3247 _16_.n13 VGND 0.021194f
C3248 net3.t0 VGND 0.067779f
C3249 net3.t7 VGND 0.019614f
C3250 net3.t4 VGND 0.031428f
C3251 net3.n0 VGND 0.061838f
C3252 net3.n1 VGND 0.008618f
C3253 net3.n2 VGND 0.005246f
C3254 net3.t2 VGND 0.029572f
C3255 net3.t3 VGND 0.018443f
C3256 net3.n3 VGND 0.059457f
C3257 net3.n4 VGND 0.019056f
C3258 net3.t6 VGND 0.030361f
C3259 net3.t5 VGND 0.055573f
C3260 net3.n5 VGND 0.744487f
C3261 net3.n6 VGND 0.124162f
C3262 net3.n7 VGND 0.092279f
C3263 net3.t1 VGND 0.037792f
C3264 net3.n8 VGND 0.040884f
C3265 net2.t2 VGND 0.015381f
C3266 net2.t5 VGND 0.026101f
C3267 net2.n0 VGND 0.037026f
C3268 net2.t6 VGND 0.015381f
C3269 net2.t10 VGND 0.026101f
C3270 net2.n1 VGND 0.033335f
C3271 net2.n2 VGND 0.017289f
C3272 net2.n3 VGND 0.0837f
C3273 net2.t7 VGND 0.026101f
C3274 net2.t8 VGND 0.016278f
C3275 net2.n4 VGND 0.052479f
C3276 net2.n5 VGND 0.259642f
C3277 net2.t9 VGND 0.013842f
C3278 net2.t3 VGND 0.011454f
C3279 net2.n6 VGND 0.060494f
C3280 net2.n7 VGND 0.03533f
C3281 net2.n8 VGND 0.650991f
C3282 net2.t11 VGND 0.017756f
C3283 net2.t4 VGND 0.028277f
C3284 net2.n9 VGND 0.038818f
C3285 net2.n10 VGND 0.03575f
C3286 net2.n11 VGND 0.11929f
C3287 net2.n12 VGND 0.278364f
C3288 net2.n13 VGND 0.037886f
C3289 net2.t0 VGND 0.08709f
C3290 net2.n14 VGND 0.10636f
C3291 net2.t1 VGND 0.032833f
C3292 _11_.t0 VGND 0.02558f
C3293 _11_.t1 VGND 0.02558f
C3294 _11_.n0 VGND 0.053419f
C3295 _11_.t17 VGND 0.042601f
C3296 _11_.t11 VGND 0.026392f
C3297 _11_.n1 VGND 0.086305f
C3298 _11_.n2 VGND 0.024278f
C3299 _11_.t6 VGND 0.027069f
C3300 _11_.t13 VGND 0.043108f
C3301 _11_.n3 VGND 0.058737f
C3302 _11_.n4 VGND 0.032841f
C3303 _11_.t14 VGND 0.023619f
C3304 _11_.t4 VGND 0.034667f
C3305 _11_.n5 VGND 0.06984f
C3306 _11_.n6 VGND 0.034707f
C3307 _11_.n7 VGND 0.494881f
C3308 _11_.t20 VGND 0.027069f
C3309 _11_.t7 VGND 0.043108f
C3310 _11_.n8 VGND 0.058739f
C3311 _11_.n9 VGND 0.133927f
C3312 _11_.n10 VGND 0.765831f
C3313 _11_.t8 VGND 0.021102f
C3314 _11_.t12 VGND 0.017461f
C3315 _11_.n11 VGND 0.092223f
C3316 _11_.n12 VGND 0.043963f
C3317 _11_.n13 VGND 0.150035f
C3318 _11_.t10 VGND 0.028052f
C3319 _11_.t21 VGND 0.019277f
C3320 _11_.n14 VGND 0.081517f
C3321 _11_.n15 VGND 0.011369f
C3322 _11_.n16 VGND 0.03744f
C3323 _11_.n17 VGND 0.156255f
C3324 _11_.t15 VGND 0.019598f
C3325 _11_.t19 VGND 0.028465f
C3326 _11_.n18 VGND 0.067767f
C3327 _11_.n19 VGND 0.143997f
C3328 _11_.n20 VGND 0.492685f
C3329 _11_.t5 VGND 0.042359f
C3330 _11_.t16 VGND 0.026451f
C3331 _11_.n21 VGND 0.080165f
C3332 _11_.n22 VGND 0.023455f
C3333 _11_.n23 VGND 0.356691f
C3334 _11_.t9 VGND 0.023619f
C3335 _11_.t18 VGND 0.034667f
C3336 _11_.n24 VGND 0.06984f
C3337 _11_.n25 VGND 0.014495f
C3338 _11_.n26 VGND 0.490885f
C3339 _11_.n27 VGND 1.19049f
C3340 _11_.n28 VGND 0.353781f
C3341 _11_.n29 VGND 0.021904f
C3342 _11_.t3 VGND 0.010743f
C3343 _11_.t2 VGND 0.010743f
C3344 _11_.n30 VGND 0.02648f
C3345 clknet_1_0__leaf_clk.t37 VGND 0.022262f
C3346 clknet_1_0__leaf_clk.t41 VGND 0.014894f
C3347 clknet_1_0__leaf_clk.n0 VGND 0.04068f
C3348 clknet_1_0__leaf_clk.n1 VGND 0.107083f
C3349 clknet_1_0__leaf_clk.t38 VGND 0.014894f
C3350 clknet_1_0__leaf_clk.t33 VGND 0.022262f
C3351 clknet_1_0__leaf_clk.n2 VGND 0.041145f
C3352 clknet_1_0__leaf_clk.n3 VGND 0.437523f
C3353 clknet_1_0__leaf_clk.t2 VGND 0.014222f
C3354 clknet_1_0__leaf_clk.t4 VGND 0.014222f
C3355 clknet_1_0__leaf_clk.n4 VGND 0.036128f
C3356 clknet_1_0__leaf_clk.t6 VGND 0.014222f
C3357 clknet_1_0__leaf_clk.t7 VGND 0.014222f
C3358 clknet_1_0__leaf_clk.n5 VGND 0.029978f
C3359 clknet_1_0__leaf_clk.n6 VGND 0.136621f
C3360 clknet_1_0__leaf_clk.t5 VGND 0.014222f
C3361 clknet_1_0__leaf_clk.t9 VGND 0.014222f
C3362 clknet_1_0__leaf_clk.n7 VGND 0.029978f
C3363 clknet_1_0__leaf_clk.n8 VGND 0.0787f
C3364 clknet_1_0__leaf_clk.t11 VGND 0.014222f
C3365 clknet_1_0__leaf_clk.t8 VGND 0.014222f
C3366 clknet_1_0__leaf_clk.n9 VGND 0.029978f
C3367 clknet_1_0__leaf_clk.n10 VGND 0.078334f
C3368 clknet_1_0__leaf_clk.t14 VGND 0.014222f
C3369 clknet_1_0__leaf_clk.t10 VGND 0.014222f
C3370 clknet_1_0__leaf_clk.n11 VGND 0.029978f
C3371 clknet_1_0__leaf_clk.n12 VGND 0.078334f
C3372 clknet_1_0__leaf_clk.t15 VGND 0.014222f
C3373 clknet_1_0__leaf_clk.t0 VGND 0.014222f
C3374 clknet_1_0__leaf_clk.n13 VGND 0.029978f
C3375 clknet_1_0__leaf_clk.t1 VGND 0.014222f
C3376 clknet_1_0__leaf_clk.t3 VGND 0.014222f
C3377 clknet_1_0__leaf_clk.n14 VGND 0.029589f
C3378 clknet_1_0__leaf_clk.t26 VGND 0.005973f
C3379 clknet_1_0__leaf_clk.t28 VGND 0.005973f
C3380 clknet_1_0__leaf_clk.n15 VGND 0.021211f
C3381 clknet_1_0__leaf_clk.t30 VGND 0.005973f
C3382 clknet_1_0__leaf_clk.t31 VGND 0.005973f
C3383 clknet_1_0__leaf_clk.n16 VGND 0.013636f
C3384 clknet_1_0__leaf_clk.n17 VGND 0.086164f
C3385 clknet_1_0__leaf_clk.t29 VGND 0.005973f
C3386 clknet_1_0__leaf_clk.t17 VGND 0.005973f
C3387 clknet_1_0__leaf_clk.n18 VGND 0.013636f
C3388 clknet_1_0__leaf_clk.n19 VGND 0.051791f
C3389 clknet_1_0__leaf_clk.t19 VGND 0.005973f
C3390 clknet_1_0__leaf_clk.t16 VGND 0.005973f
C3391 clknet_1_0__leaf_clk.n20 VGND 0.013644f
C3392 clknet_1_0__leaf_clk.n21 VGND 0.053424f
C3393 clknet_1_0__leaf_clk.t22 VGND 0.005973f
C3394 clknet_1_0__leaf_clk.t18 VGND 0.005973f
C3395 clknet_1_0__leaf_clk.n22 VGND 0.013636f
C3396 clknet_1_0__leaf_clk.n23 VGND 0.051791f
C3397 clknet_1_0__leaf_clk.t20 VGND 0.005973f
C3398 clknet_1_0__leaf_clk.t21 VGND 0.005973f
C3399 clknet_1_0__leaf_clk.n24 VGND 0.013636f
C3400 clknet_1_0__leaf_clk.n25 VGND 0.05205f
C3401 clknet_1_0__leaf_clk.t23 VGND 0.005973f
C3402 clknet_1_0__leaf_clk.t24 VGND 0.005973f
C3403 clknet_1_0__leaf_clk.n26 VGND 0.013636f
C3404 clknet_1_0__leaf_clk.n27 VGND 0.04471f
C3405 clknet_1_0__leaf_clk.t25 VGND 0.005973f
C3406 clknet_1_0__leaf_clk.t27 VGND 0.005973f
C3407 clknet_1_0__leaf_clk.n28 VGND 0.013163f
C3408 clknet_1_0__leaf_clk.n29 VGND 0.043256f
C3409 clknet_1_0__leaf_clk.n30 VGND 0.09308f
C3410 clknet_1_0__leaf_clk.n31 VGND 0.067594f
C3411 clknet_1_0__leaf_clk.n32 VGND 0.04742f
C3412 clknet_1_0__leaf_clk.t12 VGND 0.014222f
C3413 clknet_1_0__leaf_clk.t13 VGND 0.014222f
C3414 clknet_1_0__leaf_clk.n33 VGND 0.028445f
C3415 clknet_1_0__leaf_clk.n34 VGND 0.022411f
C3416 clknet_1_0__leaf_clk.n35 VGND 0.171468f
C3417 clknet_1_0__leaf_clk.t35 VGND 0.014894f
C3418 clknet_1_0__leaf_clk.t32 VGND 0.022262f
C3419 clknet_1_0__leaf_clk.n36 VGND 0.040782f
C3420 clknet_1_0__leaf_clk.n37 VGND 0.024896f
C3421 clknet_1_0__leaf_clk.t34 VGND 0.022262f
C3422 clknet_1_0__leaf_clk.t39 VGND 0.014894f
C3423 clknet_1_0__leaf_clk.n38 VGND 0.040732f
C3424 clknet_1_0__leaf_clk.n39 VGND 0.086433f
C3425 clknet_1_0__leaf_clk.n40 VGND 0.225449f
C3426 clknet_1_0__leaf_clk.t36 VGND 0.022262f
C3427 clknet_1_0__leaf_clk.t40 VGND 0.014894f
C3428 clknet_1_0__leaf_clk.n41 VGND 0.04068f
C3429 clknet_1_0__leaf_clk.n42 VGND 0.027948f
C3430 clknet_1_0__leaf_clk.n43 VGND 0.145937f
C3431 clknet_1_1__leaf_clk.t29 VGND 0.005541f
C3432 clknet_1_1__leaf_clk.t30 VGND 0.005541f
C3433 clknet_1_1__leaf_clk.n0 VGND 0.019676f
C3434 clknet_1_1__leaf_clk.t25 VGND 0.005541f
C3435 clknet_1_1__leaf_clk.t27 VGND 0.005541f
C3436 clknet_1_1__leaf_clk.n1 VGND 0.01265f
C3437 clknet_1_1__leaf_clk.n2 VGND 0.07993f
C3438 clknet_1_1__leaf_clk.t28 VGND 0.005541f
C3439 clknet_1_1__leaf_clk.t23 VGND 0.005541f
C3440 clknet_1_1__leaf_clk.n3 VGND 0.01265f
C3441 clknet_1_1__leaf_clk.n4 VGND 0.048044f
C3442 clknet_1_1__leaf_clk.t24 VGND 0.005541f
C3443 clknet_1_1__leaf_clk.t26 VGND 0.005541f
C3444 clknet_1_1__leaf_clk.n5 VGND 0.012657f
C3445 clknet_1_1__leaf_clk.n6 VGND 0.049559f
C3446 clknet_1_1__leaf_clk.t21 VGND 0.005541f
C3447 clknet_1_1__leaf_clk.t22 VGND 0.005541f
C3448 clknet_1_1__leaf_clk.n7 VGND 0.01265f
C3449 clknet_1_1__leaf_clk.n8 VGND 0.048044f
C3450 clknet_1_1__leaf_clk.t31 VGND 0.005541f
C3451 clknet_1_1__leaf_clk.t20 VGND 0.005541f
C3452 clknet_1_1__leaf_clk.n9 VGND 0.011247f
C3453 clknet_1_1__leaf_clk.t33 VGND 0.013817f
C3454 clknet_1_1__leaf_clk.t41 VGND 0.020651f
C3455 clknet_1_1__leaf_clk.n10 VGND 0.038168f
C3456 clknet_1_1__leaf_clk.t39 VGND 0.020651f
C3457 clknet_1_1__leaf_clk.t34 VGND 0.013817f
C3458 clknet_1_1__leaf_clk.n11 VGND 0.037785f
C3459 clknet_1_1__leaf_clk.n12 VGND 0.039947f
C3460 clknet_1_1__leaf_clk.t38 VGND 0.013817f
C3461 clknet_1_1__leaf_clk.t35 VGND 0.020651f
C3462 clknet_1_1__leaf_clk.n13 VGND 0.038168f
C3463 clknet_1_1__leaf_clk.n14 VGND 0.30833f
C3464 clknet_1_1__leaf_clk.t40 VGND 0.020651f
C3465 clknet_1_1__leaf_clk.t37 VGND 0.013817f
C3466 clknet_1_1__leaf_clk.n15 VGND 0.037785f
C3467 clknet_1_1__leaf_clk.n16 VGND 0.030886f
C3468 clknet_1_1__leaf_clk.n17 VGND 0.118422f
C3469 clknet_1_1__leaf_clk.t36 VGND 0.013817f
C3470 clknet_1_1__leaf_clk.t32 VGND 0.020651f
C3471 clknet_1_1__leaf_clk.n18 VGND 0.037832f
C3472 clknet_1_1__leaf_clk.n19 VGND 0.022005f
C3473 clknet_1_1__leaf_clk.n20 VGND 0.128874f
C3474 clknet_1_1__leaf_clk.n21 VGND 0.280206f
C3475 clknet_1_1__leaf_clk.n22 VGND 0.023331f
C3476 clknet_1_1__leaf_clk.n23 VGND 0.030986f
C3477 clknet_1_1__leaf_clk.t17 VGND 0.005541f
C3478 clknet_1_1__leaf_clk.t18 VGND 0.005541f
C3479 clknet_1_1__leaf_clk.n24 VGND 0.01265f
C3480 clknet_1_1__leaf_clk.n25 VGND 0.041476f
C3481 clknet_1_1__leaf_clk.t14 VGND 0.013193f
C3482 clknet_1_1__leaf_clk.t11 VGND 0.013193f
C3483 clknet_1_1__leaf_clk.n26 VGND 0.027449f
C3484 clknet_1_1__leaf_clk.t12 VGND 0.013193f
C3485 clknet_1_1__leaf_clk.t13 VGND 0.013193f
C3486 clknet_1_1__leaf_clk.n27 VGND 0.02781f
C3487 clknet_1_1__leaf_clk.t8 VGND 0.013193f
C3488 clknet_1_1__leaf_clk.t9 VGND 0.013193f
C3489 clknet_1_1__leaf_clk.n28 VGND 0.033515f
C3490 clknet_1_1__leaf_clk.t4 VGND 0.013193f
C3491 clknet_1_1__leaf_clk.t6 VGND 0.013193f
C3492 clknet_1_1__leaf_clk.n29 VGND 0.02781f
C3493 clknet_1_1__leaf_clk.n30 VGND 0.126738f
C3494 clknet_1_1__leaf_clk.t7 VGND 0.013193f
C3495 clknet_1_1__leaf_clk.t2 VGND 0.013193f
C3496 clknet_1_1__leaf_clk.n31 VGND 0.02781f
C3497 clknet_1_1__leaf_clk.n32 VGND 0.073006f
C3498 clknet_1_1__leaf_clk.t3 VGND 0.013193f
C3499 clknet_1_1__leaf_clk.t5 VGND 0.013193f
C3500 clknet_1_1__leaf_clk.n33 VGND 0.02781f
C3501 clknet_1_1__leaf_clk.n34 VGND 0.072667f
C3502 clknet_1_1__leaf_clk.t0 VGND 0.013193f
C3503 clknet_1_1__leaf_clk.t1 VGND 0.013193f
C3504 clknet_1_1__leaf_clk.n35 VGND 0.02781f
C3505 clknet_1_1__leaf_clk.n36 VGND 0.072667f
C3506 clknet_1_1__leaf_clk.t10 VGND 0.013193f
C3507 clknet_1_1__leaf_clk.t15 VGND 0.013193f
C3508 clknet_1_1__leaf_clk.n37 VGND 0.02781f
C3509 clknet_1_1__leaf_clk.n38 VGND 0.073006f
C3510 clknet_1_1__leaf_clk.n39 VGND 0.062704f
C3511 clknet_1_1__leaf_clk.n40 VGND 0.086346f
C3512 clknet_1_1__leaf_clk.n41 VGND 0.040127f
C3513 clknet_1_1__leaf_clk.t19 VGND 0.005541f
C3514 clknet_1_1__leaf_clk.t16 VGND 0.005541f
C3515 clknet_1_1__leaf_clk.n42 VGND 0.012211f
C3516 VPWR.t459 VGND 0.002088f
C3517 VPWR.t884 VGND 0.004432f
C3518 VPWR.n1 VGND 0.011362f
C3519 VPWR.t460 VGND 0.002088f
C3520 VPWR.n2 VGND 0.006189f
C3521 VPWR.n3 VGND 0.0043f
C3522 VPWR.n4 VGND 0.002447f
C3523 VPWR.t615 VGND 0.002279f
C3524 VPWR.n5 VGND 0.004063f
C3525 VPWR.n6 VGND 0.002314f
C3526 VPWR.t888 VGND 0.030181f
C3527 VPWR.t858 VGND 0.030181f
C3528 VPWR.n7 VGND 0.027762f
C3529 VPWR.n8 VGND 0.005302f
C3530 VPWR.n9 VGND 0.001225f
C3531 VPWR.n10 VGND 8.51e-19
C3532 VPWR.n11 VGND 0.001281f
C3533 VPWR.n12 VGND 8.2e-19
C3534 VPWR.n13 VGND 0.001463f
C3535 VPWR.n14 VGND 0.001414f
C3536 VPWR.n15 VGND 0.058516f
C3537 VPWR.n16 VGND 0.221149f
C3538 VPWR.n17 VGND 0.117032f
C3539 VPWR.n18 VGND 0.064545f
C3540 VPWR.n19 VGND 0.001414f
C3541 VPWR.n20 VGND 0.048231f
C3542 VPWR.n21 VGND 0.001463f
C3543 VPWR.n22 VGND 0.001146f
C3544 VPWR.n23 VGND 6.56e-19
C3545 VPWR.n24 VGND 0.001224f
C3546 VPWR.n25 VGND 0.005302f
C3547 VPWR.t609 VGND 0.002279f
C3548 VPWR.n26 VGND 0.002879f
C3549 VPWR.n27 VGND 8.51e-19
C3550 VPWR.n28 VGND 8.2e-19
C3551 VPWR.n29 VGND 0.001463f
C3552 VPWR.n30 VGND 6.56e-19
C3553 VPWR.t472 VGND 0.021641f
C3554 VPWR.t475 VGND 0.029012f
C3555 VPWR.t743 VGND 0.005881f
C3556 VPWR.t18 VGND 0.006586f
C3557 VPWR.t798 VGND 0.006586f
C3558 VPWR.t188 VGND 0.006586f
C3559 VPWR.t159 VGND 0.013016f
C3560 VPWR.t744 VGND 0.010036f
C3561 VPWR.t20 VGND 0.012389f
C3562 VPWR.t179 VGND 0.011291f
C3563 VPWR.t343 VGND 0.006586f
C3564 VPWR.t785 VGND 0.010272f
C3565 VPWR.t722 VGND 0.011761f
C3566 VPWR.t713 VGND 0.018426f
C3567 VPWR.t784 VGND 0.015525f
C3568 VPWR.t180 VGND 0.014114f
C3569 VPWR.t731 VGND 0.013722f
C3570 VPWR.t499 VGND 0.014741f
C3571 VPWR.t782 VGND 0.014271f
C3572 VPWR.t155 VGND 0.009017f
C3573 VPWR.t598 VGND 0.021641f
C3574 VPWR.n31 VGND 0.015704f
C3575 VPWR.n32 VGND 0.002501f
C3576 VPWR.t603 VGND 0.002287f
C3577 VPWR.n33 VGND 0.001522f
C3578 VPWR.t868 VGND 0.008808f
C3579 VPWR.t599 VGND 0.002071f
C3580 VPWR.n34 VGND 0.00326f
C3581 VPWR.n35 VGND 0.003332f
C3582 VPWR.t600 VGND 0.002101f
C3583 VPWR.n36 VGND 0.01479f
C3584 VPWR.n37 VGND 0.005325f
C3585 VPWR.t500 VGND 0.002286f
C3586 VPWR.n38 VGND 0.006785f
C3587 VPWR.t895 VGND 0.030181f
C3588 VPWR.t156 VGND 4.79e-19
C3589 VPWR.t783 VGND 4.79e-19
C3590 VPWR.n39 VGND 9.86e-19
C3591 VPWR.n40 VGND 0.002967f
C3592 VPWR.n41 VGND 0.002447f
C3593 VPWR.t732 VGND 0.001144f
C3594 VPWR.n42 VGND 0.002958f
C3595 VPWR.n43 VGND 0.003084f
C3596 VPWR.n44 VGND 8.51e-19
C3597 VPWR.n45 VGND 8.2e-19
C3598 VPWR.n46 VGND 0.001463f
C3599 VPWR.n47 VGND 0.048231f
C3600 VPWR.n48 VGND 0.001414f
C3601 VPWR.n49 VGND 0.058516f
C3602 VPWR.n50 VGND 0.117032f
C3603 VPWR.n51 VGND 0.001414f
C3604 VPWR.n52 VGND 0.001281f
C3605 VPWR.n53 VGND 0.001463f
C3606 VPWR.n54 VGND 8.2e-19
C3607 VPWR.n55 VGND 8.51e-19
C3608 VPWR.t476 VGND 0.002071f
C3609 VPWR.t905 VGND 0.00872f
C3610 VPWR.n57 VGND 0.015149f
C3611 VPWR.t477 VGND 0.002071f
C3612 VPWR.n58 VGND 0.008692f
C3613 VPWR.t572 VGND 0.002071f
C3614 VPWR.t878 VGND 0.00872f
C3615 VPWR.n60 VGND 0.015149f
C3616 VPWR.t573 VGND 0.002071f
C3617 VPWR.n61 VGND 0.008692f
C3618 VPWR.n62 VGND 0.00749f
C3619 VPWR.t654 VGND 0.002088f
C3620 VPWR.t841 VGND 0.004432f
C3621 VPWR.n64 VGND 0.011362f
C3622 VPWR.t655 VGND 0.002088f
C3623 VPWR.n65 VGND 0.006189f
C3624 VPWR.n66 VGND 4.71e-19
C3625 VPWR.n67 VGND 0.002447f
C3626 VPWR.t745 VGND 0.002626f
C3627 VPWR.n68 VGND 8.67e-19
C3628 VPWR.n69 VGND 9.99e-19
C3629 VPWR.t501 VGND 0.002279f
C3630 VPWR.n70 VGND 9.49e-19
C3631 VPWR.t714 VGND 0.001157f
C3632 VPWR.t723 VGND 5.61e-19
C3633 VPWR.n71 VGND 0.002356f
C3634 VPWR.n72 VGND 0.002839f
C3635 VPWR.n73 VGND 0.002363f
C3636 VPWR.n74 VGND 8.51e-19
C3637 VPWR.n75 VGND 6.56e-19
C3638 VPWR.n76 VGND 0.001197f
C3639 VPWR.n77 VGND 8.78e-19
C3640 VPWR.n78 VGND 8.2e-19
C3641 VPWR.n79 VGND 0.001463f
C3642 VPWR.n80 VGND 6.56e-19
C3643 VPWR.n81 VGND 0.001281f
C3644 VPWR.n82 VGND 8.2e-19
C3645 VPWR.n83 VGND 0.001224f
C3646 VPWR.n84 VGND 6.25e-19
C3647 VPWR.n85 VGND 0.00128f
C3648 VPWR.n86 VGND 8.2e-19
C3649 VPWR.n87 VGND 0.001995f
C3650 VPWR.n88 VGND 0.002447f
C3651 VPWR.n89 VGND 0.002447f
C3652 VPWR.n90 VGND 5.18e-19
C3653 VPWR.n91 VGND 0.001404f
C3654 VPWR.t21 VGND 0.001178f
C3655 VPWR.n92 VGND 0.00288f
C3656 VPWR.t160 VGND 7.48e-19
C3657 VPWR.t799 VGND 7.48e-19
C3658 VPWR.n93 VGND 0.001623f
C3659 VPWR.t189 VGND 7.48e-19
C3660 VPWR.t19 VGND 7.48e-19
C3661 VPWR.n94 VGND 0.001676f
C3662 VPWR.n95 VGND 0.002147f
C3663 VPWR.n96 VGND 0.001871f
C3664 VPWR.n97 VGND 3.91e-19
C3665 VPWR.n98 VGND 0.002447f
C3666 VPWR.n99 VGND 0.002447f
C3667 VPWR.n100 VGND 0.00145f
C3668 VPWR.n101 VGND 8.67e-19
C3669 VPWR.n102 VGND 7.3e-19
C3670 VPWR.n103 VGND 9.31e-19
C3671 VPWR.n104 VGND 0.003245f
C3672 VPWR.n105 VGND 3.06e-19
C3673 VPWR.n106 VGND 0.002866f
C3674 VPWR.n107 VGND 0.001281f
C3675 VPWR.n108 VGND 6.56e-19
C3676 VPWR.n109 VGND 8.2e-19
C3677 VPWR.n110 VGND 6.12e-19
C3678 VPWR.n111 VGND 0.001224f
C3679 VPWR.n112 VGND 8.51e-19
C3680 VPWR.t473 VGND 0.002088f
C3681 VPWR.t921 VGND 0.004432f
C3682 VPWR.n114 VGND 0.011362f
C3683 VPWR.t474 VGND 0.002088f
C3684 VPWR.n115 VGND 0.006189f
C3685 VPWR.n116 VGND 0.005096f
C3686 VPWR.n117 VGND 5.72e-19
C3687 VPWR.n118 VGND 0.001199f
C3688 VPWR.n119 VGND 8.78e-19
C3689 VPWR.n120 VGND 8.2e-19
C3690 VPWR.n121 VGND 6.56e-19
C3691 VPWR.n122 VGND 0.001463f
C3692 VPWR.n123 VGND 0.001414f
C3693 VPWR.n124 VGND 0.058516f
C3694 VPWR.n125 VGND 0.001414f
C3695 VPWR.n126 VGND 0.048231f
C3696 VPWR.n127 VGND 0.001281f
C3697 VPWR.n128 VGND 0.001463f
C3698 VPWR.n129 VGND 8.2e-19
C3699 VPWR.n130 VGND 8.51e-19
C3700 VPWR.n131 VGND 0.002273f
C3701 VPWR.t426 VGND 0.002088f
C3702 VPWR.t914 VGND 0.004432f
C3703 VPWR.n133 VGND 0.011362f
C3704 VPWR.t427 VGND 0.002088f
C3705 VPWR.n134 VGND 0.006189f
C3706 VPWR.n135 VGND 0.002447f
C3707 VPWR.t158 VGND 7.76e-19
C3708 VPWR.t749 VGND 8.59e-19
C3709 VPWR.n136 VGND 0.001654f
C3710 VPWR.n137 VGND 0.006836f
C3711 VPWR.t108 VGND 0.001178f
C3712 VPWR.n138 VGND 0.002692f
C3713 VPWR.t392 VGND 7.48e-19
C3714 VPWR.t110 VGND 7.48e-19
C3715 VPWR.n139 VGND 0.00168f
C3716 VPWR.n140 VGND 0.002812f
C3717 VPWR.t196 VGND 3.14e-19
C3718 VPWR.t797 VGND 3.14e-19
C3719 VPWR.n141 VGND 7.27e-19
C3720 VPWR.t747 VGND 4.65e-19
C3721 VPWR.t25 VGND -4.89e-19
C3722 VPWR.n142 VGND 0.003099f
C3723 VPWR.n143 VGND 0.00182f
C3724 VPWR.n144 VGND 0.001224f
C3725 VPWR.n145 VGND 8.2e-19
C3726 VPWR.n146 VGND 0.001463f
C3727 VPWR.n147 VGND 6.56e-19
C3728 VPWR.t777 VGND 0.001025f
C3729 VPWR.t742 VGND 7.76e-19
C3730 VPWR.n148 VGND 0.001949f
C3731 VPWR.n149 VGND 0.003882f
C3732 VPWR.n150 VGND 0.001835f
C3733 VPWR.t775 VGND 0.002616f
C3734 VPWR.t808 VGND 0.001144f
C3735 VPWR.t176 VGND 4.79e-19
C3736 VPWR.t63 VGND 4.79e-19
C3737 VPWR.n151 VGND 9.97e-19
C3738 VPWR.n152 VGND 0.002783f
C3739 VPWR.t127 VGND 0.002987f
C3740 VPWR.t597 VGND 0.002071f
C3741 VPWR.t582 VGND 0.002279f
C3742 VPWR.n153 VGND 0.004985f
C3743 VPWR.n154 VGND 0.002447f
C3744 VPWR.t842 VGND 0.008643f
C3745 VPWR.n155 VGND 0.006969f
C3746 VPWR.n156 VGND 8.51e-19
C3747 VPWR.n157 VGND 8.2e-19
C3748 VPWR.n158 VGND 0.001463f
C3749 VPWR.n159 VGND 0.048231f
C3750 VPWR.n160 VGND 0.001463f
C3751 VPWR.n161 VGND 0.001146f
C3752 VPWR.n162 VGND 6.56e-19
C3753 VPWR.n163 VGND 6.56e-19
C3754 VPWR.n164 VGND 8.2e-19
C3755 VPWR.n165 VGND 0.001224f
C3756 VPWR.t862 VGND 0.030181f
C3757 VPWR.n166 VGND 0.005302f
C3758 VPWR.n167 VGND 0.002221f
C3759 VPWR.t681 VGND 0.002279f
C3760 VPWR.n168 VGND 0.001467f
C3761 VPWR.n169 VGND 0.002447f
C3762 VPWR.t605 VGND 0.002279f
C3763 VPWR.n170 VGND 0.002879f
C3764 VPWR.t403 VGND 0.002279f
C3765 VPWR.n171 VGND 0.002879f
C3766 VPWR.n172 VGND 0.001622f
C3767 VPWR.t830 VGND 0.030181f
C3768 VPWR.n173 VGND 0.005302f
C3769 VPWR.n174 VGND 8.78e-19
C3770 VPWR.n175 VGND 8.2e-19
C3771 VPWR.n176 VGND 0.001463f
C3772 VPWR.n177 VGND 0.048231f
C3773 VPWR.n178 VGND 0.048231f
C3774 VPWR.n179 VGND 0.001463f
C3775 VPWR.n180 VGND 0.001225f
C3776 VPWR.n181 VGND 6.56e-19
C3777 VPWR.n182 VGND 0.003633f
C3778 VPWR.n183 VGND 0.002447f
C3779 VPWR.t402 VGND 0.002279f
C3780 VPWR.n184 VGND 0.004408f
C3781 VPWR.n185 VGND 0.004429f
C3782 VPWR.t412 VGND 0.002285f
C3783 VPWR.n186 VGND 0.006775f
C3784 VPWR.t563 VGND 0.027522f
C3785 VPWR.t531 VGND 0.030188f
C3786 VPWR.t592 VGND 0.045556f
C3787 VPWR.t437 VGND 0.026581f
C3788 VPWR.t566 VGND 0.045556f
C3789 VPWR.t410 VGND 0.041008f
C3790 VPWR.t425 VGND 0.021641f
C3791 VPWR.t748 VGND 0.01921f
C3792 VPWR.t157 VGND 0.013722f
C3793 VPWR.t194 VGND 0.007214f
C3794 VPWR.t569 VGND 0.002744f
C3795 VPWR.t109 VGND 0.019681f
C3796 VPWR.t391 VGND 0.015917f
C3797 VPWR.t107 VGND 0.005097f
C3798 VPWR.t796 VGND 0.008939f
C3799 VPWR.t389 VGND 0.006586f
C3800 VPWR.t195 VGND 0.006586f
C3801 VPWR.t64 VGND 0.007292f
C3802 VPWR.t746 VGND 0.007449f
C3803 VPWR.t688 VGND 0.007449f
C3804 VPWR.t24 VGND 0.01035f
C3805 VPWR.t393 VGND 0.009644f
C3806 VPWR.t741 VGND 0.00541f
C3807 VPWR.t61 VGND 0.007449f
C3808 VPWR.t776 VGND 0.007449f
C3809 VPWR.t390 VGND 0.006586f
C3810 VPWR.t774 VGND 0.006665f
C3811 VPWR.t807 VGND 0.009723f
C3812 VPWR.t733 VGND 0.005332f
C3813 VPWR.t62 VGND 0.005645f
C3814 VPWR.t126 VGND 0.006586f
C3815 VPWR.t175 VGND 0.003685f
C3816 VPWR.t595 VGND 0.030188f
C3817 VPWR.n187 VGND 0.025192f
C3818 VPWR.t580 VGND 0.041008f
C3819 VPWR.t604 VGND 0.045556f
C3820 VPWR.t679 VGND 0.041008f
C3821 VPWR.t401 VGND 0.045556f
C3822 VPWR.t496 VGND 0.036068f
C3823 VPWR.n188 VGND 0.030131f
C3824 VPWR.t568 VGND 0.002279f
C3825 VPWR.n189 VGND 0.002879f
C3826 VPWR.n190 VGND 8.51e-19
C3827 VPWR.n191 VGND 8.2e-19
C3828 VPWR.n192 VGND 0.001463f
C3829 VPWR.n193 VGND 0.048231f
C3830 VPWR.n194 VGND 0.048231f
C3831 VPWR.n195 VGND 0.001463f
C3832 VPWR.n196 VGND 0.001225f
C3833 VPWR.n197 VGND 6.56e-19
C3834 VPWR.n198 VGND 8.51e-19
C3835 VPWR.n199 VGND 0.001224f
C3836 VPWR.t903 VGND 0.030181f
C3837 VPWR.n200 VGND 0.005302f
C3838 VPWR.n201 VGND 0.002221f
C3839 VPWR.t439 VGND 0.002279f
C3840 VPWR.n202 VGND 0.002879f
C3841 VPWR.n203 VGND 0.002447f
C3842 VPWR.n204 VGND 0.003633f
C3843 VPWR.n205 VGND 0.002447f
C3844 VPWR.t894 VGND 0.030181f
C3845 VPWR.n206 VGND 0.016876f
C3846 VPWR.n207 VGND 0.001197f
C3847 VPWR.n208 VGND 8.2e-19
C3848 VPWR.n209 VGND 0.001463f
C3849 VPWR.n210 VGND 0.081008f
C3850 VPWR.n211 VGND 0.001414f
C3851 VPWR.n212 VGND 0.001463f
C3852 VPWR.n213 VGND 0.001092f
C3853 VPWR.n214 VGND 6.56e-19
C3854 VPWR.n215 VGND 0.001224f
C3855 VPWR.t892 VGND 0.015058f
C3856 VPWR.n216 VGND 0.011361f
C3857 VPWR.t453 VGND 0.002279f
C3858 VPWR.t514 VGND 0.002071f
C3859 VPWR.n217 VGND 0.004985f
C3860 VPWR.t485 VGND 0.002088f
C3861 VPWR.t902 VGND 0.004432f
C3862 VPWR.n219 VGND 0.011362f
C3863 VPWR.t486 VGND 0.002088f
C3864 VPWR.n220 VGND 0.006189f
C3865 VPWR.t585 VGND 0.002088f
C3866 VPWR.t875 VGND 0.004432f
C3867 VPWR.n222 VGND 0.011362f
C3868 VPWR.t586 VGND 0.002088f
C3869 VPWR.n223 VGND 0.006189f
C3870 VPWR.n224 VGND 0.005099f
C3871 VPWR.t441 VGND 0.002088f
C3872 VPWR.t911 VGND 0.004432f
C3873 VPWR.n226 VGND 0.011362f
C3874 VPWR.t442 VGND 0.002088f
C3875 VPWR.n227 VGND 0.006189f
C3876 VPWR.n228 VGND 0.001597f
C3877 VPWR.n229 VGND 0.00206f
C3878 VPWR.t549 VGND 0.002088f
C3879 VPWR.t886 VGND 0.004432f
C3880 VPWR.n231 VGND 0.011362f
C3881 VPWR.t550 VGND 0.002088f
C3882 VPWR.n232 VGND 0.006189f
C3883 VPWR.n233 VGND 0.005594f
C3884 VPWR.n234 VGND 0.001376f
C3885 VPWR.n235 VGND 0.001597f
C3886 VPWR.n236 VGND 0.001835f
C3887 VPWR.n237 VGND 0.001463f
C3888 VPWR.n238 VGND 0.00634f
C3889 VPWR.n239 VGND 0.010674f
C3890 VPWR.t926 VGND 0.030181f
C3891 VPWR.n240 VGND 0.016876f
C3892 VPWR.n241 VGND 0.002447f
C3893 VPWR.t515 VGND 0.002071f
C3894 VPWR.n242 VGND 0.004756f
C3895 VPWR.t488 VGND 0.002279f
C3896 VPWR.n243 VGND 0.002879f
C3897 VPWR.n244 VGND 0.002447f
C3898 VPWR.t901 VGND 0.030753f
C3899 VPWR.n245 VGND 0.014263f
C3900 VPWR.n246 VGND 0.002447f
C3901 VPWR.n247 VGND 0.004063f
C3902 VPWR.n248 VGND 8.51e-19
C3903 VPWR.n249 VGND 8.2e-19
C3904 VPWR.n250 VGND 0.001463f
C3905 VPWR.n251 VGND 0.001414f
C3906 VPWR.n252 VGND 0.001463f
C3907 VPWR.n253 VGND 0.001225f
C3908 VPWR.n254 VGND 6.56e-19
C3909 VPWR.n255 VGND 8.51e-19
C3910 VPWR.n256 VGND 8.51e-19
C3911 VPWR.n257 VGND 0.001281f
C3912 VPWR.n258 VGND 0.001225f
C3913 VPWR.t856 VGND 0.030181f
C3914 VPWR.n259 VGND 0.005302f
C3915 VPWR.n260 VGND 0.002221f
C3916 VPWR.t931 VGND 0.030753f
C3917 VPWR.t644 VGND 0.002279f
C3918 VPWR.n261 VGND 0.002879f
C3919 VPWR.n262 VGND 0.002447f
C3920 VPWR.n263 VGND 0.003633f
C3921 VPWR.n264 VGND 0.002447f
C3922 VPWR.t849 VGND 0.030181f
C3923 VPWR.n265 VGND 0.016876f
C3924 VPWR.n266 VGND 0.001197f
C3925 VPWR.n267 VGND 8.2e-19
C3926 VPWR.n268 VGND 0.001463f
C3927 VPWR.n269 VGND 0.001463f
C3928 VPWR.n270 VGND 0.001092f
C3929 VPWR.n271 VGND 6.56e-19
C3930 VPWR.n272 VGND 6.56e-19
C3931 VPWR.n273 VGND 8.2e-19
C3932 VPWR.n274 VGND 0.001224f
C3933 VPWR.t923 VGND 0.015058f
C3934 VPWR.n275 VGND 0.011361f
C3935 VPWR.t643 VGND 0.002279f
C3936 VPWR.t646 VGND 0.002071f
C3937 VPWR.n276 VGND 0.004985f
C3938 VPWR.t625 VGND 0.002088f
C3939 VPWR.t932 VGND 0.004432f
C3940 VPWR.n278 VGND 0.011362f
C3941 VPWR.t626 VGND 0.002088f
C3942 VPWR.n279 VGND 0.006189f
C3943 VPWR.t491 VGND 0.002088f
C3944 VPWR.t904 VGND 0.004432f
C3945 VPWR.n281 VGND 0.011362f
C3946 VPWR.t492 VGND 0.002088f
C3947 VPWR.n282 VGND 0.006189f
C3948 VPWR.n283 VGND 0.005099f
C3949 VPWR.t590 VGND 0.002088f
C3950 VPWR.t837 VGND 0.004432f
C3951 VPWR.n285 VGND 0.011362f
C3952 VPWR.t591 VGND 0.002088f
C3953 VPWR.n286 VGND 0.006189f
C3954 VPWR.n287 VGND 0.001597f
C3955 VPWR.n288 VGND 0.00206f
C3956 VPWR.t465 VGND 0.002088f
C3957 VPWR.t917 VGND 0.004432f
C3958 VPWR.n290 VGND 0.011362f
C3959 VPWR.t466 VGND 0.002088f
C3960 VPWR.n291 VGND 0.006189f
C3961 VPWR.n292 VGND 0.005594f
C3962 VPWR.n293 VGND 0.001376f
C3963 VPWR.n294 VGND 0.001597f
C3964 VPWR.n295 VGND 0.001835f
C3965 VPWR.n296 VGND 0.001463f
C3966 VPWR.n297 VGND 0.00634f
C3967 VPWR.n298 VGND 0.010674f
C3968 VPWR.n299 VGND 8.51e-19
C3969 VPWR.n300 VGND 0.006622f
C3970 VPWR.n301 VGND 0.00634f
C3971 VPWR.n302 VGND 8.51e-19
C3972 VPWR.n303 VGND 9.84e-19
C3973 VPWR.n304 VGND 8.2e-19
C3974 VPWR.n305 VGND 0.001281f
C3975 VPWR.n306 VGND 0.001414f
C3976 VPWR.n307 VGND 0.064545f
C3977 VPWR.n308 VGND 0.001414f
C3978 VPWR.n309 VGND 0.001281f
C3979 VPWR.n310 VGND 8.8e-19
C3980 VPWR.n311 VGND 0.00125f
C3981 VPWR.n312 VGND 0.00634f
C3982 VPWR.n313 VGND 0.008641f
C3983 VPWR.t647 VGND 0.002071f
C3984 VPWR.n314 VGND 0.004756f
C3985 VPWR.n315 VGND 0.008359f
C3986 VPWR.n316 VGND 0.002447f
C3987 VPWR.n317 VGND 0.00145f
C3988 VPWR.n318 VGND 0.001835f
C3989 VPWR.n319 VGND 0.002332f
C3990 VPWR.t628 VGND 0.002279f
C3991 VPWR.n320 VGND 0.002879f
C3992 VPWR.n321 VGND 0.005129f
C3993 VPWR.n322 VGND 0.005129f
C3994 VPWR.n323 VGND 0.002447f
C3995 VPWR.n324 VGND 0.00145f
C3996 VPWR.n325 VGND 0.001334f
C3997 VPWR.n326 VGND 0.014263f
C3998 VPWR.n327 VGND 0.001191f
C3999 VPWR.t618 VGND 0.002279f
C4000 VPWR.n328 VGND 0.002879f
C4001 VPWR.n329 VGND 0.005129f
C4002 VPWR.n330 VGND 0.002447f
C4003 VPWR.n331 VGND 0.002447f
C4004 VPWR.n332 VGND 0.001888f
C4005 VPWR.n333 VGND 0.004063f
C4006 VPWR.n334 VGND 0.015206f
C4007 VPWR.n335 VGND 0.00389f
C4008 VPWR.n336 VGND 0.005302f
C4009 VPWR.t619 VGND 0.002285f
C4010 VPWR.n337 VGND 0.006775f
C4011 VPWR.t490 VGND 0.027522f
C4012 VPWR.t464 VGND 0.030188f
C4013 VPWR.t645 VGND 0.045556f
C4014 VPWR.t642 VGND 0.026581f
C4015 VPWR.t627 VGND 0.045556f
C4016 VPWR.t617 VGND 0.041008f
C4017 VPWR.n338 VGND 0.001882f
C4018 VPWR.n339 VGND 8.51e-19
C4019 VPWR.n340 VGND 8.2e-19
C4020 VPWR.n341 VGND 0.001463f
C4021 VPWR.n342 VGND 6.56e-19
C4022 VPWR.n343 VGND 8.51e-19
C4023 VPWR.n344 VGND 0.001224f
C4024 VPWR.n345 VGND 0.005302f
C4025 VPWR.n346 VGND 0.002447f
C4026 VPWR.t927 VGND 0.030181f
C4027 VPWR.t898 VGND 0.030181f
C4028 VPWR.n347 VGND 0.027762f
C4029 VPWR.n348 VGND 0.002447f
C4030 VPWR.t511 VGND 0.002279f
C4031 VPWR.t637 VGND 0.002279f
C4032 VPWR.n349 VGND 0.003107f
C4033 VPWR.t616 VGND 0.002279f
C4034 VPWR.t448 VGND 0.002279f
C4035 VPWR.n350 VGND 0.003107f
C4036 VPWR.n351 VGND 0.001622f
C4037 VPWR.n352 VGND 0.001197f
C4038 VPWR.n353 VGND 8.78e-19
C4039 VPWR.n354 VGND 6.56e-19
C4040 VPWR.n355 VGND 8.2e-19
C4041 VPWR.n356 VGND 0.001281f
C4042 VPWR.n357 VGND 0.001225f
C4043 VPWR.n358 VGND 8.51e-19
C4044 VPWR.n359 VGND 0.005302f
C4045 VPWR.n360 VGND 0.005302f
C4046 VPWR.n361 VGND 0.005129f
C4047 VPWR.n362 VGND 0.002447f
C4048 VPWR.n363 VGND 0.002002f
C4049 VPWR.n364 VGND 0.001958f
C4050 VPWR.n365 VGND 0.002221f
C4051 VPWR.n366 VGND 0.002447f
C4052 VPWR.n367 VGND 0.005129f
C4053 VPWR.n368 VGND 0.005302f
C4054 VPWR.n369 VGND 0.004063f
C4055 VPWR.n370 VGND 0.002447f
C4056 VPWR.n371 VGND 0.002447f
C4057 VPWR.n372 VGND 0.00389f
C4058 VPWR.n373 VGND 0.005302f
C4059 VPWR.n374 VGND 0.005302f
C4060 VPWR.n375 VGND 0.002447f
C4061 VPWR.n376 VGND 0.002447f
C4062 VPWR.n377 VGND 9.31e-19
C4063 VPWR.n378 VGND 8.2e-19
C4064 VPWR.n379 VGND 0.001414f
C4065 VPWR.n380 VGND 0.001281f
C4066 VPWR.n381 VGND 0.001146f
C4067 VPWR.n382 VGND 0.001516f
C4068 VPWR.n383 VGND 0.005302f
C4069 VPWR.n384 VGND 0.005302f
C4070 VPWR.t512 VGND 0.002279f
C4071 VPWR.t638 VGND 0.002279f
C4072 VPWR.n385 VGND 0.003107f
C4073 VPWR.n386 VGND 0.005129f
C4074 VPWR.n387 VGND 8.51e-19
C4075 VPWR.n388 VGND 0.001224f
C4076 VPWR.n389 VGND 8.2e-19
C4077 VPWR.n390 VGND 6.56e-19
C4078 VPWR.n391 VGND 0.001463f
C4079 VPWR.n392 VGND 0.001414f
C4080 VPWR.n393 VGND 0.001281f
C4081 VPWR.n394 VGND 2.28e-19
C4082 VPWR.n395 VGND 0.001317f
C4083 VPWR.n396 VGND 0.001256f
C4084 VPWR.n397 VGND 0.002447f
C4085 VPWR.t508 VGND 0.002279f
C4086 VPWR.n398 VGND 0.00164f
C4087 VPWR.t887 VGND 0.015325f
C4088 VPWR.t900 VGND 0.030181f
C4089 VPWR.n399 VGND 0.016876f
C4090 VPWR.n400 VGND 0.002447f
C4091 VPWR.n401 VGND 0.008359f
C4092 VPWR.t451 VGND 0.002071f
C4093 VPWR.n402 VGND 0.004756f
C4094 VPWR.t168 VGND 6.35e-19
C4095 VPWR.t314 VGND 6.35e-19
C4096 VPWR.n403 VGND 0.00138f
C4097 VPWR.n404 VGND 0.005652f
C4098 VPWR.n405 VGND 6.14e-19
C4099 VPWR.n406 VGND 8.78e-19
C4100 VPWR.n407 VGND 0.001281f
C4101 VPWR.n408 VGND 8.2e-19
C4102 VPWR.n409 VGND 0.001463f
C4103 VPWR.n410 VGND 6.56e-19
C4104 VPWR.n411 VGND 8.2e-19
C4105 VPWR.n412 VGND 0.002447f
C4106 VPWR.t509 VGND 0.002279f
C4107 VPWR.n413 VGND 0.00177f
C4108 VPWR.n414 VGND 8.51e-19
C4109 VPWR.n415 VGND 0.001224f
C4110 VPWR.n416 VGND 6.25e-19
C4111 VPWR.n417 VGND 0.001219f
C4112 VPWR.t482 VGND 0.002279f
C4113 VPWR.n418 VGND 0.004063f
C4114 VPWR.n419 VGND 0.002447f
C4115 VPWR.t834 VGND 0.030181f
C4116 VPWR.t908 VGND 0.030181f
C4117 VPWR.n420 VGND 0.027762f
C4118 VPWR.n421 VGND 0.005302f
C4119 VPWR.n422 VGND 0.002447f
C4120 VPWR.t483 VGND 0.002279f
C4121 VPWR.t611 VGND 0.002279f
C4122 VPWR.n423 VGND 0.003107f
C4123 VPWR.n424 VGND 3.06e-19
C4124 VPWR.n425 VGND 8.2e-19
C4125 VPWR.n426 VGND 0.001463f
C4126 VPWR.n427 VGND 0.001281f
C4127 VPWR.n428 VGND 6.56e-19
C4128 VPWR.n429 VGND 8.2e-19
C4129 VPWR.n430 VGND 8.51e-19
C4130 VPWR.n431 VGND 0.001882f
C4131 VPWR.t503 VGND 0.002088f
C4132 VPWR.t867 VGND 0.004432f
C4133 VPWR.n433 VGND 0.011362f
C4134 VPWR.t504 VGND 0.002088f
C4135 VPWR.n434 VGND 0.006189f
C4136 VPWR.n435 VGND 9.97e-19
C4137 VPWR.n436 VGND 0.001224f
C4138 VPWR.n437 VGND 8.51e-19
C4139 VPWR.t661 VGND 0.002088f
C4140 VPWR.t845 VGND 0.004432f
C4141 VPWR.n439 VGND 0.011362f
C4142 VPWR.t662 VGND 0.002088f
C4143 VPWR.n440 VGND 0.006189f
C4144 VPWR.n441 VGND 0.005218f
C4145 VPWR.n442 VGND 5.72e-19
C4146 VPWR.n443 VGND 0.001199f
C4147 VPWR.n444 VGND 8.78e-19
C4148 VPWR.n445 VGND 8.2e-19
C4149 VPWR.n446 VGND 6.56e-19
C4150 VPWR.n447 VGND 0.001463f
C4151 VPWR.n448 VGND 0.001414f
C4152 VPWR.n449 VGND 0.06951f
C4153 VPWR.n450 VGND 0.048231f
C4154 VPWR.n451 VGND 0.064545f
C4155 VPWR.n452 VGND 0.001414f
C4156 VPWR.n453 VGND 0.001281f
C4157 VPWR.n454 VGND 0.001225f
C4158 VPWR.n455 VGND 0.002367f
C4159 VPWR.n456 VGND 0.005129f
C4160 VPWR.n457 VGND 0.005302f
C4161 VPWR.n458 VGND 0.005302f
C4162 VPWR.n459 VGND 0.002447f
C4163 VPWR.n460 VGND 0.002447f
C4164 VPWR.n461 VGND 0.002447f
C4165 VPWR.n462 VGND 0.005302f
C4166 VPWR.n463 VGND 0.005302f
C4167 VPWR.n464 VGND 0.00389f
C4168 VPWR.n465 VGND 0.002447f
C4169 VPWR.n466 VGND 0.002447f
C4170 VPWR.n467 VGND 0.002447f
C4171 VPWR.n468 VGND 0.005302f
C4172 VPWR.n469 VGND 0.005129f
C4173 VPWR.t610 VGND 0.002279f
C4174 VPWR.n470 VGND 0.003107f
C4175 VPWR.n471 VGND 0.001969f
C4176 VPWR.n472 VGND 0.001835f
C4177 VPWR.n473 VGND 3.88e-19
C4178 VPWR.n474 VGND 0.001281f
C4179 VPWR.n475 VGND 0.001414f
C4180 VPWR.n476 VGND 0.064545f
C4181 VPWR.n477 VGND 0.001414f
C4182 VPWR.n478 VGND 0.001463f
C4183 VPWR.n479 VGND 6.56e-19
C4184 VPWR.n480 VGND 8.2e-19
C4185 VPWR.n481 VGND 9.71e-19
C4186 VPWR.n482 VGND 7.31e-19
C4187 VPWR.n483 VGND 0.002939f
C4188 VPWR.n484 VGND 0.00372f
C4189 VPWR.n485 VGND 0.00145f
C4190 VPWR.n486 VGND 0.002447f
C4191 VPWR.n487 VGND 0.002447f
C4192 VPWR.n488 VGND 0.008641f
C4193 VPWR.n489 VGND 0.008641f
C4194 VPWR.n490 VGND 0.00634f
C4195 VPWR.n491 VGND 0.002447f
C4196 VPWR.n492 VGND 0.002447f
C4197 VPWR.n493 VGND 0.004367f
C4198 VPWR.n494 VGND 0.021777f
C4199 VPWR.n495 VGND 0.006293f
C4200 VPWR.t450 VGND 0.002071f
C4201 VPWR.n496 VGND 0.004756f
C4202 VPWR.n497 VGND 0.003605f
C4203 VPWR.n498 VGND 0.001835f
C4204 VPWR.n499 VGND 9.44e-19
C4205 VPWR.n500 VGND 9.31e-19
C4206 VPWR.n501 VGND 6.83e-19
C4207 VPWR.n502 VGND 0.009208f
C4208 VPWR.t502 VGND 0.021641f
C4209 VPWR.t481 VGND 0.086564f
C4210 VPWR.t313 VGND 0.011997f
C4211 VPWR.t167 VGND 0.009331f
C4212 VPWR.t507 VGND 0.026581f
C4213 VPWR.t449 VGND 0.038264f
C4214 VPWR.n503 VGND 0.016974f
C4215 VPWR.t510 VGND 0.086564f
C4216 VPWR.t446 VGND 0.086564f
C4217 VPWR.t458 VGND 0.022974f
C4218 VPWR.n504 VGND 0.021585f
C4219 VPWR.n505 VGND 0.006627f
C4220 VPWR.n506 VGND 0.001317f
C4221 VPWR.n507 VGND 0.001051f
C4222 VPWR.n508 VGND 0.002501f
C4223 VPWR.t629 VGND 0.002279f
C4224 VPWR.n509 VGND 0.002879f
C4225 VPWR.n510 VGND 0.005129f
C4226 VPWR.n511 VGND 8.51e-19
C4227 VPWR.n512 VGND 0.001224f
C4228 VPWR.n513 VGND 8.2e-19
C4229 VPWR.n514 VGND 0.001463f
C4230 VPWR.n515 VGND 6.56e-19
C4231 VPWR.n516 VGND 8.2e-19
C4232 VPWR.n517 VGND 9.31e-19
C4233 VPWR.n518 VGND 0.001144f
C4234 VPWR.n519 VGND 8.2e-19
C4235 VPWR.n520 VGND 0.001281f
C4236 VPWR.n521 VGND 0.001414f
C4237 VPWR.n522 VGND 0.064545f
C4238 VPWR.n523 VGND 0.048231f
C4239 VPWR.n524 VGND 0.001463f
C4240 VPWR.n525 VGND 8.2e-19
C4241 VPWR.n526 VGND 8.51e-19
C4242 VPWR.t832 VGND 0.030181f
C4243 VPWR.n527 VGND 0.015206f
C4244 VPWR.n528 VGND 0.00389f
C4245 VPWR.n529 VGND 0.001144f
C4246 VPWR.n530 VGND 6.56e-19
C4247 VPWR.n531 VGND 6.56e-19
C4248 VPWR.n532 VGND 8.2e-19
C4249 VPWR.n533 VGND 9.31e-19
C4250 VPWR.n534 VGND 0.001224f
C4251 VPWR.n535 VGND 8.51e-19
C4252 VPWR.n536 VGND 0.005302f
C4253 VPWR.n537 VGND 0.005129f
C4254 VPWR.t489 VGND 0.002279f
C4255 VPWR.n538 VGND 0.002879f
C4256 VPWR.t484 VGND 0.027522f
C4257 VPWR.t440 VGND 0.030188f
C4258 VPWR.t513 VGND 0.045556f
C4259 VPWR.t452 VGND 0.026581f
C4260 VPWR.t487 VGND 0.045556f
C4261 VPWR.t416 VGND 0.041008f
C4262 VPWR.t601 VGND 0.041008f
C4263 VPWR.t607 VGND 0.045556f
C4264 VPWR.t634 VGND 0.041008f
C4265 VPWR.t407 VGND 0.045556f
C4266 VPWR.t422 VGND 0.014427f
C4267 VPWR.n539 VGND 0.015547f
C4268 VPWR.n540 VGND 0.002598f
C4269 VPWR.n541 VGND 0.001766f
C4270 VPWR.t408 VGND 0.002286f
C4271 VPWR.t635 VGND 0.002279f
C4272 VPWR.n542 VGND 0.002879f
C4273 VPWR.n543 VGND 0.002447f
C4274 VPWR.t835 VGND 0.030181f
C4275 VPWR.t847 VGND 0.030181f
C4276 VPWR.n544 VGND 0.015206f
C4277 VPWR.n545 VGND 8.51e-19
C4278 VPWR.n546 VGND 8.2e-19
C4279 VPWR.n547 VGND 6.56e-19
C4280 VPWR.n548 VGND 6.56e-19
C4281 VPWR.n549 VGND 8.2e-19
C4282 VPWR.n550 VGND 8.51e-19
C4283 VPWR.n551 VGND 0.002447f
C4284 VPWR.n552 VGND 0.00389f
C4285 VPWR.n553 VGND 0.001224f
C4286 VPWR.n554 VGND 8.78e-19
C4287 VPWR.n555 VGND 8.2e-19
C4288 VPWR.n556 VGND 0.001197f
C4289 VPWR.n557 VGND 8.51e-19
C4290 VPWR.n558 VGND 0.005302f
C4291 VPWR.n559 VGND 0.005302f
C4292 VPWR.t636 VGND 0.002286f
C4293 VPWR.n560 VGND 0.004675f
C4294 VPWR.t608 VGND 0.002286f
C4295 VPWR.t602 VGND 0.002279f
C4296 VPWR.n561 VGND 0.002879f
C4297 VPWR.n562 VGND 0.002447f
C4298 VPWR.t866 VGND 0.030181f
C4299 VPWR.t854 VGND 0.030181f
C4300 VPWR.n563 VGND 0.015206f
C4301 VPWR.n564 VGND 0.001516f
C4302 VPWR.n565 VGND 0.002447f
C4303 VPWR.n566 VGND 0.005302f
C4304 VPWR.n567 VGND 0.00389f
C4305 VPWR.n568 VGND 0.002447f
C4306 VPWR.n569 VGND 0.002447f
C4307 VPWR.n570 VGND 0.004063f
C4308 VPWR.n571 VGND 0.00389f
C4309 VPWR.n572 VGND 0.015206f
C4310 VPWR.n573 VGND 0.00389f
C4311 VPWR.n574 VGND 0.002447f
C4312 VPWR.n575 VGND 0.002221f
C4313 VPWR.n576 VGND 0.001931f
C4314 VPWR.n577 VGND 0.004635f
C4315 VPWR.n578 VGND 0.001796f
C4316 VPWR.n579 VGND 0.001766f
C4317 VPWR.n580 VGND 0.00145f
C4318 VPWR.n581 VGND 0.001968f
C4319 VPWR.t409 VGND 0.002279f
C4320 VPWR.n582 VGND 0.002879f
C4321 VPWR.n583 VGND 0.005129f
C4322 VPWR.n584 VGND 0.005302f
C4323 VPWR.n585 VGND 0.001622f
C4324 VPWR.n586 VGND 0.001225f
C4325 VPWR.n587 VGND 0.001281f
C4326 VPWR.n588 VGND 0.001414f
C4327 VPWR.n589 VGND 0.001463f
C4328 VPWR.n590 VGND 0.001463f
C4329 VPWR.n591 VGND 0.001414f
C4330 VPWR.n592 VGND 0.001281f
C4331 VPWR.n593 VGND 0.001225f
C4332 VPWR.n594 VGND 0.002314f
C4333 VPWR.n595 VGND 0.004063f
C4334 VPWR.n596 VGND 0.00389f
C4335 VPWR.n597 VGND 0.015206f
C4336 VPWR.n598 VGND 0.00389f
C4337 VPWR.n599 VGND 0.002447f
C4338 VPWR.n600 VGND 0.001835f
C4339 VPWR.n601 VGND 0.001931f
C4340 VPWR.n602 VGND 0.004635f
C4341 VPWR.n603 VGND 0.002929f
C4342 VPWR.t424 VGND 0.002102f
C4343 VPWR.n604 VGND 0.006134f
C4344 VPWR.n605 VGND 0.006514f
C4345 VPWR.t915 VGND 0.008778f
C4346 VPWR.n606 VGND 0.008691f
C4347 VPWR.t423 VGND 0.002071f
C4348 VPWR.n607 VGND 0.002493f
C4349 VPWR.t418 VGND 0.002286f
C4350 VPWR.n608 VGND 0.004685f
C4351 VPWR.n609 VGND 0.002494f
C4352 VPWR.n610 VGND 0.001307f
C4353 VPWR.n611 VGND 9.31e-19
C4354 VPWR.n612 VGND 0.001317f
C4355 VPWR.n613 VGND 0.007114f
C4356 VPWR.n614 VGND 0.002501f
C4357 VPWR.n615 VGND 0.001051f
C4358 VPWR.n616 VGND 0.001225f
C4359 VPWR.n617 VGND 0.001281f
C4360 VPWR.n618 VGND 0.001414f
C4361 VPWR.n619 VGND 0.058516f
C4362 VPWR.n620 VGND 0.001414f
C4363 VPWR.n621 VGND 0.001281f
C4364 VPWR.n622 VGND 0.001225f
C4365 VPWR.n623 VGND 0.001888f
C4366 VPWR.n624 VGND 0.002447f
C4367 VPWR.n625 VGND 0.005302f
C4368 VPWR.n626 VGND 0.005129f
C4369 VPWR.t417 VGND 0.002279f
C4370 VPWR.n627 VGND 0.002879f
C4371 VPWR.n628 VGND 0.001191f
C4372 VPWR.n629 VGND 0.002221f
C4373 VPWR.n630 VGND 0.00145f
C4374 VPWR.n631 VGND 0.001334f
C4375 VPWR.t454 VGND 0.002279f
C4376 VPWR.n632 VGND 0.002879f
C4377 VPWR.n633 VGND 0.005129f
C4378 VPWR.n634 VGND 0.005129f
C4379 VPWR.n635 VGND 0.002447f
C4380 VPWR.n636 VGND 0.001835f
C4381 VPWR.n637 VGND 0.002332f
C4382 VPWR.n638 VGND 0.003633f
C4383 VPWR.n639 VGND 0.00145f
C4384 VPWR.n640 VGND 0.002447f
C4385 VPWR.n641 VGND 0.008359f
C4386 VPWR.n642 VGND 0.008641f
C4387 VPWR.n643 VGND 0.00634f
C4388 VPWR.n644 VGND 0.00125f
C4389 VPWR.n645 VGND 8.8e-19
C4390 VPWR.n646 VGND 8.2e-19
C4391 VPWR.n647 VGND 0.001463f
C4392 VPWR.n648 VGND 6.56e-19
C4393 VPWR.n649 VGND 0.001281f
C4394 VPWR.n650 VGND 8.2e-19
C4395 VPWR.n651 VGND 0.001197f
C4396 VPWR.n652 VGND 8.51e-19
C4397 VPWR.n653 VGND 0.006622f
C4398 VPWR.n654 VGND 0.00634f
C4399 VPWR.n655 VGND 8.51e-19
C4400 VPWR.n656 VGND 9.84e-19
C4401 VPWR.n657 VGND 8.2e-19
C4402 VPWR.n658 VGND 0.001281f
C4403 VPWR.n659 VGND 0.001414f
C4404 VPWR.n660 VGND 0.058516f
C4405 VPWR.n661 VGND 0.117032f
C4406 VPWR.n662 VGND 0.221149f
C4407 VPWR.n663 VGND 0.081008f
C4408 VPWR.n664 VGND 0.058516f
C4409 VPWR.n665 VGND 0.06951f
C4410 VPWR.n666 VGND 0.001414f
C4411 VPWR.n667 VGND 0.048231f
C4412 VPWR.n668 VGND 0.001463f
C4413 VPWR.n669 VGND 0.001225f
C4414 VPWR.n670 VGND 6.56e-19
C4415 VPWR.n671 VGND 8.51e-19
C4416 VPWR.n672 VGND 8.51e-19
C4417 VPWR.n673 VGND 0.001281f
C4418 VPWR.t576 VGND 0.002279f
C4419 VPWR.n674 VGND 0.001783f
C4420 VPWR.t545 VGND 0.002279f
C4421 VPWR.n675 VGND 0.001783f
C4422 VPWR.n676 VGND 9.99e-19
C4423 VPWR.n677 VGND 0.002447f
C4424 VPWR.t262 VGND 7.76e-19
C4425 VPWR.t266 VGND 7.76e-19
C4426 VPWR.n678 VGND 0.001601f
C4427 VPWR.t268 VGND 7.76e-19
C4428 VPWR.t272 VGND 7.76e-19
C4429 VPWR.n679 VGND 0.001601f
C4430 VPWR.n680 VGND 0.002747f
C4431 VPWR.n681 VGND 0.002447f
C4432 VPWR.t876 VGND 0.030181f
C4433 VPWR.n682 VGND 0.014093f
C4434 VPWR.t242 VGND 7.76e-19
C4435 VPWR.t244 VGND 7.76e-19
C4436 VPWR.n683 VGND 0.001602f
C4437 VPWR.t248 VGND 0.002725f
C4438 VPWR.n684 VGND 0.003983f
C4439 VPWR.t652 VGND 0.002071f
C4440 VPWR.n685 VGND 0.002596f
C4441 VPWR.n686 VGND 0.002367f
C4442 VPWR.t929 VGND 0.008643f
C4443 VPWR.n687 VGND 0.008854f
C4444 VPWR.t653 VGND 0.002071f
C4445 VPWR.t420 VGND 0.002088f
C4446 VPWR.t916 VGND 0.004432f
C4447 VPWR.n689 VGND 0.011362f
C4448 VPWR.t421 VGND 0.002088f
C4449 VPWR.n690 VGND 0.006189f
C4450 VPWR.t542 VGND 0.002088f
C4451 VPWR.t855 VGND 0.004432f
C4452 VPWR.n692 VGND 0.011362f
C4453 VPWR.t543 VGND 0.002088f
C4454 VPWR.n693 VGND 0.006189f
C4455 VPWR.n694 VGND 0.005216f
C4456 VPWR.n695 VGND 0.001225f
C4457 VPWR.n696 VGND 8.51e-19
C4458 VPWR.n697 VGND 0.001281f
C4459 VPWR.n698 VGND 8.2e-19
C4460 VPWR.n699 VGND 0.001414f
C4461 VPWR.n700 VGND 6.56e-19
C4462 VPWR.n701 VGND 8.2e-19
C4463 VPWR.n702 VGND 0.001224f
C4464 VPWR.n703 VGND 8.51e-19
C4465 VPWR.n704 VGND 8.78e-19
C4466 VPWR.n705 VGND 5.72e-19
C4467 VPWR.n706 VGND 0.001199f
C4468 VPWR.n707 VGND 0.001281f
C4469 VPWR.n708 VGND 0.053551f
C4470 VPWR.n709 VGND 0.117032f
C4471 VPWR.n710 VGND 0.058516f
C4472 VPWR.n711 VGND 0.001414f
C4473 VPWR.n712 VGND 0.053196f
C4474 VPWR.n713 VGND 0.001463f
C4475 VPWR.n714 VGND 0.001146f
C4476 VPWR.n715 VGND 6.56e-19
C4477 VPWR.n716 VGND 0.001224f
C4478 VPWR.t883 VGND 0.008643f
C4479 VPWR.n717 VGND 0.007818f
C4480 VPWR.t56 VGND 4.77e-19
C4481 VPWR.t307 VGND 3.14e-19
C4482 VPWR.n718 VGND 8.14e-19
C4483 VPWR.n719 VGND 0.004625f
C4484 VPWR.n720 VGND 8.51e-19
C4485 VPWR.n721 VGND 8.2e-19
C4486 VPWR.n722 VGND 0.001463f
C4487 VPWR.n723 VGND 6.56e-19
C4488 VPWR.t480 VGND 0.002071f
C4489 VPWR.n724 VGND 0.003578f
C4490 VPWR.n725 VGND 0.002273f
C4491 VPWR.t534 VGND 0.021641f
C4492 VPWR.t428 VGND 0.041008f
C4493 VPWR.t639 VGND 0.023993f
C4494 VPWR.t121 VGND 0.010664f
C4495 VPWR.t703 VGND 0.016544f
C4496 VPWR.t229 VGND 0.01035f
C4497 VPWR.t73 VGND 0.016544f
C4498 VPWR.t317 VGND 0.011448f
C4499 VPWR.t152 VGND 0.014114f
C4500 VPWR.t75 VGND 0.015525f
C4501 VPWR.t16 VGND 0.018426f
C4502 VPWR.t145 VGND 0.014035f
C4503 VPWR.t670 VGND 0.007449f
C4504 VPWR.t76 VGND 0.01035f
C4505 VPWR.t151 VGND 0.015525f
C4506 VPWR.t99 VGND 0.025405f
C4507 VPWR.t280 VGND 0.023052f
C4508 VPWR.t97 VGND 0.009723f
C4509 VPWR.n726 VGND 0.015857f
C4510 VPWR.n727 VGND 0.001256f
C4511 VPWR.n728 VGND 0.002447f
C4512 VPWR.t98 VGND 7.48e-19
C4513 VPWR.t281 VGND 7.48e-19
C4514 VPWR.n729 VGND 0.001676f
C4515 VPWR.t671 VGND 0.002279f
C4516 VPWR.n730 VGND 3.62e-19
C4517 VPWR.n731 VGND 0.003165f
C4518 VPWR.t100 VGND 0.001168f
C4519 VPWR.t838 VGND 0.030181f
C4520 VPWR.n732 VGND 0.014097f
C4521 VPWR.n733 VGND 0.002447f
C4522 VPWR.t146 VGND 5.61e-19
C4523 VPWR.t17 VGND 0.001157f
C4524 VPWR.n734 VGND 0.002356f
C4525 VPWR.n735 VGND 0.002939f
C4526 VPWR.n736 VGND 0.001942f
C4527 VPWR.n737 VGND 0.002984f
C4528 VPWR.n738 VGND 0.001225f
C4529 VPWR.n739 VGND 8.78e-19
C4530 VPWR.n740 VGND 0.001281f
C4531 VPWR.n741 VGND 8.2e-19
C4532 VPWR.n742 VGND 0.001463f
C4533 VPWR.n743 VGND 6.56e-19
C4534 VPWR.n744 VGND 8.2e-19
C4535 VPWR.n745 VGND 0.002447f
C4536 VPWR.t318 VGND 0.001145f
C4537 VPWR.t672 VGND 0.002279f
C4538 VPWR.n746 VGND 0.00177f
C4539 VPWR.n747 VGND 8.51e-19
C4540 VPWR.n748 VGND 0.001224f
C4541 VPWR.n749 VGND 6.25e-19
C4542 VPWR.n750 VGND 3.83e-19
C4543 VPWR.n751 VGND 0.002317f
C4544 VPWR.t74 VGND 4.79e-19
C4545 VPWR.t230 VGND 4.79e-19
C4546 VPWR.n752 VGND 9.86e-19
C4547 VPWR.n753 VGND 0.001643f
C4548 VPWR.n754 VGND 0.001436f
C4549 VPWR.t848 VGND 0.030181f
C4550 VPWR.t704 VGND 0.002929f
C4551 VPWR.n755 VGND 0.004943f
C4552 VPWR.n756 VGND 0.013997f
C4553 VPWR.t429 VGND 0.002071f
C4554 VPWR.n757 VGND 0.004756f
C4555 VPWR.n758 VGND 0.002447f
C4556 VPWR.t896 VGND 0.012177f
C4557 VPWR.n759 VGND 0.008359f
C4558 VPWR.n760 VGND 3.06e-19
C4559 VPWR.n761 VGND 8.2e-19
C4560 VPWR.n762 VGND 0.001463f
C4561 VPWR.n763 VGND 6.56e-19
C4562 VPWR.n764 VGND 6.12e-19
C4563 VPWR.n765 VGND 8.51e-19
C4564 VPWR.n766 VGND 8.78e-19
C4565 VPWR.t430 VGND 0.002071f
C4566 VPWR.t641 VGND 0.002279f
C4567 VPWR.n767 VGND 0.004985f
C4568 VPWR.n768 VGND 0.003046f
C4569 VPWR.t535 VGND 0.002088f
C4570 VPWR.t885 VGND 0.004432f
C4571 VPWR.n770 VGND 0.011362f
C4572 VPWR.t536 VGND 0.002088f
C4573 VPWR.n771 VGND 0.006189f
C4574 VPWR.t632 VGND 0.002088f
C4575 VPWR.t831 VGND 0.004432f
C4576 VPWR.n773 VGND 0.011362f
C4577 VPWR.t633 VGND 0.002088f
C4578 VPWR.n774 VGND 0.006189f
C4579 VPWR.n775 VGND 8.2e-19
C4580 VPWR.n776 VGND 0.001414f
C4581 VPWR.n777 VGND 0.001281f
C4582 VPWR.n778 VGND 0.001199f
C4583 VPWR.n779 VGND 5.72e-19
C4584 VPWR.n780 VGND 0.005216f
C4585 VPWR.n781 VGND 8.51e-19
C4586 VPWR.n782 VGND 0.001224f
C4587 VPWR.n783 VGND 8.2e-19
C4588 VPWR.n784 VGND 6.56e-19
C4589 VPWR.n785 VGND 0.001463f
C4590 VPWR.n786 VGND 0.001414f
C4591 VPWR.n787 VGND 0.001281f
C4592 VPWR.n788 VGND 0.001225f
C4593 VPWR.n789 VGND 0.002367f
C4594 VPWR.n790 VGND 0.002447f
C4595 VPWR.n791 VGND 0.008641f
C4596 VPWR.n792 VGND 0.008641f
C4597 VPWR.n793 VGND 0.018675f
C4598 VPWR.n794 VGND 0.002447f
C4599 VPWR.n795 VGND 0.001835f
C4600 VPWR.n796 VGND 0.00372f
C4601 VPWR.n797 VGND 0.002939f
C4602 VPWR.n798 VGND 0.002263f
C4603 VPWR.n799 VGND 0.002447f
C4604 VPWR.n800 VGND 0.001835f
C4605 VPWR.n801 VGND 0.00145f
C4606 VPWR.n802 VGND 0.003051f
C4607 VPWR.n803 VGND 0.003342f
C4608 VPWR.n804 VGND 0.001475f
C4609 VPWR.t640 VGND 0.002279f
C4610 VPWR.n805 VGND 0.00177f
C4611 VPWR.n806 VGND 0.001157f
C4612 VPWR.n807 VGND 0.001995f
C4613 VPWR.n808 VGND 9.99e-19
C4614 VPWR.n809 VGND 0.001281f
C4615 VPWR.n810 VGND 0.001414f
C4616 VPWR.n811 VGND 0.001414f
C4617 VPWR.n812 VGND 0.048231f
C4618 VPWR.n813 VGND 0.001463f
C4619 VPWR.n814 VGND 0.001225f
C4620 VPWR.n815 VGND 6.56e-19
C4621 VPWR.n816 VGND 8.51e-19
C4622 VPWR.n817 VGND 8.51e-19
C4623 VPWR.n818 VGND 0.001281f
C4624 VPWR.n819 VGND 0.001225f
C4625 VPWR.n820 VGND 6.64e-19
C4626 VPWR.t826 VGND 5.61e-19
C4627 VPWR.t801 VGND 0.001157f
C4628 VPWR.n821 VGND 0.002356f
C4629 VPWR.n822 VGND 0.001831f
C4630 VPWR.n823 VGND 0.002447f
C4631 VPWR.t23 VGND 0.001154f
C4632 VPWR.t822 VGND 4.79e-19
C4633 VPWR.t178 VGND 4.79e-19
C4634 VPWR.n824 VGND 9.97e-19
C4635 VPWR.n825 VGND 0.002877f
C4636 VPWR.t730 VGND 0.001154f
C4637 VPWR.t523 VGND 0.002071f
C4638 VPWR.n826 VGND 0.003648f
C4639 VPWR.n827 VGND 0.00145f
C4640 VPWR.t871 VGND 0.012177f
C4641 VPWR.t285 VGND 4.79e-19
C4642 VPWR.t132 VGND 4.79e-19
C4643 VPWR.n828 VGND 9.86e-19
C4644 VPWR.n829 VGND 0.006214f
C4645 VPWR.n830 VGND 3.06e-19
C4646 VPWR.n831 VGND 8.2e-19
C4647 VPWR.n832 VGND 0.044685f
C4648 VPWR.n833 VGND 0.117032f
C4649 VPWR.n834 VGND 0.040161f
C4650 VPWR.n835 VGND 6.56e-19
C4651 VPWR.n836 VGND 0.001269f
C4652 VPWR.n837 VGND 0.113162f
C4653 VPWR.n838 VGND 0.001269f
C4654 VPWR.n839 VGND 8.2e-19
C4655 VPWR.n840 VGND 8.51e-19
C4656 VPWR.n841 VGND 2.28e-19
C4657 VPWR.t710 VGND 0.001255f
C4658 VPWR.n842 VGND 0.002561f
C4659 VPWR.n843 VGND 9.31e-19
C4660 VPWR.t395 VGND 0.021641f
C4661 VPWR.t137 VGND 0.011997f
C4662 VPWR.t133 VGND 0.009331f
C4663 VPWR.t516 VGND 0.012153f
C4664 VPWR.t181 VGND 0.014271f
C4665 VPWR.t95 VGND 0.009331f
C4666 VPWR.t673 VGND 0.012153f
C4667 VPWR.t398 VGND 0.013094f
C4668 VPWR.t278 VGND 0.013957f
C4669 VPWR.t37 VGND 0.009488f
C4670 VPWR.t28 VGND 0.017093f
C4671 VPWR.t319 VGND 0.0069f
C4672 VPWR.t705 VGND 0.004391f
C4673 VPWR.t8 VGND 0.007214f
C4674 VPWR.t233 VGND 0.022974f
C4675 VPWR.t186 VGND 0.025013f
C4676 VPWR.t539 VGND 0.008468f
C4677 VPWR.t692 VGND 0.011448f
C4678 VPWR.t707 VGND 0.01184f
C4679 VPWR.n844 VGND 0.015857f
C4680 VPWR.t540 VGND 0.002071f
C4681 VPWR.n845 VGND 0.003648f
C4682 VPWR.t708 VGND 0.001255f
C4683 VPWR.t861 VGND 0.015325f
C4684 VPWR.n846 VGND 0.004957f
C4685 VPWR.n847 VGND 0.001835f
C4686 VPWR.t187 VGND 2.34e-19
C4687 VPWR.t693 VGND 6.29e-19
C4688 VPWR.n848 VGND 0.002869f
C4689 VPWR.n849 VGND 0.005804f
C4690 VPWR.t234 VGND 0.003122f
C4691 VPWR.n850 VGND 0.007007f
C4692 VPWR.t541 VGND 0.002071f
C4693 VPWR.n851 VGND 0.002007f
C4694 VPWR.t706 VGND 6.35e-19
C4695 VPWR.t29 VGND 6.35e-19
C4696 VPWR.n852 VGND 0.00138f
C4697 VPWR.n853 VGND 0.003248f
C4698 VPWR.n854 VGND 8.51e-19
C4699 VPWR.n855 VGND 8.2e-19
C4700 VPWR.n856 VGND 6.56e-19
C4701 VPWR.n857 VGND 0.177644f
C4702 VPWR.n858 VGND 0.001269f
C4703 VPWR.n859 VGND 6.12e-19
C4704 VPWR.t320 VGND 0.003047f
C4705 VPWR.n860 VGND 0.002247f
C4706 VPWR.n861 VGND 7.21e-19
C4707 VPWR.t399 VGND 0.002071f
C4708 VPWR.n862 VGND 0.003648f
C4709 VPWR.n863 VGND 8.2e-19
C4710 VPWR.n864 VGND 6.12e-19
C4711 VPWR.t912 VGND 0.012177f
C4712 VPWR.t674 VGND 0.002088f
C4713 VPWR.t918 VGND 0.004432f
C4714 VPWR.n866 VGND 0.011362f
C4715 VPWR.t675 VGND 0.002088f
C4716 VPWR.n867 VGND 0.005619f
C4717 VPWR.n868 VGND 0.008401f
C4718 VPWR.t517 VGND 0.002086f
C4719 VPWR.n869 VGND 9.69e-19
C4720 VPWR.t865 VGND 0.015742f
C4721 VPWR.n870 VGND 0.026863f
C4722 VPWR.n871 VGND 0.008305f
C4723 VPWR.t134 VGND 6.35e-19
C4724 VPWR.t138 VGND 6.35e-19
C4725 VPWR.n872 VGND 0.00138f
C4726 VPWR.n873 VGND 0.008883f
C4727 VPWR.n874 VGND 3.06e-19
C4728 VPWR.n875 VGND 8.2e-19
C4729 VPWR.n876 VGND 0.001269f
C4730 VPWR.n877 VGND 6.56e-19
C4731 VPWR.n878 VGND 6.12e-19
C4732 VPWR.n879 VGND 8.51e-19
C4733 VPWR.n880 VGND 8.2e-19
C4734 VPWR.n881 VGND 8.78e-19
C4735 VPWR.t518 VGND 0.002071f
C4736 VPWR.n882 VGND 0.003648f
C4737 VPWR.n883 VGND 0.002273f
C4738 VPWR.t396 VGND 0.002088f
C4739 VPWR.t907 VGND 0.004432f
C4740 VPWR.n885 VGND 0.011362f
C4741 VPWR.t397 VGND 0.002088f
C4742 VPWR.n886 VGND 0.006189f
C4743 VPWR.t505 VGND 0.002088f
C4744 VPWR.t879 VGND 0.004432f
C4745 VPWR.n888 VGND 0.011362f
C4746 VPWR.t506 VGND 0.002088f
C4747 VPWR.n889 VGND 0.006189f
C4748 VPWR.n890 VGND 0.001199f
C4749 VPWR.n891 VGND 5.72e-19
C4750 VPWR.n892 VGND 0.005217f
C4751 VPWR.n893 VGND 8.51e-19
C4752 VPWR.n894 VGND 0.001224f
C4753 VPWR.n895 VGND 8.2e-19
C4754 VPWR.n896 VGND 6.56e-19
C4755 VPWR.n897 VGND 0.100438f
C4756 VPWR.n898 VGND 0.001269f
C4757 VPWR.n899 VGND 0.001225f
C4758 VPWR.n900 VGND 0.002141f
C4759 VPWR.n901 VGND 8.38e-19
C4760 VPWR.n902 VGND 0.006423f
C4761 VPWR.n903 VGND 0.005271f
C4762 VPWR.n904 VGND 9.31e-19
C4763 VPWR.n905 VGND 0.002292f
C4764 VPWR.t96 VGND 6.35e-19
C4765 VPWR.t182 VGND 6.35e-19
C4766 VPWR.n906 VGND 0.001389f
C4767 VPWR.n907 VGND 0.008207f
C4768 VPWR.n908 VGND 8.38e-19
C4769 VPWR.n909 VGND 8.38e-19
C4770 VPWR.n910 VGND 0.001974f
C4771 VPWR.t400 VGND 0.002104f
C4772 VPWR.n911 VGND 0.003119f
C4773 VPWR.n912 VGND 0.00786f
C4774 VPWR.n913 VGND 0.00145f
C4775 VPWR.n914 VGND 0.002447f
C4776 VPWR.n915 VGND 0.001835f
C4777 VPWR.n916 VGND 0.006423f
C4778 VPWR.n917 VGND 0.016529f
C4779 VPWR.n918 VGND 9.97e-19
C4780 VPWR.n919 VGND 0.001225f
C4781 VPWR.n920 VGND 8.51e-19
C4782 VPWR.n921 VGND 0.001176f
C4783 VPWR.t38 VGND 5.7e-19
C4784 VPWR.t279 VGND 9.42e-19
C4785 VPWR.n922 VGND 0.002604f
C4786 VPWR.n923 VGND 0.003375f
C4787 VPWR.n924 VGND 6.65e-19
C4788 VPWR.n925 VGND 3.46e-19
C4789 VPWR.n926 VGND 6.12e-19
C4790 VPWR.n927 VGND 8.2e-19
C4791 VPWR.n928 VGND 6.56e-19
C4792 VPWR.n929 VGND 0.117032f
C4793 VPWR.n930 VGND 0.040161f
C4794 VPWR.n931 VGND 0.02498f
C4795 VPWR.n932 VGND 0.091099f
C4796 VPWR.n933 VGND 0.177799f
C4797 VPWR.n934 VGND 6.56e-19
C4798 VPWR.n935 VGND 0.001269f
C4799 VPWR.n936 VGND 0.001269f
C4800 VPWR.n937 VGND 6.56e-19
C4801 VPWR.n938 VGND 0.048231f
C4802 VPWR.n939 VGND 0.058067f
C4803 VPWR.n940 VGND 0.048231f
C4804 VPWR.n941 VGND 6.56e-19
C4805 VPWR.n942 VGND 0.001269f
C4806 VPWR.n943 VGND 0.001269f
C4807 VPWR.n944 VGND 8.2e-19
C4808 VPWR.n945 VGND 0.001225f
C4809 VPWR.t816 VGND 6.35e-19
C4810 VPWR.t118 VGND 6.35e-19
C4811 VPWR.n946 VGND 0.00138f
C4812 VPWR.t70 VGND 0.001631f
C4813 VPWR.t720 VGND 0.001191f
C4814 VPWR.n947 VGND 0.004218f
C4815 VPWR.n948 VGND 0.002454f
C4816 VPWR.n949 VGND 0.002221f
C4817 VPWR.t274 VGND 0.001139f
C4818 VPWR.t933 VGND 0.012177f
C4819 VPWR.n950 VGND 0.016529f
C4820 VPWR.t299 VGND 9.14e-19
C4821 VPWR.t84 VGND 9.14e-19
C4822 VPWR.n951 VGND 0.001864f
C4823 VPWR.n952 VGND 0.002706f
C4824 VPWR.t728 VGND 6.35e-19
C4825 VPWR.t354 VGND 6.35e-19
C4826 VPWR.n953 VGND 0.00141f
C4827 VPWR.t795 VGND 9.42e-19
C4828 VPWR.t68 VGND 9.7e-19
C4829 VPWR.n954 VGND 0.002279f
C4830 VPWR.n955 VGND 8.38e-19
C4831 VPWR.t495 VGND 0.002071f
C4832 VPWR.n956 VGND 0.003648f
C4833 VPWR.n957 VGND 0.00125f
C4834 VPWR.t882 VGND 0.008643f
C4835 VPWR.t340 VGND 0.002626f
C4836 VPWR.n958 VGND 0.002545f
C4837 VPWR.n959 VGND 6.12e-19
C4838 VPWR.n960 VGND 8.8e-19
C4839 VPWR.n961 VGND 6.56e-19
C4840 VPWR.n962 VGND 8.2e-19
C4841 VPWR.n963 VGND 6.56e-19
C4842 VPWR.n964 VGND 0.001092f
C4843 VPWR.t104 VGND 7.48e-19
C4844 VPWR.t102 VGND 7.48e-19
C4845 VPWR.n965 VGND 0.001639f
C4846 VPWR.n966 VGND 0.001463f
C4847 VPWR.t694 VGND 6.35e-19
C4848 VPWR.t106 VGND 6.35e-19
C4849 VPWR.n967 VGND 0.00141f
C4850 VPWR.n968 VGND 7.11e-19
C4851 VPWR.n969 VGND 0.001835f
C4852 VPWR.t276 VGND 6.35e-19
C4853 VPWR.t35 VGND 6.35e-19
C4854 VPWR.n970 VGND 0.00141f
C4855 VPWR.t529 VGND 0.002088f
C4856 VPWR.t860 VGND 0.004432f
C4857 VPWR.n972 VGND 0.011362f
C4858 VPWR.t530 VGND 0.002088f
C4859 VPWR.n973 VGND 0.006189f
C4860 VPWR.n974 VGND 0.001597f
C4861 VPWR.t630 VGND 0.002088f
C4862 VPWR.t839 VGND 0.004432f
C4863 VPWR.n976 VGND 0.011362f
C4864 VPWR.t631 VGND 0.002088f
C4865 VPWR.n977 VGND 0.006189f
C4866 VPWR.n978 VGND 0.005236f
C4867 VPWR.n979 VGND 3.77e-19
C4868 VPWR.n980 VGND 0.003736f
C4869 VPWR.n981 VGND 0.001556f
C4870 VPWR.n982 VGND 8.38e-19
C4871 VPWR.n983 VGND 0.001835f
C4872 VPWR.n984 VGND 7.11e-19
C4873 VPWR.n985 VGND 0.005275f
C4874 VPWR.n986 VGND 5.94e-19
C4875 VPWR.n987 VGND 3.59e-19
C4876 VPWR.n988 VGND 9.84e-19
C4877 VPWR.n989 VGND 8.2e-19
C4878 VPWR.n990 VGND 0.001269f
C4879 VPWR.n991 VGND 0.053551f
C4880 VPWR.n992 VGND 0.001414f
C4881 VPWR.n993 VGND 0.001463f
C4882 VPWR.n994 VGND 0.001092f
C4883 VPWR.n995 VGND 6.56e-19
C4884 VPWR.n996 VGND 0.001224f
C4885 VPWR.t578 VGND 0.002071f
C4886 VPWR.t872 VGND 0.00872f
C4887 VPWR.n998 VGND 0.015149f
C4888 VPWR.t579 VGND 0.002071f
C4889 VPWR.n999 VGND 0.008692f
C4890 VPWR.t668 VGND 0.002071f
C4891 VPWR.t930 VGND 0.00872f
C4892 VPWR.n1001 VGND 0.015149f
C4893 VPWR.t669 VGND 0.002071f
C4894 VPWR.n1002 VGND 0.008692f
C4895 VPWR.n1003 VGND 0.00749f
C4896 VPWR.t435 VGND 0.002088f
C4897 VPWR.t919 VGND 0.004432f
C4898 VPWR.n1005 VGND 0.011362f
C4899 VPWR.t436 VGND 0.002088f
C4900 VPWR.n1006 VGND 0.006189f
C4901 VPWR.t537 VGND 0.002088f
C4902 VPWR.t864 VGND 0.004432f
C4903 VPWR.n1008 VGND 0.011362f
C4904 VPWR.t538 VGND 0.002088f
C4905 VPWR.n1009 VGND 0.006189f
C4906 VPWR.n1010 VGND 0.005099f
C4907 VPWR.n1011 VGND 0.001597f
C4908 VPWR.n1012 VGND 0.002868f
C4909 VPWR.n1013 VGND 8.51e-19
C4910 VPWR.n1014 VGND 7.3e-19
C4911 VPWR.t240 VGND 7.48e-19
C4912 VPWR.t740 VGND 7.48e-19
C4913 VPWR.n1015 VGND 0.001676f
C4914 VPWR.t58 VGND 7.48e-19
C4915 VPWR.t112 VGND 7.48e-19
C4916 VPWR.n1016 VGND 0.001676f
C4917 VPWR.t239 VGND 0.001178f
C4918 VPWR.t60 VGND 0.001178f
C4919 VPWR.n1017 VGND 0.004766f
C4920 VPWR.n1018 VGND 0.002447f
C4921 VPWR.n1019 VGND 6.36e-19
C4922 VPWR.n1020 VGND 0.002447f
C4923 VPWR.t54 VGND 5.61e-19
C4924 VPWR.t719 VGND 0.001157f
C4925 VPWR.n1021 VGND 0.002356f
C4926 VPWR.t752 VGND 5.61e-19
C4927 VPWR.t712 VGND 0.001157f
C4928 VPWR.n1022 VGND 0.002356f
C4929 VPWR.n1023 VGND 0.003228f
C4930 VPWR.n1024 VGND 7.77e-19
C4931 VPWR.n1025 VGND 0.002447f
C4932 VPWR.t144 VGND 0.001154f
C4933 VPWR.t721 VGND 0.001154f
C4934 VPWR.t185 VGND 4.79e-19
C4935 VPWR.t94 VGND 4.79e-19
C4936 VPWR.n1026 VGND 9.97e-19
C4937 VPWR.n1027 VGND 0.001888f
C4938 VPWR.t2 VGND 4.79e-19
C4939 VPWR.t130 VGND 4.79e-19
C4940 VPWR.n1028 VGND 9.97e-19
C4941 VPWR.t432 VGND 0.002088f
C4942 VPWR.t920 VGND 0.004432f
C4943 VPWR.n1030 VGND 0.011362f
C4944 VPWR.t433 VGND 0.002088f
C4945 VPWR.n1031 VGND 0.006189f
C4946 VPWR.t779 VGND 7.48e-19
C4947 VPWR.t702 VGND 7.48e-19
C4948 VPWR.n1032 VGND 0.001682f
C4949 VPWR.n1033 VGND 0.005999f
C4950 VPWR.n1034 VGND 0.001225f
C4951 VPWR.n1035 VGND 0.001281f
C4952 VPWR.n1036 VGND 8.2e-19
C4953 VPWR.n1037 VGND 0.001463f
C4954 VPWR.n1038 VGND 0.053551f
C4955 VPWR.n1039 VGND 6.56e-19
C4956 VPWR.n1040 VGND 8.2e-19
C4957 VPWR.n1041 VGND 6.12e-19
C4958 VPWR.n1042 VGND 8.51e-19
C4959 VPWR.n1043 VGND 0.001224f
C4960 VPWR.n1044 VGND 8.51e-19
C4961 VPWR.t781 VGND 0.001168f
C4962 VPWR.n1045 VGND 0.002245f
C4963 VPWR.t434 VGND 0.031129f
C4964 VPWR.t577 VGND 0.037401f
C4965 VPWR.t57 VGND 0.017015f
C4966 VPWR.t111 VGND 0.023052f
C4967 VPWR.t59 VGND 0.025405f
C4968 VPWR.t142 VGND 0.015525f
C4969 VPWR.t3 VGND 0.014035f
C4970 VPWR.t53 VGND 0.017799f
C4971 VPWR.t711 VGND 0.018426f
C4972 VPWR.t0 VGND 0.015525f
C4973 VPWR.t141 VGND 0.014114f
C4974 VPWR.t143 VGND 0.021406f
C4975 VPWR.t1 VGND 0.021327f
C4976 VPWR.t93 VGND 0.01035f
C4977 VPWR.t778 VGND 0.013094f
C4978 VPWR.t431 VGND 0.006586f
C4979 VPWR.t701 VGND 0.008547f
C4980 VPWR.n1046 VGND 0.002273f
C4981 VPWR.n1047 VGND 8.51e-19
C4982 VPWR.n1048 VGND 8.2e-19
C4983 VPWR.n1049 VGND 0.001463f
C4984 VPWR.n1050 VGND 6.56e-19
C4985 VPWR.n1051 VGND 8.51e-19
C4986 VPWR.n1052 VGND 0.001224f
C4987 VPWR.t910 VGND 0.008643f
C4988 VPWR.t301 VGND 6.29e-19
C4989 VPWR.t5 VGND 2.34e-19
C4990 VPWR.n1053 VGND 0.002869f
C4991 VPWR.n1054 VGND 6.7e-19
C4992 VPWR.n1055 VGND 0.003264f
C4993 VPWR.t305 VGND 9.7e-19
C4994 VPWR.t166 VGND 9.42e-19
C4995 VPWR.n1056 VGND 0.002247f
C4996 VPWR.t328 VGND 9.14e-19
C4997 VPWR.t148 VGND 9.14e-19
C4998 VPWR.n1057 VGND 0.001864f
C4999 VPWR.n1058 VGND 0.002447f
C5000 VPWR.t696 VGND 4.65e-19
C5001 VPWR.t42 VGND -4.89e-19
C5002 VPWR.n1059 VGND 0.003109f
C5003 VPWR.n1060 VGND 7.16e-19
C5004 VPWR.n1061 VGND 0.002447f
C5005 VPWR.t818 VGND 4.65e-19
C5006 VPWR.t193 VGND -4.89e-19
C5007 VPWR.n1062 VGND 0.003109f
C5008 VPWR.t334 VGND 4.79e-19
C5009 VPWR.t86 VGND 4.79e-19
C5010 VPWR.n1063 VGND 9.97e-19
C5011 VPWR.t174 VGND 0.001149f
C5012 VPWR.n1064 VGND 0.002221f
C5013 VPWR.n1065 VGND 6.25e-19
C5014 VPWR.t162 VGND 3.14e-19
C5015 VPWR.t347 VGND 3.14e-19
C5016 VPWR.n1066 VGND 7.27e-19
C5017 VPWR.t46 VGND 4.79e-19
C5018 VPWR.t129 VGND 4.79e-19
C5019 VPWR.n1067 VGND 9.97e-19
C5020 VPWR.n1068 VGND 0.002967f
C5021 VPWR.n1069 VGND 8.78e-19
C5022 VPWR.n1070 VGND 8.2e-19
C5023 VPWR.n1071 VGND 0.001463f
C5024 VPWR.n1072 VGND 0.001414f
C5025 VPWR.n1073 VGND 0.001463f
C5026 VPWR.n1074 VGND 0.001225f
C5027 VPWR.n1075 VGND 6.56e-19
C5028 VPWR.n1076 VGND 8.51e-19
C5029 VPWR.n1077 VGND 0.001197f
C5030 VPWR.t372 VGND 7.76e-19
C5031 VPWR.t376 VGND 7.76e-19
C5032 VPWR.n1078 VGND 0.001602f
C5033 VPWR.n1079 VGND 0.003594f
C5034 VPWR.t380 VGND 7.76e-19
C5035 VPWR.t384 VGND 7.76e-19
C5036 VPWR.n1080 VGND 0.001602f
C5037 VPWR.n1081 VGND 0.003594f
C5038 VPWR.n1082 VGND 8.78e-19
C5039 VPWR.n1083 VGND 0.002447f
C5040 VPWR.t356 VGND 7.76e-19
C5041 VPWR.t360 VGND 7.48e-19
C5042 VPWR.n1084 VGND 0.001574f
C5043 VPWR.n1085 VGND 0.001775f
C5044 VPWR.t364 VGND 7.76e-19
C5045 VPWR.t368 VGND 7.76e-19
C5046 VPWR.n1086 VGND 0.001601f
C5047 VPWR.n1087 VGND 0.003372f
C5048 VPWR.t406 VGND 0.002279f
C5049 VPWR.n1088 VGND 0.001563f
C5050 VPWR.t358 VGND 7.76e-19
C5051 VPWR.t362 VGND 7.76e-19
C5052 VPWR.n1089 VGND 0.001601f
C5053 VPWR.n1090 VGND 0.00202f
C5054 VPWR.n1091 VGND 0.002447f
C5055 VPWR.t677 VGND 0.002279f
C5056 VPWR.n1092 VGND 0.001766f
C5057 VPWR.t366 VGND 7.76e-19
C5058 VPWR.t370 VGND 7.76e-19
C5059 VPWR.n1093 VGND 0.001602f
C5060 VPWR.t833 VGND 0.030181f
C5061 VPWR.n1094 VGND 0.013829f
C5062 VPWR.t374 VGND 0.002725f
C5063 VPWR.n1095 VGND 0.003161f
C5064 VPWR.n1096 VGND 0.00372f
C5065 VPWR.n1097 VGND 9.31e-19
C5066 VPWR.n1098 VGND 8.2e-19
C5067 VPWR.n1099 VGND 6.56e-19
C5068 VPWR.n1100 VGND 6.56e-19
C5069 VPWR.n1101 VGND 8.2e-19
C5070 VPWR.n1102 VGND 8.51e-19
C5071 VPWR.t554 VGND 0.027522f
C5072 VPWR.t525 VGND 0.023052f
C5073 VPWR.t587 VGND 0.038342f
C5074 VPWR.t663 VGND 0.026581f
C5075 VPWR.t557 VGND 0.045556f
C5076 VPWR.t551 VGND 0.041008f
C5077 VPWR.n1103 VGND 0.002501f
C5078 VPWR.n1104 VGND 0.002598f
C5079 VPWR.n1105 VGND 8.51e-19
C5080 VPWR.n1106 VGND 8.2e-19
C5081 VPWR.n1107 VGND 0.001463f
C5082 VPWR.n1108 VGND 0.081008f
C5083 VPWR.n1109 VGND 0.221149f
C5084 VPWR.n1110 VGND 0.048231f
C5085 VPWR.n1111 VGND 0.001463f
C5086 VPWR.n1112 VGND 0.001225f
C5087 VPWR.n1113 VGND 6.56e-19
C5088 VPWR.n1114 VGND 8.51e-19
C5089 VPWR.n1115 VGND 0.001224f
C5090 VPWR.t851 VGND 0.030181f
C5091 VPWR.n1116 VGND 0.015206f
C5092 VPWR.n1117 VGND 0.002447f
C5093 VPWR.t873 VGND 0.030181f
C5094 VPWR.n1118 VGND 0.015033f
C5095 VPWR.t665 VGND 0.002279f
C5096 VPWR.n1119 VGND 0.002879f
C5097 VPWR.n1120 VGND 0.001835f
C5098 VPWR.t589 VGND 0.002071f
C5099 VPWR.n1121 VGND 0.004756f
C5100 VPWR.n1122 VGND 0.002447f
C5101 VPWR.n1123 VGND 0.00634f
C5102 VPWR.n1124 VGND 0.001197f
C5103 VPWR.n1125 VGND 8.2e-19
C5104 VPWR.n1126 VGND 0.001463f
C5105 VPWR.n1127 VGND 6.56e-19
C5106 VPWR.n1128 VGND 9.84e-19
C5107 VPWR.t859 VGND 0.015325f
C5108 VPWR.t588 VGND 0.002071f
C5109 VPWR.n1129 VGND 0.004756f
C5110 VPWR.t527 VGND 0.00212f
C5111 VPWR.n1130 VGND 8.89e-19
C5112 VPWR.n1131 VGND 0.004844f
C5113 VPWR.t881 VGND 0.004446f
C5114 VPWR.n1132 VGND 0.00855f
C5115 VPWR.t526 VGND 0.002088f
C5116 VPWR.n1133 VGND 0.003022f
C5117 VPWR.n1134 VGND 0.002979f
C5118 VPWR.t555 VGND 0.002088f
C5119 VPWR.t874 VGND 0.004432f
C5120 VPWR.n1136 VGND 0.011362f
C5121 VPWR.t556 VGND 0.002088f
C5122 VPWR.n1137 VGND 0.006189f
C5123 VPWR.t666 VGND 0.002088f
C5124 VPWR.t924 VGND 0.004432f
C5125 VPWR.n1139 VGND 0.011362f
C5126 VPWR.t667 VGND 0.002088f
C5127 VPWR.n1140 VGND 0.006189f
C5128 VPWR.n1141 VGND 0.005099f
C5129 VPWR.n1142 VGND 0.001597f
C5130 VPWR.n1143 VGND 0.001464f
C5131 VPWR.n1144 VGND 8.38e-19
C5132 VPWR.n1145 VGND 0.001148f
C5133 VPWR.t664 VGND 0.002287f
C5134 VPWR.n1146 VGND 0.002536f
C5135 VPWR.n1147 VGND 0.003124f
C5136 VPWR.n1148 VGND 0.001835f
C5137 VPWR.n1149 VGND 8.2e-19
C5138 VPWR.n1150 VGND 0.001414f
C5139 VPWR.n1151 VGND 0.001281f
C5140 VPWR.n1152 VGND 0.001092f
C5141 VPWR.n1153 VGND 0.001463f
C5142 VPWR.n1154 VGND 0.006293f
C5143 VPWR.n1155 VGND 0.021777f
C5144 VPWR.t925 VGND 0.030181f
C5145 VPWR.n1156 VGND 0.016876f
C5146 VPWR.n1157 VGND 0.004367f
C5147 VPWR.n1158 VGND 8.51e-19
C5148 VPWR.n1159 VGND 8.51e-19
C5149 VPWR.n1160 VGND 0.001224f
C5150 VPWR.n1161 VGND 8.2e-19
C5151 VPWR.n1162 VGND 6.56e-19
C5152 VPWR.n1163 VGND 0.001463f
C5153 VPWR.n1164 VGND 0.001414f
C5154 VPWR.n1165 VGND 0.001281f
C5155 VPWR.n1166 VGND 8.8e-19
C5156 VPWR.n1167 VGND 0.00125f
C5157 VPWR.n1168 VGND 0.008641f
C5158 VPWR.n1169 VGND 0.008641f
C5159 VPWR.n1170 VGND 0.008359f
C5160 VPWR.n1171 VGND 0.002447f
C5161 VPWR.n1172 VGND 0.00145f
C5162 VPWR.n1173 VGND 0.003633f
C5163 VPWR.n1174 VGND 0.002332f
C5164 VPWR.t558 VGND 0.002279f
C5165 VPWR.n1175 VGND 0.002879f
C5166 VPWR.n1176 VGND 0.004956f
C5167 VPWR.n1177 VGND 0.002447f
C5168 VPWR.n1178 VGND 0.00145f
C5169 VPWR.n1179 VGND 0.002412f
C5170 VPWR.t552 VGND 0.002279f
C5171 VPWR.n1180 VGND 0.00164f
C5172 VPWR.n1181 VGND 0.002392f
C5173 VPWR.n1182 VGND 0.002221f
C5174 VPWR.n1183 VGND 0.002447f
C5175 VPWR.n1184 VGND 0.00389f
C5176 VPWR.n1185 VGND 0.005302f
C5177 VPWR.n1186 VGND 0.004063f
C5178 VPWR.n1187 VGND 0.002447f
C5179 VPWR.n1188 VGND 0.001888f
C5180 VPWR.n1189 VGND 0.00389f
C5181 VPWR.n1190 VGND 0.005302f
C5182 VPWR.t559 VGND 0.002279f
C5183 VPWR.n1191 VGND 0.002879f
C5184 VPWR.n1192 VGND 0.005129f
C5185 VPWR.n1193 VGND 0.005302f
C5186 VPWR.n1194 VGND 8.51e-19
C5187 VPWR.n1195 VGND 6.56e-19
C5188 VPWR.n1196 VGND 8.2e-19
C5189 VPWR.n1197 VGND 9.31e-19
C5190 VPWR.n1198 VGND 0.001144f
C5191 VPWR.n1199 VGND 8.2e-19
C5192 VPWR.n1200 VGND 0.001281f
C5193 VPWR.n1201 VGND 0.001414f
C5194 VPWR.n1202 VGND 0.058516f
C5195 VPWR.n1203 VGND 0.001414f
C5196 VPWR.n1204 VGND 0.001281f
C5197 VPWR.n1205 VGND 0.001225f
C5198 VPWR.n1206 VGND 0.001051f
C5199 VPWR.n1207 VGND 0.002425f
C5200 VPWR.t889 VGND 0.008576f
C5201 VPWR.t72 VGND 0.002867f
C5202 VPWR.n1208 VGND 0.00593f
C5203 VPWR.n1209 VGND 0.00145f
C5204 VPWR.t322 VGND 7.76e-19
C5205 VPWR.t15 VGND 7.76e-19
C5206 VPWR.n1210 VGND 0.001667f
C5207 VPWR.t405 VGND 0.002279f
C5208 VPWR.n1211 VGND 0.001468f
C5209 VPWR.n1212 VGND 0.002447f
C5210 VPWR.t751 VGND 7.76e-19
C5211 VPWR.t386 VGND 7.76e-19
C5212 VPWR.n1213 VGND 0.001663f
C5213 VPWR.n1214 VGND 0.003631f
C5214 VPWR.t378 VGND 7.76e-19
C5215 VPWR.t382 VGND 7.76e-19
C5216 VPWR.n1215 VGND 0.001602f
C5217 VPWR.t928 VGND 0.030181f
C5218 VPWR.n1216 VGND 0.001572f
C5219 VPWR.n1217 VGND 0.01411f
C5220 VPWR.n1218 VGND 0.002314f
C5221 VPWR.n1219 VGND 0.001335f
C5222 VPWR.n1220 VGND 0.003594f
C5223 VPWR.n1221 VGND 0.002603f
C5224 VPWR.n1222 VGND 0.001859f
C5225 VPWR.n1223 VGND 0.002447f
C5226 VPWR.n1224 VGND 0.001835f
C5227 VPWR.n1225 VGND 0.001196f
C5228 VPWR.n1226 VGND 0.002407f
C5229 VPWR.t521 VGND 0.002071f
C5230 VPWR.n1227 VGND 0.005866f
C5231 VPWR.n1228 VGND 0.006109f
C5232 VPWR.n1229 VGND 0.002221f
C5233 VPWR.n1230 VGND 0.001224f
C5234 VPWR.n1231 VGND 6.98e-19
C5235 VPWR.n1232 VGND 0.002862f
C5236 VPWR.n1233 VGND 0.00426f
C5237 VPWR.n1234 VGND 0.001638f
C5238 VPWR.t520 VGND 0.002071f
C5239 VPWR.n1235 VGND 0.001104f
C5240 VPWR.t553 VGND 0.002287f
C5241 VPWR.n1236 VGND 0.002594f
C5242 VPWR.n1237 VGND 9.64e-19
C5243 VPWR.n1238 VGND 8.38e-19
C5244 VPWR.n1239 VGND 9.31e-19
C5245 VPWR.n1240 VGND 0.001317f
C5246 VPWR.n1241 VGND 0.007114f
C5247 VPWR.n1242 VGND 0.015547f
C5248 VPWR.t519 VGND 0.002509f
C5249 VPWR.t71 VGND 0.006978f
C5250 VPWR.t321 VGND 0.011918f
C5251 VPWR.t14 VGND 0.008311f
C5252 VPWR.t750 VGND 0.013486f
C5253 VPWR.t385 VGND 0.013486f
C5254 VPWR.t377 VGND 0.013486f
C5255 VPWR.t381 VGND 0.013486f
C5256 VPWR.t371 VGND 0.013486f
C5257 VPWR.t375 VGND 0.010272f
C5258 VPWR.t404 VGND 0.006743f
C5259 VPWR.t379 VGND 0.009958f
C5260 VPWR.t383 VGND 0.013486f
C5261 VPWR.t355 VGND 0.013408f
C5262 VPWR.t359 VGND 0.013408f
C5263 VPWR.t363 VGND 0.013486f
C5264 VPWR.t367 VGND 0.010899f
C5265 VPWR.t357 VGND 0.009331f
C5266 VPWR.t361 VGND 0.013486f
C5267 VPWR.t365 VGND 0.013486f
C5268 VPWR.t369 VGND 0.013486f
C5269 VPWR.t373 VGND 0.020308f
C5270 VPWR.t676 VGND 0.016858f
C5271 VPWR.t682 VGND 0.026581f
C5272 VPWR.t419 VGND 0.021641f
C5273 VPWR.t651 VGND 0.035363f
C5274 VPWR.t247 VGND 0.028855f
C5275 VPWR.t544 VGND 0.006743f
C5276 VPWR.t243 VGND 0.007841f
C5277 VPWR.t241 VGND 0.013486f
C5278 VPWR.t271 VGND 0.013486f
C5279 VPWR.t267 VGND 0.013486f
C5280 VPWR.t265 VGND 0.013486f
C5281 VPWR.t261 VGND 0.013486f
C5282 VPWR.t269 VGND 0.010742f
C5283 VPWR.t257 VGND 0.009409f
C5284 VPWR.t263 VGND 0.013486f
C5285 VPWR.t259 VGND 0.013486f
C5286 VPWR.t251 VGND 0.013486f
C5287 VPWR.t255 VGND 0.013486f
C5288 VPWR.t253 VGND 0.011369f
C5289 VPWR.t574 VGND 0.006743f
C5290 VPWR.t249 VGND 0.00886f
C5291 VPWR.t245 VGND 0.013486f
C5292 VPWR.t754 VGND 0.013486f
C5293 VPWR.t758 VGND 0.013486f
C5294 VPWR.t768 VGND 0.013486f
C5295 VPWR.t756 VGND 0.009252f
C5296 VPWR.n1243 VGND 0.015547f
C5297 VPWR.t913 VGND 0.008643f
C5298 VPWR.t683 VGND 0.002071f
C5299 VPWR.n1244 VGND 0.002596f
C5300 VPWR.n1245 VGND 0.008854f
C5301 VPWR.n1246 VGND 0.006481f
C5302 VPWR.n1247 VGND 8.51e-19
C5303 VPWR.n1248 VGND 8.2e-19
C5304 VPWR.n1249 VGND 0.001224f
C5305 VPWR.n1250 VGND 0.001224f
C5306 VPWR.n1251 VGND 8.51e-19
C5307 VPWR.n1252 VGND 0.008359f
C5308 VPWR.t684 VGND 0.002071f
C5309 VPWR.n1253 VGND 0.004756f
C5310 VPWR.n1254 VGND 0.00372f
C5311 VPWR.n1255 VGND 0.00116f
C5312 VPWR.n1256 VGND 0.002447f
C5313 VPWR.t757 VGND 0.002867f
C5314 VPWR.n1257 VGND 0.002819f
C5315 VPWR.t575 VGND 0.002279f
C5316 VPWR.n1258 VGND 0.00172f
C5317 VPWR.t769 VGND 7.76e-19
C5318 VPWR.t759 VGND 7.76e-19
C5319 VPWR.n1259 VGND 0.001667f
C5320 VPWR.t863 VGND 0.030535f
C5321 VPWR.n1260 VGND 0.012522f
C5322 VPWR.n1261 VGND 0.002447f
C5323 VPWR.t755 VGND 7.76e-19
C5324 VPWR.t246 VGND 7.76e-19
C5325 VPWR.n1262 VGND 0.001663f
C5326 VPWR.n1263 VGND 0.003526f
C5327 VPWR.t250 VGND 7.76e-19
C5328 VPWR.t254 VGND 7.76e-19
C5329 VPWR.n1264 VGND 0.001602f
C5330 VPWR.n1265 VGND 0.0024f
C5331 VPWR.t256 VGND 7.76e-19
C5332 VPWR.t252 VGND 7.76e-19
C5333 VPWR.n1266 VGND 0.001602f
C5334 VPWR.n1267 VGND 0.003594f
C5335 VPWR.t260 VGND 7.76e-19
C5336 VPWR.t264 VGND 7.76e-19
C5337 VPWR.n1268 VGND 0.001602f
C5338 VPWR.n1269 VGND 0.002366f
C5339 VPWR.n1270 VGND 0.003594f
C5340 VPWR.n1271 VGND 0.002197f
C5341 VPWR.n1272 VGND 0.002265f
C5342 VPWR.n1273 VGND 0.001942f
C5343 VPWR.n1274 VGND 0.002447f
C5344 VPWR.n1275 VGND 0.002447f
C5345 VPWR.n1276 VGND 0.002062f
C5346 VPWR.n1277 VGND 0.003594f
C5347 VPWR.n1278 VGND 0.002603f
C5348 VPWR.n1279 VGND 0.001859f
C5349 VPWR.n1280 VGND 0.002447f
C5350 VPWR.n1281 VGND 0.002447f
C5351 VPWR.n1282 VGND 0.002667f
C5352 VPWR.n1283 VGND 0.001643f
C5353 VPWR.n1284 VGND 0.003761f
C5354 VPWR.n1285 VGND 0.002883f
C5355 VPWR.n1286 VGND 0.002221f
C5356 VPWR.n1287 VGND 8.38e-19
C5357 VPWR.n1288 VGND 8.38e-19
C5358 VPWR.n1289 VGND 0.001231f
C5359 VPWR.t678 VGND 0.002279f
C5360 VPWR.n1290 VGND 0.00177f
C5361 VPWR.n1291 VGND 0.006955f
C5362 VPWR.n1292 VGND 9.31e-19
C5363 VPWR.n1293 VGND 2.28e-19
C5364 VPWR.n1294 VGND 0.001281f
C5365 VPWR.n1295 VGND 0.001414f
C5366 VPWR.n1296 VGND 0.001463f
C5367 VPWR.n1297 VGND 0.001463f
C5368 VPWR.n1298 VGND 0.001414f
C5369 VPWR.n1299 VGND 0.001281f
C5370 VPWR.n1300 VGND 0.001146f
C5371 VPWR.n1301 VGND 9.04e-19
C5372 VPWR.n1302 VGND 9.31e-19
C5373 VPWR.n1303 VGND 0.002939f
C5374 VPWR.n1304 VGND 0.00181f
C5375 VPWR.n1305 VGND 0.001835f
C5376 VPWR.n1306 VGND 0.002447f
C5377 VPWR.n1307 VGND 0.002362f
C5378 VPWR.n1308 VGND 0.001717f
C5379 VPWR.n1309 VGND 0.003554f
C5380 VPWR.n1310 VGND 0.002839f
C5381 VPWR.n1311 VGND 0.002447f
C5382 VPWR.n1312 VGND 0.002221f
C5383 VPWR.n1313 VGND 0.001139f
C5384 VPWR.n1314 VGND 0.001245f
C5385 VPWR.n1315 VGND 0.00145f
C5386 VPWR.n1316 VGND 0.002447f
C5387 VPWR.n1317 VGND 0.002447f
C5388 VPWR.n1318 VGND 0.002687f
C5389 VPWR.n1319 VGND 0.003474f
C5390 VPWR.n1320 VGND 0.001977f
C5391 VPWR.n1321 VGND 0.002468f
C5392 VPWR.n1322 VGND 0.001622f
C5393 VPWR.n1323 VGND 8.2e-19
C5394 VPWR.n1324 VGND 0.001463f
C5395 VPWR.n1325 VGND 6.56e-19
C5396 VPWR.n1326 VGND 8.2e-19
C5397 VPWR.n1327 VGND 0.001281f
C5398 VPWR.n1328 VGND 0.001225f
C5399 VPWR.n1329 VGND 8.51e-19
C5400 VPWR.n1330 VGND 0.002197f
C5401 VPWR.n1331 VGND 0.002265f
C5402 VPWR.n1332 VGND 8.51e-19
C5403 VPWR.n1333 VGND 0.001224f
C5404 VPWR.n1334 VGND 8.2e-19
C5405 VPWR.n1335 VGND 0.001281f
C5406 VPWR.n1336 VGND 0.001414f
C5407 VPWR.n1337 VGND 0.058516f
C5408 VPWR.n1338 VGND 0.048231f
C5409 VPWR.n1339 VGND 0.001414f
C5410 VPWR.n1340 VGND 0.001463f
C5411 VPWR.n1341 VGND 0.001225f
C5412 VPWR.n1342 VGND 6.56e-19
C5413 VPWR.n1343 VGND 8.51e-19
C5414 VPWR.n1344 VGND 0.001197f
C5415 VPWR.t88 VGND 4.77e-19
C5416 VPWR.t170 VGND -3.03e-19
C5417 VPWR.n1345 VGND 0.003045f
C5418 VPWR.n1346 VGND 0.002345f
C5419 VPWR.t332 VGND 0.001154f
C5420 VPWR.n1347 VGND 5.61e-19
C5421 VPWR.n1348 VGND 4.78e-19
C5422 VPWR.t210 VGND 7.76e-19
C5423 VPWR.t214 VGND 7.76e-19
C5424 VPWR.n1349 VGND 0.001602f
C5425 VPWR.n1350 VGND 4.7e-19
C5426 VPWR.n1351 VGND 8.51e-19
C5427 VPWR.n1352 VGND 8.2e-19
C5428 VPWR.n1353 VGND 0.001463f
C5429 VPWR.n1354 VGND 6.56e-19
C5430 VPWR.n1355 VGND 0.001144f
C5431 VPWR.n1356 VGND 0.001224f
C5432 VPWR.t691 VGND 4.31e-19
C5433 VPWR.t345 VGND 4.31e-19
C5434 VPWR.n1357 VGND 9.01e-19
C5435 VPWR.t208 VGND 7.76e-19
C5436 VPWR.t212 VGND 7.76e-19
C5437 VPWR.n1358 VGND 0.001602f
C5438 VPWR.n1359 VGND 5.62e-19
C5439 VPWR.n1360 VGND 0.001842f
C5440 VPWR.t224 VGND 7.76e-19
C5441 VPWR.t218 VGND 7.76e-19
C5442 VPWR.n1361 VGND 0.001613f
C5443 VPWR.n1362 VGND 0.002799f
C5444 VPWR.n1363 VGND 0.002447f
C5445 VPWR.t226 VGND 0.002739f
C5446 VPWR.n1364 VGND 0.003481f
C5447 VPWR.n1365 VGND 0.002221f
C5448 VPWR.t805 VGND 6.35e-19
C5449 VPWR.t125 VGND 6.35e-19
C5450 VPWR.n1366 VGND 0.00138f
C5451 VPWR.n1367 VGND 0.008219f
C5452 VPWR.n1368 VGND 8.2e-19
C5453 VPWR.n1369 VGND 0.001463f
C5454 VPWR.n1370 VGND 6.56e-19
C5455 VPWR.n1371 VGND 8.51e-19
C5456 VPWR.n1372 VGND 3.86e-19
C5457 VPWR.n1373 VGND 0.006661f
C5458 VPWR.t836 VGND 0.015624f
C5459 VPWR.n1374 VGND 0.028164f
C5460 VPWR.t621 VGND 0.002071f
C5461 VPWR.n1375 VGND 0.006661f
C5462 VPWR.t659 VGND 0.002088f
C5463 VPWR.t844 VGND 0.004432f
C5464 VPWR.n1377 VGND 0.011362f
C5465 VPWR.t660 VGND 0.002088f
C5466 VPWR.n1378 VGND 0.006189f
C5467 VPWR.t462 VGND 0.002088f
C5468 VPWR.t893 VGND 0.004432f
C5469 VPWR.n1380 VGND 0.011362f
C5470 VPWR.t463 VGND 0.002088f
C5471 VPWR.n1381 VGND 0.006189f
C5472 VPWR.n1382 VGND 0.005236f
C5473 VPWR.n1383 VGND 0.001597f
C5474 VPWR.n1384 VGND 9.31e-19
C5475 VPWR.n1385 VGND 5.93e-19
C5476 VPWR.n1386 VGND 0.00732f
C5477 VPWR.t562 VGND 0.002071f
C5478 VPWR.n1387 VGND 0.012535f
C5479 VPWR.t877 VGND 0.011968f
C5480 VPWR.n1388 VGND 0.008075f
C5481 VPWR.n1389 VGND 0.003462f
C5482 VPWR.t561 VGND 0.002071f
C5483 VPWR.n1390 VGND 0.001617f
C5484 VPWR.n1391 VGND 0.001699f
C5485 VPWR.n1392 VGND 9.44e-19
C5486 VPWR.n1393 VGND 9.84e-19
C5487 VPWR.n1394 VGND 8.2e-19
C5488 VPWR.n1395 VGND 0.001414f
C5489 VPWR.n1396 VGND 0.001281f
C5490 VPWR.n1397 VGND 0.002997f
C5491 VPWR.n1398 VGND 0.002078f
C5492 VPWR.n1399 VGND 0.00897f
C5493 VPWR.n1400 VGND 7.31e-19
C5494 VPWR.n1401 VGND 0.001224f
C5495 VPWR.n1402 VGND 8.2e-19
C5496 VPWR.n1403 VGND 6.56e-19
C5497 VPWR.n1404 VGND 0.001463f
C5498 VPWR.n1405 VGND 0.001414f
C5499 VPWR.n1406 VGND 0.001281f
C5500 VPWR.n1407 VGND 6.14e-19
C5501 VPWR.n1408 VGND 2.53e-19
C5502 VPWR.n1409 VGND 0.005411f
C5503 VPWR.n1410 VGND 0.008883f
C5504 VPWR.t622 VGND 0.002071f
C5505 VPWR.n1411 VGND 0.003648f
C5506 VPWR.n1412 VGND 0.002391f
C5507 VPWR.n1413 VGND 0.00145f
C5508 VPWR.n1414 VGND 0.001835f
C5509 VPWR.n1415 VGND 0.002447f
C5510 VPWR.n1416 VGND 0.001018f
C5511 VPWR.n1417 VGND 0.001365f
C5512 VPWR.t698 VGND 0.00177f
C5513 VPWR.n1418 VGND 0.001629f
C5514 VPWR.t33 VGND 4.31e-19
C5515 VPWR.n1419 VGND 0.001225f
C5516 VPWR.n1420 VGND 0.002402f
C5517 VPWR.t220 VGND 7.76e-19
C5518 VPWR.t222 VGND 7.76e-19
C5519 VPWR.n1421 VGND 0.001616f
C5520 VPWR.n1422 VGND 0.002503f
C5521 VPWR.n1423 VGND 5.67e-19
C5522 VPWR.n1424 VGND 0.002447f
C5523 VPWR.t316 VGND 4.77e-19
C5524 VPWR.t342 VGND 3.14e-19
C5525 VPWR.n1425 VGND 8.24e-19
C5526 VPWR.n1426 VGND 0.001933f
C5527 VPWR.n1427 VGND 0.002447f
C5528 VPWR.n1428 VGND 0.00145f
C5529 VPWR.n1429 VGND 5.43e-19
C5530 VPWR.t228 VGND 7.76e-19
C5531 VPWR.t198 VGND 7.76e-19
C5532 VPWR.n1430 VGND 0.001616f
C5533 VPWR.n1431 VGND 0.003026f
C5534 VPWR.t283 VGND 0.001191f
C5535 VPWR.t297 VGND 0.001631f
C5536 VPWR.n1432 VGND 0.004218f
C5537 VPWR.t200 VGND 7.48e-19
C5538 VPWR.t204 VGND 7.76e-19
C5539 VPWR.n1433 VGND 0.001574f
C5540 VPWR.n1434 VGND 0.002297f
C5541 VPWR.n1435 VGND 0.003141f
C5542 VPWR.n1436 VGND 4.55e-19
C5543 VPWR.n1437 VGND 0.002447f
C5544 VPWR.n1438 VGND 0.001888f
C5545 VPWR.n1439 VGND 8.2e-19
C5546 VPWR.n1440 VGND 0.001414f
C5547 VPWR.n1441 VGND 0.001281f
C5548 VPWR.n1442 VGND 0.001225f
C5549 VPWR.n1443 VGND 8.51e-19
C5550 VPWR.n1444 VGND 7.08e-19
C5551 VPWR.n1445 VGND 0.002408f
C5552 VPWR.n1446 VGND 0.002777f
C5553 VPWR.t202 VGND 7.76e-19
C5554 VPWR.t206 VGND 7.76e-19
C5555 VPWR.n1447 VGND 0.001602f
C5556 VPWR.t136 VGND 0.001139f
C5557 VPWR.n1448 VGND 0.001724f
C5558 VPWR.n1449 VGND 0.002461f
C5559 VPWR.n1450 VGND 6.5e-19
C5560 VPWR.n1451 VGND 5.23e-19
C5561 VPWR.n1452 VGND 8.51e-19
C5562 VPWR.n1453 VGND 9.31e-19
C5563 VPWR.n1454 VGND 8.2e-19
C5564 VPWR.n1455 VGND 6.56e-19
C5565 VPWR.n1456 VGND 0.001463f
C5566 VPWR.n1457 VGND 0.001414f
C5567 VPWR.n1458 VGND 0.001281f
C5568 VPWR.n1459 VGND 0.001225f
C5569 VPWR.n1460 VGND 0.001051f
C5570 VPWR.n1461 VGND 9.31e-19
C5571 VPWR.t461 VGND 0.021484f
C5572 VPWR.t560 VGND 0.03105f
C5573 VPWR.t620 VGND 0.019367f
C5574 VPWR.t804 VGND 0.009331f
C5575 VPWR.t124 VGND 0.011997f
C5576 VPWR.t697 VGND 0.011056f
C5577 VPWR.t225 VGND 0.008155f
C5578 VPWR.t219 VGND 0.012545f
C5579 VPWR.t32 VGND 0.006743f
C5580 VPWR.t221 VGND 0.0069f
C5581 VPWR.t315 VGND 0.006743f
C5582 VPWR.t223 VGND 0.007527f
C5583 VPWR.t217 VGND 0.0069f
C5584 VPWR.t341 VGND 0.005253f
C5585 VPWR.t227 VGND 0.008233f
C5586 VPWR.t197 VGND 0.008155f
C5587 VPWR.t282 VGND 0.006743f
C5588 VPWR.t199 VGND 0.011997f
C5589 VPWR.t203 VGND 0.007684f
C5590 VPWR.t296 VGND 0.006743f
C5591 VPWR.t207 VGND 0.006743f
C5592 VPWR.t690 VGND 0.006743f
C5593 VPWR.t211 VGND 0.008155f
C5594 VPWR.t344 VGND 0.006743f
C5595 VPWR.t201 VGND 0.007841f
C5596 VPWR.t135 VGND 0.006743f
C5597 VPWR.t205 VGND 0.005097f
C5598 VPWR.t209 VGND 0.005881f
C5599 VPWR.t306 VGND 0.012153f
C5600 VPWR.t478 VGND 0.007684f
C5601 VPWR.t55 VGND 0.007527f
C5602 VPWR.t770 VGND 0.016231f
C5603 VPWR.t792 VGND 0.015368f
C5604 VPWR.t813 VGND 0.015525f
C5605 VPWR.t113 VGND 0.005645f
C5606 VPWR.t308 VGND 0.006586f
C5607 VPWR.t30 VGND 0.007527f
C5608 VPWR.t51 VGND 0.016466f
C5609 VPWR.t115 VGND 0.017721f
C5610 VPWR.t715 VGND 0.008939f
C5611 VPWR.t172 VGND 0.00886f
C5612 VPWR.t290 VGND 0.00541f
C5613 VPWR.t739 VGND 0.008625f
C5614 VPWR.t91 VGND 0.011134f
C5615 VPWR.t717 VGND 0.009331f
C5616 VPWR.t724 VGND 0.006665f
C5617 VPWR.t288 VGND 0.00737f
C5618 VPWR.t786 VGND 0.008076f
C5619 VPWR.t736 VGND 0.009174f
C5620 VPWR.t171 VGND 0.011997f
C5621 VPWR.t65 VGND 0.006665f
C5622 VPWR.t331 VGND 0.008625f
C5623 VPWR.t87 VGND 0.014114f
C5624 VPWR.t169 VGND 0.008233f
C5625 VPWR.t737 VGND 0.002352f
C5626 VPWR.t827 VGND 0.007292f
C5627 VPWR.t764 VGND 0.010585f
C5628 VPWR.t762 VGND 0.007135f
C5629 VPWR.t811 VGND 0.006743f
C5630 VPWR.t766 VGND 0.0069f
C5631 VPWR.t802 VGND 0.00298f
C5632 VPWR.t760 VGND 0.007135f
C5633 VPWR.t215 VGND 0.010115f
C5634 VPWR.t213 VGND 0.012467f
C5635 VPWR.n1462 VGND 0.00802f
C5636 VPWR.n1463 VGND 0.004707f
C5637 VPWR.n1464 VGND 0.002485f
C5638 VPWR.t216 VGND 7.76e-19
C5639 VPWR.t761 VGND 7.76e-19
C5640 VPWR.n1465 VGND 0.001694f
C5641 VPWR.n1466 VGND 0.002808f
C5642 VPWR.n1467 VGND 7.08e-19
C5643 VPWR.n1468 VGND 0.001835f
C5644 VPWR.n1469 VGND 0.001556f
C5645 VPWR.n1470 VGND 8.38e-19
C5646 VPWR.n1471 VGND 5.04e-19
C5647 VPWR.t803 VGND 6.35e-19
C5648 VPWR.t812 VGND 6.35e-19
C5649 VPWR.n1472 VGND 0.00141f
C5650 VPWR.t767 VGND 7.76e-19
C5651 VPWR.t763 VGND 7.76e-19
C5652 VPWR.n1473 VGND 0.001692f
C5653 VPWR.n1474 VGND 0.00601f
C5654 VPWR.n1475 VGND 0.002221f
C5655 VPWR.n1476 VGND 0.001835f
C5656 VPWR.n1477 VGND 8.38e-19
C5657 VPWR.t765 VGND 0.002898f
C5658 VPWR.n1478 VGND 0.003667f
C5659 VPWR.t828 VGND 4.79e-19
C5660 VPWR.t738 VGND 4.79e-19
C5661 VPWR.n1479 VGND 9.97e-19
C5662 VPWR.n1480 VGND 0.002675f
C5663 VPWR.n1481 VGND 8.51e-19
C5664 VPWR.n1482 VGND 0.002208f
C5665 VPWR.n1483 VGND 0.002314f
C5666 VPWR.n1484 VGND 0.002378f
C5667 VPWR.n1485 VGND 7.07e-19
C5668 VPWR.t66 VGND 9.12e-19
C5669 VPWR.t787 VGND 0.001104f
C5670 VPWR.n1486 VGND 0.002621f
C5671 VPWR.n1487 VGND 0.001587f
C5672 VPWR.n1488 VGND 6.64e-19
C5673 VPWR.n1489 VGND 8.78e-19
C5674 VPWR.t718 VGND 0.00119f
C5675 VPWR.t289 VGND 0.001157f
C5676 VPWR.t92 VGND 5.61e-19
C5677 VPWR.n1490 VGND 0.002356f
C5678 VPWR.n1491 VGND 0.001807f
C5679 VPWR.n1492 VGND 0.003357f
C5680 VPWR.t716 VGND 5.7e-19
C5681 VPWR.t291 VGND 9.42e-19
C5682 VPWR.n1493 VGND 0.002611f
C5683 VPWR.n1494 VGND 0.003201f
C5684 VPWR.n1495 VGND 0.002447f
C5685 VPWR.t116 VGND 0.001178f
C5686 VPWR.n1496 VGND 0.002447f
C5687 VPWR.t52 VGND 0.003055f
C5688 VPWR.t31 VGND 7.48e-19
C5689 VPWR.t114 VGND 7.48e-19
C5690 VPWR.n1497 VGND 0.001676f
C5691 VPWR.n1498 VGND 4.9e-19
C5692 VPWR.t814 VGND 0.003177f
C5693 VPWR.n1499 VGND 0.004693f
C5694 VPWR.n1500 VGND 0.001117f
C5695 VPWR.t793 VGND 0.00177f
C5696 VPWR.n1501 VGND 0.001629f
C5697 VPWR.t771 VGND 4.31e-19
C5698 VPWR.n1502 VGND 0.001225f
C5699 VPWR.n1503 VGND 0.002968f
C5700 VPWR.t479 VGND 0.002071f
C5701 VPWR.n1504 VGND 0.002042f
C5702 VPWR.n1505 VGND 0.001539f
C5703 VPWR.n1506 VGND 9.04e-19
C5704 VPWR.n1507 VGND 9.31e-19
C5705 VPWR.n1508 VGND 0.001249f
C5706 VPWR.n1509 VGND 4.53e-19
C5707 VPWR.n1510 VGND 0.001224f
C5708 VPWR.n1511 VGND 0.001835f
C5709 VPWR.n1512 VGND 0.002447f
C5710 VPWR.n1513 VGND 4.71e-19
C5711 VPWR.n1514 VGND 0.002147f
C5712 VPWR.n1515 VGND 0.002894f
C5713 VPWR.n1516 VGND 0.002663f
C5714 VPWR.n1517 VGND 3.25e-19
C5715 VPWR.n1518 VGND 0.002447f
C5716 VPWR.n1519 VGND 0.002221f
C5717 VPWR.n1520 VGND 8.38e-19
C5718 VPWR.n1521 VGND 7.77e-19
C5719 VPWR.n1522 VGND 4.57e-19
C5720 VPWR.n1523 VGND 0.001835f
C5721 VPWR.n1524 VGND 0.001622f
C5722 VPWR.n1525 VGND 8.2e-19
C5723 VPWR.n1526 VGND 0.001463f
C5724 VPWR.n1527 VGND 6.56e-19
C5725 VPWR.n1528 VGND 8.2e-19
C5726 VPWR.n1529 VGND 0.001281f
C5727 VPWR.n1530 VGND 0.001225f
C5728 VPWR.n1531 VGND 8.51e-19
C5729 VPWR.n1532 VGND 8.41e-19
C5730 VPWR.n1533 VGND 0.001148f
C5731 VPWR.n1534 VGND 8.51e-19
C5732 VPWR.n1535 VGND 0.001224f
C5733 VPWR.n1536 VGND 8.2e-19
C5734 VPWR.n1537 VGND 0.001281f
C5735 VPWR.n1538 VGND 0.001414f
C5736 VPWR.n1539 VGND 0.053551f
C5737 VPWR.n1541 VGND 0.001463f
C5738 VPWR.n1542 VGND 0.001225f
C5739 VPWR.n1543 VGND 6.56e-19
C5740 VPWR.n1544 VGND 0.002314f
C5741 VPWR.t773 VGND 0.001154f
C5742 VPWR.t78 VGND 5.61e-19
C5743 VPWR.t810 VGND 0.001157f
C5744 VPWR.n1545 VGND 0.002356f
C5745 VPWR.n1546 VGND 8.67e-19
C5746 VPWR.n1547 VGND 0.002447f
C5747 VPWR.t40 VGND 5.61e-19
C5748 VPWR.t7 VGND 0.001157f
C5749 VPWR.n1548 VGND 0.002356f
C5750 VPWR.t48 VGND 0.001168f
C5751 VPWR.n1549 VGND 8.29e-19
C5752 VPWR.n1550 VGND 0.001835f
C5753 VPWR.n1551 VGND 7.68e-19
C5754 VPWR.t50 VGND 7.48e-19
C5755 VPWR.t154 VGND 7.48e-19
C5756 VPWR.n1552 VGND 0.001676f
C5757 VPWR.n1553 VGND 0.002157f
C5758 VPWR.n1554 VGND 4.71e-19
C5759 VPWR.n1555 VGND 0.002447f
C5760 VPWR.n1556 VGND 0.002447f
C5761 VPWR.n1557 VGND 0.002447f
C5762 VPWR.n1558 VGND 5.32e-19
C5763 VPWR.n1559 VGND 0.002014f
C5764 VPWR.n1560 VGND 0.001732f
C5765 VPWR.n1561 VGND 6.64e-19
C5766 VPWR.n1562 VGND 8.67e-19
C5767 VPWR.n1563 VGND 0.002447f
C5768 VPWR.n1564 VGND 0.002447f
C5769 VPWR.n1565 VGND 0.002447f
C5770 VPWR.n1566 VGND 6.36e-19
C5771 VPWR.n1567 VGND 0.001741f
C5772 VPWR.n1568 VGND 0.002321f
C5773 VPWR.n1569 VGND 5.61e-19
C5774 VPWR.n1570 VGND 8.51e-19
C5775 VPWR.n1571 VGND 6.56e-19
C5776 VPWR.n1572 VGND 8.2e-19
C5777 VPWR.n1573 VGND 0.001197f
C5778 VPWR.n1574 VGND 8.51e-19
C5779 VPWR.n1575 VGND 0.001224f
C5780 VPWR.n1576 VGND 8.2e-19
C5781 VPWR.n1577 VGND 0.001269f
C5782 VPWR.n1578 VGND 0.001426f
C5783 VPWR.n1579 VGND 0.053196f
C5784 VPWR.n1580 VGND 0.001426f
C5785 VPWR.n1581 VGND 0.001269f
C5786 VPWR.n1582 VGND 6.14e-19
C5787 VPWR.n1583 VGND 2.53e-19
C5788 VPWR.n1584 VGND 5.65e-19
C5789 VPWR.n1585 VGND 0.008386f
C5790 VPWR.n1586 VGND 0.002877f
C5791 VPWR.n1587 VGND 0.00255f
C5792 VPWR.n1588 VGND 0.00145f
C5793 VPWR.n1589 VGND 0.001224f
C5794 VPWR.n1590 VGND 0.001835f
C5795 VPWR.n1591 VGND 7.16e-19
C5796 VPWR.n1592 VGND 0.002493f
C5797 VPWR.n1593 VGND 0.002772f
C5798 VPWR.t295 VGND 3.14e-19
C5799 VPWR.t150 VGND 3.14e-19
C5800 VPWR.n1594 VGND 7.27e-19
C5801 VPWR.n1595 VGND 0.009854f
C5802 VPWR.n1596 VGND 0.002021f
C5803 VPWR.n1597 VGND 8.25e-19
C5804 VPWR.n1598 VGND 9.31e-19
C5805 VPWR.n1599 VGND 8.2e-19
C5806 VPWR.n1600 VGND 0.001414f
C5807 VPWR.n1601 VGND 0.001281f
C5808 VPWR.n1602 VGND 0.001146f
C5809 VPWR.n1603 VGND 9.04e-19
C5810 VPWR.n1604 VGND 0.002454f
C5811 VPWR.t470 VGND 0.002071f
C5812 VPWR.n1605 VGND 0.001902f
C5813 VPWR.n1606 VGND 0.003989f
C5814 VPWR.n1607 VGND 0.006561f
C5815 VPWR.n1608 VGND 0.004818f
C5816 VPWR.t326 VGND 0.001255f
C5817 VPWR.t471 VGND 0.002071f
C5818 VPWR.n1609 VGND 0.001797f
C5819 VPWR.n1610 VGND 0.00513f
C5820 VPWR.n1611 VGND 0.005062f
C5821 VPWR.n1612 VGND 8.51e-19
C5822 VPWR.n1613 VGND 0.001224f
C5823 VPWR.n1614 VGND 8.2e-19
C5824 VPWR.n1615 VGND 6.56e-19
C5825 VPWR.n1616 VGND 0.001463f
C5826 VPWR.n1617 VGND 0.001414f
C5827 VPWR.n1618 VGND 0.001281f
C5828 VPWR.n1619 VGND 2.28e-19
C5829 VPWR.n1620 VGND 8.38e-19
C5830 VPWR.t330 VGND 7.48e-19
C5831 VPWR.t82 VGND 7.48e-19
C5832 VPWR.n1621 VGND 0.001628f
C5833 VPWR.n1622 VGND 0.00206f
C5834 VPWR.t686 VGND 0.002088f
C5835 VPWR.t922 VGND 0.004432f
C5836 VPWR.n1624 VGND 0.011362f
C5837 VPWR.t687 VGND 0.002088f
C5838 VPWR.n1625 VGND 0.006189f
C5839 VPWR.t90 VGND 0.002626f
C5840 VPWR.n1626 VGND 4.71e-19
C5841 VPWR.t789 VGND 7.48e-19
C5842 VPWR.t293 VGND 7.48e-19
C5843 VPWR.n1627 VGND 0.001676f
C5844 VPWR.n1628 VGND 0.002157f
C5845 VPWR.n1629 VGND 0.001835f
C5846 VPWR.t791 VGND 0.001178f
C5847 VPWR.t13 VGND 7.48e-19
C5848 VPWR.t337 VGND 7.48e-19
C5849 VPWR.n1630 VGND 0.001676f
C5850 VPWR.n1631 VGND 0.002157f
C5851 VPWR.n1632 VGND 0.001942f
C5852 VPWR.t11 VGND 0.001178f
C5853 VPWR.t191 VGND 5.61e-19
C5854 VPWR.t184 VGND 0.001157f
C5855 VPWR.n1633 VGND 0.002356f
C5856 VPWR.n1634 VGND 0.001831f
C5857 VPWR.n1635 VGND 3.91e-19
C5858 VPWR.n1636 VGND 0.002965f
C5859 VPWR.n1637 VGND 7.77e-19
C5860 VPWR.n1638 VGND 0.002447f
C5861 VPWR.n1639 VGND 0.002447f
C5862 VPWR.n1640 VGND 2.26e-19
C5863 VPWR.n1641 VGND 0.002965f
C5864 VPWR.n1642 VGND 7.77e-19
C5865 VPWR.n1643 VGND 0.001835f
C5866 VPWR.n1644 VGND 0.002447f
C5867 VPWR.n1645 VGND 0.001835f
C5868 VPWR.n1646 VGND 5.18e-19
C5869 VPWR.n1647 VGND 0.001513f
C5870 VPWR.n1648 VGND 0.005529f
C5871 VPWR.n1649 VGND 0.005029f
C5872 VPWR.t413 VGND 0.021641f
C5873 VPWR.t122 VGND 0.011997f
C5874 VPWR.t9 VGND 0.007998f
C5875 VPWR.t522 VGND 0.007292f
C5876 VPWR.t131 VGND 0.01035f
C5877 VPWR.t284 VGND 0.016544f
C5878 VPWR.t729 VGND 0.003764f
C5879 VPWR.t177 VGND 0.006665f
C5880 VPWR.t140 VGND 0.006586f
C5881 VPWR.t821 VGND 0.007449f
C5882 VPWR.t287 VGND 0.014741f
C5883 VPWR.t22 VGND 0.008076f
C5884 VPWR.t800 VGND 0.006665f
C5885 VPWR.t231 VGND 0.01035f
C5886 VPWR.t825 VGND 0.007449f
C5887 VPWR.t823 VGND 0.007449f
C5888 VPWR.t286 VGND 0.008076f
C5889 VPWR.t183 VGND 0.006586f
C5890 VPWR.t139 VGND 0.01035f
C5891 VPWR.t190 VGND 0.008939f
C5892 VPWR.t10 VGND 0.007449f
C5893 VPWR.t824 VGND 0.012702f
C5894 VPWR.t232 VGND 0.01035f
C5895 VPWR.t336 VGND 0.008939f
C5896 VPWR.t790 VGND 0.006586f
C5897 VPWR.t12 VGND 0.016466f
C5898 VPWR.t292 VGND 0.016152f
C5899 VPWR.t753 VGND 0.006586f
C5900 VPWR.t788 VGND 0.014741f
C5901 VPWR.t89 VGND 0.010429f
C5902 VPWR.t81 VGND 0.008547f
C5903 VPWR.t685 VGND 0.006586f
C5904 VPWR.t329 VGND 0.010036f
C5905 VPWR.t36 VGND 0.009644f
C5906 VPWR.n1650 VGND 0.008565f
C5907 VPWR.t325 VGND 0.012153f
C5908 VPWR.t469 VGND 0.006586f
C5909 VPWR.t300 VGND 0.010821f
C5910 VPWR.t4 VGND 0.014427f
C5911 VPWR.t165 VGND 0.007135f
C5912 VPWR.t149 VGND 0.005724f
C5913 VPWR.t304 VGND 0.006586f
C5914 VPWR.t294 VGND 0.00737f
C5915 VPWR.t147 VGND 0.007292f
C5916 VPWR.t695 VGND 0.007527f
C5917 VPWR.t327 VGND 0.007449f
C5918 VPWR.t41 VGND 0.007527f
C5919 VPWR.t348 VGND 0.014741f
C5920 VPWR.t192 VGND 0.015133f
C5921 VPWR.t85 VGND 0.003999f
C5922 VPWR.t817 VGND 0.006586f
C5923 VPWR.t333 VGND 0.007292f
C5924 VPWR.t346 VGND 0.007527f
C5925 VPWR.t161 VGND 0.009017f
C5926 VPWR.t173 VGND 0.007214f
C5927 VPWR.t324 VGND 0.003764f
C5928 VPWR.t128 VGND 0.007449f
C5929 VPWR.t45 VGND 0.014663f
C5930 VPWR.t809 VGND 0.014741f
C5931 VPWR.t772 VGND 0.01035f
C5932 VPWR.t77 VGND 0.006665f
C5933 VPWR.t735 VGND 0.007449f
C5934 VPWR.t335 VGND 0.007449f
C5935 VPWR.t44 VGND 0.006586f
C5936 VPWR.t323 VGND 0.008076f
C5937 VPWR.t6 VGND 0.008939f
C5938 VPWR.t47 VGND 0.01035f
C5939 VPWR.t39 VGND 0.01333f
C5940 VPWR.t43 VGND 0.010585f
C5941 VPWR.t153 VGND 0.006586f
C5942 VPWR.t734 VGND 0.006586f
C5943 VPWR.t49 VGND 0.008939f
C5944 VPWR.t780 VGND 0.011761f
C5945 VPWR.n1651 VGND 0.013116f
C5946 VPWR.n1652 VGND 0.004512f
C5947 VPWR.n1653 VGND 9.31e-19
C5948 VPWR.n1654 VGND 0.001051f
C5949 VPWR.n1655 VGND 0.001225f
C5950 VPWR.n1656 VGND 0.001281f
C5951 VPWR.n1657 VGND 0.001414f
C5952 VPWR.n1658 VGND 0.053196f
C5953 VPWR.n1659 VGND 0.001414f
C5954 VPWR.n1660 VGND 0.001463f
C5955 VPWR.n1661 VGND 6.56e-19
C5956 VPWR.n1662 VGND 8.2e-19
C5957 VPWR.n1663 VGND 3.86e-19
C5958 VPWR.n1664 VGND 7.85e-19
C5959 VPWR.n1665 VGND 5.65e-19
C5960 VPWR.n1666 VGND 0.004756f
C5961 VPWR.n1667 VGND 5.61e-19
C5962 VPWR.n1668 VGND 0.003931f
C5963 VPWR.n1669 VGND 0.002447f
C5964 VPWR.n1670 VGND 0.002447f
C5965 VPWR.n1671 VGND 0.002447f
C5966 VPWR.n1672 VGND 8.67e-19
C5967 VPWR.n1673 VGND 8.67e-19
C5968 VPWR.n1674 VGND 6.64e-19
C5969 VPWR.n1675 VGND 0.002447f
C5970 VPWR.n1676 VGND 0.002447f
C5971 VPWR.n1677 VGND 0.002447f
C5972 VPWR.n1678 VGND 8.67e-19
C5973 VPWR.n1679 VGND 8.67e-19
C5974 VPWR.n1680 VGND 6.22e-19
C5975 VPWR.n1681 VGND 0.002447f
C5976 VPWR.n1682 VGND 0.00125f
C5977 VPWR.n1683 VGND 8.8e-19
C5978 VPWR.n1684 VGND 8.2e-19
C5979 VPWR.n1685 VGND 0.001463f
C5980 VPWR.n1686 VGND 6.56e-19
C5981 VPWR.n1687 VGND 0.001281f
C5982 VPWR.n1688 VGND 8.2e-19
C5983 VPWR.n1689 VGND 0.001197f
C5984 VPWR.n1690 VGND 8.51e-19
C5985 VPWR.n1691 VGND 7.77e-19
C5986 VPWR.n1692 VGND 0.00388f
C5987 VPWR.n1693 VGND 4.71e-19
C5988 VPWR.n1694 VGND 8.51e-19
C5989 VPWR.n1695 VGND 9.84e-19
C5990 VPWR.n1696 VGND 8.2e-19
C5991 VPWR.n1697 VGND 0.001281f
C5992 VPWR.n1698 VGND 0.001414f
C5993 VPWR.n1699 VGND 0.053196f
C5994 VPWR.n1700 VGND 0.221149f
C5995 VPWR.n1701 VGND 0.081008f
C5996 VPWR.n1702 VGND 0.040334f
C5997 VPWR.n1703 VGND 0.044685f
C5998 VPWR.n1704 VGND 0.10196f
C5999 VPWR.n1705 VGND 0.001269f
C6000 VPWR.n1706 VGND 8.2e-19
C6001 VPWR.n1707 VGND 0.001197f
C6002 VPWR.n1708 VGND 8.51e-19
C6003 VPWR.n1709 VGND 0.001183f
C6004 VPWR.t494 VGND 0.002071f
C6005 VPWR.n1710 VGND 0.002042f
C6006 VPWR.n1711 VGND 0.007818f
C6007 VPWR.n1712 VGND 0.004818f
C6008 VPWR.n1713 VGND 0.006214f
C6009 VPWR.n1714 VGND 0.001835f
C6010 VPWR.n1715 VGND 8.38e-19
C6011 VPWR.n1716 VGND 0.002342f
C6012 VPWR.n1717 VGND 0.003701f
C6013 VPWR.n1718 VGND 0.003581f
C6014 VPWR.n1719 VGND 0.002221f
C6015 VPWR.n1720 VGND 0.001835f
C6016 VPWR.n1721 VGND 9.31e-19
C6017 VPWR.n1722 VGND 5.85e-19
C6018 VPWR.t657 VGND 0.002071f
C6019 VPWR.n1723 VGND 0.003648f
C6020 VPWR.n1724 VGND 0.002454f
C6021 VPWR.n1725 VGND 0.001835f
C6022 VPWR.n1726 VGND 0.001835f
C6023 VPWR.n1727 VGND 8.38e-19
C6024 VPWR.n1728 VGND 0.003421f
C6025 VPWR.n1729 VGND 0.004694f
C6026 VPWR.n1730 VGND 0.006214f
C6027 VPWR.t120 VGND 4.31e-19
C6028 VPWR.t303 VGND 4.31e-19
C6029 VPWR.n1731 VGND 9.01e-19
C6030 VPWR.t658 VGND 0.002071f
C6031 VPWR.n1732 VGND 0.003089f
C6032 VPWR.n1733 VGND 0.005595f
C6033 VPWR.n1734 VGND 0.00377f
C6034 VPWR.n1735 VGND 0.001888f
C6035 VPWR.n1736 VGND 0.001225f
C6036 VPWR.n1737 VGND 7.85e-19
C6037 VPWR.n1738 VGND 8.2e-19
C6038 VPWR.n1739 VGND 3.86e-19
C6039 VPWR.n1740 VGND 6.12e-19
C6040 VPWR.n1741 VGND 3.06e-19
C6041 VPWR.n1742 VGND 7.41e-19
C6042 VPWR.n1743 VGND 0.003244f
C6043 VPWR.t528 VGND 0.021641f
C6044 VPWR.t275 VGND 0.007292f
C6045 VPWR.t34 VGND 0.007135f
C6046 VPWR.t338 VGND 0.009644f
C6047 VPWR.t103 VGND 0.013173f
C6048 VPWR.t101 VGND 0.0069f
C6049 VPWR.t105 VGND 0.00541f
C6050 VPWR.t339 VGND 0.015917f
C6051 VPWR.t806 VGND 0.015525f
C6052 VPWR.t493 VGND 0.012938f
C6053 VPWR.t794 VGND 0.007135f
C6054 VPWR.t727 VGND 0.003058f
C6055 VPWR.t67 VGND 0.0069f
C6056 VPWR.t353 VGND 0.00737f
C6057 VPWR.t298 VGND 0.008625f
C6058 VPWR.t83 VGND 0.011056f
C6059 VPWR.t277 VGND 0.021798f
C6060 VPWR.t656 VGND 0.002431f
C6061 VPWR.t273 VGND 0.007998f
C6062 VPWR.t119 VGND 0.015995f
C6063 VPWR.t302 VGND 0.011369f
C6064 VPWR.t69 VGND 0.007214f
C6065 VPWR.t815 VGND 0.009331f
C6066 VPWR.t117 VGND 0.017877f
C6067 VPWR.t387 VGND 0.007919f
C6068 VPWR.t709 VGND 0.0069f
C6069 VPWR.t237 VGND 0.006508f
C6070 VPWR.t235 VGND 0.007214f
C6071 VPWR.t311 VGND 0.012153f
C6072 VPWR.t648 VGND 0.013094f
C6073 VPWR.t699 VGND 0.019054f
C6074 VPWR.t26 VGND 0.009331f
C6075 VPWR.t455 VGND 0.007214f
C6076 VPWR.t612 VGND 0.043204f
C6077 VPWR.t163 VGND 0.019054f
C6078 VPWR.t349 VGND 0.007214f
C6079 VPWR.t309 VGND 0.002431f
C6080 VPWR.t725 VGND 0.010429f
C6081 VPWR.t819 VGND 0.014898f
C6082 VPWR.t351 VGND 0.008939f
C6083 VPWR.t443 VGND 0.007841f
C6084 VPWR.t79 VGND 0.009488f
C6085 VPWR.n1744 VGND 0.02207f
C6086 VPWR.n1745 VGND 0.009207f
C6087 VPWR.t899 VGND 0.012177f
C6088 VPWR.t80 VGND 0.001139f
C6089 VPWR.n1746 VGND 0.004694f
C6090 VPWR.n1747 VGND 0.002447f
C6091 VPWR.t352 VGND 4.31e-19
C6092 VPWR.t820 VGND 4.31e-19
C6093 VPWR.n1748 VGND 9.01e-19
C6094 VPWR.t445 VGND 0.002071f
C6095 VPWR.n1749 VGND 0.003648f
C6096 VPWR.t726 VGND 0.001631f
C6097 VPWR.t310 VGND 0.001191f
C6098 VPWR.n1750 VGND 0.00425f
C6099 VPWR.n1751 VGND 8.38e-19
C6100 VPWR.n1752 VGND 0.001609f
C6101 VPWR.t350 VGND 6.35e-19
C6102 VPWR.t164 VGND 6.35e-19
C6103 VPWR.n1753 VGND 0.00141f
C6104 VPWR.n1754 VGND 0.001041f
C6105 VPWR.n1755 VGND 8.2e-19
C6106 VPWR.n1756 VGND 0.001197f
C6107 VPWR.n1757 VGND 0.001369f
C6108 VPWR.t613 VGND 0.002071f
C6109 VPWR.t843 VGND 0.012096f
C6110 VPWR.n1758 VGND 0.006349f
C6111 VPWR.n1759 VGND 0.008368f
C6112 VPWR.n1760 VGND 8.2e-19
C6113 VPWR.n1761 VGND 8.78e-19
C6114 VPWR.n1762 VGND 0.002447f
C6115 VPWR.t891 VGND 0.030181f
C6116 VPWR.t614 VGND 0.002071f
C6117 VPWR.n1763 VGND 0.004756f
C6118 VPWR.t27 VGND 6.35e-19
C6119 VPWR.t700 VGND 6.35e-19
C6120 VPWR.n1764 VGND 0.00138f
C6121 VPWR.n1765 VGND 0.005753f
C6122 VPWR.t457 VGND 0.002286f
C6123 VPWR.n1766 VGND 0.004705f
C6124 VPWR.n1767 VGND 0.001766f
C6125 VPWR.t236 VGND 6.29e-19
C6126 VPWR.t312 VGND 2.34e-19
C6127 VPWR.n1768 VGND 0.002889f
C6128 VPWR.t238 VGND 6.35e-19
C6129 VPWR.t388 VGND 6.35e-19
C6130 VPWR.n1769 VGND 0.00138f
C6131 VPWR.n1770 VGND 0.003352f
C6132 VPWR.n1771 VGND 3.88e-19
C6133 VPWR.n1772 VGND 8.2e-19
C6134 VPWR.n1773 VGND 6.12e-19
C6135 VPWR.n1774 VGND 9.97e-19
C6136 VPWR.n1775 VGND 3.06e-19
C6137 VPWR.n1776 VGND 5.13e-19
C6138 VPWR.n1777 VGND 0.006439f
C6139 VPWR.t650 VGND 0.002102f
C6140 VPWR.n1778 VGND 0.002457f
C6141 VPWR.n1779 VGND 0.009561f
C6142 VPWR.t829 VGND 0.008778f
C6143 VPWR.n1780 VGND 0.008691f
C6144 VPWR.t649 VGND 0.002071f
C6145 VPWR.n1781 VGND 0.002493f
C6146 VPWR.n1782 VGND 0.002473f
C6147 VPWR.n1783 VGND 0.001307f
C6148 VPWR.n1784 VGND 9.31e-19
C6149 VPWR.n1785 VGND 0.002598f
C6150 VPWR.n1786 VGND 0.003084f
C6151 VPWR.n1787 VGND 0.001835f
C6152 VPWR.n1788 VGND 0.002221f
C6153 VPWR.n1789 VGND 8.38e-19
C6154 VPWR.n1790 VGND 0.002939f
C6155 VPWR.n1791 VGND 0.00372f
C6156 VPWR.n1792 VGND 0.00145f
C6157 VPWR.n1793 VGND 0.002447f
C6158 VPWR.n1794 VGND 0.006058f
C6159 VPWR.n1795 VGND 0.016876f
C6160 VPWR.n1796 VGND 0.006622f
C6161 VPWR.n1797 VGND 0.008594f
C6162 VPWR.n1798 VGND 0.001622f
C6163 VPWR.n1799 VGND 0.001225f
C6164 VPWR.n1800 VGND 8.51e-19
C6165 VPWR.n1801 VGND 0.004086f
C6166 VPWR.t456 VGND 0.002279f
C6167 VPWR.n1802 VGND 0.004985f
C6168 VPWR.n1803 VGND 0.001597f
C6169 VPWR.n1804 VGND 8.51e-19
C6170 VPWR.n1805 VGND 8.2e-19
C6171 VPWR.n1806 VGND 6.12e-19
C6172 VPWR.n1807 VGND 4.52e-19
C6173 VPWR.n1808 VGND 6.14e-19
C6174 VPWR.n1809 VGND 0.001224f
C6175 VPWR.n1810 VGND 7.11e-19
C6176 VPWR.n1811 VGND 0.003727f
C6177 VPWR.n1812 VGND 0.003879f
C6178 VPWR.n1813 VGND 0.002096f
C6179 VPWR.n1814 VGND 0.00145f
C6180 VPWR.n1815 VGND 0.002447f
C6181 VPWR.n1816 VGND 0.005655f
C6182 VPWR.n1817 VGND 0.005805f
C6183 VPWR.n1818 VGND 0.00377f
C6184 VPWR.n1819 VGND 0.006214f
C6185 VPWR.n1820 VGND 0.002221f
C6186 VPWR.n1821 VGND 8.38e-19
C6187 VPWR.n1822 VGND 0.013527f
C6188 VPWR.t444 VGND 0.002071f
C6189 VPWR.n1823 VGND 0.003648f
C6190 VPWR.n1824 VGND 0.002273f
C6191 VPWR.n1825 VGND 9.31e-19
C6192 VPWR.n1826 VGND 9.31e-19
C6193 VPWR.n1827 VGND 0.001436f
C6194 VPWR.n1828 VGND 7.3e-19
C6195 VPWR.n1829 VGND 0.003168f
C6196 VPWR.n1830 VGND 8.51e-19
C6197 VPWR.n1831 VGND 9.97e-19
C6198 VPWR.n1832 VGND 8.2e-19
C6199 VPWR.n1833 VGND 6.56e-19
C6200 VPWR.n1834 VGND 0.033802f
C6201 VPWR.n1835 VGND 0.044685f
C6202 VPWR.n1836 VGND 0.040593f
C6203 VPWR.n1837 VGND 0.122046f
C6204 VPWR.n1838 VGND 0.025756f
C6205 VPWR.n1839 VGND 0.221149f
C6206 VPWR.n1840 VGND 0.117032f
C6207 VPWR.n1841 VGND 0.026244f
C6208 VPWR.n1842 VGND 0.058516f
C6209 VPWR.n1843 VGND 0.032796f
C6210 VPWR.n1844 VGND 0.117014f
C6211 VPWR.n1845 VGND 0.057872f
C6212 VPWR.n1846 VGND 0.057872f
C6213 VPWR.n1847 VGND 0.087246f
C6214 VPWR.n1848 VGND 0.12165f
C6215 VPWR.n1849 VGND 0.02498f
C6216 VPWR.n1850 VGND 0.06951f
C6217 VPWR.n1851 VGND 0.117032f
C6218 VPWR.n1852 VGND 0.02498f
C6219 VPWR.n1853 VGND 0.040161f
C6220 VPWR.n1854 VGND 0.044685f
C6221 VPWR.n1855 VGND 0.032759f
C6222 VPWR.n1856 VGND 0.001269f
C6223 VPWR.n1857 VGND 0.001225f
C6224 VPWR.n1858 VGND 0.001716f
C6225 VPWR.n1859 VGND 8.38e-19
C6226 VPWR.n1860 VGND 8.07e-19
C6227 VPWR.n1861 VGND 0.002454f
C6228 VPWR.n1862 VGND 0.00145f
C6229 VPWR.n1863 VGND 0.001835f
C6230 VPWR.n1864 VGND 0.004853f
C6231 VPWR.n1865 VGND 0.006423f
C6232 VPWR.n1866 VGND 0.004678f
C6233 VPWR.n1867 VGND 0.002447f
C6234 VPWR.n1868 VGND 0.002447f
C6235 VPWR.n1869 VGND 0.002221f
C6236 VPWR.n1870 VGND 0.004748f
C6237 VPWR.n1871 VGND 0.019307f
C6238 VPWR.n1872 VGND 0.003804f
C6239 VPWR.n1873 VGND 0.004364f
C6240 VPWR.n1874 VGND 8.38e-19
C6241 VPWR.n1875 VGND 9.44e-19
C6242 VPWR.n1876 VGND 0.002273f
C6243 VPWR.n1877 VGND 0.005166f
C6244 VPWR.n1878 VGND 4.8e-19
C6245 VPWR.n1879 VGND 8.51e-19
C6246 VPWR.n1880 VGND 0.001224f
C6247 VPWR.n1881 VGND 8.2e-19
C6248 VPWR.n1882 VGND 6.56e-19
C6249 VPWR.n1883 VGND 0.032584f
C6250 VPWR.n1884 VGND 0.044685f
C6251 VPWR.n1885 VGND 0.048231f
C6252 VPWR.n1886 VGND 0.117032f
C6253 VPWR.n1887 VGND 0.117032f
C6254 VPWR.n1888 VGND 0.06951f
C6255 VPWR.n1889 VGND 0.048231f
C6256 VPWR.n1890 VGND 0.053196f
C6257 VPWR.n1891 VGND 0.001463f
C6258 VPWR.n1892 VGND 6.56e-19
C6259 VPWR.n1893 VGND 6.12e-19
C6260 VPWR.n1894 VGND 8.51e-19
C6261 VPWR.n1895 VGND 8.78e-19
C6262 VPWR.t123 VGND 0.002929f
C6263 VPWR.t524 VGND 0.002071f
C6264 VPWR.n1896 VGND 0.00777f
C6265 VPWR.n1897 VGND 0.002273f
C6266 VPWR.t623 VGND 0.002088f
C6267 VPWR.t852 VGND 0.004432f
C6268 VPWR.n1899 VGND 0.011362f
C6269 VPWR.t624 VGND 0.002088f
C6270 VPWR.n1900 VGND 0.006189f
C6271 VPWR.t414 VGND 0.002088f
C6272 VPWR.t909 VGND 0.004432f
C6273 VPWR.n1902 VGND 0.011362f
C6274 VPWR.t415 VGND 0.002088f
C6275 VPWR.n1903 VGND 0.006189f
C6276 VPWR.n1904 VGND 8.2e-19
C6277 VPWR.n1905 VGND 0.001414f
C6278 VPWR.n1906 VGND 0.001281f
C6279 VPWR.n1907 VGND 0.001199f
C6280 VPWR.n1908 VGND 5.72e-19
C6281 VPWR.n1909 VGND 0.005217f
C6282 VPWR.n1910 VGND 8.51e-19
C6283 VPWR.n1911 VGND 0.001224f
C6284 VPWR.n1912 VGND 8.2e-19
C6285 VPWR.n1913 VGND 6.56e-19
C6286 VPWR.n1914 VGND 0.001463f
C6287 VPWR.n1915 VGND 0.001414f
C6288 VPWR.n1916 VGND 0.001281f
C6289 VPWR.n1917 VGND 0.001225f
C6290 VPWR.n1918 VGND 0.002128f
C6291 VPWR.n1919 VGND 8.51e-19
C6292 VPWR.n1920 VGND 0.006423f
C6293 VPWR.n1921 VGND 0.006354f
C6294 VPWR.n1922 VGND 0.005012f
C6295 VPWR.n1923 VGND 0.013387f
C6296 VPWR.n1924 VGND 0.002447f
C6297 VPWR.n1925 VGND 0.001835f
C6298 VPWR.n1926 VGND 0.002234f
C6299 VPWR.n1927 VGND 0.002359f
C6300 VPWR.n1928 VGND 0.00145f
C6301 VPWR.n1929 VGND 0.002447f
C6302 VPWR.n1930 VGND 0.002447f
C6303 VPWR.n1931 VGND 5.61e-19
C6304 VPWR.n1932 VGND 0.002524f
C6305 VPWR.n1933 VGND 5.75e-19
C6306 VPWR.n1934 VGND 0.002447f
C6307 VPWR.n1935 VGND 0.001995f
C6308 VPWR.n1936 VGND 6.36e-19
C6309 VPWR.n1937 VGND 8.67e-19
C6310 VPWR.n1938 VGND 8.51e-19
C6311 VPWR.n1939 VGND 0.001224f
C6312 VPWR.n1940 VGND 8.2e-19
C6313 VPWR.n1941 VGND 0.001463f
C6314 VPWR.n1942 VGND 6.56e-19
C6315 VPWR.n1943 VGND 8.2e-19
C6316 VPWR.n1944 VGND 8.78e-19
C6317 VPWR.n1945 VGND 0.001197f
C6318 VPWR.n1946 VGND 8.2e-19
C6319 VPWR.n1947 VGND 0.001281f
C6320 VPWR.n1948 VGND 0.001414f
C6321 VPWR.n1949 VGND 0.053196f
C6322 VPWR.n1950 VGND 0.053551f
C6323 VPWR.n1951 VGND 0.001414f
C6324 VPWR.n1952 VGND 0.001463f
C6325 VPWR.n1953 VGND 6.56e-19
C6326 VPWR.n1954 VGND 8.2e-19
C6327 VPWR.n1955 VGND 0.001197f
C6328 VPWR.n1956 VGND 8.51e-19
C6329 VPWR.n1957 VGND 0.003084f
C6330 VPWR.n1958 VGND 0.003084f
C6331 VPWR.n1959 VGND 0.002363f
C6332 VPWR.n1960 VGND 0.002447f
C6333 VPWR.n1961 VGND 0.002447f
C6334 VPWR.n1962 VGND 0.002263f
C6335 VPWR.n1963 VGND 0.003084f
C6336 VPWR.n1964 VGND 0.002263f
C6337 VPWR.n1965 VGND 0.002447f
C6338 VPWR.n1966 VGND 0.002447f
C6339 VPWR.n1967 VGND 0.002011f
C6340 VPWR.n1968 VGND 0.003353f
C6341 VPWR.n1969 VGND 0.001894f
C6342 VPWR.n1970 VGND 0.00295f
C6343 VPWR.n1971 VGND 0.002447f
C6344 VPWR.n1972 VGND 0.001835f
C6345 VPWR.n1973 VGND 9.44e-19
C6346 VPWR.n1974 VGND 6.83e-19
C6347 VPWR.n1975 VGND 0.005166f
C6348 VPWR.n1976 VGND 9.31e-19
C6349 VPWR.n1977 VGND 2.28e-19
C6350 VPWR.n1978 VGND 0.001281f
C6351 VPWR.n1979 VGND 8.2e-19
C6352 VPWR.n1980 VGND 0.001224f
C6353 VPWR.n1981 VGND 8.51e-19
C6354 VPWR.n1982 VGND 0.003282f
C6355 VPWR.n1983 VGND 0.004818f
C6356 VPWR.n1984 VGND 8.51e-19
C6357 VPWR.n1985 VGND 9.31e-19
C6358 VPWR.n1986 VGND 8.2e-19
C6359 VPWR.n1987 VGND 0.001281f
C6360 VPWR.n1988 VGND 0.001414f
C6361 VPWR.n1989 VGND 0.053551f
C6362 VPWR.n1990 VGND 0.048231f
C6363 VPWR.n1991 VGND 0.117032f
C6364 VPWR.n1992 VGND 0.117032f
C6365 VPWR.n1993 VGND 0.06951f
C6366 VPWR.n1994 VGND 0.048231f
C6367 VPWR.n1995 VGND 0.058516f
C6368 VPWR.n1996 VGND 0.001414f
C6369 VPWR.n1997 VGND 0.001463f
C6370 VPWR.n1998 VGND 0.001463f
C6371 VPWR.n1999 VGND 6.56e-19
C6372 VPWR.n2000 VGND 8.2e-19
C6373 VPWR.n2001 VGND 6.12e-19
C6374 VPWR.n2002 VGND 3.06e-19
C6375 VPWR.n2003 VGND 0.003046f
C6376 VPWR.t546 VGND 0.002279f
C6377 VPWR.n2004 VGND 0.004985f
C6378 VPWR.n2005 VGND 0.008359f
C6379 VPWR.n2006 VGND 0.006481f
C6380 VPWR.n2007 VGND 0.002447f
C6381 VPWR.n2008 VGND 0.001835f
C6382 VPWR.n2009 VGND 0.00372f
C6383 VPWR.n2010 VGND 0.001665f
C6384 VPWR.n2011 VGND 0.001835f
C6385 VPWR.n2012 VGND 0.002447f
C6386 VPWR.n2013 VGND 0.002815f
C6387 VPWR.n2014 VGND 0.001717f
C6388 VPWR.n2015 VGND 0.003554f
C6389 VPWR.n2016 VGND 0.002113f
C6390 VPWR.n2017 VGND 0.002447f
C6391 VPWR.n2018 VGND 0.002447f
C6392 VPWR.n2019 VGND 0.001572f
C6393 VPWR.n2020 VGND 0.00289f
C6394 VPWR.n2021 VGND 0.003474f
C6395 VPWR.n2022 VGND 0.001673f
C6396 VPWR.n2023 VGND 0.002447f
C6397 VPWR.n2024 VGND 0.001995f
C6398 VPWR.n2025 VGND 0.001014f
C6399 VPWR.t258 VGND 7.76e-19
C6400 VPWR.t270 VGND 7.48e-19
C6401 VPWR.n2026 VGND 0.001578f
C6402 VPWR.n2027 VGND 0.002819f
C6403 VPWR.n2028 VGND 5.49e-19
C6404 VPWR.n2029 VGND 6.25e-19
C6405 VPWR.n2030 VGND 0.001224f
C6406 VPWR.n2031 VGND 8.2e-19
C6407 VPWR.n2032 VGND 0.001463f
C6408 VPWR.n2033 VGND 6.56e-19
C6409 VPWR.n2034 VGND 8.2e-19
C6410 VPWR.n2035 VGND 8.78e-19
C6411 VPWR.n2036 VGND 0.001197f
C6412 VPWR.n2037 VGND 8.2e-19
C6413 VPWR.n2038 VGND 0.001281f
C6414 VPWR.n2039 VGND 0.001414f
C6415 VPWR.n2040 VGND 0.058516f
C6416 VPWR.n2041 VGND 0.048231f
C6417 VPWR.n2042 VGND 0.117032f
C6418 VPWR.n2043 VGND 0.117032f
C6419 VPWR.n2044 VGND 0.117032f
C6420 VPWR.n2045 VGND 0.221149f
C6421 VPWR.n2046 VGND 0.081008f
C6422 VPWR.n2047 VGND 0.001463f
C6423 VPWR.n2048 VGND 0.001092f
C6424 VPWR.n2049 VGND 6.56e-19
C6425 VPWR.n2050 VGND 6.56e-19
C6426 VPWR.n2051 VGND 8.2e-19
C6427 VPWR.n2052 VGND 0.001224f
C6428 VPWR.n2053 VGND 0.00634f
C6429 VPWR.t438 VGND 0.002279f
C6430 VPWR.t593 VGND 0.002071f
C6431 VPWR.n2054 VGND 0.004985f
C6432 VPWR.n2055 VGND 0.001597f
C6433 VPWR.t532 VGND 0.002088f
C6434 VPWR.t880 VGND 0.004432f
C6435 VPWR.n2057 VGND 0.011362f
C6436 VPWR.t533 VGND 0.002088f
C6437 VPWR.n2058 VGND 0.006189f
C6438 VPWR.n2059 VGND 0.001463f
C6439 VPWR.n2060 VGND 0.001835f
C6440 VPWR.n2061 VGND 0.00206f
C6441 VPWR.t547 VGND 0.002088f
C6442 VPWR.t853 VGND 0.004432f
C6443 VPWR.n2063 VGND 0.011362f
C6444 VPWR.t548 VGND 0.002088f
C6445 VPWR.n2064 VGND 0.006189f
C6446 VPWR.t564 VGND 0.002088f
C6447 VPWR.t870 VGND 0.004432f
C6448 VPWR.n2066 VGND 0.011362f
C6449 VPWR.t565 VGND 0.002088f
C6450 VPWR.n2067 VGND 0.006189f
C6451 VPWR.n2068 VGND 0.001597f
C6452 VPWR.t583 VGND 0.002088f
C6453 VPWR.t846 VGND 0.004432f
C6454 VPWR.n2070 VGND 0.011362f
C6455 VPWR.t584 VGND 0.002088f
C6456 VPWR.n2071 VGND 0.006189f
C6457 VPWR.n2072 VGND 0.005099f
C6458 VPWR.n2073 VGND 0.005594f
C6459 VPWR.n2074 VGND 0.001376f
C6460 VPWR.t857 VGND 0.015058f
C6461 VPWR.n2075 VGND 0.011361f
C6462 VPWR.n2076 VGND 0.010674f
C6463 VPWR.n2077 VGND 8.51e-19
C6464 VPWR.n2078 VGND 0.006622f
C6465 VPWR.n2079 VGND 0.00634f
C6466 VPWR.n2080 VGND 8.51e-19
C6467 VPWR.n2081 VGND 9.84e-19
C6468 VPWR.n2082 VGND 8.2e-19
C6469 VPWR.n2083 VGND 0.001281f
C6470 VPWR.n2084 VGND 0.001414f
C6471 VPWR.n2085 VGND 0.058516f
C6472 VPWR.n2086 VGND 0.001414f
C6473 VPWR.n2087 VGND 0.001281f
C6474 VPWR.n2088 VGND 8.8e-19
C6475 VPWR.n2089 VGND 0.00125f
C6476 VPWR.n2090 VGND 0.00634f
C6477 VPWR.n2091 VGND 0.008641f
C6478 VPWR.t594 VGND 0.002071f
C6479 VPWR.n2092 VGND 0.004756f
C6480 VPWR.n2093 VGND 0.008359f
C6481 VPWR.n2094 VGND 0.002447f
C6482 VPWR.n2095 VGND 0.00145f
C6483 VPWR.n2096 VGND 0.001835f
C6484 VPWR.n2097 VGND 0.002332f
C6485 VPWR.t567 VGND 0.002279f
C6486 VPWR.n2098 VGND 0.002879f
C6487 VPWR.n2099 VGND 0.005129f
C6488 VPWR.n2100 VGND 0.005129f
C6489 VPWR.n2101 VGND 0.002447f
C6490 VPWR.n2102 VGND 0.00145f
C6491 VPWR.n2103 VGND 0.001334f
C6492 VPWR.t869 VGND 0.030753f
C6493 VPWR.n2104 VGND 0.014263f
C6494 VPWR.n2105 VGND 0.001191f
C6495 VPWR.t411 VGND 0.002279f
C6496 VPWR.n2106 VGND 0.002879f
C6497 VPWR.n2107 VGND 0.005129f
C6498 VPWR.n2108 VGND 0.002447f
C6499 VPWR.n2109 VGND 0.002447f
C6500 VPWR.n2110 VGND 0.001888f
C6501 VPWR.n2111 VGND 0.004063f
C6502 VPWR.n2112 VGND 0.015206f
C6503 VPWR.n2113 VGND 0.00389f
C6504 VPWR.n2114 VGND 0.005129f
C6505 VPWR.n2115 VGND 0.005302f
C6506 VPWR.n2116 VGND 8.51e-19
C6507 VPWR.n2117 VGND 6.56e-19
C6508 VPWR.n2118 VGND 8.2e-19
C6509 VPWR.n2119 VGND 9.31e-19
C6510 VPWR.n2120 VGND 0.001144f
C6511 VPWR.n2121 VGND 8.2e-19
C6512 VPWR.n2122 VGND 0.001281f
C6513 VPWR.n2123 VGND 0.001414f
C6514 VPWR.n2124 VGND 0.058516f
C6515 VPWR.n2125 VGND 0.001414f
C6516 VPWR.n2126 VGND 0.001281f
C6517 VPWR.n2127 VGND 0.001225f
C6518 VPWR.n2128 VGND 0.001051f
C6519 VPWR.n2129 VGND 0.002501f
C6520 VPWR.n2130 VGND 0.006627f
C6521 VPWR.n2131 VGND 0.001317f
C6522 VPWR.n2132 VGND 0.002058f
C6523 VPWR.n2133 VGND 0.004023f
C6524 VPWR.n2134 VGND 0.005626f
C6525 VPWR.t497 VGND 0.002071f
C6526 VPWR.n2135 VGND 0.012426f
C6527 VPWR.t897 VGND 0.007283f
C6528 VPWR.n2136 VGND 0.014117f
C6529 VPWR.n2137 VGND 0.003221f
C6530 VPWR.n2138 VGND 7.21e-19
C6531 VPWR.n2139 VGND 0.004098f
C6532 VPWR.n2140 VGND 0.002221f
C6533 VPWR.n2141 VGND 0.002447f
C6534 VPWR.n2142 VGND 0.008359f
C6535 VPWR.n2143 VGND 0.008641f
C6536 VPWR.t906 VGND 0.030181f
C6537 VPWR.t498 VGND 0.002071f
C6538 VPWR.n2144 VGND 0.002455f
C6539 VPWR.n2145 VGND 0.016594f
C6540 VPWR.n2146 VGND 0.006622f
C6541 VPWR.n2147 VGND 0.002447f
C6542 VPWR.n2148 VGND 0.00145f
C6543 VPWR.n2149 VGND 0.001702f
C6544 VPWR.n2150 VGND 0.002332f
C6545 VPWR.t680 VGND 0.002279f
C6546 VPWR.n2151 VGND 0.002879f
C6547 VPWR.n2152 VGND 0.005129f
C6548 VPWR.n2153 VGND 8.51e-19
C6549 VPWR.n2154 VGND 6.56e-19
C6550 VPWR.n2155 VGND 8.2e-19
C6551 VPWR.n2156 VGND 0.001197f
C6552 VPWR.n2157 VGND 8.51e-19
C6553 VPWR.n2158 VGND 0.001224f
C6554 VPWR.n2159 VGND 8.2e-19
C6555 VPWR.n2160 VGND 0.001281f
C6556 VPWR.n2161 VGND 0.001414f
C6557 VPWR.n2162 VGND 0.058516f
C6558 VPWR.n2163 VGND 0.001414f
C6559 VPWR.n2164 VGND 0.001281f
C6560 VPWR.n2165 VGND 0.001225f
C6561 VPWR.n2166 VGND 8.51e-19
C6562 VPWR.n2167 VGND 0.004063f
C6563 VPWR.n2168 VGND 0.015206f
C6564 VPWR.n2169 VGND 0.00389f
C6565 VPWR.n2170 VGND 0.005129f
C6566 VPWR.n2171 VGND 0.002447f
C6567 VPWR.n2172 VGND 0.00145f
C6568 VPWR.n2173 VGND 0.002412f
C6569 VPWR.n2174 VGND 0.002392f
C6570 VPWR.n2175 VGND 0.002221f
C6571 VPWR.n2176 VGND 0.002447f
C6572 VPWR.n2177 VGND 0.005129f
C6573 VPWR.n2178 VGND 0.005302f
C6574 VPWR.t840 VGND 0.030181f
C6575 VPWR.n2179 VGND 0.015033f
C6576 VPWR.n2180 VGND 0.004063f
C6577 VPWR.n2181 VGND 0.002447f
C6578 VPWR.n2182 VGND 0.00145f
C6579 VPWR.n2183 VGND 0.002412f
C6580 VPWR.n2184 VGND 0.002392f
C6581 VPWR.t581 VGND 0.002279f
C6582 VPWR.n2185 VGND 0.002879f
C6583 VPWR.n2186 VGND 0.005129f
C6584 VPWR.n2187 VGND 0.002447f
C6585 VPWR.n2188 VGND 0.002447f
C6586 VPWR.n2189 VGND 0.001516f
C6587 VPWR.n2190 VGND 0.004063f
C6588 VPWR.n2191 VGND 0.015206f
C6589 VPWR.n2192 VGND 0.002501f
C6590 VPWR.t606 VGND 0.002279f
C6591 VPWR.n2193 VGND 0.002879f
C6592 VPWR.n2194 VGND 0.001224f
C6593 VPWR.n2195 VGND 8.51e-19
C6594 VPWR.n2196 VGND 0.005129f
C6595 VPWR.n2197 VGND 0.00389f
C6596 VPWR.n2198 VGND 8.51e-19
C6597 VPWR.n2199 VGND 9.31e-19
C6598 VPWR.n2200 VGND 8.2e-19
C6599 VPWR.n2201 VGND 0.001281f
C6600 VPWR.n2202 VGND 0.001414f
C6601 VPWR.n2203 VGND 0.058516f
C6602 VPWR.n2204 VGND 0.001414f
C6603 VPWR.n2205 VGND 0.001281f
C6604 VPWR.n2206 VGND 2.28e-19
C6605 VPWR.n2207 VGND 0.001317f
C6606 VPWR.n2208 VGND 0.001835f
C6607 VPWR.n2209 VGND 0.00372f
C6608 VPWR.t596 VGND 0.002071f
C6609 VPWR.n2210 VGND 0.002596f
C6610 VPWR.n2211 VGND 0.008854f
C6611 VPWR.n2212 VGND 0.006481f
C6612 VPWR.n2213 VGND 0.008359f
C6613 VPWR.n2214 VGND 0.002447f
C6614 VPWR.n2215 VGND 0.00145f
C6615 VPWR.n2216 VGND 0.00306f
C6616 VPWR.n2217 VGND 0.005055f
C6617 VPWR.n2218 VGND 8.38e-19
C6618 VPWR.n2219 VGND 0.002221f
C6619 VPWR.n2220 VGND 0.001436f
C6620 VPWR.n2221 VGND 6.88e-19
C6621 VPWR.n2222 VGND 0.00185f
C6622 VPWR.n2223 VGND 6.12e-20
C6623 VPWR.n2224 VGND 0.002277f
C6624 VPWR.n2225 VGND 6.83e-19
C6625 VPWR.n2226 VGND 0.002447f
C6626 VPWR.n2227 VGND 0.001942f
C6627 VPWR.n2228 VGND 0.001225f
C6628 VPWR.n2229 VGND 0.001414f
C6629 VPWR.n2230 VGND 0.001281f
C6630 VPWR.n2231 VGND 8.2e-19
C6631 VPWR.n2232 VGND 3.86e-19
C6632 VPWR.n2233 VGND 7.11e-19
C6633 VPWR.t394 VGND 0.001157f
C6634 VPWR.t689 VGND 5.61e-19
C6635 VPWR.n2234 VGND 0.002356f
C6636 VPWR.n2235 VGND 0.001803f
C6637 VPWR.n2236 VGND 6.64e-19
C6638 VPWR.n2237 VGND 8.51e-19
C6639 VPWR.n2238 VGND 6.12e-19
C6640 VPWR.n2239 VGND 8.2e-19
C6641 VPWR.n2240 VGND 6.56e-19
C6642 VPWR.n2241 VGND 0.001463f
C6643 VPWR.n2242 VGND 0.001414f
C6644 VPWR.n2243 VGND 0.001281f
C6645 VPWR.n2244 VGND 0.001225f
C6646 VPWR.n2245 VGND 8.51e-19
C6647 VPWR.n2246 VGND 4.62e-19
C6648 VPWR.n2247 VGND 8.67e-19
C6649 VPWR.n2248 VGND 0.006875f
C6650 VPWR.n2249 VGND 0.002021f
C6651 VPWR.n2250 VGND 9.31e-19
C6652 VPWR.n2251 VGND 0.002591f
C6653 VPWR.t850 VGND 0.015539f
C6654 VPWR.n2252 VGND 0.026019f
C6655 VPWR.t570 VGND 0.002071f
C6656 VPWR.n2253 VGND 0.005332f
C6657 VPWR.n2254 VGND 0.007114f
C6658 VPWR.n2255 VGND 8.38e-19
C6659 VPWR.n2256 VGND 0.002221f
C6660 VPWR.n2257 VGND 0.005202f
C6661 VPWR.n2258 VGND 0.004143f
C6662 VPWR.n2259 VGND 0.003282f
C6663 VPWR.t571 VGND 0.002071f
C6664 VPWR.n2260 VGND 0.003648f
C6665 VPWR.n2261 VGND 0.006214f
C6666 VPWR.n2262 VGND 0.001835f
C6667 VPWR.n2263 VGND 3.06e-19
C6668 VPWR.n2264 VGND 6.14e-19
C6669 VPWR.n2265 VGND 0.001281f
C6670 VPWR.n2266 VGND 6.56e-19
C6671 VPWR.n2267 VGND 8.2e-19
C6672 VPWR.n2268 VGND 6.12e-19
C6673 VPWR.n2269 VGND 0.001224f
C6674 VPWR.n2270 VGND 8.51e-19
C6675 VPWR.t467 VGND 0.002088f
C6676 VPWR.t890 VGND 0.004432f
C6677 VPWR.n2272 VGND 0.011362f
C6678 VPWR.t468 VGND 0.002088f
C6679 VPWR.n2273 VGND 0.006189f
C6680 VPWR.n2274 VGND 0.005217f
C6681 VPWR.n2275 VGND 5.72e-19
C6682 VPWR.n2276 VGND 0.001199f
C6683 VPWR.n2277 VGND 8.78e-19
C6684 VPWR.n2278 VGND 8.2e-19
C6685 VPWR.n2279 VGND 6.56e-19
C6686 VPWR.n2280 VGND 0.001463f
C6687 VPWR.n2281 VGND 0.001414f
C6688 VPWR.n2282 VGND 0.058516f
C6689 VPWR.n2283 VGND 0.048231f
C6690 VPWR.n2284 VGND 0.06951f
C6691 VPWR.n2285 VGND 0.117032f
C6692 VPWR.n2286 VGND 0.048231f
C6693 VPWR.n2287 VGND 0.058516f
C6694 VPWR.n2288 VGND 0.001414f
C6695 VPWR.n2289 VGND 0.001281f
C6696 VPWR.n2290 VGND 0.001225f
C6697 VPWR.n2291 VGND 0.001942f
C6698 VPWR.n2292 VGND 0.003084f
C6699 VPWR.n2293 VGND 0.003084f
C6700 VPWR.n2294 VGND 0.001659f
C6701 VPWR.n2295 VGND 0.002447f
C6702 VPWR.n2296 VGND 0.002447f
C6703 VPWR.n2297 VGND 0.002221f
C6704 VPWR.n2298 VGND 0.001576f
C6705 VPWR.n2299 VGND 0.002521f
C6706 VPWR.n2300 VGND 0.014064f
C6707 VPWR.n2301 VGND 0.001877f
C6708 VPWR.n2302 VGND 8.38e-19
C6709 VPWR.n2303 VGND 0.002538f
C6710 VPWR.n2304 VGND 8.38e-19
C6711 VPWR.n2305 VGND 9.56e-19
C6712 VPWR.n2306 VGND 0.002601f
C6713 VPWR.n2307 VGND 0.006627f
C6714 VPWR.n2308 VGND 0.001317f
C6715 VPWR.n2309 VGND 2.28e-19
C6716 VPWR.n2310 VGND 0.001281f
C6717 VPWR.n2311 VGND 8.2e-19
C6718 VPWR.n2312 VGND 0.001224f
C6719 VPWR.n2313 VGND 8.51e-19
C6720 VPWR.n2314 VGND 0.005129f
C6721 VPWR.n2315 VGND 0.005302f
C6722 VPWR.n2316 VGND 8.51e-19
C6723 VPWR.n2317 VGND 9.31e-19
C6724 VPWR.n2318 VGND 8.2e-19
C6725 VPWR.n2319 VGND 0.001281f
C6726 VPWR.n2320 VGND 0.001414f
C6727 VPWR.n2321 VGND 0.058516f
C6728 VPWR.n2322 VGND 0.048231f
C6729 VPWR.n2323 VGND 0.117032f
C6730 VPWR.n2324 VGND 0.117032f
C6731 VPWR.n2325 VGND 0.048231f
C6732 VPWR.n2326 VGND 0.064545f
C6733 VPWR.n2327 VGND 0.001414f
C6734 VPWR.n2328 VGND 0.001463f
C6735 VPWR.n2329 VGND 6.56e-19
C6736 VPWR.n2330 VGND 8.2e-19
C6737 VPWR.n2331 VGND 0.001224f
C6738 VPWR.n2332 VGND 8.51e-19
C6739 VPWR.n2333 VGND 0.005302f
C6740 VPWR.n2334 VGND 0.005302f
C6741 VPWR.n2335 VGND 0.00389f
C6742 VPWR.n2336 VGND 0.002447f
C6743 VPWR.n2337 VGND 0.002447f
C6744 VPWR.n2338 VGND 0.002447f
C6745 VPWR.n2339 VGND 0.005302f
C6746 VPWR.n2340 VGND 0.005129f
C6747 VPWR.t447 VGND 0.002279f
C6748 VPWR.n2341 VGND 0.003107f
C6749 VPWR.n2342 VGND 0.001839f
C6750 VPWR.n2343 VGND 0.001835f
C6751 VPWR.n2344 VGND 0.002058f
C6752 clknet_0_clk.t38 VGND 0.015823f
C6753 clknet_0_clk.t47 VGND 0.0074f
C6754 clknet_0_clk.t40 VGND 0.015823f
C6755 clknet_0_clk.t32 VGND 0.0074f
C6756 clknet_0_clk.t36 VGND 0.015823f
C6757 clknet_0_clk.t44 VGND 0.0074f
C6758 clknet_0_clk.t42 VGND 0.015823f
C6759 clknet_0_clk.t34 VGND 0.0074f
C6760 clknet_0_clk.n0 VGND 0.036121f
C6761 clknet_0_clk.n1 VGND 0.047576f
C6762 clknet_0_clk.n2 VGND 0.047576f
C6763 clknet_0_clk.n3 VGND 0.057784f
C6764 clknet_0_clk.n4 VGND 0.075138f
C6765 clknet_0_clk.t45 VGND 0.015823f
C6766 clknet_0_clk.t37 VGND 0.0074f
C6767 clknet_0_clk.t33 VGND 0.015823f
C6768 clknet_0_clk.t41 VGND 0.0074f
C6769 clknet_0_clk.t43 VGND 0.015823f
C6770 clknet_0_clk.t35 VGND 0.0074f
C6771 clknet_0_clk.t46 VGND 0.015823f
C6772 clknet_0_clk.t39 VGND 0.0074f
C6773 clknet_0_clk.n5 VGND 0.036121f
C6774 clknet_0_clk.n6 VGND 0.047576f
C6775 clknet_0_clk.n7 VGND 0.047576f
C6776 clknet_0_clk.n8 VGND 0.057941f
C6777 clknet_0_clk.n9 VGND 0.038186f
C6778 clknet_0_clk.t15 VGND 0.01123f
C6779 clknet_0_clk.t2 VGND 0.01123f
C6780 clknet_0_clk.n10 VGND 0.028528f
C6781 clknet_0_clk.t13 VGND 0.01123f
C6782 clknet_0_clk.t8 VGND 0.01123f
C6783 clknet_0_clk.n11 VGND 0.023672f
C6784 clknet_0_clk.n12 VGND 0.107879f
C6785 clknet_0_clk.t1 VGND 0.01123f
C6786 clknet_0_clk.t3 VGND 0.01123f
C6787 clknet_0_clk.n13 VGND 0.023672f
C6788 clknet_0_clk.n14 VGND 0.062143f
C6789 clknet_0_clk.t14 VGND 0.01123f
C6790 clknet_0_clk.t9 VGND 0.01123f
C6791 clknet_0_clk.n15 VGND 0.023672f
C6792 clknet_0_clk.n16 VGND 0.061854f
C6793 clknet_0_clk.t11 VGND 0.01123f
C6794 clknet_0_clk.t4 VGND 0.01123f
C6795 clknet_0_clk.n17 VGND 0.023672f
C6796 clknet_0_clk.n18 VGND 0.061854f
C6797 clknet_0_clk.t6 VGND 0.01123f
C6798 clknet_0_clk.t10 VGND 0.01123f
C6799 clknet_0_clk.n19 VGND 0.023672f
C6800 clknet_0_clk.n20 VGND 0.062143f
C6801 clknet_0_clk.t12 VGND 0.01123f
C6802 clknet_0_clk.t5 VGND 0.01123f
C6803 clknet_0_clk.n21 VGND 0.023672f
C6804 clknet_0_clk.n22 VGND 0.053374f
C6805 clknet_0_clk.t7 VGND 0.01123f
C6806 clknet_0_clk.t0 VGND 0.01123f
C6807 clknet_0_clk.n23 VGND 0.023364f
C6808 clknet_0_clk.n24 VGND 0.073498f
C6809 clknet_0_clk.t18 VGND 0.004717f
C6810 clknet_0_clk.t20 VGND 0.004717f
C6811 clknet_0_clk.n25 VGND 0.010394f
C6812 clknet_0_clk.n26 VGND 0.034156f
C6813 clknet_0_clk.t30 VGND 0.004717f
C6814 clknet_0_clk.t16 VGND 0.004717f
C6815 clknet_0_clk.n27 VGND 0.010767f
C6816 clknet_0_clk.n28 VGND 0.035304f
C6817 clknet_0_clk.t26 VGND 0.004717f
C6818 clknet_0_clk.t22 VGND 0.004717f
C6819 clknet_0_clk.n29 VGND 0.016749f
C6820 clknet_0_clk.t24 VGND 0.004717f
C6821 clknet_0_clk.t19 VGND 0.004717f
C6822 clknet_0_clk.n30 VGND 0.010767f
C6823 clknet_0_clk.n31 VGND 0.068037f
C6824 clknet_0_clk.t21 VGND 0.004717f
C6825 clknet_0_clk.t23 VGND 0.004717f
C6826 clknet_0_clk.n32 VGND 0.010767f
C6827 clknet_0_clk.n33 VGND 0.040895f
C6828 clknet_0_clk.t25 VGND 0.004717f
C6829 clknet_0_clk.t27 VGND 0.004717f
C6830 clknet_0_clk.n34 VGND 0.010774f
C6831 clknet_0_clk.n35 VGND 0.042184f
C6832 clknet_0_clk.t29 VGND 0.004717f
C6833 clknet_0_clk.t31 VGND 0.004717f
C6834 clknet_0_clk.n36 VGND 0.010767f
C6835 clknet_0_clk.n37 VGND 0.040895f
C6836 clknet_0_clk.n38 VGND 0.026375f
C6837 clknet_0_clk.t17 VGND 0.004717f
C6838 clknet_0_clk.t28 VGND 0.004717f
C6839 clknet_0_clk.n39 VGND 0.009573f
C6840 clknet_0_clk.n40 VGND 0.015919f
C6841 clknet_0_clk.n41 VGND 0.145873f
.ends

