** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tb_anamux.sch
**.subckt tb_anamux
x1 net1 net2 net3 net4 net5 net6 net7 net8 net9 net10 net11 net12 net13 net14 net15 net16 net17 net18 net19 net20 net21 net22
+ net23 net24 net25 net26 net27 net28 net29 net30 net31 net32 net33 net34 net35 net36 net37 net38 net39 net40 EN_COUNTER VRES LADOUTPX
+ RSEL1 RINGOUTPX SEL1 RSEL2 EN_RING RSEL0 MUXOUTPX SEL0 VCC VSS tt_um_patdeegan_anamux_parax
R6 RINGOUTPX VSS 100k m=1
R1 MUXOUTPX VSS 100k m=1
R2 LADOUTPX VSS 100k m=1
R3 RINGOUT VSS 100k m=1
R4 MUXOUT VSS 100k m=1
R5 LADOUT VSS 100k m=1
x2 net41 net42 net43 VRES RINGOUT MUXOUT LADOUT net44 net45 net46 net47 RSEL0 RSEL1 RSEL2 SEL0 SEL1 EN_COUNTER EN_RING net48 net49
+ net50 net51 net52 net53 net54 net55 net56 net57 net58 net59 net60 net61 net62 net63 net64 net65 net66 net67 net68 net69 net70 net71
+ net72 net73 net74 net75 net76 net77 net78 net79 net80 VCC VSS tt_um_patdeegan_anamux
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  tt_um_patdeegan_anamux.sym # of pins=53
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sch
.subckt tt_um_patdeegan_anamux clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VSS
*.ipin ena
*.ipin clk
*.ipin rst_n
*.iopin ua[4]
*.iopin ua[5]
*.iopin ua[6]
*.ipin ui_in[7]
*.ipin uio_in[0]
*.ipin uio_in[1]
*.ipin uio_in[2]
*.ipin uio_in[3]
*.ipin uio_in[4]
*.ipin uio_in[5]
*.ipin uio_in[6]
*.ipin uio_in[7]
*.opin uio_oe[0]
*.opin uio_oe[1]
*.opin uio_oe[2]
*.opin uio_oe[3]
*.opin uio_oe[4]
*.opin uio_oe[5]
*.opin uio_oe[6]
*.opin uio_oe[7]
*.iopin uio_out[0]
*.iopin uio_out[1]
*.iopin uio_out[2]
*.iopin uio_out[3]
*.iopin uio_out[4]
*.iopin uio_out[5]
*.iopin uio_out[6]
*.iopin uio_out[7]
*.opin uo_out[0]
*.opin uo_out[1]
*.opin uo_out[2]
*.opin uo_out[3]
*.opin uo_out[4]
*.opin uo_out[5]
*.opin uo_out[6]
*.opin uo_out[7]
*.ipin ui_in[0]
*.ipin ui_in[1]
*.ipin ui_in[2]
*.ipin ui_in[3]
*.ipin ui_in[4]
*.ipin ui_in[5]
*.ipin ui_in[6]
*.iopin ua[0]
*.iopin ua[1]
*.iopin ua[2]
*.iopin ua[3]
*.ipin VSS
*.ipin VDPWR
*.iopin ua[7]
x1 ua[0] ui_in[3] VDPWR ui_in[4] ua[1] VSS ui_in[0] ui_in[1] ua[2] ui_in[2] ua[3] ui_in[6] ui_in[5] fulltest_userarea
.ends


* expanding   symbol:  tt_um_patdeegan_anamux_parax.sym # of pins=53
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sym
.include /home/ttuser/vmswap/tt09-analogmux/xschem/extracted/tt_um_patdeegan_anamux_parax.spice

* expanding   symbol:  fulltest_userarea.sym # of pins=13
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sch
.subckt fulltest_userarea VRES select0 VDD select1 ring_out VSS rsel0 rsel1 muxtest_out rsel2 ladderout enable_ring enable_counter
*.ipin VDD
*.ipin VSS
*.ipin select0
*.ipin select1
*.ipin rsel0
*.ipin rsel1
*.ipin rsel2
*.ipin enable_ring
*.ipin enable_counter
*.opin ring_out
*.opin muxtest_out
*.opin ladderout
*.ipin VRES
x1 VSS VDD select0 select1 VRES rsel0 rsel1 rsel2 muxtest_out ladderout muxtest
x2 VDD VSS enable_ring select0 select1 enable_counter ring_out ringtest
.ends


* expanding   symbol:  muxtest.sym # of pins=10
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sch
.subckt muxtest VSS VDD SELECT0 SELECT1 VRES RSEL0 RSEL1 RSEL2 OUT LADDEROUT
*.ipin VSS
*.ipin VDD
*.ipin SELECT0
*.ipin SELECT1
*.ipin VRES
*.ipin RSEL0
*.ipin RSEL1
*.ipin RSEL2
*.opin OUT
*.opin LADDEROUT
x1 RSEL0 RSEL1 RSEL2 A1 A2 A3 A4 A5 A6 A7 VRES LADDEROUT VDD VSS mux8onehot
x2 SELECT0 SELECT1 VDD LADDEROUT VRES A5 A1 OUT OUT OUT OUT net1 VDD VSS mux4onehot_b
XR1 A7 VRES VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR2 A6 A7 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR3 A5 A6 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR4 A4 A5 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR5 A3 A4 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR6 A2 A3 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR7 A1 A2 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR8 VSS A1 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
.ends


* expanding   symbol:  ringtest.sym # of pins=7
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sch
.subckt ringtest VDD VSS enable_ring select0 select1 enable_counter mux_out
*.ipin VDD
*.ipin VSS
*.ipin enable_ring
*.ipin select0
*.ipin select1
*.ipin enable_counter
*.opin mux_out
x3 select0 select1 VDD ring_out drv_out counter3 counter7 mux_out mux_out mux_out mux_out net1 VDD VSS mux4onehot_b
x4 VSS VDD drv_out enable_counter net2 net3 counter7 net4 net5 net6 counter3 net7 net8 net9 simplecounter
x1 VDD VSS enable_ring ring_out ring
x2 VDD VSS ring_out drv_out driver
.ends


* expanding   symbol:  mux8onehot.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sch
.subckt mux8onehot select0 select1 select2 A1 A2 A3 A4 A5 A6 A7 A8 Z VDD VSS
*.ipin select0
*.ipin select1
*.ipin select2
*.ipin VDD
*.ipin VSS
*.iopin Z
*.iopin A1
*.iopin A2
*.iopin A3
*.iopin A4
*.iopin A5
*.iopin A6
*.iopin A7
*.iopin A8
x4 OUT_HIGH select2 nSEL2 Z VDD VSS passgate
x5 OUT_LOW nSEL2 select2 Z VDD VSS passgate
x2 A1 gno0 gpo0 OUT_LOW A2 gno1 gpo1 OUT_LOW A3 gno2 gpo2 OUT_LOW A4 gno3 gpo3 OUT_LOW VDD VSS passgatex4
x1 select0 select1 select2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nSEL2 VDD VSS passgatesCtrlManual
x3 A5 gno0 gpo0 OUT_HIGH A6 gno1 gpo1 OUT_HIGH A7 gno2 gpo2 OUT_HIGH A8 gno3 gpo3 OUT_HIGH VDD VSS passgatex4
.ends


* expanding   symbol:  mux4onehot_b.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sch
.subckt mux4onehot_b select0 select1 select2 A1 A2 A3 A4 Z1 Z2 Z3 Z4 nselect2 VDD VSS
*.ipin select0
*.ipin select1
*.ipin select2
*.iopin A1
*.iopin A2
*.iopin A3
*.iopin A4
*.iopin Z1
*.iopin Z2
*.iopin Z3
*.iopin Z4
*.opin nselect2
*.ipin VDD
*.ipin VSS
x2 A1 gno0 gpo0 Z1 A2 gno1 gpo1 Z2 A3 gno2 gpo2 Z3 A4 gno3 gpo3 Z4 VDD VSS passgatex4
x1 select0 select1 select2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nselect2 VDD VSS passgatesCtrlManual
.ends


* expanding   symbol:  ring.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ring.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ring.sch
.subckt ring VDD VSS enable out
*.iopin VDD
*.ipin enable
*.iopin VSS
*.opin out
x2 enable net18 VSS VSS VDD VDD out sky130_fd_sc_hd__nand2_2
x1 VDD VSS out net1 inverter
x3 VDD VSS net1 net2 inverter
x4 VDD VSS net2 net3 inverter
x5 VDD VSS net3 net4 inverter
x6 VDD VSS net4 net5 inverter
x7 VDD VSS net5 net6 inverter
x8 VDD VSS net6 net7 inverter
x9 VDD VSS net7 net8 inverter
x10 VDD VSS net8 net9 inverter
x11 VDD VSS net9 net10 inverter
x12 VDD VSS net10 net11 inverter
x13 VDD VSS net11 net12 inverter
x14 VDD VSS net12 net13 inverter
x15 VDD VSS net13 net14 inverter
x16 VDD VSS net14 net15 inverter
x17 VDD VSS net15 net16 inverter
x18 VDD VSS net16 net17 inverter
x19 VDD VSS net17 net18 inverter
.ends


* expanding   symbol:  driver.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/driver.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/driver.sch
.subckt driver VDD VSS in out
*.iopin VDD
*.iopin VSS
*.opin out
*.ipin in
XM9 net1 in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net1 in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=72 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=24 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  passgate.sym # of pins=6
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sch
.subckt passgate A GN GP Z VDD VSS
*.ipin GN
*.ipin VDD
*.ipin VSS
*.ipin GP
*.iopin A
*.iopin Z
XM1 Z GN A VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 Z GP A VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  passgatex4.sym # of pins=18
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sch
.subckt passgatex4 A1 GN1 GP1 Z1 A2 GN2 GP2 Z2 A3 GN3 GP3 Z3 A4 GN4 GP4 Z4 VDD VSS
*.ipin VDD
*.ipin VSS
*.ipin GP1
*.ipin GN1
*.iopin A1
*.iopin Z1
*.ipin GP2
*.ipin GN2
*.iopin A2
*.iopin Z2
*.ipin GP3
*.ipin GN3
*.iopin A3
*.iopin Z3
*.ipin GP4
*.ipin GN4
*.iopin A4
*.iopin Z4
x1 A1 GN1 GP1 Z1 VDD VSS passgate
x2 A2 GN2 GP2 Z2 VDD VSS passgate
x3 A3 GN3 GP3 Z3 VDD VSS passgate
x4 A4 GN4 GP4 Z4 VDD VSS passgate
.ends


* expanding   symbol:  passgatesCtrlManual.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sch
.subckt passgatesCtrlManual SEL0 SEL1 SEL2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nSEL2 VPWR VGND
*.ipin SEL0
*.ipin SEL1
*.ipin SEL2
*.opin gno0
*.opin gpo0
*.opin gno1
*.opin gpo1
*.opin gno2
*.opin gpo2
*.opin gno3
*.opin gpo3
*.opin nSEL2
*.ipin VPWR
*.ipin VGND
x1 SEL0 VGND VGND VPWR VPWR nSEL0 sky130_fd_sc_hd__inv_2
x2 SEL1 VGND VGND VPWR VPWR nSEL1 sky130_fd_sc_hd__inv_2
x7 nSEL0 nSEL1 VGND VGND VPWR VPWR gno0 sky130_fd_sc_hd__and2_1
x10 SEL1 SEL0 VGND VGND VPWR VPWR gno3 sky130_fd_sc_hd__and2_1
x11 gno0 VGND VGND VPWR VPWR gpo0 sky130_fd_sc_hd__inv_2
x12 gno1 VGND VGND VPWR VPWR gpo1 sky130_fd_sc_hd__inv_2
x13 gno2 VGND VGND VPWR VPWR gpo2 sky130_fd_sc_hd__inv_2
x14 gno3 VGND VGND VPWR VPWR gpo3 sky130_fd_sc_hd__inv_2
x15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x8 SEL1 SEL0 VGND VGND VPWR VPWR gno1 sky130_fd_sc_hd__and2b_1
x9 SEL0 SEL1 VGND VGND VPWR VPWR gno2 sky130_fd_sc_hd__and2b_1
x18 SEL2 VGND VGND VPWR VPWR nSEL2 sky130_fd_sc_hd__inv_2
x19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/inverter.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/inverter.sch
.subckt inverter VDD VSS in out
*.opin out
*.iopin VDD
*.iopin VSS
*.ipin in
x1 in VSS VSS VDD VDD out sky130_fd_sc_hd__inv_2
.ends

**** begin user architecture code


* ngspice commands
* .options savecurrents

.param VCC = 1.8
.param SRCRES = 1k
* need this for matt's weird inverter and add
.include /home/ttuser/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
* don't want to deal with verilog, so:
.include ../extracted/simplecounter_parax.spice
.include stimuli_tb_anamux.cir
.control
save all
* op
* write tb_anamux.raw
* set appendwrite
tran 1n 185n uic
write tb_anamux.raw
* quit 0
.endc



**** end user architecture code
.end
