magic
tech sky130A
magscale 1 2
timestamp 1725652981
<< metal1 >>
rect 2810 -336 2820 -204
rect 2928 -336 2938 -204
rect 3892 -328 3902 -198
rect 4010 -328 4020 -198
rect 4910 -336 4920 -194
rect 5022 -336 5032 -194
rect 6012 -318 6022 -184
rect 6094 -318 6104 -184
<< via1 >>
rect 2820 -336 2928 -204
rect 3902 -328 4010 -198
rect 4920 -336 5022 -194
rect 6022 -318 6094 -184
<< metal2 >>
rect 568 1134 6082 1190
rect 758 889 814 892
rect 758 839 5825 889
rect 758 198 814 839
rect 1310 632 4994 688
rect 1310 -722 1366 632
rect 1472 426 4760 482
rect 1472 -1586 1528 426
rect 1284 -1642 1528 -1586
rect 1684 202 3982 258
rect 1684 -2506 1740 202
rect 1292 -2562 1740 -2506
rect 1838 72 3716 128
rect 1838 -3426 1894 72
rect 1306 -3482 1894 -3426
rect 1964 -84 2902 -28
rect 1964 -4346 2020 -84
rect 1272 -4402 2020 -4346
rect 2097 -198 2687 -139
rect 2846 -194 2902 -84
rect 2097 -5266 2156 -198
rect 2578 -272 2687 -198
rect 2628 -278 2687 -272
rect 2575 -337 2687 -278
rect 2820 -204 2928 -194
rect 3660 -334 3716 72
rect 3926 -188 3982 202
rect 3902 -198 4010 -188
rect 4704 -322 4760 426
rect 4938 -184 4994 632
rect 4920 -194 5022 -184
rect 2820 -346 2928 -336
rect 3902 -338 4010 -328
rect 5775 -303 5825 839
rect 6026 -174 6082 1134
rect 6022 -184 6094 -174
rect 6022 -328 6094 -318
rect 4920 -346 5022 -336
rect 1278 -5322 2156 -5266
rect 2097 -5323 2156 -5322
use passgatesdigital  passgatesdigital_0
timestamp 1725652498
transform 0 -1 2512 1 0 -6078
box 750 1142 7254 6332
use passgatex4  passgatex4_0
timestamp 1725644236
transform 1 0 -9124 0 1 -4842
box 11366 -356 15589 4682
<< end >>
