* NGSPICE file created from tt_um_patdeegan_anamux.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.102877 pd=0.95413 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.244946 ps=2.271739 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.087768 pd=0.816449 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.102877 ps=0.95413 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.135832 ps=1.263551 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111244 pd=0.929204 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.264867 ps=2.212389 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13602 ps=1.457047 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.111244 ps=0.929204 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111244 pd=0.929204 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08789 pd=0.941476 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08789 ps=0.941476 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=1.05
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.05
**devattr d=5720,324
.ends

.subckt passgatesCtrlManual SEL0 SEL1 SEL2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3
+ nSEL2 VPWR VGND
Xx1 SEL0 VGND VGND VPWR VPWR nSEL0 sky130_fd_sc_hd__inv_2
Xx2 SEL1 VGND VGND VPWR VPWR nSEL1 sky130_fd_sc_hd__inv_2
Xx7 nSEL0 nSEL1 VGND VGND VPWR VPWR gno0 sky130_fd_sc_hd__and2_1
Xx8 SEL1 SEL0 VGND VGND VPWR VPWR gno1 sky130_fd_sc_hd__and2b_1
Xx9 SEL0 SEL1 VGND VGND VPWR VPWR gno2 sky130_fd_sc_hd__and2b_1
Xx10 SEL1 SEL0 VGND VGND VPWR VPWR gno3 sky130_fd_sc_hd__and2_1
Xx11 gno0 VGND VGND VPWR VPWR gpo0 sky130_fd_sc_hd__inv_2
Xx12 gno1 VGND VGND VPWR VPWR gpo1 sky130_fd_sc_hd__inv_2
Xx13 gno2 VGND VGND VPWR VPWR gpo2 sky130_fd_sc_hd__inv_2
Xx15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xx14 gno3 VGND VGND VPWR VPWR gpo3 sky130_fd_sc_hd__inv_2
Xx16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xx17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xx18 SEL2 VGND VGND VPWR VPWR nSEL2 sky130_fd_sc_hd__inv_2
Xx19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_PEJ72P a_n35_21# a_35_109# a_n195_n1883# a_n35_n1797#
+ a_n93_n1709# a_n93_109# a_35_n1709#
X0 a_35_n1709# a_n35_n1797# a_n93_n1709# a_n195_n1883# sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
X1 a_35_109# a_n35_21# a_n93_109# a_n195_n1883# sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
**devattr s=92800,3316 d=92800,3316
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4QFMR3 a_n35_21# a_n93_118# a_n35_n2215# a_n93_n2118#
+ a_35_118# a_35_n2118# w_n231_n2337#
X0 a_35_n2118# a_n35_n2215# a_n93_n2118# w_n231_n2337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
X1 a_35_118# a_n35_21# a_n93_118# w_n231_n2337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
**devattr s=116000,4116 d=116000,4116
.ends

.subckt passgate A GN GP Z VSS VDD
XXM1 GN Z VSS GN A A Z sky130_fd_pr__nfet_01v8_lvt_PEJ72P
XXM3 GP Z GP Z A A VDD sky130_fd_pr__pfet_01v8_lvt_4QFMR3
.ends

.subckt passgatex4 A1 GN1 A2 GN2 GP2 Z2 A3 GN3 GP3 Z3 A4 GN4 GP4 Z4 GP1 Z1 VSS VDD
Xx1 A1 GN1 GP1 Z1 VSS VDD passgate
Xx2 A2 GN2 GP2 Z2 VSS VDD passgate
Xx3 A3 GN3 GP3 Z3 VSS VDD passgate
Xx4 A4 GN4 GP4 Z4 VSS VDD passgate
.ends

.subckt mux8onehot select0 select1 select2 A1 A2 A3 A4 A5 A6 A7 A8 Z VDD VSS
Xx1 select0 select1 select2 x3/GN1 x3/GP1 x3/GN2 x3/GP2 x3/GN3 x3/GP3 x3/GN4 x3/GP4
+ x5/GN VDD VSS passgatesCtrlManual
Xx2 A1 x3/GN1 A2 x3/GN2 x3/GP2 x5/A A3 x3/GN3 x3/GP3 x5/A A4 x3/GN4 x3/GP4 x5/A x3/GP1
+ x5/A VSS VDD passgatex4
Xx3 A5 x3/GN1 A6 x3/GN2 x3/GP2 x4/A A7 x3/GN3 x3/GP3 x4/A A8 x3/GN4 x3/GP4 x4/A x3/GP1
+ x4/A VSS VDD passgatex4
Xx4 x4/A select2 x5/GN Z VSS VDD passgate
Xx5 x5/A x5/GN select2 Z VSS VDD passgate
.ends

.subckt mux4onehot_b select0 select1 select2 A1 A2 A3 A4 Z1 Z2 Z3 Z4 nselect2 VDD
+ m3_8196_n3226# VSS
Xx1 select0 select1 select2 x2/GN1 x2/GP1 x2/GN2 x2/GP2 x2/GN3 x2/GP3 x2/GN4 x2/GP4
+ nselect2 VDD VSS passgatesCtrlManual
Xx2 A1 x2/GN1 A2 x2/GN2 x2/GP2 Z2 A3 x2/GN3 x2/GP3 Z3 A4 x2/GN4 x2/GP4 Z4 x2/GP1 Z1
+ VSS VDD passgatex4
.ends

.subckt sky130_fd_pr__res_high_po_1p41_DV8LAQ a_n141_n591# a_n141_159# a_n271_n721#
X0 a_n141_159# a_n141_n591# a_n271_n721# sky130_fd_pr__res_high_po_1p41 l=1.75
.ends

.subckt muxtest SELECT0 SELECT1 VRES RSEL0 RSEL1 RSEL2 LADDEROUT OUT VDD VSS
Xx1 RSEL0 RSEL1 RSEL2 R7R8 R6R7 R5R6 R4R5 R3R4 R2R3 R1R2 VRES LADDEROUT VDD VSS mux8onehot
Xx2 SELECT0 SELECT1 VDD LADDEROUT VRES R3R4 R7R8 OUT OUT OUT OUT x2/nselect2 VDD VRES
+ VSS mux4onehot_b
XXR1 VRES R1R2 VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
XXR2 R1R2 R2R3 VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
XXR3 R2R3 R3R4 VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
XXR5 R4R5 R5R6 VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
XXR4 R3R4 R4R5 VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
XXR6 R5R6 R6R7 VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
XXR7 R6R7 R7R8 VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
XXR8 R7R8 VSS VSS sky130_fd_pr__res_high_po_1p41_DV8LAQ
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1975 pd=1.895 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.128375 pd=1.37 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1975 ps=1.895 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.128375 ps=1.37 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt ring VDD enable out VSS
Xsky130_fd_sc_hd__inv_2_10 out VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_11/A sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_11 sky130_fd_sc_hd__inv_2_11/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_12/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nand2_2_0 enable sky130_fd_sc_hd__inv_2_9/Y VSS VSS VDD VDD out
+ sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_12 sky130_fd_sc_hd__inv_2_12/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_13/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_13 sky130_fd_sc_hd__inv_2_13/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_14/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_14 sky130_fd_sc_hd__inv_2_14/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_15/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_7/Y VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_9/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_15 sky130_fd_sc_hd__inv_2_15/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_16/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 sky130_fd_sc_hd__inv_2_8/Y VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_2/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_16 sky130_fd_sc_hd__inv_2_16/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_17/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_2 sky130_fd_sc_hd__inv_2_2/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_3/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_17 sky130_fd_sc_hd__inv_2_17/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_8/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_3 sky130_fd_sc_hd__inv_2_3/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_4/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_4 sky130_fd_sc_hd__inv_2_4/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_5/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_5 sky130_fd_sc_hd__inv_2_5/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_6/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_6 sky130_fd_sc_hd__inv_2_6/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_7/A
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_7 sky130_fd_sc_hd__inv_2_7/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_7/Y
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_8 sky130_fd_sc_hd__inv_2_8/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_8/Y
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_9 sky130_fd_sc_hd__inv_2_9/A VSS VSS VDD VDD sky130_fd_sc_hd__inv_2_9/Y
+ sky130_fd_sc_hd__inv_2
.ends

.subckt sky130_fd_pr__nfet_01v8_F5PS5H a_n33_n300# a_n369_n388# a_303_322# a_15_n388#
+ a_n81_322# a_n177_n388# a_159_n300# a_n515_n474# a_n273_322# a_n413_n300# a_255_n300#
+ a_351_n300# a_n129_n300# a_63_n300# a_n225_n300# a_n321_n300# a_111_322# a_207_n388#
X0 a_255_n300# a_207_n388# a_159_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X1 a_n321_n300# a_n369_n388# a_n413_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
**devattr s=37200,1324 d=19800,666
X2 a_159_n300# a_111_322# a_63_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X3 a_n225_n300# a_n273_322# a_n321_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X4 a_63_n300# a_15_n388# a_n33_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X5 a_n129_n300# a_n177_n388# a_n225_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X6 a_n33_n300# a_n81_322# a_n129_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
**devattr s=19800,666 d=19800,666
X7 a_351_n300# a_303_322# a_255_n300# a_n515_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
**devattr s=19800,666 d=37200,1324
.ends

.subckt sky130_fd_pr__pfet_01v8_XGSFBL a_n33_n997# a_n73_n900# a_15_n900# w_n211_n1119#
X0 a_15_n900# a_n33_n997# a_n73_n900# w_n211_n1119# sky130_fd_pr__pfet_01v8 ad=2.61 pd=18.58 as=2.61 ps=18.58 w=9 l=0.15
**devattr s=104400,3716 d=104400,3716
.ends

.subckt sky130_fd_pr__nfet_01v8_J2SMEF a_n175_n474# a_n73_n300# a_n33_n388# a_15_n300#
X0 a_15_n300# a_n33_n388# a_n73_n300# a_n175_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
**devattr s=34800,1316 d=34800,1316
.ends

.subckt sky130_fd_pr__pfet_01v8_UG67RG a_n33_n900# a_159_n900# a_n413_n900# a_111_931#
+ a_255_n900# a_207_n997# a_351_n900# a_n369_n997# a_303_931# a_n129_n900# a_63_n900#
+ w_n551_n1119# a_n225_n900# a_15_n997# a_n81_931# a_n177_n997# a_n273_931# a_n321_n900#
X0 a_255_n900# a_207_n997# a_159_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X1 a_n321_n900# a_n369_n997# a_n413_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=2.79 ps=18.62 w=9 l=0.15
**devattr s=111600,3724 d=59400,1866
X2 a_159_n900# a_111_931# a_63_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X3 a_n225_n900# a_n273_931# a_n321_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X4 a_63_n900# a_15_n997# a_n33_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X5 a_n129_n900# a_n177_n997# a_n225_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X6 a_n33_n900# a_n81_931# a_n129_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
**devattr s=59400,1866 d=59400,1866
X7 a_351_n900# a_303_931# a_255_n900# w_n551_n1119# sky130_fd_pr__pfet_01v8 ad=2.79 pd=18.62 as=1.485 ps=9.33 w=9 l=0.15
**devattr s=59400,1866 d=111600,3724
.ends

.subckt driver VDD in out VSS
XXM12 VSS m1_3340_n180# m1_3340_n180# m1_3340_n180# m1_3340_n180# m1_3340_n180# VSS
+ VSS m1_3340_n180# VSS out VSS out out VSS out m1_3340_n180# m1_3340_n180# sky130_fd_pr__nfet_01v8_F5PS5H
XXM9 in VDD m1_3340_n180# VDD sky130_fd_pr__pfet_01v8_XGSFBL
XXM10 VSS VSS in m1_3340_n180# sky130_fd_pr__nfet_01v8_J2SMEF
XXM11 VDD VDD VDD m1_3340_n180# out m1_3340_n180# VDD m1_3340_n180# m1_3340_n180#
+ out out VDD VDD m1_3340_n180# m1_3340_n180# m1_3340_n180# m1_3340_n180# out sky130_fd_pr__pfet_01v8_UG67RG
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=4.73
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=4.73
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=0.59
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=0.59
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.3375 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6900,269
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.16875 ps=1.3375 w=1 l=0.15
**devattr s=6900,269 d=6400,264
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
**devattr s=4160,194 d=4290,196
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.144083 ps=1.31 w=0.65 l=0.15
**devattr s=4485,199 d=4160,194
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.144083 pd=1.31 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=4485,199
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.144083 pd=1.31 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=8320,388
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
**devattr s=4290,196 d=4290,196
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16875 pd=1.3375 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6400,264 d=6600,266
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.1625 ps=1.325 w=1 l=0.15
**devattr s=6600,266 d=12800,528
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.16875 ps=1.3375 w=1 l=0.15
**devattr s=6600,266 d=6600,266
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.139399 ps=0.987313 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.331903 ps=2.350746 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.139399 ps=0.987313 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139399 pd=0.987313 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.154085 pd=1.044112 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139399 pd=0.987313 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.238465 ps=1.615888 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.128382 ps=1.053134 w=0.42 l=0.15
**devattr s=5830,267 d=5160,236
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2646,147 d=4368,272
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06831 pd=0.73445 as=0.0742 ps=0.913333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
**devattr s=2688,148 d=1764,126
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.913333 as=0.06831 ps=0.73445 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128382 pd=1.053134 as=0.129 ps=1.18 w=0.42 l=0.15
**devattr s=5160,236 d=8370,269
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.128382 ps=1.053134 w=0.42 l=0.15
**devattr s=8370,269 d=2688,148
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.06831 ps=0.73445 w=0.42 l=0.15
**devattr s=3945,196 d=2646,147
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305672 pd=2.507463 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5830,267
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128382 pd=1.053134 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=4368,272
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.105719 pd=1.136649 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3945,196
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=3835,189
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.1475 ps=1.295 w=1 l=0.15
**devattr s=5900,259 d=10600,506
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
**devattr s=6890,366 d=3640,186
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.181667 ps=1.696667 w=1 l=0.15
**devattr s=5600,256 d=5900,259
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.181667 pd=1.696667 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
**devattr s=3835,189 d=6890,366
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.723333 as=0.265 ps=2.53 w=1 l=0.15
**devattr s=10600,506 d=6500,265
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.723333 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
**devattr s=4452,274 d=2730,149
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.723333 w=1 l=0.15
**devattr s=6500,265 d=5400,254
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0819 ps=0.95 w=0.42 l=0.15
**devattr s=2730,149 d=2268,138
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.95 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12054 ps=1.304827 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.071208 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12353 pd=1.162647 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.193015 ps=1.816635 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.081066 ps=0.762987 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.074954 ps=0.823846 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193015 pd=1.816635 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.081066 pd=0.762987 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.126592 pd=1.2736 as=0.118685 ps=1.284752 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.140385 pd=1.378205 as=0.144761 ps=1.362476 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.071077 ps=0.802308 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.077887 ps=0.843119 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.078615 ps=0.771795 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.064246 pd=0.706154 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.060923 pd=0.687692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.081066 pd=0.762987 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.075046 ps=0.766154 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12353 ps=1.162647 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.12054 pd=1.304827 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.087554 pd=0.893846 as=0.077887 ps=0.843119 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077887 pd=0.843119 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066633 ps=0.67519 w=0.42 l=0.15
**devattr s=4010,197 d=4368,272
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.278216 pd=2.336257 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=11200,512
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.103122 pd=1.044937 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4010,197
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.116851 ps=0.981228 w=0.42 l=0.15
**devattr s=7430,283 d=4704,280
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103122 pd=1.044937 as=0.128917 ps=1.263333 w=0.65 l=0.15
**devattr s=4290,196 d=3510,184
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4290,196
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.278216 ps=2.336257 w=1 l=0.15
**devattr s=12000,520 d=6600,266
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
**devattr s=6600,266 d=4200,242
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128917 pd=1.263333 as=0.103122 ps=1.044937 w=0.65 l=0.15
**devattr s=3510,184 d=6890,366
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.278216 pd=2.336257 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=7430,283
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073937 pd=0.752655 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.073937 pd=0.752655 as=0.0805 ps=0.943333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103351 pd=0.894953 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.943333 as=0.073937 ps=0.752655 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.17604 ps=1.792035 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.159949 ps=1.385047 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138125 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.4 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.4 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.176667 ps=1.686667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176667 pd=1.686667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.138125 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=2.89
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=2.89
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=10600,506 d=5600,256
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2310,139
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5500,255
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.063945 pd=0.7665 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15225 pd=1.4045 as=0.14 ps=1.28 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15225 ps=1.4045 w=1 l=0.15
**devattr s=5600,256 d=5600,256
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.063945 ps=0.7665 w=0.42 l=0.15
**devattr s=2310,139 d=2352,140
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.2262 ps=2.26 w=0.87 l=1.97
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.97
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=4200,242
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
.ends

.subckt simplecounter VPWR clk enable counter[0] counter[1] counter[2] counter[3]
+ counter[4] counter[5] counter[6] counter[7] counter[8] counter[9] VGND
X_49_ _23_ _24_ VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput7 net7 VGND VGND VPWR VPWR counter[5] sky130_fd_sc_hd__buf_1
XFILLER_0_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_48_ _11_ _15_ _22_ net10 VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_12_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR counter[8] sky130_fd_sc_hd__buf_1
Xoutput8 net8 VGND VGND VPWR VPWR counter[6] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_47_ net10 _11_ _15_ _22_ VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput11 net11 VGND VGND VPWR VPWR counter[9] sky130_fd_sc_hd__buf_1
Xoutput9 net9 VGND VGND VPWR VPWR counter[7] sky130_fd_sc_hd__buf_1
X_46_ _16_ _22_ _21_ net9 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29_ net2 net1 net3 VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28_ _10_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__clkbuf_2
X_45_ net6 net7 net8 net9 VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__and4_1
X_61_ clknet_1_1__leaf_clk _09_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
X_44_ net8 _17_ _21_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_4_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27_ net2 net3 net1 VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_60_ clknet_1_1__leaf_clk _08_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
X_26_ net2 net1 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__xor2_1
X_43_ _11_ _15_ _20_ VGND VGND VPWR VPWR _21_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_42_ net6 net7 net8 VGND VGND VPWR VPWR _20_ sky130_fd_sc_hd__and3_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_41_ _19_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_40_ _17_ _18_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 enable VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_59_ clknet_1_1__leaf_clk _07_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_58_ clknet_1_1__leaf_clk _06_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_57_ clknet_1_1__leaf_clk _05_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_56_ clknet_1_0__leaf_clk _04_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_1
X_39_ net6 _11_ _15_ net7 VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__a31o_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_55_ clknet_1_0__leaf_clk _03_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_38_ net6 net7 _11_ _15_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_54_ clknet_1_0__leaf_clk _02_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_2_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_37_ net6 _16_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_53_ clknet_1_0__leaf_clk _01_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfxtp_1
X_36_ net5 _14_ _16_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_52_ clknet_1_0__leaf_clk _00_ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dfxtp_1
X_35_ _11_ _15_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_51_ net11 _23_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_34_ net4 net5 VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33_ _13_ _14_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__nor2_1
X_50_ _25_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_32_ net4 _11_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31_ net4 _11_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30_ _11_ _12_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput2 net2 VGND VGND VPWR VPWR counter[0] sky130_fd_sc_hd__buf_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput3 net3 VGND VGND VPWR VPWR counter[1] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_8_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR counter[2] sky130_fd_sc_hd__buf_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR counter[3] sky130_fd_sc_hd__buf_1
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput6 net6 VGND VGND VPWR VPWR counter[4] sky130_fd_sc_hd__buf_1
.ends

.subckt ringtest enable_ring select0 select1 enable_counter mux_out VDD VSS
Xx1 VDD enable_ring ring_out VSS ring
Xx2 VDD ring_out drv_out VSS driver
Xx3 select0 select1 VDD ring_out drv_out counter3 counter7 mux_out mux_out mux_out
+ mux_out x3/nselect2 VDD x3/m3_8196_n3226# VSS mux4onehot_b
Xx4 VDD drv_out enable_counter x4/counter[0] x4/counter[1] x4/counter[2] counter3
+ x4/counter[4] x4/counter[5] x4/counter[6] counter7 x4/counter[8] x4/counter[9] VSS
+ simplecounter
.ends

.subckt tt_um_patdeegan_anamux clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VSS
Xmuxtest_0 ui_in[3] ui_in[4] ua[0] ui_in[0] ui_in[1] ui_in[2] ua[3] ua[2] VDPWR VSS
+ muxtest
Xringtest_0 ui_in[6] ui_in[3] ui_in[4] ui_in[5] ua[1] VDPWR VSS ringtest
R0 VSS uio_oe[7] 0.000000
R1 VSS uo_out[2] 0.000000
R2 VSS uio_oe[6] 0.000000
R3 VSS uo_out[1] 0.000000
R4 VSS uio_oe[5] 0.000000
R5 VSS uo_out[0] 0.000000
R6 VSS uio_oe[4] 0.000000
R7 VSS uio_out[7] 0.000000
R8 VSS uio_oe[3] 0.000000
R9 VSS uio_out[6] 0.000000
R10 VSS uio_oe[1] 0.000000
R11 VSS uio_oe[2] 0.000000
R12 VSS uio_out[4] 0.000000
R13 VSS uio_out[5] 0.000000
R14 VSS uo_out[7] 0.000000
R15 VSS uio_out[3] 0.000000
R16 VSS uo_out[6] 0.000000
R17 VSS uo_out[5] 0.000000
R18 VSS uio_oe[0] 0.000000
R19 VSS uio_out[2] 0.000000
R20 VSS uio_out[1] 0.000000
R21 VSS uo_out[4] 0.000000
R22 VSS uio_out[0] 0.000000
R23 VSS uo_out[3] 0.000000
.ends

