magic
tech sky130A
magscale 1 2
timestamp 1728327329
<< metal1 >>
rect 4798 -2878 4926 -2784
rect 4798 -2958 4840 -2878
rect 7146 -3218 7334 -3030
rect 7630 -3186 7640 -3098
rect 7758 -3186 7768 -3098
rect 8196 -3226 8396 -3026
rect 8690 -3178 8700 -3030
rect 8842 -3178 8852 -3030
rect 9240 -3230 9440 -3030
rect 9720 -3162 9730 -3056
rect 9884 -3162 9894 -3056
rect 10270 -3216 10470 -3016
rect 10766 -3172 10776 -3038
rect 10910 -3172 10920 -3038
rect 4852 -4981 4918 -4786
rect 4982 -4985 5048 -4790
rect 5096 -4985 5162 -4785
rect 7112 -7960 7312 -7596
rect 8180 -7956 8380 -7756
rect 9250 -7992 9450 -7792
rect 10308 -7994 10508 -7592
<< via1 >>
rect 7640 -3186 7758 -3098
rect 8700 -3178 8842 -3030
rect 9730 -3162 9884 -3056
rect 10776 -3172 10910 -3038
<< metal2 >>
rect 6430 -2452 10861 -2405
rect 6430 -3270 6477 -2452
rect 6526 -2522 10628 -2482
rect 6526 -3319 6566 -2522
rect 6431 -3359 6566 -3319
rect 6602 -2596 9816 -2556
rect 6602 -3511 6642 -2596
rect 6454 -3551 6642 -3511
rect 6679 -2679 9586 -2638
rect 6679 -3609 6720 -2679
rect 6458 -3650 6720 -3609
rect 6758 -2758 8787 -2719
rect 6758 -3881 6797 -2758
rect 6453 -3920 6797 -3881
rect 6838 -2839 8535 -2801
rect 6838 -4083 6876 -2839
rect 7671 -2879 7714 -2876
rect 6462 -4116 6876 -4083
rect 6838 -4118 6876 -4116
rect 6911 -2917 7714 -2879
rect 6911 -4164 6949 -2917
rect 6471 -4194 6949 -4164
rect 6911 -4198 6949 -4194
rect 6985 -2984 7483 -2949
rect 6985 -4776 7020 -2984
rect 7448 -3181 7483 -2984
rect 7671 -3088 7714 -2917
rect 7640 -3098 7758 -3088
rect 8497 -3131 8535 -2839
rect 8748 -3020 8787 -2758
rect 8700 -3030 8842 -3020
rect 8497 -3169 8567 -3131
rect 7640 -3196 7758 -3186
rect 8700 -3188 8842 -3178
rect 9545 -3182 9586 -2679
rect 9776 -3046 9816 -2596
rect 9730 -3056 9884 -3046
rect 9730 -3172 9884 -3162
rect 10588 -3170 10628 -2522
rect 10814 -3028 10861 -2452
rect 10776 -3038 10910 -3028
rect 9776 -3182 9816 -3172
rect 10776 -3182 10910 -3172
rect 6465 -4806 7020 -4776
rect 6985 -4808 7020 -4806
rect 5750 -4877 6864 -4872
rect 5746 -4963 5755 -4877
rect 5841 -4963 6864 -4877
rect 5750 -4968 6864 -4963
rect 6960 -4968 6969 -4872
rect 6864 -7651 7556 -7646
rect 6860 -7737 6869 -7651
rect 6955 -7737 7556 -7651
rect 6864 -7742 7556 -7737
rect 7398 -7848 7494 -7742
<< via2 >>
rect 5755 -4963 5841 -4877
rect 6864 -4968 6960 -4872
rect 6869 -7737 6955 -7651
<< metal3 >>
rect 6281 -2799 6451 -2527
rect 6281 -2969 8112 -2799
rect 6281 -2971 6451 -2969
rect 7942 -3447 8112 -2969
rect 8196 -3226 8396 -3026
rect 9240 -3230 9440 -3030
rect 10270 -3216 10470 -3016
rect 5750 -4870 5846 -4672
rect 5742 -4877 5864 -4870
rect 5742 -4963 5755 -4877
rect 5841 -4963 5864 -4877
rect 5742 -4980 5864 -4963
rect 6859 -4872 6965 -4867
rect 6859 -4968 6864 -4872
rect 6960 -4968 6965 -4872
rect 6859 -4973 6965 -4968
rect 6864 -7651 6960 -4973
rect 6864 -7737 6869 -7651
rect 6955 -7737 6960 -7651
rect 6864 -7742 6960 -7737
use passgatesCtrlManual  x1
timestamp 1728289486
transform 0 -1 1696 1 0 -5526
box 666 -4798 2906 -2962
use passgatex4  x2
timestamp 1728255086
transform 1 0 -4302 0 1 -7698
box 11366 -356 15589 4682
<< labels >>
flabel metal1 4984 -4980 5046 -4918 0 FreeSans 640 0 0 0 select0
port 0 nsew
flabel metal1 4854 -4976 4916 -4914 0 FreeSans 640 0 0 0 select1
port 1 nsew
flabel metal1 5098 -4980 5160 -4918 0 FreeSans 640 0 0 0 select2
port 2 nsew
flabel metal1 8196 -3226 8396 -3026 0 FreeSans 640 0 0 0 A2
port 4 nsew
flabel metal1 9240 -3230 9440 -3030 0 FreeSans 640 0 0 0 A3
port 5 nsew
flabel metal1 10270 -3216 10470 -3016 0 FreeSans 640 0 0 0 A4
port 6 nsew
flabel metal1 7112 -7960 7312 -7596 0 FreeSans 640 0 0 0 Z1
port 7 nsew
flabel metal1 8180 -7956 8380 -7756 0 FreeSans 640 0 0 0 Z2
port 8 nsew
flabel metal1 9250 -7992 9450 -7792 0 FreeSans 640 0 0 0 Z3
port 9 nsew
flabel metal1 10308 -7994 10508 -7592 0 FreeSans 640 0 0 0 Z4
port 10 nsew
flabel metal1 4798 -2878 4926 -2784 0 FreeSans 640 0 0 0 nselect2
port 11 nsew
flabel metal3 5742 -4980 5864 -4870 0 FreeSans 800 0 0 0 VDD
port 12 nsew
flabel metal3 6281 -2695 6451 -2525 0 FreeSans 800 0 0 0 VSS
port 13 nsew
flabel metal1 7146 -3218 7334 -3030 0 FreeSans 1600 0 0 0 A1
port 3 nsew
<< end >>
