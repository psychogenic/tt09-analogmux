magic
tech sky130A
magscale 1 2
timestamp 1728370683
<< metal1 >>
rect 26516 44628 26522 44761
rect 26655 44628 26661 44761
rect 27071 44649 27077 44776
rect 27204 44649 27210 44776
rect 27629 44655 27635 44769
rect 27749 44655 27755 44769
rect 25414 42326 25614 42332
rect 10916 42126 10922 42326
rect 11122 42126 25414 42326
rect 25414 42120 25614 42126
rect 10388 41688 10394 41864
rect 10570 41688 25948 41864
rect 26124 41688 26130 41864
rect 17921 35009 18068 35016
rect 17921 34876 17928 35009
rect 18061 34876 18068 35009
rect 17921 33145 18068 34876
rect 26522 35009 26655 44628
rect 26522 34870 26655 34876
rect 18185 34507 18307 34513
rect 18185 34346 18307 34385
rect 27077 34510 27204 44649
rect 27077 34377 27204 34383
rect 18184 34263 18307 34346
rect 18184 33160 18305 34263
rect 18450 34085 18583 34091
rect 27635 34075 27749 44655
rect 27629 33961 27635 34075
rect 27749 33961 27755 34075
rect 18450 33864 18583 33952
rect 18445 33274 18583 33864
rect 18445 33203 18571 33274
rect 21616 30836 22914 30864
rect 21616 30296 22338 30836
rect 22878 30296 22914 30836
rect 21616 30262 22914 30296
rect 6874 25260 7090 25268
rect 6874 25060 11440 25260
rect 6874 698 7090 25060
rect 7880 24691 7886 24891
rect 8086 24691 10922 24891
rect 11122 24691 11680 24891
rect 7438 24297 7444 24497
rect 7644 24297 10390 24497
rect 10590 24297 11448 24497
rect 21404 20702 30357 21024
rect 7318 19117 7539 19128
rect 7318 18917 8392 19117
rect 7318 1233 7539 18917
rect 7881 17599 7887 17798
rect 8086 17797 12169 17798
rect 8086 17599 12897 17797
rect 13095 17599 13101 17797
rect 7730 17330 7930 17336
rect 7930 17130 12638 17330
rect 12838 17130 12844 17330
rect 17648 17206 23838 17486
rect 24118 17206 24124 17486
rect 7730 17124 7930 17130
rect 17648 15982 17928 17206
rect 11884 1812 12084 7280
rect 11884 1612 26698 1812
rect 7318 1012 22798 1233
rect 22577 817 22798 1012
rect 26498 949 26698 1612
rect 30035 1086 30357 20702
rect 30035 1065 30611 1086
rect 18741 698 18747 703
rect 6874 482 18747 698
rect 18741 477 18747 482
rect 18973 477 18979 703
rect 22577 578 22599 817
rect 22593 566 22599 578
rect 22850 566 22856 817
rect 26469 753 26708 949
rect 30035 875 30315 1065
rect 30037 790 30315 875
rect 30590 790 30611 1065
rect 30037 768 30611 790
rect 26463 514 26469 753
rect 26708 514 26714 753
<< via1 >>
rect 26522 44628 26655 44761
rect 27077 44649 27204 44776
rect 27635 44655 27749 44769
rect 10922 42126 11122 42326
rect 25414 42126 25614 42326
rect 10394 41688 10570 41864
rect 25948 41688 26124 41864
rect 17928 34876 18061 35009
rect 26522 34876 26655 35009
rect 18185 34385 18307 34507
rect 27077 34383 27204 34510
rect 18450 33952 18583 34085
rect 27635 33961 27749 34075
rect 22338 30296 22878 30836
rect 7886 24691 8086 24891
rect 10922 24691 11122 24891
rect 7444 24297 7644 24497
rect 10390 24297 10590 24497
rect 7887 17599 8086 17798
rect 12897 17599 13095 17797
rect 7730 17130 7930 17330
rect 12638 17130 12838 17330
rect 23838 17206 24118 17486
rect 18747 477 18973 703
rect 22599 566 22850 817
rect 30315 790 30590 1065
rect 26469 514 26708 753
<< metal2 >>
rect 27077 44864 27204 44882
rect 25414 44834 25610 44858
rect 25414 44743 25439 44834
rect 25530 44743 25610 44834
rect 25414 44604 25610 44743
rect 25954 44817 26118 44844
rect 25954 44708 25982 44817
rect 26091 44708 26118 44817
rect 25954 44704 26118 44708
rect 26522 44818 26655 44843
rect 26522 44761 26547 44818
rect 26630 44761 26655 44818
rect 10922 42326 11122 42332
rect 25414 42326 25614 44604
rect 25408 42126 25414 42326
rect 25614 42126 25620 42326
rect 10394 41864 10570 41870
rect 10394 26551 10570 41688
rect 7886 24891 8086 24897
rect 7886 24685 8086 24691
rect 7444 24497 7644 24503
rect 7444 17330 7644 24297
rect 7887 17798 8086 24685
rect 10394 24503 10571 26551
rect 10922 24891 11122 42126
rect 25948 41864 26124 44704
rect 27077 44776 27094 44864
rect 27186 44776 27204 44864
rect 27635 44859 27749 44875
rect 27635 44777 27651 44859
rect 27733 44777 27749 44859
rect 27635 44769 27749 44777
rect 27635 44649 27749 44655
rect 27077 44643 27204 44649
rect 26522 44622 26655 44628
rect 25948 41682 26124 41688
rect 17922 34876 17928 35009
rect 18061 34876 26522 35009
rect 26655 34876 26661 35009
rect 27071 34507 27077 34510
rect 18179 34385 18185 34507
rect 18307 34385 27077 34507
rect 27071 34383 27077 34385
rect 27204 34383 27210 34510
rect 18444 33952 18450 34085
rect 18583 34075 27759 34085
rect 18583 33961 27635 34075
rect 27749 33961 27759 34075
rect 18583 33952 27759 33961
rect 23838 33472 24118 33481
rect 22294 30853 23566 30892
rect 22294 30836 22973 30853
rect 22294 30296 22338 30836
rect 22878 30296 22973 30836
rect 22294 30280 22973 30296
rect 23546 30280 23566 30853
rect 22294 30248 23566 30280
rect 10922 24685 11122 24691
rect 10390 24497 10590 24503
rect 10390 24291 10590 24297
rect 7887 17593 8086 17599
rect 12897 17800 13095 17803
rect 12897 17797 13097 17800
rect 13095 17599 13097 17797
rect 12897 17593 13097 17599
rect 12638 17330 12838 17336
rect 7444 17130 7730 17330
rect 7930 17130 7936 17330
rect 12638 17124 12838 17130
rect 12715 15905 12833 17124
rect 12960 15875 13097 17593
rect 23838 17486 24118 33192
rect 23838 17200 24118 17206
rect 24306 33344 24498 33353
rect 24306 16648 24498 33152
rect 21892 16456 24498 16648
rect 11959 13050 11968 13306
rect 12224 13050 12554 13306
rect 30315 1065 30590 1071
rect 22599 817 22850 823
rect 18747 703 18973 709
rect 18747 299 18761 477
rect 18959 299 18973 477
rect 22599 358 22618 566
rect 22830 358 22850 566
rect 22599 339 22850 358
rect 26469 753 26708 759
rect 26469 328 26483 514
rect 26694 328 26708 514
rect 30315 700 30590 790
rect 30315 464 30334 700
rect 30570 464 30590 700
rect 30315 445 30590 464
rect 26469 314 26708 328
rect 18747 285 18973 299
<< via2 >>
rect 25439 44743 25530 44834
rect 25982 44708 26091 44817
rect 26547 44761 26630 44818
rect 26547 44735 26630 44761
rect 27094 44776 27186 44864
rect 27094 44772 27186 44776
rect 27651 44777 27733 44859
rect 23838 33192 24118 33472
rect 22973 30280 23546 30853
rect 24306 33152 24498 33344
rect 11968 13050 12224 13306
rect 18761 477 18959 497
rect 18761 299 18959 477
rect 22618 566 22830 570
rect 22618 358 22830 566
rect 26483 514 26694 539
rect 26483 328 26694 514
rect 30334 464 30570 700
<< metal3 >>
rect 25434 44904 25535 44923
rect 24890 44891 24976 44892
rect 24257 44834 24475 44869
rect 24257 44743 24335 44834
rect 24426 44743 24475 44834
rect 23838 43883 24118 43884
rect 24257 43883 24475 44743
rect 23838 43665 24475 43883
rect 24836 44807 24891 44891
rect 24975 44807 25031 44891
rect 23838 33477 24118 43665
rect 24836 43493 25031 44807
rect 25434 44840 25452 44904
rect 25516 44840 25535 44904
rect 25434 44834 25535 44840
rect 25434 44743 25439 44834
rect 25530 44743 25535 44834
rect 25434 44738 25535 44743
rect 25977 44916 26096 44944
rect 25977 44852 26004 44916
rect 26068 44852 26096 44916
rect 25977 44817 26096 44852
rect 25977 44708 25982 44817
rect 26091 44708 26096 44817
rect 26542 44916 26635 44931
rect 26542 44852 26556 44916
rect 26620 44852 26635 44916
rect 26542 44818 26635 44852
rect 26542 44735 26547 44818
rect 26630 44735 26635 44818
rect 27089 44918 27191 44937
rect 27089 44864 27108 44918
rect 27172 44864 27191 44918
rect 27089 44772 27094 44864
rect 27186 44772 27191 44864
rect 27646 44918 27738 44932
rect 27646 44859 27660 44918
rect 27724 44859 27738 44918
rect 27646 44777 27651 44859
rect 27733 44777 27738 44859
rect 27646 44772 27738 44777
rect 27089 44767 27191 44772
rect 26542 44730 26635 44735
rect 25977 44703 26096 44708
rect 24305 43298 25031 43493
rect 23833 33472 24123 33477
rect 23833 33192 23838 33472
rect 24118 33192 24123 33472
rect 24305 33349 24500 43298
rect 23833 33187 24123 33192
rect 24301 33344 24503 33349
rect 24301 33152 24306 33344
rect 24498 33152 24503 33344
rect 24301 33147 24503 33152
rect 5454 32660 5464 32664
rect 5359 32154 5464 32660
rect 5454 32126 5464 32154
rect 6168 32660 6178 32664
rect 6168 32154 17902 32660
rect 29916 32563 29926 32646
rect 20452 32394 29926 32563
rect 29916 32338 29926 32394
rect 30720 32563 30730 32646
rect 30720 32394 30852 32563
rect 30720 32338 30730 32394
rect 6168 32126 6178 32154
rect 5384 31118 12145 31133
rect 5384 30900 5464 31118
rect 5454 30896 5464 30900
rect 6080 30900 12145 31118
rect 6080 30896 6090 30900
rect 22916 30853 30818 30904
rect 22916 30280 22973 30853
rect 23546 30834 30818 30853
rect 23546 30302 29836 30834
rect 30720 30302 30818 30834
rect 23546 30280 30818 30302
rect 22916 30212 30818 30280
rect 5318 22410 5328 22616
rect 6258 22588 6268 22616
rect 6258 22561 8905 22588
rect 6258 22465 9010 22561
rect 6258 22438 8905 22465
rect 6258 22410 6268 22438
rect 17651 21343 18033 21529
rect 18219 21343 18225 21529
rect 17952 20136 30742 20188
rect 17952 20078 29864 20136
rect 17952 19570 17986 20078
rect 18270 19570 29864 20078
rect 17952 19536 29864 19570
rect 30692 19536 30742 20136
rect 5378 16765 5388 16824
rect 5330 16393 5388 16765
rect 5378 16310 5388 16393
rect 6198 16765 6208 16824
rect 6198 16393 13138 16765
rect 6198 16310 6208 16393
rect 5418 13342 5428 13424
rect 5322 13014 5428 13342
rect 5418 12926 5428 13014
rect 6270 13342 6280 13424
rect 6270 13306 12260 13342
rect 6270 13050 11968 13306
rect 12224 13050 12260 13306
rect 6270 13014 12260 13050
rect 6270 12926 6280 13014
rect 28192 11764 30836 11784
rect 28192 11738 29852 11764
rect 28124 11426 29852 11738
rect 28192 11400 29852 11426
rect 30790 11400 30836 11764
rect 28192 11380 30836 11400
rect 5380 10727 5390 10768
rect 5315 10521 5390 10727
rect 5380 10462 5390 10521
rect 6240 10727 6250 10768
rect 6240 10521 12762 10727
rect 6240 10462 6250 10521
rect 27956 10348 30798 10378
rect 27956 9958 29874 10348
rect 30698 9958 30798 10348
rect 27956 9924 30798 9958
rect 27946 7146 30788 7174
rect 27946 6756 29878 7146
rect 30702 6756 30788 7146
rect 27946 6720 30788 6756
rect 27950 4908 30792 4948
rect 27950 4518 29888 4908
rect 30712 4518 30792 4908
rect 27950 4494 30792 4518
rect 5348 3620 5358 3656
rect 5328 3118 5358 3620
rect 5348 3054 5358 3118
rect 6264 3620 6274 3656
rect 6264 3118 20901 3620
rect 6264 3054 6274 3118
rect 30329 700 30575 705
rect 22613 570 22835 575
rect 18756 497 18964 502
rect 18756 299 18761 497
rect 18959 299 18964 497
rect 18756 173 18771 299
rect 18949 173 18964 299
rect 22613 358 22618 570
rect 22830 358 22835 570
rect 22613 219 22635 358
rect 22813 219 22835 358
rect 22613 197 22835 219
rect 26478 539 26699 544
rect 26478 328 26483 539
rect 26694 328 26699 539
rect 18756 158 18964 173
rect 26478 179 26499 328
rect 26677 179 26699 328
rect 30329 464 30334 700
rect 30570 464 30575 700
rect 30329 459 30575 464
rect 30329 281 30363 459
rect 30541 281 30575 459
rect 30329 247 30575 281
rect 26478 158 26699 179
<< via3 >>
rect 24335 44743 24426 44834
rect 24891 44807 24975 44891
rect 25452 44840 25516 44904
rect 26004 44852 26068 44916
rect 26556 44852 26620 44916
rect 27108 44864 27172 44918
rect 27108 44854 27172 44864
rect 27660 44859 27724 44918
rect 27660 44854 27724 44859
rect 5464 32126 6168 32664
rect 29926 32338 30720 32646
rect 5464 30896 6080 31118
rect 29836 30302 30720 30834
rect 5328 22410 6258 22616
rect 18033 21343 18219 21529
rect 17986 19570 18270 20078
rect 29864 19536 30692 20136
rect 5388 16310 6198 16824
rect 5428 12926 6270 13424
rect 29852 11400 30790 11764
rect 5390 10462 6240 10768
rect 29874 9958 30698 10348
rect 29878 6756 30702 7146
rect 29888 4518 30712 4908
rect 5358 3054 6264 3656
rect 18771 299 18949 351
rect 18771 173 18949 299
rect 22635 358 22813 397
rect 22635 219 22813 358
rect 26499 328 26677 357
rect 26499 179 26677 328
rect 30363 281 30541 459
<< metal4 >>
rect 6134 44532 6194 45152
rect 6686 44532 6746 45152
rect 7238 44532 7298 45152
rect 7790 44532 7850 45152
rect 8342 44532 8402 45152
rect 8894 44532 8954 45152
rect 9446 44532 9506 45152
rect 9998 44532 10058 45152
rect 10550 44532 10610 45152
rect 11102 44532 11162 45152
rect 11654 44532 11714 45152
rect 12206 44532 12266 45152
rect 12758 44532 12818 45152
rect 13310 44532 13370 45152
rect 13862 44532 13922 45152
rect 14414 44532 14474 45152
rect 14966 44532 15026 45152
rect 15518 44532 15578 45152
rect 16070 44532 16130 45152
rect 16622 44532 16682 45152
rect 17174 44532 17234 45152
rect 17726 44532 17786 45152
rect 18278 44532 18338 45152
rect 18830 44532 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44936 22754 45152
rect 23246 44936 23306 45152
rect 23798 44952 23858 45152
rect 24350 44951 24410 45152
rect 24902 45047 24962 45152
rect 24334 44834 24427 44951
rect 24902 44892 24963 45047
rect 25454 44905 25514 45152
rect 26006 44917 26066 45152
rect 26558 44917 26618 45152
rect 27110 44919 27170 45152
rect 27662 44919 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27107 44918 27173 44919
rect 26003 44916 26069 44917
rect 25451 44904 25517 44905
rect 24334 44743 24335 44834
rect 24426 44743 24427 44834
rect 24890 44891 24976 44892
rect 24890 44807 24891 44891
rect 24975 44807 24976 44891
rect 25451 44840 25452 44904
rect 25516 44840 25517 44904
rect 26003 44852 26004 44916
rect 26068 44852 26069 44916
rect 26003 44851 26069 44852
rect 26555 44916 26621 44917
rect 26555 44852 26556 44916
rect 26620 44852 26621 44916
rect 27107 44854 27108 44918
rect 27172 44854 27173 44918
rect 27107 44853 27173 44854
rect 27659 44918 27725 44919
rect 27659 44854 27660 44918
rect 27724 44854 27725 44918
rect 27659 44853 27725 44854
rect 26555 44851 26621 44852
rect 25451 44839 25517 44840
rect 24890 44806 24976 44807
rect 24334 44742 24427 44743
rect 6106 44176 30826 44532
rect 6106 43912 30846 44176
rect 5280 32664 6346 43338
rect 5280 32126 5464 32664
rect 6168 32126 6346 32664
rect 5280 31118 6346 32126
rect 5280 30896 5464 31118
rect 6080 30896 6346 31118
rect 5280 22616 6346 30896
rect 5280 22410 5328 22616
rect 6258 22410 6346 22616
rect 5280 16824 6346 22410
rect 29780 32646 30846 43912
rect 29780 32338 29926 32646
rect 30720 32338 30846 32646
rect 29780 30834 30846 32338
rect 29780 30302 29836 30834
rect 30720 30302 30846 30834
rect 17988 21529 18264 21574
rect 17988 21343 18033 21529
rect 18219 21343 18264 21529
rect 17988 20079 18264 21343
rect 29780 20136 30846 30302
rect 17985 20078 18271 20079
rect 17985 19570 17986 20078
rect 18270 19570 18271 20078
rect 17985 19569 18271 19570
rect 17988 19542 18264 19569
rect 5280 16310 5388 16824
rect 6198 16310 6346 16824
rect 5280 13424 6346 16310
rect 5280 12926 5428 13424
rect 6270 12926 6346 13424
rect 5280 10768 6346 12926
rect 5280 10462 5390 10768
rect 6240 10462 6346 10768
rect 5280 3656 6346 10462
rect 5280 3054 5358 3656
rect 6264 3054 6346 3656
rect 5280 748 6346 3054
rect 29780 19536 29864 20136
rect 30692 19536 30846 20136
rect 29780 11764 30846 19536
rect 29780 11400 29852 11764
rect 30790 11400 30846 11764
rect 29780 10348 30846 11400
rect 29780 9958 29874 10348
rect 30698 9958 30846 10348
rect 29780 7146 30846 9958
rect 29780 6756 29878 7146
rect 30702 6756 30846 7146
rect 29780 4908 30846 6756
rect 29780 4518 29888 4908
rect 30712 4518 30846 4908
rect 29780 1408 30846 4518
rect 30362 459 30542 460
rect 22634 397 22814 398
rect 18770 351 18950 352
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 173 18771 351
rect 18949 173 18950 351
rect 18770 0 18950 173
rect 22634 219 22635 397
rect 22813 219 22814 397
rect 22634 0 22814 219
rect 26498 357 26678 358
rect 26498 179 26499 357
rect 26677 179 26678 357
rect 26498 0 26678 179
rect 30362 281 30363 459
rect 30541 281 30542 459
rect 30362 0 30542 281
use muxtest  muxtest_0
timestamp 1728362514
transform 0 1 23718 -1 0 37419
box 4086 -15558 19281 -1352
use ringtest  ringtest_0
timestamp 1728347809
transform 1 0 -1830 0 1 14049
box 13714 -11825 30474 2702
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 5330 37948 6284 39026 0 FreeSans 1600 0 0 0 VDPWR
port 51 nsew
flabel metal4 29780 38563 30846 39629 0 FreeSans 1600 0 0 0 VSS
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
