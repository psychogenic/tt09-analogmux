magic
tech sky130A
magscale 1 2
timestamp 1728360080
<< metal1 >>
rect 11365 7381 11466 7398
rect 11365 7314 11382 7381
rect 11449 7314 11466 7381
rect 11129 7262 11216 7278
rect 11129 7206 11144 7262
rect 11200 7206 11216 7262
rect 10317 7140 10395 7153
rect 5168 7088 5210 7111
rect 10317 7088 10330 7140
rect 10382 7088 10395 7140
rect 5157 7036 5163 7088
rect 5215 7036 5221 7088
rect 10091 7036 10158 7044
rect 10091 6984 10098 7036
rect 10150 6984 10158 7036
rect 9294 6905 9346 6908
rect 9291 6902 9349 6905
rect 9291 6850 9294 6902
rect 9346 6850 9349 6902
rect 9050 6783 9102 6788
rect 9049 6782 9103 6783
rect 9049 6730 9050 6782
rect 9102 6730 9103 6782
rect 8236 6642 8288 6648
rect 8236 6584 8288 6590
rect 7694 6150 7894 6350
rect 8239 6209 8286 6584
rect 8750 6148 8950 6348
rect 9049 6185 9103 6730
rect 9291 6199 9349 6850
rect 9794 6144 9994 6344
rect 10091 6173 10158 6984
rect 10317 6157 10395 7088
rect 10824 6158 11024 6358
rect 11129 6189 11216 7206
rect 11365 6200 11466 7314
rect 12008 6152 12208 6352
rect 12490 6204 12500 6336
rect 12640 6204 12650 6336
rect 13064 6150 13264 6350
rect 13550 6198 13560 6330
rect 13700 6198 13710 6330
rect 14108 6146 14308 6346
rect 14592 6198 14602 6330
rect 14742 6198 14752 6330
rect 15138 6160 15338 6360
rect 15624 6212 15634 6344
rect 15774 6212 15784 6344
rect 5222 5149 5288 5358
rect 5352 5251 5418 5357
rect 5352 5179 5418 5185
rect 5047 5083 5053 5149
rect 5119 5083 5288 5149
rect 5466 5049 5532 5355
rect 5466 4977 5532 4983
rect 7694 1254 7801 1601
rect 8776 1254 8883 1589
rect 9849 1254 9956 1637
rect 10902 1254 11023 1541
rect 7513 1172 11023 1254
rect 12019 1259 12126 1553
rect 12593 1259 12743 1280
rect 13095 1259 13202 1525
rect 14154 1259 14261 1511
rect 15270 1259 15377 1495
rect 12019 1181 15377 1259
rect 7513 1147 11016 1172
rect 12019 1152 12593 1181
rect 7513 332 7620 1147
rect 12743 1152 15377 1181
rect 12593 1025 12743 1031
rect 12111 581 12261 587
rect 7682 420 7692 574
rect 7846 420 7856 574
rect 7942 432 7952 544
rect 8088 432 8098 544
rect 12111 425 12261 431
rect 7513 225 7815 332
rect 7910 220 7920 346
rect 8114 220 8124 346
rect 11998 158 13042 358
rect 12149 -486 12299 -480
rect 7462 -530 7538 -524
rect 7538 -606 7852 -530
rect 7462 -612 7538 -606
rect 7974 -628 7984 -510
rect 8130 -628 8140 -510
rect 12149 -642 12299 -636
rect 7729 -991 7879 -705
rect 7952 -828 7962 -700
rect 8150 -828 8160 -700
rect 12842 -710 13042 158
rect 12030 -910 13042 -710
rect 7729 -1141 12593 -991
rect 12743 -1141 12749 -991
<< via1 >>
rect 11382 7314 11449 7381
rect 11144 7206 11200 7262
rect 10330 7088 10382 7140
rect 5163 7036 5215 7088
rect 10098 6984 10150 7036
rect 9294 6850 9346 6902
rect 9050 6730 9102 6782
rect 8236 6590 8288 6642
rect 12500 6204 12640 6336
rect 13560 6198 13700 6330
rect 14602 6198 14742 6330
rect 15634 6212 15774 6344
rect 5352 5185 5418 5251
rect 5053 5083 5119 5149
rect 5466 4983 5532 5049
rect 12593 1031 12743 1181
rect 7692 420 7846 574
rect 7952 432 8088 544
rect 12111 431 12261 581
rect 7920 220 8114 346
rect 7462 -606 7538 -530
rect 7984 -628 8130 -510
rect 12149 -636 12299 -486
rect 7962 -828 8150 -700
rect 12593 -1141 12743 -991
<< metal2 >>
rect 6793 7314 11382 7381
rect 11449 7314 15739 7381
rect 5225 7104 5339 7119
rect 5197 7094 5339 7104
rect 5163 7088 5339 7094
rect 5215 7059 5339 7088
rect 5215 7036 5225 7059
rect 5163 7030 5225 7036
rect 5197 7020 5225 7030
rect 5225 6936 5339 6945
rect 6793 6863 6860 7314
rect 6934 7206 11144 7262
rect 11200 7206 15510 7262
rect 6934 6832 6990 7206
rect 10324 7138 10330 7140
rect 6782 6776 6990 6832
rect 7050 7090 10330 7138
rect 7050 6637 7098 7090
rect 10324 7088 10330 7090
rect 10382 7138 10388 7140
rect 10382 7090 14672 7138
rect 10382 7088 10388 7090
rect 10092 7034 10098 7036
rect 6808 6589 7098 6637
rect 7141 6985 10098 7034
rect 7141 6539 7190 6985
rect 10092 6984 10098 6985
rect 10150 7034 10156 7036
rect 10150 6985 14462 7034
rect 10150 6984 10156 6985
rect 6794 6490 7190 6539
rect 7264 6898 7654 6902
rect 9288 6898 9294 6902
rect 7264 6858 9294 6898
rect 7264 6265 7308 6858
rect 7578 6854 9294 6858
rect 9288 6850 9294 6854
rect 9346 6898 9352 6902
rect 9346 6854 13656 6898
rect 9346 6850 9352 6854
rect 6794 6221 7308 6265
rect 7351 6776 7696 6778
rect 9044 6776 9050 6782
rect 7351 6737 9050 6776
rect 7351 6065 7392 6737
rect 7578 6735 9050 6737
rect 9044 6730 9050 6735
rect 9102 6776 9108 6782
rect 9102 6735 13410 6776
rect 9102 6730 9108 6735
rect 8230 6639 8236 6642
rect 7578 6636 8236 6639
rect 7432 6592 8236 6636
rect 7432 6586 7649 6592
rect 8230 6590 8236 6592
rect 8288 6639 8294 6642
rect 8288 6592 12579 6639
rect 8288 6590 8294 6592
rect 6796 6024 7392 6065
rect 7434 5989 7481 6586
rect 6787 5942 7481 5989
rect 7539 6471 12357 6513
rect 7539 5374 7581 6471
rect 8003 6195 8045 6471
rect 12315 6203 12357 6471
rect 12532 6346 12579 6592
rect 12500 6336 12640 6346
rect 12500 6194 12640 6204
rect 13369 6235 13410 6735
rect 13612 6340 13656 6854
rect 13560 6330 13700 6340
rect 13369 6194 13444 6235
rect 14413 6253 14462 6985
rect 14624 6340 14672 7090
rect 14602 6330 14742 6340
rect 14413 6204 14504 6253
rect 13560 6188 13700 6198
rect 14429 6195 14471 6204
rect 14602 6188 14742 6198
rect 14624 6182 14702 6188
rect 15454 6184 15510 7206
rect 15672 6354 15739 7314
rect 15634 6344 15774 6354
rect 15634 6202 15774 6212
rect 15672 6193 15739 6202
rect 6857 5332 7581 5374
rect 4995 5185 5352 5251
rect 5418 5185 5424 5251
rect 5655 5198 5721 5202
rect 5650 5193 7462 5198
rect 5053 5149 5119 5155
rect 4991 5083 5053 5149
rect 5650 5127 5655 5193
rect 5721 5127 7462 5193
rect 5650 5122 7462 5127
rect 7538 5122 7547 5198
rect 5655 5118 5721 5122
rect 5053 5077 5119 5083
rect 7186 5049 7250 5064
rect 4993 4983 5466 5049
rect 5532 4983 7250 5049
rect 7186 4968 7250 4983
rect 7346 4968 7355 5064
rect 6989 1498 6998 1674
rect 7174 1498 8456 1674
rect 11126 1426 12834 1612
rect 7692 574 7846 584
rect 12364 581 12514 1426
rect 12587 1031 12593 1181
rect 12743 1031 12749 1181
rect 7952 544 8088 554
rect 7952 422 8088 432
rect 12105 431 12111 581
rect 12261 431 12514 581
rect 7692 410 7846 420
rect 7928 360 8108 370
rect 7920 346 7928 356
rect 8108 346 8114 356
rect 7920 210 8114 220
rect 12364 -486 12514 431
rect 7984 -509 8130 -500
rect 7984 -510 8019 -509
rect 8121 -510 8130 -509
rect 7456 -606 7462 -530
rect 7538 -606 7544 -530
rect 7984 -638 8130 -628
rect 12143 -636 12149 -486
rect 12299 -636 12514 -486
rect 7962 -690 8148 -684
rect 7962 -694 8150 -690
rect 8148 -700 8150 -694
rect 8148 -836 8150 -828
rect 7962 -838 8150 -836
rect 7962 -846 8148 -838
rect 12593 -991 12743 1031
rect 12593 -1147 12743 -1141
<< via2 >>
rect 5225 6945 5339 7059
rect 5655 5127 5721 5193
rect 7462 5122 7538 5198
rect 7250 4968 7346 5064
rect 6998 1498 7174 1674
rect 7692 420 7846 574
rect 7952 432 8088 544
rect 7928 346 8108 360
rect 7928 224 8108 346
rect 8019 -510 8121 -509
rect 7467 -601 7533 -535
rect 8019 -611 8121 -510
rect 7962 -700 8148 -694
rect 7962 -828 8148 -700
rect 7962 -836 8148 -828
<< metal3 >>
rect 6655 7419 6841 7425
rect 6655 7227 6841 7233
rect 8492 7420 8680 7426
rect 5220 7059 5344 7064
rect 5220 6945 5225 7059
rect 5339 6945 5344 7059
rect 5220 6940 5344 6945
rect 5244 5748 5320 6940
rect 8492 6576 8680 7232
rect 8492 6388 12989 6576
rect 8497 5967 8675 6388
rect 12810 5921 12980 6388
rect 5244 5672 5508 5748
rect 5432 5198 5508 5672
rect 5432 5193 5726 5198
rect 5432 5127 5655 5193
rect 5721 5127 5726 5193
rect 5432 5122 5726 5127
rect 6120 4771 6216 5596
rect 7457 5198 7543 5203
rect 7457 5122 7462 5198
rect 7538 5122 7543 5198
rect 7457 5117 7543 5122
rect 7245 5064 7351 5069
rect 7245 4968 7250 5064
rect 7346 4968 7351 5064
rect 7245 4963 7351 4968
rect 6057 4765 6231 4771
rect 6057 4585 6231 4591
rect 6998 4766 7174 4794
rect 6998 1679 7174 4590
rect 6993 1674 7179 1679
rect 6993 1498 6998 1674
rect 7174 1498 7179 1674
rect 6993 1493 7179 1498
rect 7254 824 7343 4963
rect 7254 818 7356 824
rect 7254 718 7256 818
rect 7254 712 7356 718
rect 7254 -303 7343 712
rect 7254 -398 7343 -392
rect 7462 514 7538 5117
rect 7714 819 7816 825
rect 7706 717 7714 774
rect 7816 717 7824 774
rect 7706 579 7824 717
rect 7462 -535 7538 438
rect 7682 574 7856 579
rect 7682 420 7692 574
rect 7846 420 7856 574
rect 7942 544 8098 549
rect 7942 432 7952 544
rect 8088 432 8098 544
rect 7942 427 8098 432
rect 7682 415 7856 420
rect 8496 367 8666 5719
rect 7930 365 8666 367
rect 7918 360 8666 365
rect 7918 224 7928 360
rect 8108 238 8666 360
rect 8108 224 8118 238
rect 7918 219 8118 224
rect 7945 -290 8055 -285
rect 7944 -291 8126 -290
rect 7944 -401 7945 -291
rect 8055 -401 8126 -291
rect 7944 -402 8126 -401
rect 7945 -407 8126 -402
rect 7462 -601 7467 -535
rect 7533 -601 7538 -535
rect 7462 -606 7538 -601
rect 8014 -509 8126 -407
rect 8014 -611 8019 -509
rect 8121 -611 8126 -509
rect 8014 -616 8126 -611
rect 8496 -681 8666 238
rect 7947 -694 8666 -681
rect 7947 -827 7962 -694
rect 7952 -836 7962 -827
rect 8148 -827 8666 -694
rect 8148 -836 8158 -827
rect 7952 -841 8158 -836
rect 8496 -839 8666 -827
<< via3 >>
rect 6655 7233 6841 7419
rect 8492 7232 8680 7420
rect 6057 4591 6231 4765
rect 6998 4590 7174 4766
rect 7256 718 7356 818
rect 7254 -392 7343 -303
rect 7714 717 7816 819
rect 7462 438 7538 514
rect 7952 432 8088 544
rect 7945 -401 8055 -291
<< metal4 >>
rect 8491 7420 8681 7421
rect 6654 7419 8492 7420
rect 6654 7233 6655 7419
rect 6841 7233 8492 7419
rect 6654 7232 8492 7233
rect 8680 7232 8681 7420
rect 8491 7231 8681 7232
rect 6997 4766 7175 4767
rect 6056 4765 6998 4766
rect 6056 4591 6057 4765
rect 6231 4591 6998 4765
rect 6056 4590 6998 4591
rect 7174 4590 7175 4766
rect 6997 4589 7175 4590
rect 7713 819 7817 820
rect 7255 818 7714 819
rect 7255 718 7256 818
rect 7356 718 7714 818
rect 7255 717 7714 718
rect 7816 717 7817 819
rect 7713 716 7817 717
rect 7951 544 8089 545
rect 7461 514 7539 515
rect 7951 514 7952 544
rect 7461 438 7462 514
rect 7538 438 7952 514
rect 7461 437 7539 438
rect 7951 432 7952 438
rect 8088 432 8089 544
rect 7951 431 8089 432
rect 7944 -291 8119 -290
rect 7944 -302 7945 -291
rect 7253 -303 7945 -302
rect 7253 -392 7254 -303
rect 7343 -391 7945 -303
rect 7343 -392 7344 -391
rect 7253 -393 7344 -392
rect 7944 -401 7945 -391
rect 8055 -401 8119 -291
rect 7944 -402 8119 -401
use passgatesCtrlManual  x1
timestamp 1728289486
transform 0 -1 2066 1 0 4618
box 666 -4798 2906 -2962
use passgatex4  x2
timestamp 1728255086
transform 1 0 -3748 0 1 1676
box 11366 -356 15589 4682
use passgatex4  x3
timestamp 1728255086
transform 1 0 566 0 1 1678
box 11366 -356 15589 4682
use passgate  x4
timestamp 1725640011
transform 1 0 4272 0 1 -58
box 3356 -890 8072 137
use passgate  x5
timestamp 1725640011
transform 1 0 4234 0 1 1000
box 3356 -890 8072 137
<< labels >>
flabel metal2 5000 5186 5060 5248 0 FreeSans 640 0 0 0 select0
port 0 nsew
flabel metal2 5000 5084 5060 5146 0 FreeSans 640 0 0 0 select1
port 1 nsew
flabel metal2 5002 4984 5062 5046 0 FreeSans 640 0 0 0 select2
port 2 nsew
flabel metal4 6242 4596 6446 4756 0 FreeSans 640 0 0 0 VDD
port 3 nsew
flabel metal4 6822 7248 7026 7408 0 FreeSans 640 0 0 0 VSS
port 4 nsew
flabel metal1 12846 -378 13034 -198 0 FreeSans 640 0 0 0 Z
port 5 nsew
flabel metal1 7694 6150 7894 6350 0 FreeSans 640 0 0 0 A1
port 6 nsew
flabel metal1 8750 6148 8950 6348 0 FreeSans 640 0 0 0 A2
port 7 nsew
flabel metal1 9794 6144 9994 6344 0 FreeSans 640 0 0 0 A3
port 8 nsew
flabel metal1 10824 6158 11024 6358 0 FreeSans 640 0 0 0 A4
port 9 nsew
flabel metal1 12008 6152 12208 6352 0 FreeSans 640 0 0 0 A5
port 10 nsew
flabel metal1 13064 6150 13264 6350 0 FreeSans 640 0 0 0 A6
port 11 nsew
flabel metal1 14108 6146 14308 6346 0 FreeSans 640 0 0 0 A7
port 12 nsew
flabel metal1 15138 6160 15338 6360 0 FreeSans 640 0 0 0 A8
port 13 nsew
<< end >>
