* NGSPICE file created from passgatesCtrl_parax.ext - technology: sky130A

.subckt passgatesCtrl gno0 gno2 gpo0 gpo1 gpo2 gpo3 select0 VDD gno1 select1
+ gno3 VSS
X0 VSS.t57 select0.t0 a_2822_3855# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X1 VSS.t74 VDD.t88 VSS.t73 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X2 VDD.t46 a_2101_3476# gpo0.t1 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X3 net6 a_2879_2223# VDD.t38 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X4 a_2463_3073# net1 VDD.t7 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=4368,272
X5 VSS.t34 net2 a_2235_4215# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=6300,234
X6 _02_ a_1448_2473# VDD.t37 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X7 gpo3.t1 a_3431_2223# VDD.t2 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X8 VSS.t8 net1 a_1448_2473# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X9 VSS.t61 a_2101_3476# gpo0.t0 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X10 net3 net1 VSS.t5 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X11 VDD.t21 a_2835_2986# net8 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X12 VSS.t52 a_2007_4074# net4 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X13 net6 a_2879_2223# VSS.t54 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X14 a_1587_3855# a_1407_3855# VDD.t48 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=2856,152 d=2436,142
X15 net3 net2 a_1873_3561# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
**devattr s=4200,242 d=10400,504
X16 VDD.t0 a_3123_2999# _03_ _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.475 ps=2.95 w=1 l=0.15
**devattr s=19000,590 d=6662,278
X17 VDD.t39 _02_ a_1499_3311# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X18 net10 net1 a_2689_2223# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X19 gno1.t1 a_1407_2767# VDD.t15 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X20 gpo3.t0 a_3431_2223# VSS.t2 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X21 a_2427_3971# a_2235_4215# VSS.t51 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6300,234 d=2268,138
X22 VSS.t39 a_2838_4551# a_2787_4399# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3880,195
X23 a_3318_3855# a_3141_3855# VSS.t81 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X24 gno2.t1 a_2327_2223# VDD.t84 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X25 gno3.t1 a_3155_2223# VDD.t57 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X26 a_1683_3127# net1 VDD.t9 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=4704,280
X27 VDD.t83 VSS.t88 VDD.t82 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X28 a_2838_4551# a_2934_4373# VSS.t78 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=3880,195 d=4368,272
X29 a_2287_2741# net2 VDD.t28 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0 ps=0 w=0.42 l=0.15
**devattr s=9116,348 d=2436,142
X30 a_3297_3105# net2 VSS.t37 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4472,208 d=2268,138
X31 VSS.t55 _02_ a_1499_3311# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X32 VSS.t76 VDD.t89 VSS.t75 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X33 VDD.t81 VSS.t89 VDD.t80 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X34 _00_ a_2427_3971# VSS.t64 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X35 a_2287_2741# a_2463_3073# a_2415_3133# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4368,272
X36 VSS.t80 a_2287_2741# _04_ PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4052,198
X37 VSS.t28 a_2835_2986# net8 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X38 gno2.t0 a_2327_2223# VSS.t84 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X39 net1 a_2822_3855# VDD.t20 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5630,265 d=10400,504
X40 gno3.t0 a_3155_2223# VSS.t83 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X41 net10 net2 VDD.t27 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X42 VSS.t70 VDD.t90 VSS.t69 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X43 VSS.t10 net1 a_3141_3855# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X44 VDD.t17 a_3440_4551# net2 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5630,265
X45 gno1.t0 a_1407_2767# VSS.t12 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X46 VDD.t8 net1 a_2509_3971# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5930,268
X47 a_3123_2999# net2 VDD.t22 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6662,278 d=2268,138
X48 _05_ a_1587_3855# VDD.t45 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=9116,348 d=10400,504
X49 VDD.t35 a_3121_4551# a_2934_4373# FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5630,265
X50 _02_ a_1448_2473# VSS.t53 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X51 VSS.t30 net2 a_1875_2883# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X52 a_2653_3476# net3 VDD.t3 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X53 VDD.t79 VSS.t90 VDD.t78 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X54 VDD.t40 net6 a_3155_2223# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X55 a_3481_3476# net9 VDD.t53 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X56 VSS.t77 a_3318_3855# a_3424_3855# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X57 a_2415_3133# net2 VSS.t32 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0 ps=0 w=0.42 l=0.15
**devattr s=4052,198 d=2016,132
X58 a_1407_3855# net2 VSS.t36 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X59 VDD.t5 _03_ a_2879_2223# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X60 a_1530_2473# net2 a_1448_2473# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X61 a_2838_4551# a_2934_4373# VDD.t52 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=5630,265 d=4368,272
X62 VSS.t29 net2 net3 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X63 _01_ a_1875_2883# VSS.t38 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X64 a_2653_3476# net3 VSS.t3 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X65 VSS.t56 net6 a_3155_2223# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X66 a_3481_3476# net9 VSS.t79 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X67 net7 a_1499_3311# VDD.t47 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X68 a_2377_3476# net8 VDD.t1 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X69 VSS.t72 VDD.t91 VSS.t71 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X70 net9 a_3155_3311# VDD.t85 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X71 VSS.t4 _03_ a_2879_2223# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X72 VDD.t41 select0.t1 a_2822_3855# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5630,265
X73 a_1448_2473# net2 VSS.t35 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X74 VSS.t45 VDD.t92 VSS.t44 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X75 a_1957_2883# a_1683_3127# a_1875_2883# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X76 VSS.t47 VDD.t93 VSS.t46 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X77 VDD.t49 net10 a_3431_2223# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X78 a_3318_3855# a_3141_3855# VDD.t55 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5630,265 d=10400,504
X79 net7 a_1499_3311# VSS.t62 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X80 a_3601_3855# a_3424_3855# VSS.t87 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X81 a_2377_3476# net8 VSS.t1 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X82 VSS.t66 VDD.t94 VSS.t65 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X83 net5 a_2051_2223# VDD.t44 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X84 net9 a_3155_3311# VSS.t85 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X85 a_2007_4074# _05_ VDD.t32 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X86 a_2689_2223# net2 VSS.t31 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0 ps=0 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X87 VSS.t6 net1 a_2463_3073# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X88 VSS.t11 net1 a_1677_4221# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0504 ps=0.66 w=0.42 l=0.15
**devattr s=2016,132 d=4052,198
X89 a_3440_4551# select1.t0 VSS.t41 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=3880,195 d=4368,272
X90 VDD.t42 net4 a_1407_2767# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X91 a_2235_4215# net2 VDD.t25 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
**devattr s=4368,272 d=4704,280
X92 _00_ a_2427_3971# VDD.t50 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X93 VSS.t63 net10 a_3431_2223# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X94 VDD.t54 a_2287_2741# _04_ _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=9116,348
X95 VDD.t33 net5 a_2327_2223# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X96 net5 a_2051_2223# VSS.t59 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X97 VDD.t77 VSS.t91 VDD.t76 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X98 VDD.t75 VSS.t92 VDD.t74 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X99 VDD.t30 a_2838_4551# a_2787_4399# FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5630,265
X100 VSS.t68 VDD.t95 VSS.t67 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
**devattr d=5720,324
X101 VDD.t19 _00_ a_3155_3311# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X102 a_3121_4551# net2 VSS.t33 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=3880,195 d=4368,272
X103 VSS.t7 net1 a_1683_3127# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=6300,234
X104 VDD.t73 VSS.t93 VDD.t72 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X105 a_2007_4074# _05_ VSS.t43 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X106 VSS.t48 net5 a_2327_2223# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X107 a_2835_2986# _01_ VDD.t86 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X108 VDD.t11 net1 a_1587_3855# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=9116,348
X109 a_1677_4221# a_1407_3855# a_1587_3855# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2016,132
X110 VSS.t58 net4 a_1407_2767# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X111 VDD.t18 _04_ a_2051_2223# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X112 VSS.t16 _00_ a_3155_3311# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X113 VDD.t71 VSS.t94 VDD.t70 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X114 VSS.t24 VDD.t96 VSS.t23 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X115 VDD.t14 net1 a_3141_3855# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5630,265
X116 VSS.t26 VDD.t97 VSS.t25 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X117 VSS.t18 VDD.t98 VSS.t17 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X118 VSS.t9 net1 a_2427_3971# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X119 a_3440_4551# select1.t1 VDD.t43 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=5630,265 d=4368,272
X120 a_1875_2883# a_1683_3127# VSS.t40 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0 ps=0 w=0.42 l=0.15
**devattr s=6300,234 d=2268,138
X121 VSS.t0 a_3123_2999# _03_ PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
**devattr s=7280,372 d=4472,208
X122 _01_ a_1875_2883# VDD.t29 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X123 VSS.t20 VDD.t99 VSS.t19 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X124 VDD.t4 a_2463_3073# a_2287_2741# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=2856,152
X125 VDD.t56 a_2653_3476# gno0.t1 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X126 VDD.t10 net1 a_1530_2473# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X127 VDD.t34 a_3481_3476# gpo2.t1 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X128 VSS.t15 _04_ a_2051_2223# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X129 a_3123_2999# net1 a_3297_3105# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X130 VSS.t14 a_3440_4551# net2 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3880,195
X131 a_2835_2986# _01_ VSS.t86 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X132 a_2101_3476# net7 VDD.t31 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X133 VDD.t69 VSS.t95 VDD.t68 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
**devattr d=9048,452
X134 a_3121_4551# net2 VDD.t23 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
**devattr s=5630,265 d=4368,272
X135 VDD.t51 a_3318_3855# a_3424_3855# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5630,265
X136 VDD.t13 net1 net10 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X137 VDD.t26 net2 a_1407_3855# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2856,152
X138 VSS.t82 a_2653_3476# gno0.t0 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X139 VSS.t49 a_3481_3476# gpo2.t0 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X140 VSS.t50 a_3121_4551# a_2934_4373# PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3880,195
X141 a_3601_3855# a_3424_3855# VDD.t87 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
**devattr s=5630,265 d=10400,504
X142 VDD.t24 net2 a_1957_2883# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5930,268
X143 VDD.t67 VSS.t96 VDD.t66 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X144 VDD.t16 a_2377_3476# gpo1.t1 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X145 a_2509_3971# a_2235_4215# a_2427_3971# _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X146 VDD.t6 net1 a_3123_2999# _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4704,280
X147 a_2101_3476# net7 VSS.t42 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X148 net1 a_2822_3855# VSS.t27 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X149 VDD.t65 VSS.t97 VDD.t64 FILLER_0_4_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X150 VDD.t63 VSS.t98 VDD.t62 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X151 VDD.t61 VSS.t99 VDD.t60 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X152 VDD.t59 VSS.t100 VDD.t58 _09_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
**devattr d=9048,452
X153 VSS.t13 a_2377_3476# gpo1.t0 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
X154 _05_ a_1587_3855# VSS.t60 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
**devattr s=4052,198 d=6760,364
X155 VSS.t22 VDD.t100 VSS.t21 PHY_EDGE_ROW_4_Right_4.VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
**devattr d=5720,324
X156 VDD.t36 a_2007_4074# net4 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X157 a_1873_3561# net1 VDD.t12 _12_.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=4200,242
R0 select0.n0 select0.t1 323.55
R1 select0.n0 select0.t0 195.017
R2 select0.n1 select0.n0 152.792
R3 select0 select0.n1 9.4552
R4 select0.n1 select0 2.2438
R5 VSS.n200 VSS.t92 262.784
R6 VSS.n201 VSS.t93 262.784
R7 VSS.n262 VSS.t98 262.784
R8 VSS.n263 VSS.t100 262.784
R9 VSS.n45 VSS.t97 262.784
R10 VSS.n46 VSS.t99 262.784
R11 VSS.n301 VSS.t88 262.784
R12 VSS.n302 VSS.t89 262.784
R13 VSS.n311 VSS.t95 262.719
R14 VSS.n229 VSS.t96 259.082
R15 VSS.n95 VSS.t90 259.082
R16 VSS.n150 VSS.t91 259.082
R17 VSS.n335 VSS.t94 259.082
R18 VSS.n146 VSS.t35 246.506
R19 VSS.n238 VSS.t6 237.327
R20 VSS.n300 VSS.t36 237.327
R21 VSS.n7 VSS.t67 218.203
R22 VSS.n230 VSS.t18 214.456
R23 VSS.n26 VSS.t17 214.456
R24 VSS.n200 VSS.t47 214.456
R25 VSS.n200 VSS.t46 214.456
R26 VSS.n201 VSS.t72 214.456
R27 VSS.n201 VSS.t71 214.456
R28 VSS.n262 VSS.t20 214.456
R29 VSS.n262 VSS.t19 214.456
R30 VSS.n263 VSS.t26 214.456
R31 VSS.n263 VSS.t25 214.456
R32 VSS.n149 VSS.t45 214.456
R33 VSS.n147 VSS.t44 214.456
R34 VSS.n99 VSS.t76 214.456
R35 VSS.n96 VSS.t75 214.456
R36 VSS.n299 VSS.t68 214.456
R37 VSS.n334 VSS.t66 214.456
R38 VSS.n338 VSS.t65 214.456
R39 VSS.n45 VSS.t24 214.456
R40 VSS.n45 VSS.t23 214.456
R41 VSS.n46 VSS.t22 214.456
R42 VSS.n46 VSS.t21 214.456
R43 VSS.n301 VSS.t74 214.456
R44 VSS.n301 VSS.t73 214.456
R45 VSS.n302 VSS.t70 214.456
R46 VSS.n302 VSS.t69 214.456
R47 VSS.n160 VSS.n144 210.601
R48 VSS.n247 VSS.n246 200.231
R49 VSS.n29 VSS.n28 200.105
R50 VSS.n198 VSS.n197 199.739
R51 VSS.n245 VSS.n244 199.739
R52 VSS.n251 VSS.n21 199.739
R53 VSS.n269 VSS.n258 199.739
R54 VSS.n268 VSS.n261 199.739
R55 VSS.n93 VSS.n92 199.739
R56 VSS.n90 VSS.n89 199.739
R57 VSS.n185 VSS.n120 199.739
R58 VSS.n124 VSS.n123 199.739
R59 VSS.n126 VSS.n125 199.739
R60 VSS.n253 VSS.n252 198.475
R61 VSS.n312 VSS.n297 197.476
R62 VSS.n239 VSS.n24 196.442
R63 VSS.n209 VSS.n208 196.442
R64 VSS.n9 VSS.n8 196.442
R65 VSS.n336 VSS.n3 195.612
R66 VSS.n44 VSS.n43 194.809
R67 VSS.n52 VSS.n51 194.809
R68 VSS.n60 VSS.n41 194.809
R69 VSS.n59 VSS.n42 194.809
R70 VSS.n65 VSS.n62 194.809
R71 VSS.n64 VSS.n63 194.809
R72 VSS.n232 VSS.n231 189.335
R73 VSS.n232 VSS.n25 176
R74 VSS.n281 VSS.t29 156.915
R75 VSS.n179 VSS.t31 150.922
R76 VSS.n271 VSS.t5 150.101
R77 VSS.n333 VSS.n5 100.331
R78 VSS.n254 VSS.t7 89.3033
R79 VSS.n254 VSS.t40 88.8109
R80 VSS.n4 VSS.t51 88.6006
R81 VSS.n4 VSS.t34 88.6006
R82 VSS.n28 VSS.t37 72.8576
R83 VSS.n255 VSS.n254 70.457
R84 VSS.n5 VSS.n4 70.4126
R85 VSS.n246 VSS.t32 58.5719
R86 VSS.n297 VSS.t11 58.5719
R87 VSS.n144 VSS.t8 55.7148
R88 VSS.n252 VSS.t30 52.8576
R89 VSS.n3 VSS.t9 52.8576
R90 VSS.n43 VSS.t41 45.7148
R91 VSS.n51 VSS.t77 45.7148
R92 VSS.n41 VSS.t33 45.7148
R93 VSS.n42 VSS.t10 45.7148
R94 VSS.n62 VSS.t78 45.7148
R95 VSS.n63 VSS.t57 45.7148
R96 VSS.n210 VSS.n209 34.6358
R97 VSS.n239 VSS.n237 34.6358
R98 VSS.n53 VSS.n50 34.6358
R99 VSS.n66 VSS.n2 34.6358
R100 VSS.n210 VSS.n207 34.6358
R101 VSS.n243 VSS.n23 34.6358
R102 VSS.n271 VSS.n270 34.6358
R103 VSS.n106 VSS.n105 34.6358
R104 VSS.n186 VSS.n119 34.6358
R105 VSS.n184 VSS.n121 34.6358
R106 VSS.n180 VSS.n121 34.6358
R107 VSS.n174 VSS.n173 34.6358
R108 VSS.n134 VSS.n133 34.6358
R109 VSS.n143 VSS.n134 34.6358
R110 VSS.n162 VSS.n143 34.6358
R111 VSS.n162 VSS.n161 34.6358
R112 VSS.n159 VSS.n145 34.6358
R113 VSS.n57 VSS.n56 34.6358
R114 VSS.n58 VSS.n57 34.6358
R115 VSS.n71 VSS.n70 34.6358
R116 VSS.n70 VSS.n61 34.6358
R117 VSS.n43 VSS.t14 34.506
R118 VSS.n51 VSS.t87 34.506
R119 VSS.n41 VSS.t50 34.506
R120 VSS.n42 VSS.t81 34.506
R121 VSS.n62 VSS.t39 34.506
R122 VSS.n63 VSS.t27 34.506
R123 VSS.n24 VSS.t3 33.462
R124 VSS.n24 VSS.t82 33.462
R125 VSS.n208 VSS.t85 33.462
R126 VSS.n208 VSS.t16 33.462
R127 VSS.n231 VSS.t86 33.462
R128 VSS.n231 VSS.t28 33.462
R129 VSS.n197 VSS.t79 33.462
R130 VSS.n197 VSS.t49 33.462
R131 VSS.n244 VSS.t1 33.462
R132 VSS.n244 VSS.t13 33.462
R133 VSS.n21 VSS.t42 33.462
R134 VSS.n21 VSS.t61 33.462
R135 VSS.n258 VSS.t62 33.462
R136 VSS.n258 VSS.t55 33.462
R137 VSS.n261 VSS.t12 33.462
R138 VSS.n261 VSS.t58 33.462
R139 VSS.n92 VSS.t2 33.462
R140 VSS.n92 VSS.t63 33.462
R141 VSS.n89 VSS.t83 33.462
R142 VSS.n89 VSS.t56 33.462
R143 VSS.n120 VSS.t54 33.462
R144 VSS.n120 VSS.t4 33.462
R145 VSS.n123 VSS.t84 33.462
R146 VSS.n123 VSS.t48 33.462
R147 VSS.n125 VSS.t59 33.462
R148 VSS.n125 VSS.t15 33.462
R149 VSS.n8 VSS.t43 33.462
R150 VSS.n8 VSS.t52 33.462
R151 VSS.n238 VSS.n23 32.377
R152 VSS.n252 VSS.t38 27.5691
R153 VSS.n3 VSS.t64 27.5691
R154 VSS.n144 VSS.t53 26.8576
R155 VSS.n60 VSS.n59 26.7299
R156 VSS.n281 VSS.n280 25.977
R157 VSS.n225 VSS.n224 25.7355
R158 VSS.n101 VSS.n100 25.7355
R159 VSS.n155 VSS.n154 25.7355
R160 VSS.n339 VSS.n2 25.7355
R161 VSS.n246 VSS.t80 25.4291
R162 VSS.n297 VSS.t60 25.4291
R163 VSS.n203 VSS.n202 23.7181
R164 VSS.n267 VSS.n264 23.7181
R165 VSS.n179 VSS.n178 23.7181
R166 VSS.n50 VSS.n47 23.7181
R167 VSS.n28 VSS.t0 22.3257
R168 VSS.n203 VSS.n198 22.2123
R169 VSS.n207 VSS.n198 22.2123
R170 VSS.n237 VSS.n25 22.2123
R171 VSS.n245 VSS.n243 22.2123
R172 VSS.n251 VSS.n20 22.2123
R173 VSS.n270 VSS.n269 22.2123
R174 VSS.n268 VSS.n267 22.2123
R175 VSS.n101 VSS.n93 22.2123
R176 VSS.n105 VSS.n93 22.2123
R177 VSS.n106 VSS.n90 22.2123
R178 VSS.n119 VSS.n90 22.2123
R179 VSS.n186 VSS.n185 22.2123
R180 VSS.n185 VSS.n184 22.2123
R181 VSS.n180 VSS.n179 22.2123
R182 VSS.n178 VSS.n124 22.2123
R183 VSS.n174 VSS.n124 22.2123
R184 VSS.n173 VSS.n126 22.2123
R185 VSS.n133 VSS.n126 22.2123
R186 VSS.n247 VSS.n20 21.4593
R187 VSS.n64 VSS.n61 20.3299
R188 VSS.n271 VSS.n255 19.9534
R189 VSS.n56 VSS.n44 19.9534
R190 VSS.n224 VSS.n29 18.824
R191 VSS.n161 VSS.n160 16.1887
R192 VSS.n209 VSS.n29 15.8123
R193 VSS.n305 VSS.n304 15.3963
R194 VSS.n146 VSS.n145 15.0593
R195 VSS.n280 VSS.n255 14.6829
R196 VSS.n52 VSS.n44 13.177
R197 VSS.n65 VSS.n64 13.177
R198 VSS.n253 VSS.n251 11.2946
R199 VSS.n269 VSS.n268 9.78874
R200 VSS VSS.n96 9.74003
R201 VSS.n149 VSS.n148 9.71789
R202 VSS.n204 VSS.n203 9.3005
R203 VSS.n205 VSS.n198 9.3005
R204 VSS.n207 VSS.n206 9.3005
R205 VSS.n211 VSS.n210 9.3005
R206 VSS.n209 VSS.n30 9.3005
R207 VSS.n224 VSS.n223 9.3005
R208 VSS.n226 VSS.n225 9.3005
R209 VSS.n228 VSS.n227 9.3005
R210 VSS.n235 VSS.n234 9.3005
R211 VSS.n237 VSS.n236 9.3005
R212 VSS.n240 VSS.n239 9.3005
R213 VSS.n241 VSS.n23 9.3005
R214 VSS.n243 VSS.n242 9.3005
R215 VSS.n245 VSS.n22 9.3005
R216 VSS.n248 VSS.n247 9.3005
R217 VSS.n249 VSS.n20 9.3005
R218 VSS.n251 VSS.n250 9.3005
R219 VSS.n253 VSS.n18 9.3005
R220 VSS.n282 VSS.n281 9.3005
R221 VSS.n280 VSS.n279 9.3005
R222 VSS.n272 VSS.n271 9.3005
R223 VSS.n270 VSS.n257 9.3005
R224 VSS.n269 VSS.n259 9.3005
R225 VSS.n268 VSS.n260 9.3005
R226 VSS.n267 VSS.n266 9.3005
R227 VSS.n152 VSS.n151 9.3005
R228 VSS.n154 VSS.n153 9.3005
R229 VSS.n98 VSS.n97 9.3005
R230 VSS.n100 VSS.n94 9.3005
R231 VSS.n102 VSS.n101 9.3005
R232 VSS.n103 VSS.n93 9.3005
R233 VSS.n105 VSS.n104 9.3005
R234 VSS.n107 VSS.n106 9.3005
R235 VSS.n116 VSS.n90 9.3005
R236 VSS.n119 VSS.n118 9.3005
R237 VSS.n187 VSS.n186 9.3005
R238 VSS.n185 VSS.n88 9.3005
R239 VSS.n184 VSS.n183 9.3005
R240 VSS.n182 VSS.n121 9.3005
R241 VSS.n181 VSS.n180 9.3005
R242 VSS.n179 VSS.n122 9.3005
R243 VSS.n178 VSS.n177 9.3005
R244 VSS.n176 VSS.n124 9.3005
R245 VSS.n175 VSS.n174 9.3005
R246 VSS.n173 VSS.n172 9.3005
R247 VSS.n171 VSS.n126 9.3005
R248 VSS.n133 VSS.n127 9.3005
R249 VSS.n136 VSS.n134 9.3005
R250 VSS.n143 VSS.n142 9.3005
R251 VSS.n163 VSS.n162 9.3005
R252 VSS.n161 VSS.n132 9.3005
R253 VSS.n159 VSS.n158 9.3005
R254 VSS.n157 VSS.n145 9.3005
R255 VSS.n156 VSS.n155 9.3005
R256 VSS.n306 VSS.n305 9.3005
R257 VSS.n307 VSS.n298 9.3005
R258 VSS.n309 VSS.n308 9.3005
R259 VSS.n310 VSS.n294 9.3005
R260 VSS.n314 VSS.n313 9.3005
R261 VSS.n296 VSS.n293 9.3005
R262 VSS.n295 VSS.n292 9.3005
R263 VSS.n10 VSS.n9 9.3005
R264 VSS.n329 VSS.n328 9.3005
R265 VSS.n331 VSS.n330 9.3005
R266 VSS.n50 VSS.n49 9.3005
R267 VSS.n54 VSS.n53 9.3005
R268 VSS.n56 VSS.n55 9.3005
R269 VSS.n57 VSS.n37 9.3005
R270 VSS.n58 VSS.n38 9.3005
R271 VSS.n72 VSS.n71 9.3005
R272 VSS.n70 VSS.n69 9.3005
R273 VSS.n68 VSS.n61 9.3005
R274 VSS.n67 VSS.n66 9.3005
R275 VSS.n2 VSS.n0 9.3005
R276 VSS.n340 VSS.n339 9.3005
R277 VSS.n337 VSS.n1 9.3005
R278 VSS.n333 VSS 9.3005
R279 VSS.n330 VSS.n329 8.23546
R280 VSS.n329 VSS.n9 8.23546
R281 VSS.n295 VSS.n9 8.23546
R282 VSS.n296 VSS.n295 8.23546
R283 VSS.n313 VSS.n296 8.23546
R284 VSS.n310 VSS.n309 8.23546
R285 VSS.n309 VSS.n298 8.23546
R286 VSS.n233 VSS.n232 7.84566
R287 VSS.n299 VSS.n298 7.6984
R288 VSS.n281 VSS.n253 7.52991
R289 VSS.n330 VSS.n7 6.44526
R290 VSS.n228 VSS.n26 5.98311
R291 VSS.n99 VSS.n98 5.98311
R292 VSS.n151 VSS.n147 5.98311
R293 VSS.n338 VSS.n337 5.98311
R294 VSS.n247 VSS.n245 5.64756
R295 VSS.n202 VSS.n200 5.13108
R296 VSS.n202 VSS.n201 5.13108
R297 VSS.n264 VSS.n262 5.13108
R298 VSS.n264 VSS.n263 5.13108
R299 VSS.n47 VSS.n45 5.13108
R300 VSS.n47 VSS.n46 5.13108
R301 VSS.n304 VSS.n301 5.13108
R302 VSS.n304 VSS.n302 5.13108
R303 VSS.n7 VSS.n6 4.93764
R304 VSS.n229 VSS.n228 4.8005
R305 VSS.n98 VSS.n95 4.8005
R306 VSS.n151 VSS.n150 4.8005
R307 VSS.n332 VSS.n6 4.62124
R308 VSS.n81 VSS.n35 4.51401
R309 VSS.n40 VSS.n39 4.51401
R310 VSS.n285 VSS.n16 4.51401
R311 VSS.n278 VSS.n277 4.51401
R312 VSS.n216 VSS.n195 4.51401
R313 VSS.n220 VSS.n27 4.51401
R314 VSS.n109 VSS.n108 4.51401
R315 VSS.n189 VSS.n188 4.51401
R316 VSS.n170 VSS.n169 4.51401
R317 VSS.n165 VSS.n164 4.51401
R318 VSS.n327 VSS.n326 4.51401
R319 VSS.n318 VSS.n315 4.51401
R320 VSS.n276 VSS.n256 4.5005
R321 VSS.n284 VSS.n283 4.5005
R322 VSS.n273 VSS.n19 4.5005
R323 VSS.n215 VSS.n214 4.5005
R324 VSS.n213 VSS.n212 4.5005
R325 VSS.n222 VSS.n221 4.5005
R326 VSS.n110 VSS.n91 4.5005
R327 VSS.n115 VSS.n114 4.5005
R328 VSS.n117 VSS.n87 4.5005
R329 VSS.n141 VSS.n131 4.5005
R330 VSS.n135 VSS.n128 4.5005
R331 VSS.n140 VSS.n139 4.5005
R332 VSS.n291 VSS.n11 4.5005
R333 VSS.n322 VSS.n321 4.5005
R334 VSS.n320 VSS.n319 4.5005
R335 VSS.n80 VSS.n79 4.5005
R336 VSS.n78 VSS.n77 4.5005
R337 VSS.n74 VSS.n73 4.5005
R338 VSS.n6 VSS.n5 4.38907
R339 VSS.n336 VSS.n335 4.17441
R340 VSS.n59 VSS.n58 4.14168
R341 VSS.n311 VSS.n310 4.11798
R342 VSS.n71 VSS.n60 3.76521
R343 VSS.n312 VSS.n311 3.67043
R344 VSS.n39 VSS.n33 3.43925
R345 VSS.n82 VSS.n81 3.43925
R346 VSS.n277 VSS.n13 3.43925
R347 VSS.n286 VSS.n285 3.43925
R348 VSS.n220 VSS.n219 3.43925
R349 VSS.n217 VSS.n216 3.43925
R350 VSS.n166 VSS.n165 3.43925
R351 VSS.n169 VSS.n168 3.43925
R352 VSS.n36 VSS.n34 3.4105
R353 VSS.n76 VSS.n75 3.4105
R354 VSS.n17 VSS.n15 3.4105
R355 VSS.n275 VSS.n274 3.4105
R356 VSS.n196 VSS.n194 3.4105
R357 VSS.n32 VSS.n31 3.4105
R358 VSS.n191 VSS.n190 3.4105
R359 VSS.n191 VSS.n85 3.4105
R360 VSS.n190 VSS.n189 3.4105
R361 VSS.n109 VSS.n85 3.4105
R362 VSS.n112 VSS.n111 3.4105
R363 VSS.n113 VSS.n86 3.4105
R364 VSS.n137 VSS.n129 3.4105
R365 VSS.n138 VSS.n130 3.4105
R366 VSS.n317 VSS.n288 3.4105
R367 VSS.n325 VSS.n288 3.4105
R368 VSS.n318 VSS.n317 3.4105
R369 VSS.n326 VSS.n325 3.4105
R370 VSS.n324 VSS.n323 3.4105
R371 VSS.n316 VSS.n290 3.4105
R372 VSS.n202 VSS.n199 3.05586
R373 VSS.n48 VSS.n47 3.05586
R374 VSS.n265 VSS.n264 3.04861
R375 VSS.n304 VSS.n303 3.04861
R376 VSS.n239 VSS.n238 2.25932
R377 VSS.n160 VSS.n159 2.25932
R378 VSS.n234 VSS.n25 2.01789
R379 VSS.n219 VSS.n218 1.69188
R380 VSS.n218 VSS.n217 1.69188
R381 VSS.n83 VSS.n33 1.69188
R382 VSS.n83 VSS.n82 1.69188
R383 VSS.n191 VSS.n84 1.69188
R384 VSS.n167 VSS.n166 1.69188
R385 VSS.n168 VSS.n167 1.69188
R386 VSS.n287 VSS.n13 1.69188
R387 VSS.n287 VSS.n286 1.69188
R388 VSS.n289 VSS.n288 1.69188
R389 VSS.n155 VSS.n146 1.50638
R390 VSS.n53 VSS.n52 1.50638
R391 VSS.n230 VSS.n229 1.18311
R392 VSS.n96 VSS.n95 1.18311
R393 VSS.n150 VSS.n149 1.18311
R394 VSS.n335 VSS.n334 1.18311
R395 VSS.n66 VSS.n65 1.12991
R396 VSS.n337 VSS.n336 0.626587
R397 VSS.n83 VSS.n12 0.500712
R398 VSS.n193 VSS.n192 0.500125
R399 VSS.n313 VSS.n312 0.448052
R400 VSS.n305 VSS.n300 0.448052
R401 VSS.n225 VSS.n26 0.417891
R402 VSS.n100 VSS.n99 0.417891
R403 VSS.n154 VSS.n147 0.417891
R404 VSS.n339 VSS.n338 0.417891
R405 VSS.n334 VSS.n333 0.417891
R406 VSS.n288 VSS.n12 0.381087
R407 VSS.n192 VSS.n14 0.3805
R408 VSS.n233 VSS.n230 0.278761
R409 VSS.n204 VSS.n199 0.232472
R410 VSS.n49 VSS.n48 0.232472
R411 VSS.n303 VSS 0.217246
R412 VSS VSS.n265 0.208476
R413 VSS.n332 VSS.n331 0.180304
R414 VSS.n218 VSS.n83 0.1603
R415 VSS.n288 VSS.n287 0.1603
R416 VSS VSS.n332 0.158169
R417 VSS.n303 VSS 0.14207
R418 VSS.n265 VSS 0.141725
R419 VSS.n234 VSS.n233 0.13963
R420 VSS.n193 VSS.n191 0.126812
R421 VSS.n167 VSS.n14 0.126812
R422 VSS.n227 VSS.n226 0.120292
R423 VSS.n242 VSS.n241 0.120292
R424 VSS.n248 VSS.n22 0.120292
R425 VSS.n249 VSS.n248 0.120292
R426 VSS.n272 VSS.n257 0.120292
R427 VSS.n260 VSS.n259 0.120292
R428 VSS.n97 VSS.n94 0.120292
R429 VSS.n102 VSS.n94 0.120292
R430 VSS.n103 VSS.n102 0.120292
R431 VSS.n104 VSS.n103 0.120292
R432 VSS.n187 VSS.n88 0.120292
R433 VSS.n183 VSS.n88 0.120292
R434 VSS.n182 VSS.n181 0.120292
R435 VSS.n181 VSS.n122 0.120292
R436 VSS.n177 VSS.n176 0.120292
R437 VSS.n176 VSS.n175 0.120292
R438 VSS.n172 VSS.n171 0.120292
R439 VSS.n163 VSS.n132 0.120292
R440 VSS.n158 VSS.n132 0.120292
R441 VSS.n158 VSS.n157 0.120292
R442 VSS.n157 VSS.n156 0.120292
R443 VSS.n153 VSS.n152 0.120292
R444 VSS.n152 VSS.n148 0.120292
R445 VSS.n55 VSS.n54 0.120292
R446 VSS.n69 VSS.n68 0.120292
R447 VSS.n68 VSS.n67 0.120292
R448 VSS.n67 VSS.n0 0.120292
R449 VSS.n340 VSS.n1 0.120292
R450 VSS VSS.n1 0.120292
R451 VSS.n314 VSS.n294 0.120292
R452 VSS.n308 VSS.n294 0.120292
R453 VSS.n308 VSS.n307 0.120292
R454 VSS.n307 VSS.n306 0.120292
R455 VSS.n199 VSS 0.105238
R456 VSS.n48 VSS 0.105238
R457 VSS.n54 VSS 0.104667
R458 VSS.n172 VSS 0.10076
R459 VSS.n259 VSS 0.0994583
R460 VSS.n328 VSS 0.0994583
R461 VSS.n235 VSS 0.0981562
R462 VSS.n236 VSS 0.0981562
R463 VSS.n241 VSS 0.0981562
R464 VSS.n266 VSS 0.0981562
R465 VSS.n97 VSS 0.0981562
R466 VSS VSS.n182 0.0981562
R467 VSS.n153 VSS 0.0981562
R468 VSS.n226 VSS.n27 0.0968542
R469 VSS.n188 VSS.n187 0.0968542
R470 VSS.n177 VSS 0.0968542
R471 VSS.n69 VSS.n40 0.0968542
R472 VSS.n205 VSS 0.0955521
R473 VSS.n240 VSS 0.0955521
R474 VSS VSS.n22 0.0955521
R475 VSS.n250 VSS 0.0955521
R476 VSS.n81 VSS.n80 0.0950946
R477 VSS.n74 VSS.n39 0.0950946
R478 VSS.n285 VSS.n284 0.0950946
R479 VSS.n277 VSS.n276 0.0950946
R480 VSS.n216 VSS.n215 0.0950946
R481 VSS.n221 VSS.n220 0.0950946
R482 VSS.n110 VSS.n109 0.0950946
R483 VSS.n189 VSS.n87 0.0950946
R484 VSS.n169 VSS.n128 0.0950946
R485 VSS.n165 VSS.n131 0.0950946
R486 VSS.n326 VSS.n11 0.0950946
R487 VSS.n319 VSS.n318 0.0950946
R488 VSS.n250 VSS.n16 0.0916458
R489 VSS.n171 VSS.n170 0.0916458
R490 VSS VSS.n340 0.0916458
R491 VSS.n300 VSS.n299 0.0900105
R492 VSS.n206 VSS 0.0864375
R493 VSS.n214 VSS.n213 0.0838333
R494 VSS.n115 VSS.n91 0.0838333
R495 VSS.n141 VSS.n140 0.0838333
R496 VSS.n79 VSS.n78 0.0838333
R497 VSS.n321 VSS.n320 0.0838333
R498 VSS.n12 VSS 0.0827875
R499 VSS.n192 VSS 0.0827875
R500 VSS.n256 VSS 0.078625
R501 VSS.n211 VSS.n195 0.0708125
R502 VSS.n108 VSS.n107 0.0708125
R503 VSS.n37 VSS.n35 0.0708125
R504 VSS VSS.n327 0.0695104
R505 VSS.n77 VSS.n36 0.0680676
R506 VSS.n77 VSS.n76 0.0680676
R507 VSS.n273 VSS.n17 0.0680676
R508 VSS.n275 VSS.n273 0.0680676
R509 VSS.n212 VSS.n196 0.0680676
R510 VSS.n212 VSS.n31 0.0680676
R511 VSS.n114 VSS.n112 0.0680676
R512 VSS.n114 VSS.n113 0.0680676
R513 VSS.n139 VSS.n137 0.0680676
R514 VSS.n139 VSS.n138 0.0680676
R515 VSS.n323 VSS.n322 0.0680676
R516 VSS.n322 VSS.n290 0.0680676
R517 VSS.n283 VSS.n282 0.0656042
R518 VSS.n279 VSS.n278 0.0656042
R519 VSS.n136 VSS.n135 0.0656042
R520 VSS.n292 VSS.n291 0.0656042
R521 VSS.n315 VSS.n293 0.0656042
R522 VSS.n222 VSS.n30 0.0603958
R523 VSS.n223 VSS.n222 0.0603958
R524 VSS.n117 VSS.n116 0.0603958
R525 VSS.n118 VSS.n117 0.0603958
R526 VSS.n73 VSS.n38 0.0603958
R527 VSS.n73 VSS.n72 0.0603958
R528 VSS.n75 VSS.n34 0.0574697
R529 VSS.n274 VSS.n15 0.0574697
R530 VSS.n194 VSS.n32 0.0574697
R531 VSS.n111 VSS.n85 0.0574697
R532 VSS.n190 VSS.n86 0.0574697
R533 VSS.n130 VSS.n129 0.0574697
R534 VSS.n325 VSS.n324 0.0574697
R535 VSS.n317 VSS.n316 0.0574697
R536 VSS.n283 VSS.n18 0.0551875
R537 VSS.n278 VSS.n272 0.0551875
R538 VSS.n164 VSS.n163 0.0551875
R539 VSS.n291 VSS.n10 0.0551875
R540 VSS.n315 VSS.n314 0.0551875
R541 VSS.n55 VSS.n35 0.0499792
R542 VSS.n80 VSS.n36 0.0410405
R543 VSS.n76 VSS.n74 0.0410405
R544 VSS.n284 VSS.n17 0.0410405
R545 VSS.n276 VSS.n275 0.0410405
R546 VSS.n215 VSS.n196 0.0410405
R547 VSS.n221 VSS.n31 0.0410405
R548 VSS.n112 VSS.n110 0.0410405
R549 VSS.n113 VSS.n87 0.0410405
R550 VSS.n137 VSS.n128 0.0410405
R551 VSS.n138 VSS.n131 0.0410405
R552 VSS.n323 VSS.n11 0.0410405
R553 VSS.n319 VSS.n290 0.0410405
R554 VSS VSS.n205 0.0343542
R555 VSS.n142 VSS 0.0343542
R556 VSS.n218 VSS.n193 0.0339875
R557 VSS.n287 VSS.n14 0.0339875
R558 VSS.n135 VSS 0.0330521
R559 VSS.n164 VSS 0.03175
R560 VSS.n108 VSS 0.0304479
R561 VSS.n217 VSS.n194 0.0292489
R562 VSS.n219 VSS.n32 0.0292489
R563 VSS.n82 VSS.n34 0.0292489
R564 VSS.n75 VSS.n33 0.0292489
R565 VSS.n86 VSS.n84 0.0292489
R566 VSS.n111 VSS.n84 0.0292489
R567 VSS.n168 VSS.n129 0.0292489
R568 VSS.n166 VSS.n130 0.0292489
R569 VSS.n286 VSS.n15 0.0292489
R570 VSS.n274 VSS.n13 0.0292489
R571 VSS.n316 VSS.n289 0.0292489
R572 VSS.n324 VSS.n289 0.0292489
R573 VSS.n18 VSS.n16 0.0291458
R574 VSS.n170 VSS.n127 0.0291458
R575 VSS VSS.n0 0.0291458
R576 VSS.n327 VSS.n10 0.0291458
R577 VSS VSS.n195 0.0278438
R578 VSS VSS.n204 0.0252396
R579 VSS.n236 VSS 0.0252396
R580 VSS.n242 VSS 0.0252396
R581 VSS VSS.n249 0.0252396
R582 VSS.n213 VSS.n30 0.0239375
R583 VSS.n116 VSS.n115 0.0239375
R584 VSS VSS.n122 0.0239375
R585 VSS.n78 VSS.n38 0.0239375
R586 VSS.n72 VSS.n40 0.0239375
R587 VSS.n206 VSS 0.0226354
R588 VSS.n223 VSS 0.0226354
R589 VSS.n227 VSS 0.0226354
R590 VSS VSS.n235 0.0226354
R591 VSS VSS.n240 0.0226354
R592 VSS VSS.n260 0.0226354
R593 VSS.n183 VSS 0.0226354
R594 VSS VSS.n127 0.0226354
R595 VSS.n156 VSS 0.0226354
R596 VSS.n148 VSS 0.0226354
R597 VSS.n328 VSS 0.0226354
R598 VSS.n306 VSS 0.0226354
R599 VSS VSS.n257 0.0213333
R600 VSS.n331 VSS 0.0213333
R601 VSS.n266 VSS 0.0200312
R602 VSS.n104 VSS 0.0200312
R603 VSS.n118 VSS 0.0200312
R604 VSS.n175 VSS 0.0200312
R605 VSS.n282 VSS.n19 0.0187292
R606 VSS.n279 VSS.n256 0.0187292
R607 VSS.n140 VSS.n136 0.0187292
R608 VSS.n142 VSS.n141 0.0187292
R609 VSS.n321 VSS.n292 0.0187292
R610 VSS.n320 VSS.n293 0.0187292
R611 VSS.n49 VSS 0.016125
R612 VSS.n214 VSS.n211 0.0135208
R613 VSS.n107 VSS.n91 0.0135208
R614 VSS.n79 VSS.n37 0.0135208
R615 VSS.n191 VSS 0.00755
R616 VSS.n167 VSS 0.00755
R617 VSS VSS.n19 0.00570833
R618 VSS.n188 VSS 0.00440625
R619 VSS VSS.n27 0.00180208
R620 VDD.n13 VDD.t61 804.731
R621 VDD.n18 VDD.t75 804.731
R622 VDD.n30 VDD.t67 804.731
R623 VDD.n58 VDD.t81 804.731
R624 VDD.n61 VDD.t63 804.731
R625 VDD.n208 VDD.t73 804.731
R626 VDD.n232 VDD.t79 804.731
R627 VDD.n276 VDD.t59 804.731
R628 VDD.n284 VDD.t77 804.731
R629 VDD.n167 VDD.t69 804.731
R630 VDD.n148 VDD.t68 804.731
R631 VDD.t61 VDD.n12 725.173
R632 VDD.t75 VDD.n17 725.173
R633 VDD.t67 VDD.n29 725.173
R634 VDD.t81 VDD.n57 725.173
R635 VDD.t63 VDD.n60 725.173
R636 VDD.t73 VDD.n207 725.173
R637 VDD.t79 VDD.n231 725.173
R638 VDD.t59 VDD.n275 725.173
R639 VDD.t77 VDD.n283 725.173
R640 VDD.n352 VDD.t25 701.529
R641 VDD.n299 VDD.t9 697.264
R642 VDD.n239 VDD.t6 675.293
R643 VDD.n341 VDD.n54 602.456
R644 VDD.n255 VDD.n254 602.456
R645 VDD.n21 VDD.n19 596.97
R646 VDD.n374 VDD.n26 595.043
R647 VDD.n25 VDD.n24 594.144
R648 VDD.n124 VDD.n123 585
R649 VDD.n101 VDD.n100 585
R650 VDD.n104 VDD.n103 585
R651 VDD.n168 VDD.t82 381.443
R652 VDD.n132 VDD.t70 381.443
R653 VDD.n91 VDD.t71 381.443
R654 VDD.n105 VDD.t64 381.443
R655 VDD.n108 VDD.t65 381.443
R656 VDD.n181 VDD.t83 381.443
R657 VDD.n11 VDD.t60 380.193
R658 VDD.n16 VDD.t74 380.193
R659 VDD.n28 VDD.t66 380.193
R660 VDD.n56 VDD.t80 380.193
R661 VDD.n59 VDD.t62 380.193
R662 VDD.n206 VDD.t72 380.193
R663 VDD.n230 VDD.t78 380.193
R664 VDD.n274 VDD.t58 380.193
R665 VDD.n282 VDD.t76 380.193
R666 VDD.n200 VDD.n199 322.329
R667 VDD.n363 VDD.n40 315.406
R668 VDD.n306 VDD.n261 315.406
R669 VDD.n32 VDD.n31 312.053
R670 VDD.n42 VDD.n41 312.053
R671 VDD.n351 VDD.n45 312.053
R672 VDD.n342 VDD.n53 312.053
R673 VDD.n204 VDD.n203 312.053
R674 VDD.n247 VDD.n246 312.053
R675 VDD.n260 VDD.n259 312.053
R676 VDD.n350 VDD.n46 312.051
R677 VDD.n197 VDD.n196 312.051
R678 VDD.n266 VDD.n265 312.051
R679 VDD.n298 VDD.n264 312.005
R680 VDD.n21 VDD.n20 311.582
R681 VDD.n378 VDD.n23 308.755
R682 VDD.n314 VDD.n256 308.755
R683 VDD.n241 VDD.n202 308.755
R684 VDD.n155 VDD.t95 306.735
R685 VDD.n258 VDD.n257 259.697
R686 VDD.n344 VDD.n51 259.697
R687 VDD.n251 VDD.t13 249.363
R688 VDD.n255 VDD.t27 246.805
R689 VDD.n12 VDD.t100 245.667
R690 VDD.n17 VDD.t93 245.667
R691 VDD.n29 VDD.t98 245.667
R692 VDD.n57 VDD.t90 245.667
R693 VDD.n60 VDD.t99 245.667
R694 VDD.n207 VDD.t91 245.667
R695 VDD.n231 VDD.t89 245.667
R696 VDD.n275 VDD.t97 245.667
R697 VDD.n283 VDD.t92 245.667
R698 VDD.n81 VDD.t88 242.282
R699 VDD.n131 VDD.t94 242.282
R700 VDD.n107 VDD.t96 242.282
R701 VDD.n50 VDD.t12 240.215
R702 VDD.n257 VDD.t28 157.014
R703 VDD.n51 VDD.t11 156.998
R704 VDD.n51 VDD.t45 137.095
R705 VDD.n257 VDD.t54 137.079
R706 VDD.n199 VDD.t22 116.341
R707 VDD.n40 VDD.t8 96.1553
R708 VDD.n54 VDD.t48 96.1553
R709 VDD.n254 VDD.t4 96.1553
R710 VDD.n261 VDD.t24 96.1553
R711 VDD.n264 VDD.t10 96.1553
R712 VDD.n19 VDD.t51 77.3934
R713 VDD.n24 VDD.t14 77.3934
R714 VDD.n26 VDD.t41 77.3934
R715 VDD.n103 VDD.t43 77.3934
R716 VDD.n100 VDD.t23 77.3934
R717 VDD.n123 VDD.t52 77.3934
R718 VDD.n54 VDD.t26 63.3219
R719 VDD.n254 VDD.t7 63.3219
R720 VDD.n19 VDD.t87 41.0422
R721 VDD.n24 VDD.t55 41.0422
R722 VDD.n26 VDD.t20 41.0422
R723 VDD.n103 VDD.t17 41.0422
R724 VDD.n100 VDD.t35 41.0422
R725 VDD.n123 VDD.t30 41.0422
R726 VDD.n23 VDD.t85 36.1587
R727 VDD.n23 VDD.t19 36.1587
R728 VDD.n20 VDD.t53 36.1587
R729 VDD.n20 VDD.t34 36.1587
R730 VDD.n31 VDD.t3 36.1587
R731 VDD.n31 VDD.t56 36.1587
R732 VDD.n41 VDD.t1 36.1587
R733 VDD.n41 VDD.t16 36.1587
R734 VDD.n45 VDD.t31 36.1587
R735 VDD.n45 VDD.t46 36.1587
R736 VDD.n46 VDD.t32 36.1587
R737 VDD.n46 VDD.t36 36.1587
R738 VDD.n53 VDD.t47 36.1587
R739 VDD.n53 VDD.t39 36.1587
R740 VDD.n256 VDD.t84 36.1587
R741 VDD.n256 VDD.t33 36.1587
R742 VDD.n202 VDD.t57 36.1587
R743 VDD.n202 VDD.t40 36.1587
R744 VDD.n203 VDD.t2 36.1587
R745 VDD.n203 VDD.t49 36.1587
R746 VDD.n246 VDD.t38 36.1587
R747 VDD.n246 VDD.t5 36.1587
R748 VDD.n196 VDD.t86 36.1587
R749 VDD.n196 VDD.t21 36.1587
R750 VDD.n259 VDD.t44 36.1587
R751 VDD.n259 VDD.t18 36.1587
R752 VDD.n265 VDD.t15 36.1587
R753 VDD.n265 VDD.t42 36.1587
R754 VDD.n379 VDD.n378 34.6358
R755 VDD.n241 VDD.n240 34.6358
R756 VDD.n315 VDD.n314 34.6358
R757 VDD.n380 VDD.n379 34.6358
R758 VDD.n349 VDD.n48 34.6358
R759 VDD.n245 VDD.n244 34.6358
R760 VDD.n311 VDD.n310 34.6358
R761 VDD.n305 VDD.n262 34.6358
R762 VDD.n301 VDD.n262 34.6358
R763 VDD.n301 VDD.n300 34.6358
R764 VDD.n125 VDD.n122 34.6358
R765 VDD.n117 VDD.n116 34.6358
R766 VDD.n118 VDD.n117 34.6358
R767 VDD.n113 VDD.n112 34.6358
R768 VDD.n50 VDD.n48 32.377
R769 VDD.n375 VDD.n25 30.4946
R770 VDD.n199 VDD.t0 28.4453
R771 VDD.n122 VDD.n121 27.1064
R772 VDD.n40 VDD.t50 26.5955
R773 VDD.n261 VDD.t29 26.5955
R774 VDD.n353 VDD.n352 25.977
R775 VDD.n253 VDD.n251 25.977
R776 VDD.n264 VDD.t37 25.6105
R777 VDD.n129 VDD.n98 25.224
R778 VDD.n133 VDD.n129 25.1912
R779 VDD.n112 VDD.n109 25.1912
R780 VDD.n385 VDD.n384 23.7181
R781 VDD.n375 VDD.n374 23.7181
R782 VDD.n374 VDD.n373 23.7181
R783 VDD.n340 VDD.n62 23.7181
R784 VDD.n234 VDD.n233 23.7181
R785 VDD.n285 VDD.n273 23.7181
R786 VDD.n125 VDD.n124 23.019
R787 VDD.n363 VDD.n362 22.9652
R788 VDD.n315 VDD.n255 22.9652
R789 VDD.n306 VDD.n305 22.9652
R790 VDD.n373 VDD.n32 22.2123
R791 VDD.n362 VDD.n42 22.2123
R792 VDD.n353 VDD.n42 22.2123
R793 VDD.n350 VDD.n349 22.2123
R794 VDD.n343 VDD.n342 22.2123
R795 VDD.n234 VDD.n204 22.2123
R796 VDD.n238 VDD.n204 22.2123
R797 VDD.n247 VDD.n245 22.2123
R798 VDD.n310 VDD.n260 22.2123
R799 VDD.n297 VDD.n266 22.2123
R800 VDD.n273 VDD.n266 22.2123
R801 VDD.n384 VDD.n21 21.4593
R802 VDD.n341 VDD.n340 21.4593
R803 VDD.n255 VDD.n253 21.4593
R804 VDD.n299 VDD.n298 21.4593
R805 VDD.n118 VDD.n101 20.3837
R806 VDD.n380 VDD.n21 18.824
R807 VDD.n241 VDD.n200 18.824
R808 VDD.n345 VDD.n344 18.4476
R809 VDD.n311 VDD.n258 18.0711
R810 VDD.n149 VDD.n147 17.612
R811 VDD.n170 VDD.n169 17.3413
R812 VDD.n314 VDD.n258 16.5652
R813 VDD.n344 VDD.n343 16.1887
R814 VDD.n244 VDD.n200 15.8123
R815 VDD.n363 VDD.n32 12.8005
R816 VDD.n306 VDD.n260 12.8005
R817 VDD.n298 VDD.n297 12.0476
R818 VDD.n352 VDD.n351 11.6711
R819 VDD.n251 VDD.n197 11.2946
R820 VDD.n342 VDD.n341 10.5417
R821 VDD.n351 VDD.n350 9.78874
R822 VDD.n247 VDD.n197 9.78874
R823 VDD.n116 VDD.n104 9.73495
R824 VDD.n153 VDD.n89 9.73273
R825 VDD.n154 VDD.n153 9.73273
R826 VDD.n156 VDD.n87 9.73273
R827 VDD.n160 VDD.n87 9.73273
R828 VDD.n161 VDD.n160 9.73273
R829 VDD.n162 VDD.n161 9.73273
R830 VDD.n162 VDD.n85 9.73273
R831 VDD.n166 VDD.n85 9.73273
R832 VDD.n182 VDD.n181 9.60526
R833 VDD.n105 VDD.n0 9.60526
R834 VDD.n240 VDD.n239 9.41227
R835 VDD.n73 VDD.n62 9.3005
R836 VDD.n71 VDD.n62 9.3005
R837 VDD.n64 VDD.n62 9.3005
R838 VDD.n385 VDD.n15 9.3005
R839 VDD.n386 VDD.n385 9.3005
R840 VDD.n385 VDD.n14 9.3005
R841 VDD.n384 VDD.n383 9.3005
R842 VDD.n382 VDD.n21 9.3005
R843 VDD.n381 VDD.n380 9.3005
R844 VDD.n379 VDD.n22 9.3005
R845 VDD.n378 VDD.n377 9.3005
R846 VDD.n376 VDD.n375 9.3005
R847 VDD.n373 VDD.n372 9.3005
R848 VDD.n33 VDD.n32 9.3005
R849 VDD.n364 VDD.n363 9.3005
R850 VDD.n362 VDD.n361 9.3005
R851 VDD.n355 VDD.n42 9.3005
R852 VDD.n354 VDD.n353 9.3005
R853 VDD.n352 VDD.n43 9.3005
R854 VDD.n351 VDD.n44 9.3005
R855 VDD.n350 VDD.n47 9.3005
R856 VDD.n349 VDD.n348 9.3005
R857 VDD.n347 VDD.n48 9.3005
R858 VDD.n346 VDD.n345 9.3005
R859 VDD.n343 VDD.n49 9.3005
R860 VDD.n342 VDD.n52 9.3005
R861 VDD.n341 VDD.n55 9.3005
R862 VDD.n340 VDD.n339 9.3005
R863 VDD.n286 VDD.n285 9.3005
R864 VDD.n285 VDD.n281 9.3005
R865 VDD.n285 VDD.n278 9.3005
R866 VDD.n233 VDD.n229 9.3005
R867 VDD.n233 VDD.n209 9.3005
R868 VDD.n233 VDD.n205 9.3005
R869 VDD.n235 VDD.n234 9.3005
R870 VDD.n236 VDD.n204 9.3005
R871 VDD.n238 VDD.n237 9.3005
R872 VDD.n240 VDD.n201 9.3005
R873 VDD.n242 VDD.n241 9.3005
R874 VDD.n244 VDD.n243 9.3005
R875 VDD.n245 VDD.n198 9.3005
R876 VDD.n248 VDD.n247 9.3005
R877 VDD.n249 VDD.n197 9.3005
R878 VDD.n251 VDD.n250 9.3005
R879 VDD.n253 VDD.n252 9.3005
R880 VDD.n255 VDD.n193 9.3005
R881 VDD.n316 VDD.n315 9.3005
R882 VDD.n314 VDD.n313 9.3005
R883 VDD.n312 VDD.n311 9.3005
R884 VDD.n310 VDD.n309 9.3005
R885 VDD.n308 VDD.n260 9.3005
R886 VDD.n307 VDD.n306 9.3005
R887 VDD.n305 VDD.n304 9.3005
R888 VDD.n303 VDD.n262 9.3005
R889 VDD.n302 VDD.n301 9.3005
R890 VDD.n300 VDD.n263 9.3005
R891 VDD.n297 VDD.n296 9.3005
R892 VDD.n295 VDD.n266 9.3005
R893 VDD.n273 VDD.n267 9.3005
R894 VDD.n106 VDD.n1 9.3005
R895 VDD.n110 VDD.n109 9.3005
R896 VDD.n112 VDD.n111 9.3005
R897 VDD.n114 VDD.n113 9.3005
R898 VDD.n116 VDD.n115 9.3005
R899 VDD.n117 VDD.n102 9.3005
R900 VDD.n119 VDD.n118 9.3005
R901 VDD.n121 VDD.n120 9.3005
R902 VDD.n122 VDD.n99 9.3005
R903 VDD.n126 VDD.n125 9.3005
R904 VDD.n127 VDD.n98 9.3005
R905 VDD.n129 VDD.n128 9.3005
R906 VDD.n134 VDD.n133 9.3005
R907 VDD.n130 VDD.n92 9.3005
R908 VDD.n147 VDD.n146 9.3005
R909 VDD.n150 VDD.n149 9.3005
R910 VDD.n151 VDD.n89 9.3005
R911 VDD.n153 VDD.n152 9.3005
R912 VDD.n154 VDD.n88 9.3005
R913 VDD.n157 VDD.n156 9.3005
R914 VDD.n158 VDD.n87 9.3005
R915 VDD.n160 VDD.n159 9.3005
R916 VDD.n161 VDD.n86 9.3005
R917 VDD.n163 VDD.n162 9.3005
R918 VDD.n164 VDD.n85 9.3005
R919 VDD.n166 VDD.n165 9.3005
R920 VDD.n171 VDD.n170 9.3005
R921 VDD.n169 VDD.n82 9.3005
R922 VDD.n180 VDD.n179 9.3005
R923 VDD.n148 VDD.n89 9.09802
R924 VDD.n167 VDD.n166 9.09802
R925 VDD.n155 VDD.n154 5.18397
R926 VDD.n156 VDD.n155 4.54926
R927 VDD.n404 VDD.n3 4.51401
R928 VDD.n325 VDD.n191 4.51401
R929 VDD.n195 VDD.n194 4.51401
R930 VDD.n371 VDD.n370 4.51401
R931 VDD.n360 VDD.n359 4.51401
R932 VDD.n65 VDD.n63 4.51401
R933 VDD.n75 VDD.n74 4.51401
R934 VDD.n10 VDD.n9 4.51401
R935 VDD.n226 VDD.n212 4.51401
R936 VDD.n294 VDD.n293 4.51401
R937 VDD.n288 VDD.n287 4.51401
R938 VDD.n84 VDD.n83 4.51401
R939 VDD.n184 VDD.n183 4.51401
R940 VDD.n139 VDD.n96 4.51401
R941 VDD.n143 VDD.n90 4.51401
R942 VDD.n338 VDD.n337 4.5005
R943 VDD.n70 VDD.n66 4.5005
R944 VDD.n72 VDD.n69 4.5005
R945 VDD.n38 VDD.n34 4.5005
R946 VDD.n366 VDD.n365 4.5005
R947 VDD.n356 VDD.n39 4.5005
R948 VDD.n391 VDD.n8 4.5005
R949 VDD.n388 VDD.n387 4.5005
R950 VDD.n216 VDD.n210 4.5005
R951 VDD.n228 VDD.n227 4.5005
R952 VDD.n324 VDD.n323 4.5005
R953 VDD.n322 VDD.n321 4.5005
R954 VDD.n318 VDD.n317 4.5005
R955 VDD.n277 VDD.n268 4.5005
R956 VDD.n280 VDD.n279 4.5005
R957 VDD.n272 VDD.n271 4.5005
R958 VDD.n398 VDD.n397 4.5005
R959 VDD.n406 VDD.n405 4.5005
R960 VDD.n173 VDD.n172 4.5005
R961 VDD.n178 VDD.n177 4.5005
R962 VDD.n80 VDD.n79 4.5005
R963 VDD.n138 VDD.n137 4.5005
R964 VDD.n136 VDD.n135 4.5005
R965 VDD.n145 VDD.n144 4.5005
R966 VDD.n181 VDD.n180 4.36875
R967 VDD.n130 VDD.n91 4.36875
R968 VDD.n106 VDD.n105 4.36875
R969 VDD.n113 VDD.n104 4.19546
R970 VDD.n378 VDD.n25 4.14168
R971 VDD.n239 VDD.n238 4.14168
R972 VDD.n385 VDD.n13 4.02033
R973 VDD.n385 VDD.n18 4.02033
R974 VDD.n374 VDD.n30 4.02033
R975 VDD.n62 VDD.n58 4.02033
R976 VDD.n62 VDD.n61 4.02033
R977 VDD.n233 VDD.n208 4.02033
R978 VDD.n233 VDD.n232 4.02033
R979 VDD.n285 VDD.n276 4.02033
R980 VDD.n285 VDD.n284 4.02033
R981 VDD.n180 VDD.n81 3.50526
R982 VDD.n131 VDD.n130 3.50526
R983 VDD.n107 VDD.n106 3.50526
R984 VDD.n394 VDD.n393 3.48706
R985 VDD.n401 VDD.n400 3.48706
R986 VDD.n219 VDD.n218 3.45831
R987 VDD.n404 VDD.n403 3.43925
R988 VDD.n143 VDD.n142 3.43925
R989 VDD.n194 VDD.n188 3.43925
R990 VDD.n326 VDD.n325 3.43925
R991 VDD.n140 VDD.n139 3.43925
R992 VDD.n333 VDD.n75 3.43925
R993 VDD.n67 VDD.n65 3.43925
R994 VDD.n9 VDD.n5 3.43925
R995 VDD.n289 VDD.n288 3.43925
R996 VDD.n293 VDD.n292 3.43925
R997 VDD.n399 VDD.n396 3.4105
R998 VDD.n4 VDD.n2 3.4105
R999 VDD.n192 VDD.n190 3.4105
R1000 VDD.n320 VDD.n319 3.4105
R1001 VDD.n358 VDD.n35 3.4105
R1002 VDD.n369 VDD.n35 3.4105
R1003 VDD.n359 VDD.n358 3.4105
R1004 VDD.n370 VDD.n369 3.4105
R1005 VDD.n368 VDD.n367 3.4105
R1006 VDD.n357 VDD.n37 3.4105
R1007 VDD.n336 VDD.n335 3.4105
R1008 VDD.n334 VDD.n68 3.4105
R1009 VDD.n392 VDD.n7 3.4105
R1010 VDD.n390 VDD.n389 3.4105
R1011 VDD.n225 VDD.n224 3.4105
R1012 VDD.n224 VDD.n219 3.4105
R1013 VDD.n226 VDD.n225 3.4105
R1014 VDD.n217 VDD.n215 3.4105
R1015 VDD.n213 VDD.n211 3.4105
R1016 VDD.n291 VDD.n269 3.4105
R1017 VDD.n290 VDD.n270 3.4105
R1018 VDD.n186 VDD.n185 3.4105
R1019 VDD.n186 VDD.n77 3.4105
R1020 VDD.n185 VDD.n184 3.4105
R1021 VDD.n83 VDD.n77 3.4105
R1022 VDD.n175 VDD.n174 3.4105
R1023 VDD.n176 VDD.n78 3.4105
R1024 VDD.n97 VDD.n95 3.4105
R1025 VDD.n94 VDD.n93 3.4105
R1026 VDD.n374 VDD.n27 3.04861
R1027 VDD.n13 VDD.n11 2.63539
R1028 VDD.n18 VDD.n16 2.63539
R1029 VDD.n30 VDD.n28 2.63539
R1030 VDD.n58 VDD.n56 2.63539
R1031 VDD.n61 VDD.n59 2.63539
R1032 VDD.n208 VDD.n206 2.63539
R1033 VDD.n232 VDD.n230 2.63539
R1034 VDD.n276 VDD.n274 2.63539
R1035 VDD.n284 VDD.n282 2.63539
R1036 VDD.n17 VDD.n16 2.37495
R1037 VDD.n12 VDD.n11 2.37495
R1038 VDD.n29 VDD.n28 2.37495
R1039 VDD.n60 VDD.n59 2.37495
R1040 VDD.n57 VDD.n56 2.37495
R1041 VDD.n231 VDD.n230 2.37495
R1042 VDD.n207 VDD.n206 2.37495
R1043 VDD.n283 VDD.n282 2.37495
R1044 VDD.n275 VDD.n274 2.37495
R1045 VDD.n393 VDD.n8 2.33488
R1046 VDD.n218 VDD.n210 2.33488
R1047 VDD.n400 VDD.n397 2.33488
R1048 VDD.n345 VDD.n50 2.25932
R1049 VDD.n327 VDD.n188 1.69188
R1050 VDD.n327 VDD.n326 1.69188
R1051 VDD.n142 VDD.n141 1.69188
R1052 VDD.n141 VDD.n140 1.69188
R1053 VDD.n36 VDD.n35 1.69188
R1054 VDD.n395 VDD.n5 1.69188
R1055 VDD.n395 VDD.n394 1.69188
R1056 VDD.n403 VDD.n402 1.69188
R1057 VDD.n402 VDD.n401 1.69188
R1058 VDD.n224 VDD.n214 1.69188
R1059 VDD.n292 VDD.n187 1.69188
R1060 VDD.n289 VDD.n187 1.69188
R1061 VDD.n332 VDD.n67 1.69188
R1062 VDD.n333 VDD.n332 1.69188
R1063 VDD.n186 VDD.n76 1.69188
R1064 VDD.n300 VDD.n299 1.12991
R1065 VDD.n121 VDD.n101 1.07613
R1066 VDD.n168 VDD.n81 0.863992
R1067 VDD.n132 VDD.n131 0.863992
R1068 VDD.n108 VDD.n107 0.863992
R1069 VDD.n149 VDD.n148 0.635211
R1070 VDD.n170 VDD.n167 0.635211
R1071 VDD.n329 VDD.n6 0.500125
R1072 VDD.n223 VDD.n222 0.500125
R1073 VDD.n222 VDD.n189 0.3805
R1074 VDD.n329 VDD.n328 0.3805
R1075 VDD.n221 VDD.n220 0.3805
R1076 VDD.n331 VDD.n330 0.3805
R1077 VDD.n124 VDD.n98 0.323189
R1078 VDD.n169 VDD.n168 0.305262
R1079 VDD.n133 VDD.n132 0.305262
R1080 VDD.n147 VDD.n91 0.305262
R1081 VDD.n109 VDD.n108 0.305262
R1082 VDD.n27 VDD 0.217246
R1083 VDD.n141 VDD.n35 0.1603
R1084 VDD.n402 VDD.n395 0.1603
R1085 VDD.n332 VDD.n186 0.1603
R1086 VDD.n328 VDD.n327 0.14385
R1087 VDD.n224 VDD.n6 0.14385
R1088 VDD.n331 VDD.n187 0.14385
R1089 VDD VDD.n27 0.14207
R1090 VDD.n383 VDD.n14 0.120292
R1091 VDD.n382 VDD.n381 0.120292
R1092 VDD.n381 VDD.n22 0.120292
R1093 VDD.n377 VDD.n22 0.120292
R1094 VDD.n377 VDD.n376 0.120292
R1095 VDD.n355 VDD.n354 0.120292
R1096 VDD.n354 VDD.n43 0.120292
R1097 VDD.n348 VDD.n47 0.120292
R1098 VDD.n347 VDD.n346 0.120292
R1099 VDD.n346 VDD.n49 0.120292
R1100 VDD.n52 VDD.n49 0.120292
R1101 VDD.n55 VDD.n52 0.120292
R1102 VDD.n235 VDD.n205 0.120292
R1103 VDD.n236 VDD.n235 0.120292
R1104 VDD.n242 VDD.n201 0.120292
R1105 VDD.n243 VDD.n242 0.120292
R1106 VDD.n248 VDD.n198 0.120292
R1107 VDD.n313 VDD.n312 0.120292
R1108 VDD.n309 VDD.n308 0.120292
R1109 VDD.n308 VDD.n307 0.120292
R1110 VDD.n304 VDD.n303 0.120292
R1111 VDD.n302 VDD.n263 0.120292
R1112 VDD.n296 VDD.n295 0.120292
R1113 VDD.n111 VDD.n110 0.120292
R1114 VDD.n115 VDD.n114 0.120292
R1115 VDD.n115 VDD.n102 0.120292
R1116 VDD.n119 VDD.n102 0.120292
R1117 VDD.n120 VDD.n119 0.120292
R1118 VDD.n120 VDD.n99 0.120292
R1119 VDD.n126 VDD.n99 0.120292
R1120 VDD.n127 VDD.n126 0.120292
R1121 VDD.n128 VDD.n127 0.120292
R1122 VDD.n151 VDD.n150 0.120292
R1123 VDD.n152 VDD.n151 0.120292
R1124 VDD.n152 VDD.n88 0.120292
R1125 VDD.n157 VDD.n88 0.120292
R1126 VDD.n158 VDD.n157 0.120292
R1127 VDD.n159 VDD.n158 0.120292
R1128 VDD.n159 VDD.n86 0.120292
R1129 VDD.n163 VDD.n86 0.120292
R1130 VDD.n164 VDD.n163 0.120292
R1131 VDD.n165 VDD.n164 0.120292
R1132 VDD.n330 VDD.n329 0.120125
R1133 VDD.n222 VDD.n221 0.120125
R1134 VDD.n14 VDD.n10 0.117688
R1135 VDD.n212 VDD.n205 0.117688
R1136 VDD.n110 VDD.n3 0.117688
R1137 VDD.n295 VDD.n294 0.112479
R1138 VDD.n165 VDD.n84 0.112479
R1139 VDD.n114 VDD 0.104667
R1140 VDD.n296 VDD 0.0994583
R1141 VDD VDD.n382 0.0981562
R1142 VDD.n372 VDD 0.0981562
R1143 VDD.n44 VDD 0.0981562
R1144 VDD.n47 VDD 0.0981562
R1145 VDD VDD.n201 0.0981562
R1146 VDD VDD.n198 0.0981562
R1147 VDD.n249 VDD 0.0981562
R1148 VDD.n250 VDD 0.0981562
R1149 VDD.n309 VDD 0.0981562
R1150 VDD.n304 VDD 0.0981562
R1151 VDD VDD.n347 0.0968542
R1152 VDD.n405 VDD.n404 0.0950946
R1153 VDD.n325 VDD.n324 0.0950946
R1154 VDD.n318 VDD.n194 0.0950946
R1155 VDD.n370 VDD.n34 0.0950946
R1156 VDD.n359 VDD.n356 0.0950946
R1157 VDD.n337 VDD.n65 0.0950946
R1158 VDD.n75 VDD.n69 0.0950946
R1159 VDD.n388 VDD.n9 0.0950946
R1160 VDD.n227 VDD.n226 0.0950946
R1161 VDD.n293 VDD.n268 0.0950946
R1162 VDD.n288 VDD.n271 0.0950946
R1163 VDD.n173 VDD.n83 0.0950946
R1164 VDD.n184 VDD.n79 0.0950946
R1165 VDD.n139 VDD.n138 0.0950946
R1166 VDD.n144 VDD.n143 0.0950946
R1167 VDD.n63 VDD 0.0903438
R1168 VDD.n400 VDD.n399 0.0878527
R1169 VDD.n393 VDD.n392 0.0878527
R1170 VDD.n218 VDD.n217 0.0878527
R1171 VDD.n237 VDD 0.0877396
R1172 VDD VDD.n302 0.0877396
R1173 VDD.n365 VDD.n38 0.0838333
R1174 VDD.n74 VDD.n72 0.0838333
R1175 VDD.n323 VDD.n322 0.0838333
R1176 VDD.n287 VDD.n272 0.0838333
R1177 VDD.n137 VDD.n136 0.0838333
R1178 VDD.n183 VDD.n80 0.0838333
R1179 VDD.n387 VDD.n386 0.0812292
R1180 VDD.n364 VDD.n39 0.0812292
R1181 VDD.n71 VDD.n70 0.0812292
R1182 VDD.n228 VDD.n209 0.0812292
R1183 VDD.n281 VDD.n280 0.0812292
R1184 VDD.n406 VDD.n1 0.0812292
R1185 VDD.n145 VDD.n92 0.0812292
R1186 VDD.n179 VDD.n178 0.0812292
R1187 VDD.n360 VDD.n355 0.0760208
R1188 VDD.n313 VDD.n195 0.0760208
R1189 VDD.n150 VDD.n90 0.0760208
R1190 VDD.n250 VDD.n191 0.0708125
R1191 VDD.n128 VDD.n96 0.0708125
R1192 VDD.n399 VDD.n398 0.0680676
R1193 VDD.n398 VDD.n2 0.0680676
R1194 VDD.n321 VDD.n192 0.0680676
R1195 VDD.n321 VDD.n320 0.0680676
R1196 VDD.n367 VDD.n366 0.0680676
R1197 VDD.n366 VDD.n37 0.0680676
R1198 VDD.n336 VDD.n66 0.0680676
R1199 VDD.n68 VDD.n66 0.0680676
R1200 VDD.n392 VDD.n391 0.0680676
R1201 VDD.n391 VDD.n390 0.0680676
R1202 VDD.n217 VDD.n216 0.0680676
R1203 VDD.n216 VDD.n211 0.0680676
R1204 VDD.n279 VDD.n269 0.0680676
R1205 VDD.n279 VDD.n270 0.0680676
R1206 VDD.n177 VDD.n175 0.0680676
R1207 VDD.n177 VDD.n176 0.0680676
R1208 VDD.n135 VDD.n97 0.0680676
R1209 VDD.n317 VDD 0.0577917
R1210 VDD.n396 VDD.n4 0.0574697
R1211 VDD.n95 VDD.n94 0.0574697
R1212 VDD.n319 VDD.n190 0.0574697
R1213 VDD.n369 VDD.n368 0.0574697
R1214 VDD.n358 VDD.n357 0.0574697
R1215 VDD.n335 VDD.n334 0.0574697
R1216 VDD.n389 VDD.n7 0.0574697
R1217 VDD.n219 VDD.n215 0.0574697
R1218 VDD.n225 VDD.n213 0.0574697
R1219 VDD.n291 VDD.n290 0.0574697
R1220 VDD.n174 VDD.n77 0.0574697
R1221 VDD.n185 VDD.n78 0.0574697
R1222 VDD.n277 VDD 0.0538854
R1223 VDD.n172 VDD 0.0538854
R1224 VDD.n327 VDD.n189 0.051025
R1225 VDD.n224 VDD.n223 0.051025
R1226 VDD.n220 VDD.n187 0.051025
R1227 VDD.n371 VDD.n33 0.0499792
R1228 VDD.n252 VDD.n191 0.0499792
R1229 VDD.n134 VDD.n96 0.0499792
R1230 VDD.n15 VDD.n8 0.0447708
R1231 VDD VDD.n338 0.0447708
R1232 VDD.n338 VDD.n64 0.0447708
R1233 VDD.n229 VDD.n210 0.0447708
R1234 VDD.n316 VDD.n195 0.0447708
R1235 VDD.n278 VDD.n277 0.0447708
R1236 VDD.n397 VDD.n0 0.0447708
R1237 VDD.n172 VDD.n82 0.0447708
R1238 VDD VDD.n371 0.0421667
R1239 VDD.n405 VDD.n2 0.0410405
R1240 VDD.n324 VDD.n192 0.0410405
R1241 VDD.n320 VDD.n318 0.0410405
R1242 VDD.n367 VDD.n34 0.0410405
R1243 VDD.n356 VDD.n37 0.0410405
R1244 VDD.n337 VDD.n336 0.0410405
R1245 VDD.n69 VDD.n68 0.0410405
R1246 VDD.n390 VDD.n388 0.0410405
R1247 VDD.n227 VDD.n211 0.0410405
R1248 VDD.n269 VDD.n268 0.0410405
R1249 VDD.n271 VDD.n270 0.0410405
R1250 VDD.n175 VDD.n173 0.0410405
R1251 VDD.n176 VDD.n79 0.0410405
R1252 VDD.n138 VDD.n97 0.0410405
R1253 VDD.n144 VDD.n93 0.0410405
R1254 VDD.n361 VDD.n39 0.0395625
R1255 VDD.n70 VDD.n64 0.0395625
R1256 VDD.n317 VDD.n316 0.0395625
R1257 VDD.n280 VDD.n278 0.0395625
R1258 VDD.n146 VDD.n145 0.0395625
R1259 VDD.n178 VDD.n82 0.0395625
R1260 VDD.n189 VDD 0.036925
R1261 VDD.n223 VDD 0.036925
R1262 VDD.n220 VDD 0.036925
R1263 VDD.n38 VDD.n33 0.0343542
R1264 VDD.n74 VDD.n73 0.0343542
R1265 VDD.n287 VDD.n286 0.0343542
R1266 VDD.n137 VDD.n134 0.0343542
R1267 VDD.n183 VDD.n182 0.0343542
R1268 VDD.n135 VDD 0.0342838
R1269 VDD VDD.n93 0.0342838
R1270 VDD VDD.n236 0.0330521
R1271 VDD.n303 VDD 0.0330521
R1272 VDD.n140 VDD.n95 0.0292489
R1273 VDD.n326 VDD.n190 0.0292489
R1274 VDD.n319 VDD.n188 0.0292489
R1275 VDD.n142 VDD.n94 0.0292489
R1276 VDD.n357 VDD.n36 0.0292489
R1277 VDD.n368 VDD.n36 0.0292489
R1278 VDD.n335 VDD.n67 0.0292489
R1279 VDD.n334 VDD.n333 0.0292489
R1280 VDD.n394 VDD.n7 0.0292489
R1281 VDD.n389 VDD.n5 0.0292489
R1282 VDD.n401 VDD.n396 0.0292489
R1283 VDD.n403 VDD.n4 0.0292489
R1284 VDD.n214 VDD.n213 0.0292489
R1285 VDD.n215 VDD.n214 0.0292489
R1286 VDD.n292 VDD.n291 0.0292489
R1287 VDD.n290 VDD.n289 0.0292489
R1288 VDD.n78 VDD.n76 0.0292489
R1289 VDD.n174 VDD.n76 0.0292489
R1290 VDD.n348 VDD 0.0239375
R1291 VDD VDD.n193 0.0239375
R1292 VDD.n330 VDD 0.022975
R1293 VDD.n221 VDD 0.022975
R1294 VDD.n15 VDD 0.0226354
R1295 VDD.n383 VDD 0.0226354
R1296 VDD.n376 VDD 0.0226354
R1297 VDD.n372 VDD 0.0226354
R1298 VDD.n361 VDD 0.0226354
R1299 VDD VDD.n360 0.0226354
R1300 VDD VDD.n44 0.0226354
R1301 VDD VDD.n55 0.0226354
R1302 VDD.n339 VDD 0.0226354
R1303 VDD.n73 VDD 0.0226354
R1304 VDD.n229 VDD 0.0226354
R1305 VDD.n237 VDD 0.0226354
R1306 VDD.n243 VDD 0.0226354
R1307 VDD VDD.n248 0.0226354
R1308 VDD VDD.n249 0.0226354
R1309 VDD.n252 VDD 0.0226354
R1310 VDD.n312 VDD 0.0226354
R1311 VDD.n307 VDD 0.0226354
R1312 VDD VDD.n267 0.0226354
R1313 VDD.n286 VDD 0.0226354
R1314 VDD VDD.n0 0.0226354
R1315 VDD.n146 VDD 0.0226354
R1316 VDD VDD.n90 0.0226354
R1317 VDD VDD.n171 0.0226354
R1318 VDD.n182 VDD 0.0226354
R1319 VDD VDD.n43 0.0213333
R1320 VDD VDD.n263 0.0213333
R1321 VDD.n387 VDD 0.0174271
R1322 VDD VDD.n228 0.0174271
R1323 VDD VDD.n406 0.0174271
R1324 VDD.n328 VDD.n35 0.01695
R1325 VDD.n395 VDD.n6 0.01695
R1326 VDD.n332 VDD.n331 0.01695
R1327 VDD.n111 VDD 0.016125
R1328 VDD.n323 VDD 0.0122188
R1329 VDD.n339 VDD.n63 0.0083125
R1330 VDD.n294 VDD.n267 0.0083125
R1331 VDD.n171 VDD.n84 0.0083125
R1332 VDD.n386 VDD.n10 0.00310417
R1333 VDD.n365 VDD.n364 0.00310417
R1334 VDD.n72 VDD.n71 0.00310417
R1335 VDD.n212 VDD.n209 0.00310417
R1336 VDD.n322 VDD.n193 0.00310417
R1337 VDD.n281 VDD.n272 0.00310417
R1338 VDD.n3 VDD.n1 0.00310417
R1339 VDD.n136 VDD.n92 0.00310417
R1340 VDD.n179 VDD.n80 0.00310417
R1341 gpo0.n0 gpo0.t1 368.521
R1342 gpo0.n2 gpo0.t0 216.155
R1343 gpo0 gpo0.n2 78.8791
R1344 gpo0.n1 gpo0 27.368
R1345 gpo0.n1 gpo0.n0 6.52665
R1346 gpo0.n0 gpo0 5.48477
R1347 gpo0.n2 gpo0 5.16973
R1348 gpo0 gpo0.n1 4.03013
R1349 gpo3.n0 gpo3.t1 368.521
R1350 gpo3.n1 gpo3.t0 216.155
R1351 gpo3.n1 gpo3 78.8791
R1352 gpo3 gpo3.n2 19.5448
R1353 gpo3 gpo3.n0 10.5563
R1354 gpo3.n0 gpo3 5.48477
R1355 gpo3.n2 gpo3 4.18512
R1356 gpo3.n2 gpo3.n1 0.985115
R1357 gno1 gno1.t1 744.352
R1358 gno1.t1 gno1.n0 732.75
R1359 gno1 gno1.t0 219.355
R1360 gno1.n0 gno1 80.894
R1361 gno1 gno1.n1 18.0805
R1362 gno1.n1 gno1 12.0894
R1363 gno1.n1 gno1 4.03013
R1364 gno1.n0 gno1 2.84494
R1365 gno2.n0 gno2.t1 368.521
R1366 gno2.n1 gno2.t0 216.155
R1367 gno2 gno2.n1 78.8791
R1368 gno2 gno2.n2 17.9912
R1369 gno2.n2 gno2.n0 6.52665
R1370 gno2.n0 gno2 5.48477
R1371 gno2.n1 gno2 5.16973
R1372 gno2.n2 gno2 4.03013
R1373 gno3.n0 gno3.t1 368.521
R1374 gno3.n1 gno3.t0 216.155
R1375 gno3 gno3.n1 78.8791
R1376 gno3 gno3.n2 19.2233
R1377 gno3.n2 gno3.n0 6.52665
R1378 gno3.n0 gno3 5.48477
R1379 gno3.n1 gno3 5.16973
R1380 gno3.n2 gno3 4.03013
R1381 select1.n0 select1.t1 323.55
R1382 select1.n0 select1.t0 195.017
R1383 select1.n1 select1.n0 152
R1384 select1 select1.n1 7.52215
R1385 select1.n1 select1 1.45205
R1386 gno0.n2 gno0.t1 748.383
R1387 gno0.n1 gno0.t1 732.75
R1388 gno0.n0 gno0.t0 216.155
R1389 gno0 gno0.n0 78.8791
R1390 gno0 gno0.n2 29.2251
R1391 gno0 gno0.n1 10.9042
R1392 gno0.n1 gno0 5.21532
R1393 gno0.n0 gno0 5.16973
R1394 gno0.n2 gno0 4.03013
R1395 gpo2.n0 gpo2.t1 368.521
R1396 gpo2.n1 gpo2.t0 216.155
R1397 gpo2.n1 gpo2 78.8791
R1398 gpo2.n2 gpo2 22.4394
R1399 gpo2 gpo2.n0 10.5563
R1400 gpo2.n0 gpo2 5.48477
R1401 gpo2 gpo2.n2 4.18512
R1402 gpo2.n2 gpo2.n1 0.985115
R1403 gpo1.n0 gpo1.t1 368.521
R1404 gpo1.n1 gpo1.t0 216.155
R1405 gpo1.n1 gpo1 78.8791
R1406 gpo1 gpo1.n2 19.84
R1407 gpo1 gpo1.n0 10.5563
R1408 gpo1.n0 gpo1 5.48477
R1409 gpo1.n2 gpo1 4.18512
R1410 gpo1.n2 gpo1.n1 0.985115
C0 a_2835_2986# _01_ 0.205122f
C1 VSS a_1957_2883# 0.00141f
C2 a_1875_2883# a_2051_2223# 2.09e-19
C3 net2 VDD 1.8528f
C4 gpo0 gpo2 3.01e-20
C5 a_2509_3971# _05_ 1.6e-20
C6 gno0 a_2653_3476# 0.10943f
C7 VDD a_2822_3855# 0.134668f
C8 FILLER_0_4_3.VPB select1 0.126422f
C9 select0 a_1677_4221# 1.46e-19
C10 _09_.VPB gpo1 0.009846f
C11 VSS gpo3 0.366122f
C12 VSS gno2 0.209898f
C13 gpo0 net5 3.07e-20
C14 a_2835_2986# _04_ 9.57e-21
C15 _01_ a_3123_2999# 0.018831f
C16 select0 a_2934_4373# 0.010864f
C17 a_3155_2223# net10 0.075584f
C18 FILLER_0_4_3.VPB a_3440_4551# 0.050085f
C19 gpo3 _03_ 1.15e-21
C20 gno2 _03_ 0.092606f
C21 a_1875_2883# a_1407_2767# 0.001479f
C22 _00_ net1 0.31755f
C23 a_3121_4551# _09_.VPB 2.08e-21
C24 a_1448_2473# gno1 0.019861f
C25 a_2287_2741# gpo1 0.0123f
C26 VDD a_1448_2473# 0.117521f
C27 VSS net6 0.145452f
C28 a_1875_2883# gpo1 0.00954f
C29 a_2835_2986# a_2879_2223# 3.69e-20
C30 a_2463_3073# a_2427_3971# 4.61e-20
C31 net6 _03_ 0.014088f
C32 _01_ a_2327_2223# 3.88e-21
C33 a_3318_3855# a_3440_4551# 0.004336f
C34 a_2463_3073# net3 4.68e-20
C35 FILLER_0_4_3.VPB gpo1 6.96e-20
C36 _01_ net10 1.4e-20
C37 net7 net3 0.164881f
C38 VSS a_1499_3311# 0.128946f
C39 a_3431_2223# _09_.VPB 0.065768f
C40 VSS a_2377_3476# 0.105766f
C41 a_3121_4551# FILLER_0_4_3.VPB 0.044717f
C42 _09_.VPB gno1 0.031392f
C43 VDD _05_ 0.092744f
C44 _12_.VPB _04_ 9.81e-20
C45 gno3 a_2879_2223# 5.95e-19
C46 VDD a_2838_4551# 0.150291f
C47 VDD _09_.VPB 0.793352f
C48 a_3601_3855# a_3424_3855# 0.134298f
C49 VDD a_2007_4074# 0.204643f
C50 a_2934_4373# a_2787_4399# 0.003683f
C51 gno0 gpo1 0.022239f
C52 gpo3 gno2 1.12e-20
C53 net4 a_1407_2767# 0.230389f
C54 select0 a_3424_3855# 2.23e-19
C55 net2 VSS 1.49865f
C56 net7 net5 1.52e-19
C57 a_3155_3311# gpo1 1.48e-19
C58 select0 a_2835_2986# 0.001113f
C59 net2 _03_ 0.207324f
C60 VSS a_2822_3855# 0.160404f
C61 a_2287_2741# VDD 0.122209f
C62 _12_.VPB a_1407_3855# 0.083293f
C63 a_2327_2223# a_2879_2223# 8.26e-20
C64 net4 gpo1 0.024817f
C65 net3 a_3481_3476# 2e-19
C66 a_2879_2223# net10 0.084114f
C67 gpo3 net6 0.004299f
C68 VDD a_1875_2883# 0.064911f
C69 net6 gno2 0.003297f
C70 net1 a_3297_3105# 0.001645f
C71 gpo2 a_3424_3855# 0.001135f
C72 VDD FILLER_0_4_3.VPB 0.449342f
C73 gpo0 a_1530_2473# 2.71e-19
C74 a_2415_3133# net8 0.001464f
C75 a_2835_2986# gpo2 2.9e-19
C76 gpo2 a_3481_3476# 0.125542f
C77 _02_ net8 1.73e-20
C78 VSS a_1448_2473# 0.122486f
C79 _01_ a_2051_2223# 3.52e-19
C80 a_3431_2223# a_3318_3855# 2.45e-20
C81 a_3601_3855# net9 5.39e-19
C82 net2 a_1957_2883# 0.001973f
C83 a_3601_3855# _12_.VPB 0.008512f
C84 gno0 gno1 4.86e-20
C85 a_3123_2999# gpo2 0.011389f
C86 gno3 gpo2 0.175495f
C87 VDD gno0 1.09581f
C88 select0 _12_.VPB 0.119544f
C89 a_2101_3476# net1 0.001251f
C90 net1 net8 0.337544f
C91 VDD a_3318_3855# 0.090605f
C92 select0 net10 1.32e-21
C93 VDD a_3155_3311# 0.200073f
C94 _04_ a_2051_2223# 0.197541f
C95 net1 a_1587_3855# 0.197032f
C96 net2 gno2 0.131109f
C97 _12_.VPB a_2427_3971# 0.050824f
C98 net9 net3 5.04e-19
C99 gno3 net5 2.59e-20
C100 VSS _05_ 0.115038f
C101 _12_.VPB net3 0.09613f
C102 _01_ a_1407_2767# 3.94e-19
C103 _00_ net8 2.1e-19
C104 net4 gno1 0.038639f
C105 a_1683_3127# _02_ 0.001836f
C106 a_2822_3855# gno2 8.65e-20
C107 net3 net10 6.79e-21
C108 VSS a_2838_4551# 0.141222f
C109 VSS _09_.VPB 0.468673f
C110 VSS a_2007_4074# 0.123104f
C111 _00_ a_1587_3855# 1.69e-21
C112 VDD net4 0.603334f
C113 net9 gpo2 0.285364f
C114 _12_.VPB gpo2 0.010735f
C115 net1 a_3141_3855# 0.326148f
C116 _09_.VPB _03_ 0.080888f
C117 gpo2 net10 0.019855f
C118 _04_ a_1407_2767# 4.31e-19
C119 net2 net6 0.003038f
C120 _01_ gpo1 0.0373f
C121 gpo0 _02_ 0.11618f
C122 a_1683_3127# net1 0.178111f
C123 a_2287_2741# VSS 0.106771f
C124 a_2327_2223# net5 0.30312f
C125 _12_.VPB net5 1.7e-19
C126 _00_ a_3141_3855# 0.021686f
C127 net10 net5 0.005473f
C128 a_2287_2741# _03_ 8.26e-19
C129 select0 a_2235_4215# 0.002455f
C130 a_3431_2223# a_3155_2223# 5.3e-19
C131 gno2 a_1448_2473# 1.94e-21
C132 select0 a_2653_3476# 1.73e-20
C133 VSS a_1875_2883# 0.163756f
C134 _04_ gpo1 0.163792f
C135 gpo0 net1 0.049099f
C136 VSS FILLER_0_4_3.VPB 0.624348f
C137 net2 a_1499_3311# 6.78e-20
C138 net2 a_2377_3476# 0.013442f
C139 a_2235_4215# a_2427_3971# 0.101254f
C140 VDD a_3155_2223# 0.131112f
C141 a_2427_3971# a_2653_3476# 0.009254f
C142 a_2653_3476# net3 0.234265f
C143 gpo0 _00_ 4.55e-20
C144 net6 a_1448_2473# 5.53e-20
C145 a_3601_3855# select1 1.69e-19
C146 gpo2 a_2653_3476# 1.04e-20
C147 select0 select1 0.042686f
C148 VSS gno0 0.069452f
C149 gpo3 _09_.VPB 0.01539f
C150 net2 a_2822_3855# 0.069048f
C151 VSS a_3318_3855# 0.1224f
C152 gno2 _09_.VPB 0.020967f
C153 _01_ gno1 1.59e-19
C154 a_2235_4215# net5 4.27e-21
C155 VSS a_3155_3311# 0.180026f
C156 net3 a_2051_2223# 2.78e-21
C157 select0 a_3440_4551# 0.002452f
C158 VDD _01_ 0.139005f
C159 a_1499_3311# a_1448_2473# 1.02e-19
C160 a_2934_4373# net1 2.37e-19
C161 a_3297_3105# net8 3.3e-19
C162 a_1875_2883# a_1957_2883# 0.005162f
C163 net7 _02_ 0.004001f
C164 VSS net4 0.277144f
C165 _04_ gno1 0.00104f
C166 gpo2 select1 4.04e-19
C167 net6 _09_.VPB 0.072968f
C168 a_2934_4373# _00_ 1.42e-20
C169 VDD _04_ 0.158452f
C170 a_2463_3073# net1 0.231204f
C171 a_2051_2223# net5 0.150686f
C172 net2 a_1448_2473# 0.149541f
C173 gpo2 a_3440_4551# 1.87e-19
C174 net7 net1 0.084243f
C175 a_2101_3476# net8 0.001248f
C176 a_2509_3971# a_2427_3971# 0.005162f
C177 a_1407_3855# gno1 8.44e-20
C178 a_1499_3311# _09_.VPB 0.001545f
C179 _09_.VPB a_2377_3476# 2.07e-19
C180 net3 gpo1 0.045549f
C181 net7 _00_ 7.47e-20
C182 select0 a_3121_4551# 0.005848f
C183 select1 a_2787_4399# 7.82e-20
C184 VDD a_1407_3855# 0.189382f
C185 VDD a_2879_2223# 0.201027f
C186 a_2689_2223# net10 0.009374f
C187 VSS a_3155_2223# 0.14125f
C188 net2 _05_ 0.328235f
C189 gpo2 gpo1 1.09e-19
C190 a_2287_2741# a_2377_3476# 9.45e-20
C191 a_3155_2223# _03_ 2.5e-20
C192 net2 a_2007_4074# 0.055537f
C193 net2 a_2838_4551# 0.021582f
C194 a_2822_3855# _05_ 1.83e-19
C195 net2 _09_.VPB 0.54652f
C196 VDD a_1873_3561# 0.004308f
C197 a_2838_4551# a_2822_3855# 0.001939f
C198 net1 a_3424_3855# 0.002022f
C199 a_1683_3127# net8 2.05e-19
C200 gpo1 net5 0.049541f
C201 a_2835_2986# net1 0.08131f
C202 a_2287_2741# net2 0.231859f
C203 gno3 _02_ 2.38e-20
C204 _00_ a_3424_3855# 0.001777f
C205 a_3601_3855# VDD 0.190138f
C206 gpo0 a_2101_3476# 0.109539f
C207 VSS _01_ 0.070541f
C208 a_2835_2986# _00_ 5.47e-21
C209 net6 a_3155_3311# 1.19e-20
C210 _00_ a_3481_3476# 0.003847f
C211 gpo0 net8 5.92e-19
C212 select0 VDD 0.202684f
C213 net2 a_1875_2883# 0.136666f
C214 a_3123_2999# net1 0.129843f
C215 gpo0 a_1587_3855# 3.85e-20
C216 _01_ _03_ 0.048419f
C217 net2 FILLER_0_4_3.VPB 0.131622f
C218 net1 gno3 0.004575f
C219 a_1448_2473# _09_.VPB 0.067685f
C220 a_1499_3311# gno0 0.014566f
C221 VDD a_2427_3971# 0.10994f
C222 a_2327_2223# _02_ 2.74e-19
C223 gno0 a_2377_3476# 0.129898f
C224 VDD net3 0.224335f
C225 VSS _04_ 0.148265f
C226 _00_ a_3123_2999# 0.002755f
C227 _12_.VPB _02_ 0.062793f
C228 a_3431_2223# gpo2 0.023631f
C229 net10 _02_ 6.74e-20
C230 _04_ _03_ 8.06e-22
C231 gpo3 a_3155_2223# 5.97e-19
C232 gno2 a_3155_2223# 0.00194f
C233 VDD gpo2 0.29255f
C234 a_3431_2223# net5 3.42e-20
C235 net1 a_2327_2223# 0.033066f
C236 net1 net9 0.001873f
C237 net2 gno0 0.026337f
C238 gpo0 a_1683_3127# 3.69e-20
C239 a_1499_3311# net4 0.018726f
C240 net5 gno1 3.82e-19
C241 _12_.VPB net1 0.524087f
C242 net2 a_3318_3855# 0.007023f
C243 net4 a_2377_3476# 3.8e-19
C244 net1 net10 0.262465f
C245 _09_.VPB _05_ 1.28e-19
C246 a_2007_4074# _05_ 0.21089f
C247 net2 a_3155_3311# 0.006758f
C248 VDD net5 0.159348f
C249 VSS a_1407_3855# 0.094513f
C250 a_1677_4221# a_1587_3855# 0.004764f
C251 _01_ a_1957_2883# 3.82e-19
C252 a_2007_4074# _09_.VPB 1.99e-19
C253 VSS a_2879_2223# 0.103288f
C254 _00_ net9 0.019964f
C255 _12_.VPB _00_ 0.085785f
C256 net6 a_3155_2223# 0.304122f
C257 _00_ net10 2.08e-21
C258 a_2879_2223# _03_ 0.192462f
C259 net2 net4 0.08589f
C260 VDD a_2787_4399# 0.190451f
C261 a_2463_3073# net8 0.087486f
C262 VSS a_1873_3561# 0.003349f
C263 _04_ a_1957_2883# 6.78e-19
C264 _01_ gno2 1.16e-19
C265 net7 a_2101_3476# 0.22001f
C266 a_2822_3855# net4 5.16e-21
C267 a_2287_2741# _09_.VPB 0.053671f
C268 net7 net8 0.01152f
C269 a_1875_2883# _05_ 5.91e-20
C270 gno0 a_1448_2473# 1.25e-21
C271 a_1875_2883# _09_.VPB 0.049913f
C272 a_1875_2883# a_2007_4074# 4.04e-20
C273 VSS a_3601_3855# 0.11806f
C274 _04_ gno2 7.28e-21
C275 a_2838_4551# FILLER_0_4_3.VPB 0.04542f
C276 a_2689_2223# gpo1 1.31e-19
C277 net1 a_2235_4215# 0.133144f
C278 select0 VSS 0.167044f
C279 net1 a_2653_3476# 0.024925f
C280 select0 _03_ 1.64e-19
C281 _02_ a_2051_2223# 0.034234f
C282 net2 a_3155_2223# 0.001717f
C283 a_2287_2741# a_1875_2883# 0.0172f
C284 a_1448_2473# net4 5.53e-19
C285 VSS a_2427_3971# 0.131372f
C286 _00_ a_2235_4215# 1.34e-19
C287 a_3123_2999# a_3297_3105# 0.006584f
C288 VSS net3 0.325078f
C289 _00_ a_2653_3476# 2.67e-19
C290 net7 a_1683_3127# 2.21e-20
C291 gno0 _05_ 2.04e-20
C292 _04_ net6 4.96e-20
C293 a_3318_3855# _05_ 3.76e-20
C294 gno0 a_2007_4074# 1.61e-19
C295 a_2835_2986# net8 0.108906f
C296 gpo3 a_2879_2223# 2.94e-21
C297 a_3318_3855# _09_.VPB 2.25e-19
C298 net1 a_2051_2223# 0.043809f
C299 VSS gpo2 0.547934f
C300 a_2879_2223# gno2 0.007243f
C301 a_3155_3311# _09_.VPB 8.77e-19
C302 a_1407_2767# _02_ 0.032607f
C303 gpo2 _03_ 0.004978f
C304 gpo0 net7 0.070286f
C305 VSS net5 0.073283f
C306 net4 _05_ 0.19743f
C307 a_2287_2741# gno0 3.77e-20
C308 net2 _01_ 0.277698f
C309 a_2415_3133# gpo1 9.15e-19
C310 a_3123_2999# net8 4.13e-19
C311 a_1530_2473# gno1 5e-19
C312 net5 _03_ 4.04e-19
C313 net4 a_2007_4074# 0.108536f
C314 net4 _09_.VPB 0.065043f
C315 net6 a_2879_2223# 0.147004f
C316 VDD a_1530_2473# 0.001866f
C317 _02_ gpo1 0.006386f
C318 a_1875_2883# gno0 6.47e-21
C319 net1 a_1407_2767# 0.023828f
C320 VSS a_2787_4399# 0.11699f
C321 a_2689_2223# VDD 4.73e-19
C322 gno0 FILLER_0_4_3.VPB 4.93e-19
C323 a_3318_3855# FILLER_0_4_3.VPB 6.56e-19
C324 net2 _04_ 0.451777f
C325 select0 gno2 1.01e-19
C326 a_3155_3311# FILLER_0_4_3.VPB 4.76e-20
C327 a_1499_3311# a_1407_3855# 9.39e-19
C328 a_2509_3971# net1 0.002969f
C329 a_3123_2999# a_3141_3855# 4.19e-20
C330 net1 gpo1 0.077177f
C331 a_2101_3476# net9 7.03e-20
C332 _12_.VPB a_2101_3476# 0.062237f
C333 net9 net8 2.12e-19
C334 _12_.VPB net8 0.057086f
C335 a_2427_3971# gno2 3.94e-22
C336 a_1875_2883# net4 0.002118f
C337 gpo0 a_3481_3476# 4.56e-20
C338 gno2 net3 1.47e-19
C339 _12_.VPB a_1587_3855# 0.052044f
C340 a_2509_3971# _00_ 3.51e-19
C341 net4 FILLER_0_4_3.VPB 4.16e-21
C342 a_3155_2223# _09_.VPB 0.063076f
C343 net2 a_1407_3855# 0.249396f
C344 _00_ gpo1 6.23e-20
C345 a_3121_4551# net1 0.003252f
C346 gpo3 gpo2 0.016822f
C347 net2 a_2879_2223# 0.001672f
C348 gno2 gpo2 0.086952f
C349 gno0 a_3155_3311# 2.63e-19
C350 a_3155_3311# a_3318_3855# 1.14e-20
C351 _04_ a_1448_2473# 0.008052f
C352 a_3121_4551# _00_ 8.26e-21
C353 VDD a_2415_3133# 5.22e-19
C354 _12_.VPB a_3141_3855# 0.045488f
C355 gpo3 net5 1.06e-20
C356 gno2 net5 0.011106f
C357 _02_ gno1 0.123122f
C358 net2 a_1873_3561# 0.001151f
C359 _12_.VPB a_1683_3127# 8.16e-19
C360 gno0 net4 0.026243f
C361 _01_ _05_ 7.44e-20
C362 VDD _02_ 0.558073f
C363 net6 gpo2 0.005954f
C364 _01_ _09_.VPB 0.082504f
C365 a_3431_2223# net1 0.001379f
C366 net2 a_3601_3855# 0.001579f
C367 a_1499_3311# net3 0.002239f
C368 net1 gno1 0.074678f
C369 net3 a_2377_3476# 0.041368f
C370 a_2653_3476# net8 0.03577f
C371 gpo0 net9 7.39e-20
C372 net6 net5 2.93e-19
C373 gpo0 _12_.VPB 0.038917f
C374 select0 net2 0.379578f
C375 VDD net1 1.41714f
C376 VSS a_1530_2473# 2.93e-19
C377 a_2287_2741# _01_ 0.065112f
C378 _04_ a_2007_4074# 1.2e-20
C379 _04_ _09_.VPB 0.08635f
C380 select0 a_2822_3855# 0.26988f
C381 gpo2 a_2377_3476# 5.79e-21
C382 a_2689_2223# VSS 0.001907f
C383 net2 a_2427_3971# 0.060279f
C384 net2 net3 0.165605f
C385 VDD _00_ 0.604619f
C386 a_1875_2883# _01_ 0.107635f
C387 a_2101_3476# a_2051_2223# 2.33e-20
C388 a_2822_3855# a_2427_3971# 6.61e-19
C389 net5 a_2377_3476# 1.97e-19
C390 a_2822_3855# net3 3.84e-19
C391 a_3155_3311# a_3155_2223# 7.96e-19
C392 a_1407_3855# _05_ 7.03e-19
C393 a_2287_2741# _04_ 0.072473f
C394 net2 gpo2 0.034773f
C395 a_1407_3855# _09_.VPB 1.75e-19
C396 a_1875_2883# _04_ 0.027452f
C397 a_2879_2223# _09_.VPB 0.062897f
C398 _12_.VPB a_2934_4373# 6.37e-19
C399 net2 net5 0.0519f
C400 gpo0 a_2653_3476# 2.24e-19
C401 a_1407_2767# net8 1.12e-19
C402 _01_ gno0 8.78e-21
C403 a_3481_3476# a_3424_3855# 4.02e-19
C404 VSS a_2415_3133# 0.006037f
C405 a_2463_3073# a_2327_2223# 1.37e-19
C406 net2 a_2787_4399# 9.43e-19
C407 a_2463_3073# _12_.VPB 7.13e-19
C408 a_3601_3855# _05_ 5.39e-21
C409 net7 net9 0.002191f
C410 VSS _02_ 0.273082f
C411 net7 _12_.VPB 0.074567f
C412 a_2101_3476# gpo1 0.120482f
C413 gpo1 net8 0.052745f
C414 gno0 _04_ 1.07e-20
C415 select0 _05_ 0.002171f
C416 _02_ _03_ 4.68e-20
C417 _01_ net4 0.001208f
C418 a_2689_2223# gno2 2.26e-19
C419 select0 a_2007_4074# 9.32e-19
C420 select0 a_2838_4551# 0.030629f
C421 select0 _09_.VPB 1.62e-19
C422 gno3 a_3424_3855# 1.68e-21
C423 a_1448_2473# net5 8.26e-19
C424 a_2427_3971# _05_ 0.002611f
C425 gno3 a_3481_3476# 4.99e-21
C426 a_1683_3127# a_1407_2767# 7.37e-19
C427 net3 _05_ 1.96e-20
C428 VSS net1 1.53591f
C429 a_2427_3971# _09_.VPB 1.44e-19
C430 a_2007_4074# net3 8.96e-20
C431 net3 _09_.VPB 0.00188f
C432 net1 _03_ 0.414085f
C433 _04_ net4 2.68e-19
C434 a_2689_2223# net6 8.38e-20
C435 VSS _00_ 0.156785f
C436 gpo0 a_1407_2767# 0.003395f
C437 net9 a_3424_3855# 0.01148f
C438 a_1683_3127# gpo1 0.004604f
C439 gpo2 _09_.VPB 0.029009f
C440 _12_.VPB a_3424_3855# 0.045195f
C441 _00_ _03_ 2.23e-20
C442 _12_.VPB a_2835_2986# 0.001483f
C443 net9 a_3481_3476# 0.230747f
C444 net10 a_3424_3855# 1.48e-20
C445 a_2287_2741# net3 6.36e-20
C446 a_3121_4551# a_3141_3855# 0.001973f
C447 _12_.VPB a_3481_3476# 0.060474f
C448 select0 FILLER_0_4_3.VPB 0.010922f
C449 a_2835_2986# net10 1.1e-19
C450 a_1957_2883# _02_ 2.96e-19
C451 a_3481_3476# net10 8.52e-19
C452 gno0 a_1873_3561# 0.002605f
C453 net7 a_2653_3476# 5.41e-19
C454 _09_.VPB net5 0.091056f
C455 a_1407_3855# net4 0.005147f
C456 gno1 net8 7.96e-20
C457 a_1875_2883# net3 2.48e-20
C458 gpo0 gpo1 0.003113f
C459 a_2934_4373# select1 8.91e-19
C460 net3 FILLER_0_4_3.VPB 3.22e-19
C461 VDD a_2101_3476# 0.128916f
C462 _12_.VPB a_3123_2999# 6.21e-19
C463 a_1587_3855# gno1 1.01e-19
C464 VDD net8 0.173368f
C465 net9 gno3 3.17e-21
C466 a_3123_2999# net10 8.67e-20
C467 gno2 _02_ 1.22e-19
C468 net1 a_1957_2883# 7.28e-19
C469 VDD a_1587_3855# 0.115408f
C470 a_3601_3855# a_3318_3855# 0.003683f
C471 a_2838_4551# a_2787_4399# 0.134298f
C472 a_2287_2741# net5 6.56e-19
C473 net2 a_1530_2473# 8.47e-19
C474 gno3 net10 0.139448f
C475 gpo2 FILLER_0_4_3.VPB 2.09e-20
C476 select0 a_3318_3855# 6.4e-19
C477 net7 a_2051_2223# 8.9e-19
C478 net1 gno2 0.087277f
C479 gno0 a_2427_3971# 2.86e-19
C480 gno0 net3 0.204196f
C481 VDD a_3141_3855# 0.125966f
C482 net6 _02_ 1.36e-19
C483 a_1683_3127# gno1 0.060626f
C484 _12_.VPB net9 0.072855f
C485 net3 a_3155_3311# 5.16e-19
C486 select0 net4 4.06e-19
C487 a_2879_2223# a_3155_2223# 5.3e-19
C488 a_2327_2223# net10 0.002287f
C489 net9 net10 6.91e-21
C490 VDD a_1683_3127# 0.037512f
C491 _12_.VPB net10 2.04e-19
C492 gno0 gpo2 8.83e-20
C493 _00_ gno2 1.31e-20
C494 _01_ _04_ 0.251489f
C495 gpo2 a_3318_3855# 6.94e-19
C496 FILLER_0_4_3.VPB a_2787_4399# 0.008512f
C497 gpo2 a_3155_3311# 0.003329f
C498 a_1530_2473# a_1448_2473# 0.004767f
C499 a_2427_3971# net4 2.73e-21
C500 net1 net6 0.042251f
C501 gpo0 gno1 0.113014f
C502 a_1499_3311# _02_ 0.190762f
C503 net4 net3 0.002408f
C504 a_3121_4551# a_2934_4373# 0.159555f
C505 gno0 net5 1.29e-21
C506 gpo0 VDD 0.436425f
C507 a_2463_3073# gpo1 0.00386f
C508 VSS a_3297_3105# 0.007629f
C509 a_3424_3855# select1 0.004336f
C510 a_3297_3105# _03_ 5.76e-19
C511 _00_ net6 9.47e-19
C512 net7 gpo1 0.085308f
C513 net2 a_2415_3133# 3.56e-19
C514 a_3481_3476# select1 5.13e-20
C515 a_1499_3311# net1 0.035267f
C516 _01_ a_2879_2223# 4.52e-19
C517 net1 a_2377_3476# 0.0112f
C518 a_3424_3855# a_3440_4551# 0.001939f
C519 net2 _02_ 0.114417f
C520 a_3481_3476# a_3440_4551# 6.41e-20
C521 _12_.VPB a_2235_4215# 0.046227f
C522 net9 a_2653_3476# 7.47e-19
C523 VSS a_2101_3476# 0.105512f
C524 _12_.VPB a_2653_3476# 0.060778f
C525 VSS net8 0.391582f
C526 a_1677_4221# gno1 1.08e-19
C527 VSS a_1587_3855# 0.12794f
C528 net2 net1 1.88615f
C529 _03_ net8 0.006368f
C530 VDD a_1677_4221# 4.22e-19
C531 VDD a_2934_4373# 0.090121f
C532 net1 a_2822_3855# 0.217495f
C533 gpo2 a_3155_2223# 0.008614f
C534 a_2835_2986# gpo1 7.93e-19
C535 net2 _00_ 0.165646f
C536 a_3481_3476# gpo1 1.71e-21
C537 a_2327_2223# a_2051_2223# 5.3e-19
C538 select0 _01_ 3.3e-21
C539 _12_.VPB a_2051_2223# 1.02e-19
C540 a_1448_2473# _02_ 0.122755f
C541 VSS a_3141_3855# 0.172193f
C542 _00_ a_2822_3855# 0.126561f
C543 a_2463_3073# VDD 0.129236f
C544 net9 select1 3.65e-19
C545 a_3155_2223# net5 7.89e-20
C546 _12_.VPB select1 0.001606f
C547 net7 gno1 0.001213f
C548 _01_ a_2427_3971# 4.35e-21
C549 VSS a_1683_3127# 0.159059f
C550 _01_ net3 1.11e-19
C551 net7 VDD 0.194093f
C552 net9 a_3440_4551# 7.64e-20
C553 net1 a_1448_2473# 0.170339f
C554 _01_ gpo2 1.34e-19
C555 gpo0 VSS 0.341564f
C556 a_3121_4551# a_3123_2999# 1.59e-19
C557 _02_ _09_.VPB 0.063276f
C558 a_3431_2223# a_3424_3855# 1.09e-20
C559 gno2 net8 0.00314f
C560 select0 a_1407_3855# 3.09e-19
C561 a_3431_2223# a_3481_3476# 2.41e-20
C562 a_2327_2223# gpo1 0.005654f
C563 net9 gpo1 0.002226f
C564 a_2287_2741# a_2415_3133# 0.004764f
C565 _12_.VPB gpo1 0.013905f
C566 select0 a_2879_2223# 1.41e-20
C567 net1 _05_ 0.223818f
C568 net10 gpo1 0.001452f
C569 VDD a_3424_3855# 0.154511f
C570 VDD a_2835_2986# 0.127687f
C571 net1 a_2007_4074# 0.032005f
C572 a_2838_4551# net1 2.41e-20
C573 net1 _09_.VPB 0.349064f
C574 VDD a_3481_3476# 0.211597f
C575 _04_ net5 0.016958f
C576 a_1683_3127# a_1957_2883# 3.5e-20
C577 a_3121_4551# _12_.VPB 5.41e-19
C578 _00_ _05_ 2.4e-19
C579 a_3431_2223# gno3 0.148999f
C580 VSS a_1677_4221# 0.006151f
C581 a_1875_2883# _02_ 0.002397f
C582 VSS a_2934_4373# 0.09114f
C583 _00_ a_2007_4074# 5.79e-21
C584 _00_ _09_.VPB 0.001043f
C585 VDD a_3123_2999# 0.154092f
C586 a_2287_2741# net1 0.042316f
C587 a_2879_2223# gpo2 0.002285f
C588 net2 a_3297_3105# 6.66e-19
C589 net3 a_1873_3561# 0.011812f
C590 select0 a_3601_3855# 6.16e-20
C591 VDD gno3 0.470009f
C592 a_1499_3311# a_2101_3476# 0.002507f
C593 a_2101_3476# a_2377_3476# 5.3e-19
C594 a_1499_3311# net8 1.76e-19
C595 a_1875_2883# net1 0.048135f
C596 a_2377_3476# net8 0.197847f
C597 a_2463_3073# VSS 0.072214f
C598 a_2879_2223# net5 1.5e-19
C599 a_1499_3311# a_1587_3855# 3.09e-19
C600 net1 FILLER_0_4_3.VPB 0.001364f
C601 a_2509_3971# a_2235_4215# 3.5e-20
C602 a_3431_2223# net9 8.58e-19
C603 _12_.VPB a_3431_2223# 1.12e-19
C604 a_2463_3073# _03_ 0.002314f
C605 a_2235_4215# gpo1 2.73e-19
C606 net7 VSS 0.358556f
C607 a_2653_3476# gpo1 6.47e-19
C608 a_3431_2223# net10 0.200625f
C609 select0 a_2427_3971# 0.023337f
C610 select1 a_3440_4551# 0.259127f
C611 select0 net3 4.24e-19
C612 _12_.VPB gno1 1.48e-19
C613 gno0 _02_ 0.003141f
C614 VDD a_2327_2223# 0.149216f
C615 VDD net9 0.231582f
C616 net2 a_2101_3476# 0.028919f
C617 _12_.VPB VDD 0.728115f
C618 net2 net8 0.036688f
C619 VDD net10 0.391297f
C620 net2 a_1587_3855# 0.077927f
C621 a_2427_3971# net3 3.24e-20
C622 gno0 net1 0.030842f
C623 net1 a_3318_3855# 0.017767f
C624 gpo1 a_2051_2223# 0.012433f
C625 net4 _02_ 0.259598f
C626 net1 a_3155_3311# 4.89e-19
C627 gpo2 net3 9.89e-20
C628 _00_ gno0 1.65e-19
C629 net2 a_3141_3855# 0.016567f
C630 _00_ a_3318_3855# 0.003194f
C631 VSS a_3424_3855# 0.150239f
C632 VSS a_2835_2986# 0.104843f
C633 gpo0 a_1499_3311# 0.034289f
C634 VSS a_3481_3476# 0.141257f
C635 net3 net5 4.86e-21
C636 gpo0 a_2377_3476# 5.81e-19
C637 _00_ a_3155_3311# 0.19814f
C638 net2 a_1683_3127# 0.127798f
C639 select0 a_2787_4399# 0.012102f
C640 net1 net4 0.337599f
C641 a_3121_4551# select1 0.001676f
C642 a_2835_2986# _03_ 0.122289f
C643 a_1407_2767# gpo1 2.59e-19
C644 a_2463_3073# gno2 9.74e-19
C645 gpo2 net5 3.74e-21
C646 VDD a_2235_4215# 0.045634f
C647 _00_ net4 9.12e-20
C648 VDD a_2653_3476# 0.224108f
C649 net3 a_2787_4399# 1.27e-19
C650 VSS a_3123_2999# 0.159626f
C651 gpo0 net2 0.060123f
C652 a_3155_2223# _02_ 4.78e-20
C653 VSS gno3 0.19108f
C654 a_3123_2999# _03_ 0.110282f
C655 gno3 _03_ 3.12e-19
C656 a_2101_3476# _05_ 0.011082f
C657 a_2051_2223# gno1 0.002022f
C658 a_2101_3476# a_2007_4074# 1.62e-19
C659 net1 a_3155_2223# 0.006467f
C660 a_2101_3476# _09_.VPB 5.83e-19
C661 a_1587_3855# _05_ 0.07349f
C662 VDD a_2051_2223# 0.139815f
C663 _09_.VPB net8 0.012846f
C664 VSS a_2327_2223# 0.101183f
C665 VSS net9 0.181564f
C666 a_1587_3855# a_2007_4074# 0.017591f
C667 VDD select1 0.359874f
C668 VSS _12_.VPB 0.494511f
C669 VSS net10 0.227483f
C670 _00_ a_3155_2223# 1.83e-20
C671 a_2327_2223# _03_ 0.003128f
C672 _01_ _02_ 2.81e-19
C673 _12_.VPB _03_ 4.66e-20
C674 net2 a_1677_4221# 0.001503f
C675 VDD a_3440_4551# 0.210176f
C676 a_2463_3073# a_2377_3476# 4.64e-19
C677 gpo0 a_1448_2473# 0.003515f
C678 a_2287_2741# net8 0.016501f
C679 net10 _03_ 0.072824f
C680 net2 a_2934_4373# 0.07548f
C681 a_3141_3855# _05_ 3e-20
C682 a_2835_2986# gno2 1.5e-20
C683 _04_ a_2415_3133# 8.17e-20
C684 a_1407_2767# gno1 0.109859f
C685 net7 a_1499_3311# 0.115891f
C686 net7 a_2377_3476# 0.03289f
C687 a_2934_4373# a_2822_3855# 0.004336f
C688 VDD a_1407_2767# 0.221138f
C689 a_1875_2883# a_2101_3476# 0.00928f
C690 a_1683_3127# _05_ 1.33e-19
C691 a_1875_2883# net8 4.74e-19
C692 _04_ _02_ 0.01572f
C693 _01_ net1 0.53404f
C694 a_1683_3127# _09_.VPB 0.045434f
C695 a_2463_3073# net2 0.134082f
C696 gpo1 gno1 0.096064f
C697 a_2509_3971# VDD 0.001374f
C698 gpo3 gno3 0.206568f
C699 net7 net2 0.058965f
C700 gno3 gno2 0.004646f
C701 VDD gpo1 0.195934f
C702 _04_ net1 0.093539f
C703 gpo0 a_2007_4074# 4.16e-19
C704 gpo0 _09_.VPB 0.018313f
C705 a_1407_3855# _02_ 0.011074f
C706 VSS a_2235_4215# 0.146168f
C707 VSS a_2653_3476# 0.146592f
C708 a_2101_3476# gno0 0.021549f
C709 a_3121_4551# VDD 0.130745f
C710 a_3141_3855# FILLER_0_4_3.VPB 4.27e-19
C711 a_2879_2223# _02_ 8.14e-20
C712 gno0 net8 0.045623f
C713 a_3123_2999# net6 0.001999f
C714 a_1683_3127# a_1875_2883# 0.101254f
C715 gno0 a_1587_3855# 5.11e-20
C716 net9 gpo3 1.46e-19
C717 net6 gno3 0.004644f
C718 a_2327_2223# gno2 0.112838f
C719 _12_.VPB gno2 1.53e-19
C720 gpo3 net10 0.003316f
C721 a_1407_3855# net1 0.095088f
C722 gno2 net10 0.15439f
C723 a_1530_2473# net5 1.53e-19
C724 net1 a_2879_2223# 0.040234f
C725 gpo0 a_1875_2883# 3.42e-19
C726 VSS a_2051_2223# 0.1137f
C727 net2 a_3424_3855# 0.004493f
C728 a_2101_3476# net4 9.85e-19
C729 a_1677_4221# _05_ 8.17e-20
C730 net7 a_1448_2473# 7.15e-21
C731 net4 net8 0.003939f
C732 net2 a_2835_2986# 0.040447f
C733 gpo0 FILLER_0_4_3.VPB 2.6e-19
C734 VSS select1 0.126239f
C735 net2 a_3481_3476# 0.001017f
C736 net4 a_1587_3855# 0.026154f
C737 a_3141_3855# a_3318_3855# 0.159555f
C738 VDD a_3431_2223# 0.154305f
C739 net6 a_2327_2223# 3.72e-19
C740 a_2838_4551# a_2934_4373# 0.313533f
C741 a_2835_2986# a_2822_3855# 6.43e-20
C742 a_3141_3855# a_3155_3311# 0.009783f
C743 net1 a_1873_3561# 0.001139f
C744 a_1683_3127# gno0 3.03e-20
C745 VDD gno1 0.38374f
C746 VSS a_3440_4551# 0.208394f
C747 net6 net10 0.116149f
C748 net2 a_3123_2999# 0.184932f
C749 VSS a_1407_2767# 0.146177f
C750 a_3601_3855# net1 4.81e-19
C751 net7 _05_ 1.19e-20
C752 a_2463_3073# _09_.VPB 0.086969f
C753 a_3141_3855# net4 3.11e-22
C754 net3 _02_ 2.01e-19
C755 gpo0 gno0 0.790824f
C756 a_2327_2223# a_2377_3476# 3.05e-22
C757 net9 a_2377_3476# 3.68e-19
C758 _12_.VPB a_1499_3311# 0.067172f
C759 select0 net1 0.111065f
C760 _12_.VPB a_2377_3476# 0.060297f
C761 net7 a_2007_4074# 5.13e-20
C762 a_1683_3127# net4 0.005685f
C763 net7 _09_.VPB 0.001883f
C764 gpo0 a_3155_3311# 7.71e-20
C765 gno2 a_2653_3476# 5.64e-19
C766 a_3601_3855# _00_ 6.23e-19
C767 a_2934_4373# FILLER_0_4_3.VPB 0.120773f
C768 a_2287_2741# a_2463_3073# 0.185422f
C769 VSS gpo1 0.394879f
C770 net1 a_2427_3971# 0.172078f
C771 net1 net3 0.077714f
C772 select0 _00_ 0.068996f
C773 net2 a_2327_2223# 0.072764f
C774 net2 net9 0.001868f
C775 net2 _12_.VPB 0.229591f
C776 gpo0 net4 0.041458f
C777 _02_ net5 0.001552f
C778 net2 net10 0.054992f
C779 a_3121_4551# VSS 0.159248f
C780 _00_ a_2427_3971# 0.095678f
C781 net1 gpo2 0.07155f
C782 _12_.VPB a_2822_3855# 0.04928f
C783 _00_ net3 0.007445f
C784 gno2 a_2051_2223# 1.43e-20
C785 net7 a_1875_2883# 5.88e-20
C786 a_3121_4551# _03_ 5.49e-21
C787 a_3424_3855# _05_ 1.91e-20
C788 a_2101_3476# _01_ 2.04e-19
C789 _01_ net8 0.019674f
C790 a_3424_3855# _09_.VPB 1.13e-19
C791 net1 net5 0.105051f
C792 _00_ gpo2 0.003901f
C793 a_2835_2986# _09_.VPB 0.062491f
C794 a_3481_3476# _09_.VPB 0.001307f
C795 a_2653_3476# a_2377_3476# 5.3e-19
C796 net6 a_2051_2223# 1.9e-19
C797 a_2101_3476# _04_ 1.77e-19
C798 a_2463_3073# gno0 2.73e-20
C799 a_1957_2883# gpo1 9.32e-20
C800 _04_ net8 9.44e-19
C801 VSS a_3431_2223# 0.12041f
C802 _12_.VPB a_1448_2473# 3.17e-20
C803 a_3123_2999# _09_.VPB 0.064387f
C804 net7 gno0 0.019334f
C805 VSS gno1 0.200508f
C806 gno3 _09_.VPB 0.025899f
C807 net2 a_2235_4215# 0.184401f
C808 net2 a_2653_3476# 0.001333f
C809 VSS VDD 17.2463f
C810 net7 a_3155_3311# 1.25e-19
C811 a_1683_3127# _01_ 0.002557f
C812 gno2 gpo1 0.10388f
C813 VDD _03_ 0.384622f
C814 a_3481_3476# FILLER_0_4_3.VPB 1.17e-19
C815 a_1407_3855# a_1587_3855# 0.185422f
C816 net7 net4 0.020243f
C817 _12_.VPB _05_ 0.08189f
C818 gpo0 _01_ 1.78e-20
C819 a_1683_3127# _04_ 0.001331f
C820 a_2327_2223# _09_.VPB 0.061936f
C821 net9 _09_.VPB 0.001883f
C822 _12_.VPB a_2007_4074# 0.064732f
C823 net2 a_2051_2223# 0.001392f
C824 net10 _09_.VPB 0.088792f
C825 net6 gpo1 3.21e-20
C826 a_1499_3311# a_1407_2767# 1.79e-19
C827 net2 select1 0.019976f
C828 a_3318_3855# a_3424_3855# 0.313533f
C829 gno0 a_3481_3476# 1.1e-19
C830 gpo0 _04_ 8.71e-20
C831 a_3481_3476# a_3318_3855# 0.008873f
C832 a_2287_2741# a_2327_2223# 9.96e-20
C833 net2 a_3440_4551# 0.162139f
C834 a_2287_2741# _12_.VPB 0.001506f
C835 a_3155_3311# a_3481_3476# 0.024568f
C836 a_1530_2473# _02_ 0.001276f
C837 VDD a_1957_2883# 4.1e-19
C838 a_1499_3311# gpo1 1.19e-19
C839 a_3431_2223# gpo3 0.109562f
C840 gpo1 a_2377_3476# 0.110408f
C841 net2 a_1407_2767# 0.001661f
C842 a_3431_2223# gno2 4.68e-19
C843 a_3297_3105# gpo2 8.14e-19
C844 _12_.VPB a_1875_2883# 6.37e-19
C845 select0 net8 1.37e-20
C846 a_3123_2999# a_3318_3855# 2.06e-20
C847 net9 FILLER_0_4_3.VPB 1.04e-19
C848 gno2 gno1 8.34e-22
C849 select0 a_1587_3855# 4.71e-19
C850 a_3123_2999# a_3155_3311# 0.001353f
C851 gno3 a_3318_3855# 1.4e-21
C852 gpo0 a_1407_3855# 4.27e-20
C853 VDD gpo3 0.270382f
C854 VDD gno2 0.385961f
C855 a_2235_4215# _05_ 0.007197f
C856 a_2101_3476# net3 0.039065f
C857 net2 a_2509_3971# 7.19e-19
C858 a_2427_3971# net8 4.28e-21
C859 net3 net8 0.060274f
C860 a_2689_2223# net1 5.39e-19
C861 net2 gpo1 0.206314f
C862 a_2235_4215# a_2007_4074# 0.039733f
C863 a_3431_2223# net6 0.001454f
C864 a_2463_3073# _01_ 0.031901f
C865 select0 a_3141_3855# 0.001244f
C866 gpo2 net8 3.46e-20
C867 net6 gno1 1.13e-20
C868 gno0 net9 3.91e-19
C869 gpo0 a_1873_3561# 0.002686f
C870 a_3121_4551# net2 0.378668f
C871 net9 a_3318_3855# 2.84e-20
C872 _12_.VPB gno0 0.036135f
C873 net7 _01_ 1.1e-19
C874 _12_.VPB a_3318_3855# 0.120218f
C875 VDD net6 0.122191f
C876 VSS _03_ 0.136276f
C877 a_2287_2741# a_2235_4215# 3.22e-20
C878 a_1448_2473# a_1407_2767# 2.73e-19
C879 net10 a_3318_3855# 6.25e-20
C880 net9 a_3155_3311# 0.121931f
C881 a_2051_2223# _05_ 3.01e-21
C882 _12_.VPB a_3155_3311# 0.058947f
C883 a_3155_3311# net10 1.28e-21
C884 a_2463_3073# _04_ 1.87e-20
C885 a_2007_4074# a_2051_2223# 2.81e-21
C886 _09_.VPB a_2051_2223# 0.072393f
C887 a_1499_3311# gno1 4.17e-19
C888 a_1683_3127# net3 6.34e-19
C889 a_2838_4551# select1 4.21e-19
C890 a_2235_4215# FILLER_0_4_3.VPB 0.001637f
C891 net7 _04_ 8.57e-19
C892 select1 _09_.VPB 2.08e-20
C893 VDD a_1499_3311# 0.164378f
C894 _12_.VPB net4 0.027353f
C895 a_1448_2473# gpo1 1.64e-20
C896 VDD a_2377_3476# 0.140318f
C897 a_3123_2999# a_3155_2223# 0.002238f
C898 net1 a_2415_3133# 0.001719f
C899 gno3 a_3155_2223# 0.109558f
C900 gpo0 net3 0.253726f
C901 net2 gno1 0.126901f
C902 net1 _02_ 0.07032f
C903 a_1407_2767# _09_.VPB 0.068336f
C904 gpo3 PHY_EDGE_ROW_4_Right_4.VNB 0.589287f
C905 gno3 PHY_EDGE_ROW_4_Right_4.VNB 0.286728f
C906 gno2 PHY_EDGE_ROW_4_Right_4.VNB 0.214753f
C907 gno1 PHY_EDGE_ROW_4_Right_4.VNB 0.228206f
C908 gpo2 PHY_EDGE_ROW_4_Right_4.VNB 0.369825f
C909 gno0 PHY_EDGE_ROW_4_Right_4.VNB 0.985536f
C910 gpo1 PHY_EDGE_ROW_4_Right_4.VNB 0.236398f
C911 gpo0 PHY_EDGE_ROW_4_Right_4.VNB 0.435747f
C912 select0 PHY_EDGE_ROW_4_Right_4.VNB 0.522349f
C913 VDD PHY_EDGE_ROW_4_Right_4.VNB 8.659544f
C914 select1 PHY_EDGE_ROW_4_Right_4.VNB 0.70546f
C915 VSS PHY_EDGE_ROW_4_Right_4.VNB 7.90502f
C916 a_3431_2223# PHY_EDGE_ROW_4_Right_4.VNB 0.116639f
C917 net10 PHY_EDGE_ROW_4_Right_4.VNB 0.149646f
C918 a_3155_2223# PHY_EDGE_ROW_4_Right_4.VNB 0.113384f
C919 net6 PHY_EDGE_ROW_4_Right_4.VNB 0.151314f
C920 a_2879_2223# PHY_EDGE_ROW_4_Right_4.VNB 0.115927f
C921 a_2327_2223# PHY_EDGE_ROW_4_Right_4.VNB 0.114033f
C922 net5 PHY_EDGE_ROW_4_Right_4.VNB 0.137753f
C923 a_2051_2223# PHY_EDGE_ROW_4_Right_4.VNB 0.130178f
C924 a_1448_2473# PHY_EDGE_ROW_4_Right_4.VNB 0.115034f
C925 _03_ PHY_EDGE_ROW_4_Right_4.VNB 0.154061f
C926 _04_ PHY_EDGE_ROW_4_Right_4.VNB 0.161265f
C927 a_3123_2999# PHY_EDGE_ROW_4_Right_4.VNB 0.127927f
C928 _01_ PHY_EDGE_ROW_4_Right_4.VNB 0.137112f
C929 a_2835_2986# PHY_EDGE_ROW_4_Right_4.VNB 0.11472f
C930 a_2463_3073# PHY_EDGE_ROW_4_Right_4.VNB 0.149926f
C931 a_2287_2741# PHY_EDGE_ROW_4_Right_4.VNB 0.112385f
C932 a_1875_2883# PHY_EDGE_ROW_4_Right_4.VNB 0.105801f
C933 a_1683_3127# PHY_EDGE_ROW_4_Right_4.VNB 0.134526f
C934 a_1407_2767# PHY_EDGE_ROW_4_Right_4.VNB 0.108731f
C935 net9 PHY_EDGE_ROW_4_Right_4.VNB 0.154581f
C936 a_3481_3476# PHY_EDGE_ROW_4_Right_4.VNB 0.114121f
C937 a_3155_3311# PHY_EDGE_ROW_4_Right_4.VNB 0.114513f
C938 net3 PHY_EDGE_ROW_4_Right_4.VNB 0.139709f
C939 a_2653_3476# PHY_EDGE_ROW_4_Right_4.VNB 0.106568f
C940 net8 PHY_EDGE_ROW_4_Right_4.VNB 0.161889f
C941 a_2377_3476# PHY_EDGE_ROW_4_Right_4.VNB 0.106397f
C942 net7 PHY_EDGE_ROW_4_Right_4.VNB 0.16123f
C943 a_2101_3476# PHY_EDGE_ROW_4_Right_4.VNB 0.108228f
C944 a_1499_3311# PHY_EDGE_ROW_4_Right_4.VNB 0.12267f
C945 _02_ PHY_EDGE_ROW_4_Right_4.VNB 0.205905f
C946 a_3601_3855# PHY_EDGE_ROW_4_Right_4.VNB 0.013393f
C947 _00_ PHY_EDGE_ROW_4_Right_4.VNB 0.186938f
C948 a_3424_3855# PHY_EDGE_ROW_4_Right_4.VNB 0.101836f
C949 a_3318_3855# PHY_EDGE_ROW_4_Right_4.VNB 0.145879f
C950 a_3141_3855# PHY_EDGE_ROW_4_Right_4.VNB 0.100956f
C951 a_2822_3855# PHY_EDGE_ROW_4_Right_4.VNB 0.107457f
C952 a_2427_3971# PHY_EDGE_ROW_4_Right_4.VNB 0.104634f
C953 a_2235_4215# PHY_EDGE_ROW_4_Right_4.VNB 0.142236f
C954 net4 PHY_EDGE_ROW_4_Right_4.VNB 0.190518f
C955 _05_ PHY_EDGE_ROW_4_Right_4.VNB 0.121261f
C956 a_2007_4074# PHY_EDGE_ROW_4_Right_4.VNB 0.112198f
C957 a_1587_3855# PHY_EDGE_ROW_4_Right_4.VNB 0.104898f
C958 net1 PHY_EDGE_ROW_4_Right_4.VNB 1.2353f
C959 a_1407_3855# PHY_EDGE_ROW_4_Right_4.VNB 0.143524f
C960 a_2787_4399# PHY_EDGE_ROW_4_Right_4.VNB 0.013393f
C961 a_3440_4551# PHY_EDGE_ROW_4_Right_4.VNB 0.114511f
C962 net2 PHY_EDGE_ROW_4_Right_4.VNB 1.3614f
C963 a_3121_4551# PHY_EDGE_ROW_4_Right_4.VNB 0.107124f
C964 a_2934_4373# PHY_EDGE_ROW_4_Right_4.VNB 0.149918f
C965 a_2838_4551# PHY_EDGE_ROW_4_Right_4.VNB 0.107834f
C966 _09_.VPB PHY_EDGE_ROW_4_Right_4.VNB 4.97174f
C967 _12_.VPB PHY_EDGE_ROW_4_Right_4.VNB 4.97174f
C968 FILLER_0_4_3.VPB PHY_EDGE_ROW_4_Right_4.VNB 2.81966f
C969 VDD.n0 PHY_EDGE_ROW_4_Right_4.VNB 0.005554f
C970 VDD.n1 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C971 VDD.n2 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C972 VDD.n3 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C973 VDD.n4 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C974 VDD.n5 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C975 VDD.n6 PHY_EDGE_ROW_4_Right_4.VNB 0.489933f
C976 VDD.n7 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C977 VDD.n8 PHY_EDGE_ROW_4_Right_4.VNB 0.034024f
C978 VDD.n9 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C979 VDD.n10 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C980 VDD.t60 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C981 VDD.t100 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C982 VDD.n12 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C983 VDD.t61 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C984 VDD.n13 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C985 VDD.n14 PHY_EDGE_ROW_4_Right_4.VNB 0.018066f
C986 VDD.n15 PHY_EDGE_ROW_4_Right_4.VNB 0.005063f
C987 VDD.t74 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C988 VDD.t93 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C989 VDD.n17 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C990 VDD.t75 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C991 VDD.n18 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C992 VDD.t87 PHY_EDGE_ROW_4_Right_4.VNB 0.00988f
C993 VDD.t51 PHY_EDGE_ROW_4_Right_4.VNB 0.002866f
C994 VDD.n19 PHY_EDGE_ROW_4_Right_4.VNB 0.01075f
C995 VDD.t53 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C996 VDD.t34 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C997 VDD.n20 PHY_EDGE_ROW_4_Right_4.VNB 0.010496f
C998 VDD.n21 PHY_EDGE_ROW_4_Right_4.VNB 0.042225f
C999 VDD.n22 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1000 VDD.t85 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1001 VDD.t19 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1002 VDD.n23 PHY_EDGE_ROW_4_Right_4.VNB 0.010304f
C1003 VDD.t55 PHY_EDGE_ROW_4_Right_4.VNB 0.00988f
C1004 VDD.t14 PHY_EDGE_ROW_4_Right_4.VNB 0.002866f
C1005 VDD.n24 PHY_EDGE_ROW_4_Right_4.VNB 0.01068f
C1006 VDD.n25 PHY_EDGE_ROW_4_Right_4.VNB 0.016627f
C1007 VDD.t20 PHY_EDGE_ROW_4_Right_4.VNB 0.00988f
C1008 VDD.t41 PHY_EDGE_ROW_4_Right_4.VNB 0.002866f
C1009 VDD.n26 PHY_EDGE_ROW_4_Right_4.VNB 0.010707f
C1010 VDD.n27 PHY_EDGE_ROW_4_Right_4.VNB 0.018969f
C1011 VDD.t66 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1012 VDD.t98 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C1013 VDD.n29 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C1014 VDD.t67 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1015 VDD.n30 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C1016 VDD.t3 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1017 VDD.t56 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1018 VDD.n31 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1019 VDD.n32 PHY_EDGE_ROW_4_Right_4.VNB 0.027607f
C1020 VDD.n33 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1021 VDD.n34 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1022 VDD.n35 PHY_EDGE_ROW_4_Right_4.VNB 0.397065f
C1023 VDD.n37 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1024 VDD.n38 PHY_EDGE_ROW_4_Right_4.VNB 0.008934f
C1025 VDD.n39 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1026 VDD.t8 PHY_EDGE_ROW_4_Right_4.VNB 0.003561f
C1027 VDD.t50 PHY_EDGE_ROW_4_Right_4.VNB 0.005584f
C1028 VDD.n40 PHY_EDGE_ROW_4_Right_4.VNB 0.016424f
C1029 VDD.t1 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1030 VDD.t16 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1031 VDD.n41 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1032 VDD.n42 PHY_EDGE_ROW_4_Right_4.VNB 0.028485f
C1033 VDD.n43 PHY_EDGE_ROW_4_Right_4.VNB 0.010721f
C1034 VDD.t25 PHY_EDGE_ROW_4_Right_4.VNB 0.009541f
C1035 VDD.n44 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1036 VDD.t31 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1037 VDD.t46 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1038 VDD.n45 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1039 VDD.t32 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1040 VDD.t36 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1041 VDD.n46 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1042 VDD.n47 PHY_EDGE_ROW_4_Right_4.VNB 0.016578f
C1043 VDD.n48 PHY_EDGE_ROW_4_Right_4.VNB 0.006258f
C1044 VDD.n49 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1045 VDD.t12 PHY_EDGE_ROW_4_Right_4.VNB 0.02186f
C1046 VDD.n50 PHY_EDGE_ROW_4_Right_4.VNB 0.034002f
C1047 VDD.t45 PHY_EDGE_ROW_4_Right_4.VNB 0.019484f
C1048 VDD.t11 PHY_EDGE_ROW_4_Right_4.VNB 0.007327f
C1049 VDD.n51 PHY_EDGE_ROW_4_Right_4.VNB 0.011051f
C1050 VDD.n52 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1051 VDD.t47 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1052 VDD.t39 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1053 VDD.n53 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1054 VDD.t48 PHY_EDGE_ROW_4_Right_4.VNB 0.003561f
C1055 VDD.t26 PHY_EDGE_ROW_4_Right_4.VNB 0.002345f
C1056 VDD.n54 PHY_EDGE_ROW_4_Right_4.VNB 0.006152f
C1057 VDD.n55 PHY_EDGE_ROW_4_Right_4.VNB 0.01082f
C1058 VDD.t80 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1059 VDD.t90 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C1060 VDD.n57 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C1061 VDD.t81 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1062 VDD.n58 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C1063 VDD.t62 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1064 VDD.t99 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C1065 VDD.n60 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C1066 VDD.t63 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1067 VDD.n61 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C1068 VDD.n62 PHY_EDGE_ROW_4_Right_4.VNB 0.039055f
C1069 VDD.n63 PHY_EDGE_ROW_4_Right_4.VNB 0.007459f
C1070 VDD.n64 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1071 VDD.n65 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1072 VDD.n66 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1073 VDD.n67 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1074 VDD.n68 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1075 VDD.n69 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1076 VDD.n70 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1077 VDD.n71 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1078 VDD.n72 PHY_EDGE_ROW_4_Right_4.VNB 0.006552f
C1079 VDD.n73 PHY_EDGE_ROW_4_Right_4.VNB 0.004268f
C1080 VDD.n74 PHY_EDGE_ROW_4_Right_4.VNB 0.008948f
C1081 VDD.n75 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1082 VDD.n77 PHY_EDGE_ROW_4_Right_4.VNB 0.010646f
C1083 VDD.n78 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1084 VDD.n79 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1085 VDD.n80 PHY_EDGE_ROW_4_Right_4.VNB 0.006552f
C1086 VDD.t88 PHY_EDGE_ROW_4_Right_4.VNB 0.032488f
C1087 VDD.n81 PHY_EDGE_ROW_4_Right_4.VNB 0.049158f
C1088 VDD.n82 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1089 VDD.n83 PHY_EDGE_ROW_4_Right_4.VNB 0.009474f
C1090 VDD.n84 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C1091 VDD.n85 PHY_EDGE_ROW_4_Right_4.VNB 0.023022f
C1092 VDD.n86 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1093 VDD.n87 PHY_EDGE_ROW_4_Right_4.VNB 0.023022f
C1094 VDD.n88 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1095 VDD.t95 PHY_EDGE_ROW_4_Right_4.VNB 0.225277f
C1096 VDD.n89 PHY_EDGE_ROW_4_Right_4.VNB 0.022271f
C1097 VDD.n90 PHY_EDGE_ROW_4_Right_4.VNB 0.007459f
C1098 VDD.t71 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1099 VDD.n91 PHY_EDGE_ROW_4_Right_4.VNB 0.0271f
C1100 VDD.n92 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1101 VDD.n93 PHY_EDGE_ROW_4_Right_4.VNB 0.003367f
C1102 VDD.n94 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1103 VDD.n95 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1104 VDD.n96 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C1105 VDD.n97 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1106 VDD.n98 PHY_EDGE_ROW_4_Right_4.VNB 0.010042f
C1107 VDD.n99 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1108 VDD.t23 PHY_EDGE_ROW_4_Right_4.VNB 0.002866f
C1109 VDD.t35 PHY_EDGE_ROW_4_Right_4.VNB 0.00988f
C1110 VDD.n100 PHY_EDGE_ROW_4_Right_4.VNB 0.01054f
C1111 VDD.n101 PHY_EDGE_ROW_4_Right_4.VNB 0.011039f
C1112 VDD.n102 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1113 VDD.t43 PHY_EDGE_ROW_4_Right_4.VNB 0.002866f
C1114 VDD.t17 PHY_EDGE_ROW_4_Right_4.VNB 0.00988f
C1115 VDD.n103 PHY_EDGE_ROW_4_Right_4.VNB 0.01054f
C1116 VDD.n104 PHY_EDGE_ROW_4_Right_4.VNB 0.012492f
C1117 VDD.t96 PHY_EDGE_ROW_4_Right_4.VNB 0.032488f
C1118 VDD.t64 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1119 VDD.n105 PHY_EDGE_ROW_4_Right_4.VNB 0.04209f
C1120 VDD.n106 PHY_EDGE_ROW_4_Right_4.VNB 0.040389f
C1121 VDD.n107 PHY_EDGE_ROW_4_Right_4.VNB 0.049158f
C1122 VDD.t65 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1123 VDD.n108 PHY_EDGE_ROW_4_Right_4.VNB 0.00912f
C1124 VDD.n109 PHY_EDGE_ROW_4_Right_4.VNB 0.01832f
C1125 VDD.n110 PHY_EDGE_ROW_4_Right_4.VNB 0.018066f
C1126 VDD.n111 PHY_EDGE_ROW_4_Right_4.VNB 0.010324f
C1127 VDD.n112 PHY_EDGE_ROW_4_Right_4.VNB 0.006021f
C1128 VDD.n113 PHY_EDGE_ROW_4_Right_4.VNB 0.008032f
C1129 VDD.n114 PHY_EDGE_ROW_4_Right_4.VNB 0.017074f
C1130 VDD.n115 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1131 VDD.n116 PHY_EDGE_ROW_4_Right_4.VNB 0.005947f
C1132 VDD.n117 PHY_EDGE_ROW_4_Right_4.VNB 0.006469f
C1133 VDD.n118 PHY_EDGE_ROW_4_Right_4.VNB 0.006045f
C1134 VDD.n119 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1135 VDD.n120 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1136 VDD.n121 PHY_EDGE_ROW_4_Right_4.VNB 0.009738f
C1137 VDD.n122 PHY_EDGE_ROW_4_Right_4.VNB 0.006117f
C1138 VDD.t52 PHY_EDGE_ROW_4_Right_4.VNB 0.002866f
C1139 VDD.t30 PHY_EDGE_ROW_4_Right_4.VNB 0.00988f
C1140 VDD.n123 PHY_EDGE_ROW_4_Right_4.VNB 0.01054f
C1141 VDD.n124 PHY_EDGE_ROW_4_Right_4.VNB 0.010527f
C1142 VDD.n125 PHY_EDGE_ROW_4_Right_4.VNB 0.006187f
C1143 VDD.n126 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1144 VDD.n127 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1145 VDD.n128 PHY_EDGE_ROW_4_Right_4.VNB 0.014493f
C1146 VDD.n129 PHY_EDGE_ROW_4_Right_4.VNB 0.005732f
C1147 VDD.t94 PHY_EDGE_ROW_4_Right_4.VNB 0.032488f
C1148 VDD.n130 PHY_EDGE_ROW_4_Right_4.VNB 0.040389f
C1149 VDD.n131 PHY_EDGE_ROW_4_Right_4.VNB 0.049158f
C1150 VDD.t70 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1151 VDD.n132 PHY_EDGE_ROW_4_Right_4.VNB 0.00912f
C1152 VDD.n133 PHY_EDGE_ROW_4_Right_4.VNB 0.01832f
C1153 VDD.n134 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1154 VDD.n135 PHY_EDGE_ROW_4_Right_4.VNB 0.004591f
C1155 VDD.n136 PHY_EDGE_ROW_4_Right_4.VNB 0.006552f
C1156 VDD.n137 PHY_EDGE_ROW_4_Right_4.VNB 0.008934f
C1157 VDD.n138 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1158 VDD.n139 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1159 VDD.n140 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1160 VDD.n141 PHY_EDGE_ROW_4_Right_4.VNB 0.391771f
C1161 VDD.n142 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1162 VDD.n143 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1163 VDD.n144 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1164 VDD.n145 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1165 VDD.n146 PHY_EDGE_ROW_4_Right_4.VNB 0.004666f
C1166 VDD.n147 PHY_EDGE_ROW_4_Right_4.VNB 0.017968f
C1167 VDD.t68 PHY_EDGE_ROW_4_Right_4.VNB 0.017009f
C1168 VDD.n148 PHY_EDGE_ROW_4_Right_4.VNB 0.013214f
C1169 VDD.n149 PHY_EDGE_ROW_4_Right_4.VNB 0.008927f
C1170 VDD.n150 PHY_EDGE_ROW_4_Right_4.VNB 0.01489f
C1171 VDD.n151 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1172 VDD.n152 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1173 VDD.n153 PHY_EDGE_ROW_4_Right_4.VNB 0.023022f
C1174 VDD.n154 PHY_EDGE_ROW_4_Right_4.VNB 0.01764f
C1175 VDD.n155 PHY_EDGE_ROW_4_Right_4.VNB 0.105224f
C1176 VDD.n156 PHY_EDGE_ROW_4_Right_4.VNB 0.01689f
C1177 VDD.n157 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1178 VDD.n158 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1179 VDD.n159 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1180 VDD.n160 PHY_EDGE_ROW_4_Right_4.VNB 0.023022f
C1181 VDD.n161 PHY_EDGE_ROW_4_Right_4.VNB 0.023022f
C1182 VDD.n162 PHY_EDGE_ROW_4_Right_4.VNB 0.023022f
C1183 VDD.n163 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1184 VDD.n164 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1185 VDD.n165 PHY_EDGE_ROW_4_Right_4.VNB 0.017669f
C1186 VDD.n166 PHY_EDGE_ROW_4_Right_4.VNB 0.022271f
C1187 VDD.t69 PHY_EDGE_ROW_4_Right_4.VNB 0.017009f
C1188 VDD.n167 PHY_EDGE_ROW_4_Right_4.VNB 0.013214f
C1189 VDD.t82 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1190 VDD.n168 PHY_EDGE_ROW_4_Right_4.VNB 0.00912f
C1191 VDD.n169 PHY_EDGE_ROW_4_Right_4.VNB 0.017982f
C1192 VDD.n170 PHY_EDGE_ROW_4_Right_4.VNB 0.009091f
C1193 VDD.n171 PHY_EDGE_ROW_4_Right_4.VNB 0.002283f
C1194 VDD.n172 PHY_EDGE_ROW_4_Right_4.VNB 0.007445f
C1195 VDD.n173 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1196 VDD.n174 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1197 VDD.n175 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1198 VDD.n176 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1199 VDD.n177 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1200 VDD.n178 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1201 VDD.n179 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1202 VDD.n180 PHY_EDGE_ROW_4_Right_4.VNB 0.040389f
C1203 VDD.t83 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1204 VDD.n181 PHY_EDGE_ROW_4_Right_4.VNB 0.04209f
C1205 VDD.n182 PHY_EDGE_ROW_4_Right_4.VNB 0.00476f
C1206 VDD.n183 PHY_EDGE_ROW_4_Right_4.VNB 0.008948f
C1207 VDD.n184 PHY_EDGE_ROW_4_Right_4.VNB 0.009474f
C1208 VDD.n185 PHY_EDGE_ROW_4_Right_4.VNB 0.010646f
C1209 VDD.n186 PHY_EDGE_ROW_4_Right_4.VNB 0.391771f
C1210 VDD.n187 PHY_EDGE_ROW_4_Right_4.VNB 0.436772f
C1211 VDD.n188 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1212 VDD.n189 PHY_EDGE_ROW_4_Right_4.VNB 0.195885f
C1213 VDD.n190 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1214 VDD.n191 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C1215 VDD.n192 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1216 VDD.n193 PHY_EDGE_ROW_4_Right_4.VNB 0.001985f
C1217 VDD.n194 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1218 VDD.n195 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C1219 VDD.t86 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1220 VDD.t21 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1221 VDD.n196 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1222 VDD.n197 PHY_EDGE_ROW_4_Right_4.VNB 0.026306f
C1223 VDD.n198 PHY_EDGE_ROW_4_Right_4.VNB 0.016578f
C1224 VDD.t0 PHY_EDGE_ROW_4_Right_4.VNB 0.00175f
C1225 VDD.t22 PHY_EDGE_ROW_4_Right_4.VNB 0.004692f
C1226 VDD.n199 PHY_EDGE_ROW_4_Right_4.VNB 0.021417f
C1227 VDD.n200 PHY_EDGE_ROW_4_Right_4.VNB 0.022584f
C1228 VDD.n201 PHY_EDGE_ROW_4_Right_4.VNB 0.016578f
C1229 VDD.t57 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1230 VDD.t40 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1231 VDD.n202 PHY_EDGE_ROW_4_Right_4.VNB 0.010304f
C1232 VDD.t2 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1233 VDD.t49 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1234 VDD.n203 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1235 VDD.n204 PHY_EDGE_ROW_4_Right_4.VNB 0.028485f
C1236 VDD.n205 PHY_EDGE_ROW_4_Right_4.VNB 0.018066f
C1237 VDD.t72 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1238 VDD.t91 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C1239 VDD.n207 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C1240 VDD.t73 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1241 VDD.n208 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C1242 VDD.n209 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1243 VDD.n210 PHY_EDGE_ROW_4_Right_4.VNB 0.034024f
C1244 VDD.n211 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1245 VDD.n212 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C1246 VDD.n213 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1247 VDD.n215 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1248 VDD.n216 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1249 VDD.n217 PHY_EDGE_ROW_4_Right_4.VNB 0.008178f
C1250 VDD.n218 PHY_EDGE_ROW_4_Right_4.VNB 0.013311f
C1251 VDD.n219 PHY_EDGE_ROW_4_Right_4.VNB 0.010781f
C1252 VDD.n220 PHY_EDGE_ROW_4_Right_4.VNB 0.195885f
C1253 VDD.n221 PHY_EDGE_ROW_4_Right_4.VNB 0.518832f
C1254 VDD.n222 PHY_EDGE_ROW_4_Right_4.VNB 1.28627f
C1255 VDD.n223 PHY_EDGE_ROW_4_Right_4.VNB 0.325813f
C1256 VDD.n224 PHY_EDGE_ROW_4_Right_4.VNB 0.436772f
C1257 VDD.n225 PHY_EDGE_ROW_4_Right_4.VNB 0.010646f
C1258 VDD.n226 PHY_EDGE_ROW_4_Right_4.VNB 0.009474f
C1259 VDD.n227 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1260 VDD.n228 PHY_EDGE_ROW_4_Right_4.VNB 0.007445f
C1261 VDD.n229 PHY_EDGE_ROW_4_Right_4.VNB 0.005063f
C1262 VDD.t78 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1263 VDD.t89 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C1264 VDD.n231 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C1265 VDD.t79 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1266 VDD.n232 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C1267 VDD.n233 PHY_EDGE_ROW_4_Right_4.VNB 0.039055f
C1268 VDD.n234 PHY_EDGE_ROW_4_Right_4.VNB 0.004289f
C1269 VDD.n235 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1270 VDD.n236 PHY_EDGE_ROW_4_Right_4.VNB 0.011614f
C1271 VDD.n237 PHY_EDGE_ROW_4_Right_4.VNB 0.008338f
C1272 VDD.n238 PHY_EDGE_ROW_4_Right_4.VNB 0.002461f
C1273 VDD.t6 PHY_EDGE_ROW_4_Right_4.VNB 0.009461f
C1274 VDD.n239 PHY_EDGE_ROW_4_Right_4.VNB 0.020989f
C1275 VDD.n240 PHY_EDGE_ROW_4_Right_4.VNB 0.004113f
C1276 VDD.n241 PHY_EDGE_ROW_4_Right_4.VNB 0.024911f
C1277 VDD.n242 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1278 VDD.n243 PHY_EDGE_ROW_4_Right_4.VNB 0.01082f
C1279 VDD.n244 PHY_EDGE_ROW_4_Right_4.VNB 0.004711f
C1280 VDD.n245 PHY_EDGE_ROW_4_Right_4.VNB 0.005309f
C1281 VDD.t38 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1282 VDD.t5 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1283 VDD.n246 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1284 VDD.n247 PHY_EDGE_ROW_4_Right_4.VNB 0.027325f
C1285 VDD.n248 PHY_EDGE_ROW_4_Right_4.VNB 0.01082f
C1286 VDD.n249 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1287 VDD.n250 PHY_EDGE_ROW_4_Right_4.VNB 0.012805f
C1288 VDD.t13 PHY_EDGE_ROW_4_Right_4.VNB 0.022269f
C1289 VDD.n251 PHY_EDGE_ROW_4_Right_4.VNB 0.030894f
C1290 VDD.n252 PHY_EDGE_ROW_4_Right_4.VNB 0.00546f
C1291 VDD.n253 PHY_EDGE_ROW_4_Right_4.VNB 0.00443f
C1292 VDD.t7 PHY_EDGE_ROW_4_Right_4.VNB 0.002345f
C1293 VDD.t4 PHY_EDGE_ROW_4_Right_4.VNB 0.003561f
C1294 VDD.n254 PHY_EDGE_ROW_4_Right_4.VNB 0.006152f
C1295 VDD.t27 PHY_EDGE_ROW_4_Right_4.VNB 0.022216f
C1296 VDD.n255 PHY_EDGE_ROW_4_Right_4.VNB 0.046525f
C1297 VDD.t84 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1298 VDD.t33 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1299 VDD.n256 PHY_EDGE_ROW_4_Right_4.VNB 0.010304f
C1300 VDD.t28 PHY_EDGE_ROW_4_Right_4.VNB 0.007329f
C1301 VDD.t54 PHY_EDGE_ROW_4_Right_4.VNB 0.019482f
C1302 VDD.n257 PHY_EDGE_ROW_4_Right_4.VNB 0.011051f
C1303 VDD.n258 PHY_EDGE_ROW_4_Right_4.VNB 0.029709f
C1304 VDD.t44 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1305 VDD.t18 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1306 VDD.n259 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1307 VDD.n260 PHY_EDGE_ROW_4_Right_4.VNB 0.027607f
C1308 VDD.t24 PHY_EDGE_ROW_4_Right_4.VNB 0.003561f
C1309 VDD.t29 PHY_EDGE_ROW_4_Right_4.VNB 0.005584f
C1310 VDD.n261 PHY_EDGE_ROW_4_Right_4.VNB 0.016424f
C1311 VDD.n262 PHY_EDGE_ROW_4_Right_4.VNB 0.006469f
C1312 VDD.n263 PHY_EDGE_ROW_4_Right_4.VNB 0.010721f
C1313 VDD.t9 PHY_EDGE_ROW_4_Right_4.VNB 0.009392f
C1314 VDD.t10 PHY_EDGE_ROW_4_Right_4.VNB 0.003561f
C1315 VDD.t37 PHY_EDGE_ROW_4_Right_4.VNB 0.005377f
C1316 VDD.n264 PHY_EDGE_ROW_4_Right_4.VNB 0.016067f
C1317 VDD.t15 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1318 VDD.t42 PHY_EDGE_ROW_4_Right_4.VNB 0.004738f
C1319 VDD.n265 PHY_EDGE_ROW_4_Right_4.VNB 0.010526f
C1320 VDD.n266 PHY_EDGE_ROW_4_Right_4.VNB 0.028485f
C1321 VDD.n267 PHY_EDGE_ROW_4_Right_4.VNB 0.002283f
C1322 VDD.n268 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1323 VDD.n269 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1324 VDD.n270 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1325 VDD.n271 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1326 VDD.n272 PHY_EDGE_ROW_4_Right_4.VNB 0.006552f
C1327 VDD.n273 PHY_EDGE_ROW_4_Right_4.VNB 0.004289f
C1328 VDD.t58 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1329 VDD.t97 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C1330 VDD.n275 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C1331 VDD.t59 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1332 VDD.n276 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C1333 VDD.n277 PHY_EDGE_ROW_4_Right_4.VNB 0.007445f
C1334 VDD.n278 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1335 VDD.n279 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1336 VDD.n280 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1337 VDD.n281 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1338 VDD.t76 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1339 VDD.t92 PHY_EDGE_ROW_4_Right_4.VNB 0.033078f
C1340 VDD.n283 PHY_EDGE_ROW_4_Right_4.VNB 0.084809f
C1341 VDD.t77 PHY_EDGE_ROW_4_Right_4.VNB 0.015585f
C1342 VDD.n284 PHY_EDGE_ROW_4_Right_4.VNB 0.046196f
C1343 VDD.n285 PHY_EDGE_ROW_4_Right_4.VNB 0.039055f
C1344 VDD.n286 PHY_EDGE_ROW_4_Right_4.VNB 0.004268f
C1345 VDD.n287 PHY_EDGE_ROW_4_Right_4.VNB 0.008948f
C1346 VDD.n288 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1347 VDD.n289 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1348 VDD.n290 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1349 VDD.n291 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1350 VDD.n292 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1351 VDD.n293 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1352 VDD.n294 PHY_EDGE_ROW_4_Right_4.VNB 0.009146f
C1353 VDD.n295 PHY_EDGE_ROW_4_Right_4.VNB 0.017669f
C1354 VDD.n296 PHY_EDGE_ROW_4_Right_4.VNB 0.016677f
C1355 VDD.n297 PHY_EDGE_ROW_4_Right_4.VNB 0.003199f
C1356 VDD.n298 PHY_EDGE_ROW_4_Right_4.VNB 0.024076f
C1357 VDD.n299 PHY_EDGE_ROW_4_Right_4.VNB 0.025796f
C1358 VDD.n300 PHY_EDGE_ROW_4_Right_4.VNB 0.00334f
C1359 VDD.n301 PHY_EDGE_ROW_4_Right_4.VNB 0.006469f
C1360 VDD.n302 PHY_EDGE_ROW_4_Right_4.VNB 0.015783f
C1361 VDD.n303 PHY_EDGE_ROW_4_Right_4.VNB 0.011614f
C1362 VDD.n304 PHY_EDGE_ROW_4_Right_4.VNB 0.016578f
C1363 VDD.n305 PHY_EDGE_ROW_4_Right_4.VNB 0.005379f
C1364 VDD.n306 PHY_EDGE_ROW_4_Right_4.VNB 0.024765f
C1365 VDD.n307 PHY_EDGE_ROW_4_Right_4.VNB 0.01082f
C1366 VDD.n308 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1367 VDD.n309 PHY_EDGE_ROW_4_Right_4.VNB 0.016578f
C1368 VDD.n310 PHY_EDGE_ROW_4_Right_4.VNB 0.005309f
C1369 VDD.n311 PHY_EDGE_ROW_4_Right_4.VNB 0.004922f
C1370 VDD.n312 PHY_EDGE_ROW_4_Right_4.VNB 0.01082f
C1371 VDD.n313 PHY_EDGE_ROW_4_Right_4.VNB 0.01489f
C1372 VDD.n314 PHY_EDGE_ROW_4_Right_4.VNB 0.0247f
C1373 VDD.n315 PHY_EDGE_ROW_4_Right_4.VNB 0.005379f
C1374 VDD.n316 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1375 VDD.n317 PHY_EDGE_ROW_4_Right_4.VNB 0.007346f
C1376 VDD.n318 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1377 VDD.n319 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1378 VDD.n320 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1379 VDD.n321 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1380 VDD.n322 PHY_EDGE_ROW_4_Right_4.VNB 0.006552f
C1381 VDD.n323 PHY_EDGE_ROW_4_Right_4.VNB 0.007246f
C1382 VDD.n324 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1383 VDD.n325 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1384 VDD.n326 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1385 VDD.n327 PHY_EDGE_ROW_4_Right_4.VNB 0.436772f
C1386 VDD.n328 PHY_EDGE_ROW_4_Right_4.VNB 0.360006f
C1387 VDD.n329 PHY_EDGE_ROW_4_Right_4.VNB 1.28627f
C1388 VDD.n330 PHY_EDGE_ROW_4_Right_4.VNB 0.518832f
C1389 VDD.n331 PHY_EDGE_ROW_4_Right_4.VNB 0.360006f
C1390 VDD.n332 PHY_EDGE_ROW_4_Right_4.VNB 0.397065f
C1391 VDD.n333 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1392 VDD.n334 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1393 VDD.n335 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1394 VDD.n336 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1395 VDD.n337 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1396 VDD.n338 PHY_EDGE_ROW_4_Right_4.VNB 0.00675f
C1397 VDD.n339 PHY_EDGE_ROW_4_Right_4.VNB 0.002283f
C1398 VDD.n340 PHY_EDGE_ROW_4_Right_4.VNB 0.004219f
C1399 VDD.n341 PHY_EDGE_ROW_4_Right_4.VNB 0.019668f
C1400 VDD.n342 PHY_EDGE_ROW_4_Right_4.VNB 0.027396f
C1401 VDD.n343 PHY_EDGE_ROW_4_Right_4.VNB 0.003586f
C1402 VDD.n344 PHY_EDGE_ROW_4_Right_4.VNB 0.029709f
C1403 VDD.n345 PHY_EDGE_ROW_4_Right_4.VNB 0.001934f
C1404 VDD.n346 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1405 VDD.n347 PHY_EDGE_ROW_4_Right_4.VNB 0.016478f
C1406 VDD.n348 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1407 VDD.n349 PHY_EDGE_ROW_4_Right_4.VNB 0.005309f
C1408 VDD.n350 PHY_EDGE_ROW_4_Right_4.VNB 0.027325f
C1409 VDD.n351 PHY_EDGE_ROW_4_Right_4.VNB 0.026341f
C1410 VDD.n352 PHY_EDGE_ROW_4_Right_4.VNB 0.030641f
C1411 VDD.n353 PHY_EDGE_ROW_4_Right_4.VNB 0.0045f
C1412 VDD.n354 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1413 VDD.n355 PHY_EDGE_ROW_4_Right_4.VNB 0.01489f
C1414 VDD.n356 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1415 VDD.n357 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1416 VDD.n358 PHY_EDGE_ROW_4_Right_4.VNB 0.010646f
C1417 VDD.n359 PHY_EDGE_ROW_4_Right_4.VNB 0.009474f
C1418 VDD.n360 PHY_EDGE_ROW_4_Right_4.VNB 0.007459f
C1419 VDD.n361 PHY_EDGE_ROW_4_Right_4.VNB 0.004666f
C1420 VDD.n362 PHY_EDGE_ROW_4_Right_4.VNB 0.004219f
C1421 VDD.n363 PHY_EDGE_ROW_4_Right_4.VNB 0.024765f
C1422 VDD.n364 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1423 VDD.n365 PHY_EDGE_ROW_4_Right_4.VNB 0.006552f
C1424 VDD.n366 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1425 VDD.n367 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1426 VDD.n368 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1427 VDD.n369 PHY_EDGE_ROW_4_Right_4.VNB 0.010646f
C1428 VDD.n370 PHY_EDGE_ROW_4_Right_4.VNB 0.009474f
C1429 VDD.n371 PHY_EDGE_ROW_4_Right_4.VNB 0.006962f
C1430 VDD.n372 PHY_EDGE_ROW_4_Right_4.VNB 0.009132f
C1431 VDD.n373 PHY_EDGE_ROW_4_Right_4.VNB 0.004289f
C1432 VDD.n374 PHY_EDGE_ROW_4_Right_4.VNB 0.045321f
C1433 VDD.n375 PHY_EDGE_ROW_4_Right_4.VNB 0.005063f
C1434 VDD.n376 PHY_EDGE_ROW_4_Right_4.VNB 0.01082f
C1435 VDD.n377 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1436 VDD.n378 PHY_EDGE_ROW_4_Right_4.VNB 0.02354f
C1437 VDD.n379 PHY_EDGE_ROW_4_Right_4.VNB 0.006469f
C1438 VDD.n380 PHY_EDGE_ROW_4_Right_4.VNB 0.004992f
C1439 VDD.n381 PHY_EDGE_ROW_4_Right_4.VNB 0.018265f
C1440 VDD.n382 PHY_EDGE_ROW_4_Right_4.VNB 0.016578f
C1441 VDD.n383 PHY_EDGE_ROW_4_Right_4.VNB 0.01082f
C1442 VDD.n384 PHY_EDGE_ROW_4_Right_4.VNB 0.004219f
C1443 VDD.n385 PHY_EDGE_ROW_4_Right_4.VNB 0.039055f
C1444 VDD.n386 PHY_EDGE_ROW_4_Right_4.VNB 0.006353f
C1445 VDD.n387 PHY_EDGE_ROW_4_Right_4.VNB 0.007445f
C1446 VDD.n388 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1447 VDD.n389 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1448 VDD.n390 PHY_EDGE_ROW_4_Right_4.VNB 0.004897f
C1449 VDD.n391 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1450 VDD.n392 PHY_EDGE_ROW_4_Right_4.VNB 0.008178f
C1451 VDD.n393 PHY_EDGE_ROW_4_Right_4.VNB 0.0134f
C1452 VDD.n394 PHY_EDGE_ROW_4_Right_4.VNB 0.010692f
C1453 VDD.n395 PHY_EDGE_ROW_4_Right_4.VNB 0.397065f
C1454 VDD.n396 PHY_EDGE_ROW_4_Right_4.VNB 0.010919f
C1455 VDD.n397 PHY_EDGE_ROW_4_Right_4.VNB 0.034024f
C1456 VDD.n398 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1457 VDD.n399 PHY_EDGE_ROW_4_Right_4.VNB 0.008178f
C1458 VDD.n400 PHY_EDGE_ROW_4_Right_4.VNB 0.0134f
C1459 VDD.n401 PHY_EDGE_ROW_4_Right_4.VNB 0.010692f
C1460 VDD.n402 PHY_EDGE_ROW_4_Right_4.VNB 0.391771f
C1461 VDD.n403 PHY_EDGE_ROW_4_Right_4.VNB 0.010557f
C1462 VDD.n404 PHY_EDGE_ROW_4_Right_4.VNB 0.009563f
C1463 VDD.n405 PHY_EDGE_ROW_4_Right_4.VNB 0.006121f
C1464 VDD.n406 PHY_EDGE_ROW_4_Right_4.VNB 0.007445f
C1465 VSS.n0 PHY_EDGE_ROW_4_Right_4.VNB 0.013717f
C1466 VSS.n1 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1467 VSS.n2 PHY_EDGE_ROW_4_Right_4.VNB 0.00734f
C1468 VSS.t64 PHY_EDGE_ROW_4_Right_4.VNB 0.002751f
C1469 VSS.t9 PHY_EDGE_ROW_4_Right_4.VNB 0.003895f
C1470 VSS.n3 PHY_EDGE_ROW_4_Right_4.VNB 0.014283f
C1471 VSS.t94 PHY_EDGE_ROW_4_Right_4.VNB 0.057386f
C1472 VSS.t51 PHY_EDGE_ROW_4_Right_4.VNB 0.010155f
C1473 VSS.t34 PHY_EDGE_ROW_4_Right_4.VNB 0.010155f
C1474 VSS.n4 PHY_EDGE_ROW_4_Right_4.VNB 0.01199f
C1475 VSS.n5 PHY_EDGE_ROW_4_Right_4.VNB 0.032479f
C1476 VSS.n6 PHY_EDGE_ROW_4_Right_4.VNB 0.017898f
C1477 VSS.t67 PHY_EDGE_ROW_4_Right_4.VNB 0.013216f
C1478 VSS.n7 PHY_EDGE_ROW_4_Right_4.VNB 0.048771f
C1479 VSS.t43 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1480 VSS.t52 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1481 VSS.n8 PHY_EDGE_ROW_4_Right_4.VNB 0.008008f
C1482 VSS.n9 PHY_EDGE_ROW_4_Right_4.VNB 0.045105f
C1483 VSS.n10 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1484 VSS.n11 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1485 VSS.n12 PHY_EDGE_ROW_4_Right_4.VNB 1.73714f
C1486 VSS.n13 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1487 VSS.n14 PHY_EDGE_ROW_4_Right_4.VNB 0.436375f
C1488 VSS.n15 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1489 VSS.n16 PHY_EDGE_ROW_4_Right_4.VNB 0.011087f
C1490 VSS.n17 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1491 VSS.n18 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1492 VSS.n19 PHY_EDGE_ROW_4_Right_4.VNB 0.002166f
C1493 VSS.n20 PHY_EDGE_ROW_4_Right_4.VNB 0.004943f
C1494 VSS.t42 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1495 VSS.t61 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1496 VSS.n21 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1497 VSS.n22 PHY_EDGE_ROW_4_Right_4.VNB 0.019854f
C1498 VSS.n23 PHY_EDGE_ROW_4_Right_4.VNB 0.007585f
C1499 VSS.t3 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1500 VSS.t82 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1501 VSS.n24 PHY_EDGE_ROW_4_Right_4.VNB 0.008008f
C1502 VSS.n25 PHY_EDGE_ROW_4_Right_4.VNB 0.009648f
C1503 VSS.t96 PHY_EDGE_ROW_4_Right_4.VNB 0.057386f
C1504 VSS.t17 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1505 VSS.n26 PHY_EDGE_ROW_4_Right_4.VNB 0.022675f
C1506 VSS.n27 PHY_EDGE_ROW_4_Right_4.VNB 0.009041f
C1507 VSS.t37 PHY_EDGE_ROW_4_Right_4.VNB 0.005369f
C1508 VSS.t0 PHY_EDGE_ROW_4_Right_4.VNB -0.001821f
C1509 VSS.n28 PHY_EDGE_ROW_4_Right_4.VNB 0.019464f
C1510 VSS.n29 PHY_EDGE_ROW_4_Right_4.VNB 0.01486f
C1511 VSS.n30 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1512 VSS.n31 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1513 VSS.n32 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1514 VSS.n33 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1515 VSS.n34 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1516 VSS.n35 PHY_EDGE_ROW_4_Right_4.VNB 0.011087f
C1517 VSS.n36 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1518 VSS.n37 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1519 VSS.n38 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1520 VSS.n39 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1521 VSS.n40 PHY_EDGE_ROW_4_Right_4.VNB 0.011087f
C1522 VSS.t33 PHY_EDGE_ROW_4_Right_4.VNB 0.003369f
C1523 VSS.t50 PHY_EDGE_ROW_4_Right_4.VNB 0.006656f
C1524 VSS.n41 PHY_EDGE_ROW_4_Right_4.VNB 0.009918f
C1525 VSS.t81 PHY_EDGE_ROW_4_Right_4.VNB 0.006656f
C1526 VSS.t10 PHY_EDGE_ROW_4_Right_4.VNB 0.003369f
C1527 VSS.n42 PHY_EDGE_ROW_4_Right_4.VNB 0.009918f
C1528 VSS.t41 PHY_EDGE_ROW_4_Right_4.VNB 0.003369f
C1529 VSS.t14 PHY_EDGE_ROW_4_Right_4.VNB 0.006656f
C1530 VSS.n43 PHY_EDGE_ROW_4_Right_4.VNB 0.009918f
C1531 VSS.n44 PHY_EDGE_ROW_4_Right_4.VNB 0.018699f
C1532 VSS.t97 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1533 VSS.t23 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1534 VSS.t24 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1535 VSS.n45 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1536 VSS.t21 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1537 VSS.t99 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1538 VSS.t22 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1539 VSS.n46 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1540 VSS.n47 PHY_EDGE_ROW_4_Right_4.VNB 0.060111f
C1541 VSS.n48 PHY_EDGE_ROW_4_Right_4.VNB 0.02108f
C1542 VSS.n49 PHY_EDGE_ROW_4_Right_4.VNB 0.026019f
C1543 VSS.n50 PHY_EDGE_ROW_4_Right_4.VNB 0.006605f
C1544 VSS.t87 PHY_EDGE_ROW_4_Right_4.VNB 0.006656f
C1545 VSS.t77 PHY_EDGE_ROW_4_Right_4.VNB 0.003369f
C1546 VSS.n51 PHY_EDGE_ROW_4_Right_4.VNB 0.009918f
C1547 VSS.n52 PHY_EDGE_ROW_4_Right_4.VNB 0.01661f
C1548 VSS.n53 PHY_EDGE_ROW_4_Right_4.VNB 0.004091f
C1549 VSS.n54 PHY_EDGE_ROW_4_Right_4.VNB 0.020696f
C1550 VSS.n55 PHY_EDGE_ROW_4_Right_4.VNB 0.015642f
C1551 VSS.n56 PHY_EDGE_ROW_4_Right_4.VNB 0.006179f
C1552 VSS.n57 PHY_EDGE_ROW_4_Right_4.VNB 0.007841f
C1553 VSS.n58 PHY_EDGE_ROW_4_Right_4.VNB 0.004389f
C1554 VSS.n59 PHY_EDGE_ROW_4_Right_4.VNB 0.018443f
C1555 VSS.n60 PHY_EDGE_ROW_4_Right_4.VNB 0.0184f
C1556 VSS.n61 PHY_EDGE_ROW_4_Right_4.VNB 0.006222f
C1557 VSS.t78 PHY_EDGE_ROW_4_Right_4.VNB 0.003369f
C1558 VSS.t39 PHY_EDGE_ROW_4_Right_4.VNB 0.006656f
C1559 VSS.n62 PHY_EDGE_ROW_4_Right_4.VNB 0.009918f
C1560 VSS.t27 PHY_EDGE_ROW_4_Right_4.VNB 0.006656f
C1561 VSS.t57 PHY_EDGE_ROW_4_Right_4.VNB 0.003369f
C1562 VSS.n63 PHY_EDGE_ROW_4_Right_4.VNB 0.009918f
C1563 VSS.n64 PHY_EDGE_ROW_4_Right_4.VNB 0.018741f
C1564 VSS.n65 PHY_EDGE_ROW_4_Right_4.VNB 0.016568f
C1565 VSS.n66 PHY_EDGE_ROW_4_Right_4.VNB 0.004048f
C1566 VSS.n67 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1567 VSS.n68 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1568 VSS.n69 PHY_EDGE_ROW_4_Right_4.VNB 0.019974f
C1569 VSS.n70 PHY_EDGE_ROW_4_Right_4.VNB 0.007841f
C1570 VSS.n71 PHY_EDGE_ROW_4_Right_4.VNB 0.004347f
C1571 VSS.n72 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1572 VSS.n73 PHY_EDGE_ROW_4_Right_4.VNB 0.01107f
C1573 VSS.n74 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1574 VSS.n75 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1575 VSS.n76 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1576 VSS.n77 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1577 VSS.n78 PHY_EDGE_ROW_4_Right_4.VNB 0.009867f
C1578 VSS.n79 PHY_EDGE_ROW_4_Right_4.VNB 0.008904f
C1579 VSS.n80 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1580 VSS.n81 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1581 VSS.n82 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1582 VSS.n83 PHY_EDGE_ROW_4_Right_4.VNB 1.17543f
C1583 VSS.n85 PHY_EDGE_ROW_4_Right_4.VNB 0.012905f
C1584 VSS.n86 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1585 VSS.n87 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1586 VSS.n88 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1587 VSS.t83 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1588 VSS.t56 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1589 VSS.n89 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1590 VSS.n90 PHY_EDGE_ROW_4_Right_4.VNB 0.022556f
C1591 VSS.n91 PHY_EDGE_ROW_4_Right_4.VNB 0.008904f
C1592 VSS.t2 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1593 VSS.t63 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1594 VSS.n92 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1595 VSS.n93 PHY_EDGE_ROW_4_Right_4.VNB 0.022556f
C1596 VSS.n94 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1597 VSS.t90 PHY_EDGE_ROW_4_Right_4.VNB 0.057386f
C1598 VSS.n95 PHY_EDGE_ROW_4_Right_4.VNB 0.054365f
C1599 VSS.t75 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1600 VSS.n96 PHY_EDGE_ROW_4_Right_4.VNB 0.019533f
C1601 VSS.n97 PHY_EDGE_ROW_4_Right_4.VNB 0.020094f
C1602 VSS.n98 PHY_EDGE_ROW_4_Right_4.VNB 0.035746f
C1603 VSS.t76 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1604 VSS.n99 PHY_EDGE_ROW_4_Right_4.VNB 0.022675f
C1605 VSS.n100 PHY_EDGE_ROW_4_Right_4.VNB 0.01671f
C1606 VSS.n101 PHY_EDGE_ROW_4_Right_4.VNB 0.005934f
C1607 VSS.n102 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1608 VSS.n103 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1609 VSS.n104 PHY_EDGE_ROW_4_Right_4.VNB 0.012875f
C1610 VSS.n105 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1611 VSS.n106 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1612 VSS.n107 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1613 VSS.n108 PHY_EDGE_ROW_4_Right_4.VNB 0.009282f
C1614 VSS.n109 PHY_EDGE_ROW_4_Right_4.VNB 0.011484f
C1615 VSS.n110 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1616 VSS.n111 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1617 VSS.n112 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1618 VSS.n113 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1619 VSS.n114 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1620 VSS.n115 PHY_EDGE_ROW_4_Right_4.VNB 0.009867f
C1621 VSS.n116 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1622 VSS.n117 PHY_EDGE_ROW_4_Right_4.VNB 0.01107f
C1623 VSS.n118 PHY_EDGE_ROW_4_Right_4.VNB 0.00734f
C1624 VSS.n119 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1625 VSS.t54 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1626 VSS.t4 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1627 VSS.n120 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1628 VSS.n121 PHY_EDGE_ROW_4_Right_4.VNB 0.007841f
C1629 VSS.n122 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1630 VSS.t31 PHY_EDGE_ROW_4_Right_4.VNB 0.016422f
C1631 VSS.t84 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1632 VSS.t48 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1633 VSS.n123 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1634 VSS.n124 PHY_EDGE_ROW_4_Right_4.VNB 0.022556f
C1635 VSS.t59 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1636 VSS.t15 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1637 VSS.n125 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1638 VSS.n126 PHY_EDGE_ROW_4_Right_4.VNB 0.022556f
C1639 VSS.n127 PHY_EDGE_ROW_4_Right_4.VNB 0.004693f
C1640 VSS.n128 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1641 VSS.n129 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1642 VSS.n130 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1643 VSS.n131 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1644 VSS.n132 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1645 VSS.n133 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1646 VSS.n134 PHY_EDGE_ROW_4_Right_4.VNB 0.007841f
C1647 VSS.n135 PHY_EDGE_ROW_4_Right_4.VNB 0.009024f
C1648 VSS.n136 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1649 VSS.n137 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1650 VSS.n138 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1651 VSS.n139 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1652 VSS.n140 PHY_EDGE_ROW_4_Right_4.VNB 0.009385f
C1653 VSS.n141 PHY_EDGE_ROW_4_Right_4.VNB 0.009385f
C1654 VSS.n142 PHY_EDGE_ROW_4_Right_4.VNB 0.004813f
C1655 VSS.n143 PHY_EDGE_ROW_4_Right_4.VNB 0.007841f
C1656 VSS.t53 PHY_EDGE_ROW_4_Right_4.VNB 0.005028f
C1657 VSS.t8 PHY_EDGE_ROW_4_Right_4.VNB 0.004106f
C1658 VSS.n144 PHY_EDGE_ROW_4_Right_4.VNB 0.011966f
C1659 VSS.n145 PHY_EDGE_ROW_4_Right_4.VNB 0.005625f
C1660 VSS.t35 PHY_EDGE_ROW_4_Right_4.VNB 0.010532f
C1661 VSS.n146 PHY_EDGE_ROW_4_Right_4.VNB 0.018657f
C1662 VSS.t44 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1663 VSS.n147 PHY_EDGE_ROW_4_Right_4.VNB 0.022675f
C1664 VSS.n148 PHY_EDGE_ROW_4_Right_4.VNB 0.013687f
C1665 VSS.t91 PHY_EDGE_ROW_4_Right_4.VNB 0.057386f
C1666 VSS.t45 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1667 VSS.n149 PHY_EDGE_ROW_4_Right_4.VNB 0.019501f
C1668 VSS.n150 PHY_EDGE_ROW_4_Right_4.VNB 0.054365f
C1669 VSS.n151 PHY_EDGE_ROW_4_Right_4.VNB 0.035746f
C1670 VSS.n152 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1671 VSS.n153 PHY_EDGE_ROW_4_Right_4.VNB 0.020094f
C1672 VSS.n154 PHY_EDGE_ROW_4_Right_4.VNB 0.01671f
C1673 VSS.n155 PHY_EDGE_ROW_4_Right_4.VNB 0.00359f
C1674 VSS.n156 PHY_EDGE_ROW_4_Right_4.VNB 0.013115f
C1675 VSS.n157 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1676 VSS.n158 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1677 VSS.n159 PHY_EDGE_ROW_4_Right_4.VNB 0.004176f
C1678 VSS.n160 PHY_EDGE_ROW_4_Right_4.VNB 0.015752f
C1679 VSS.n161 PHY_EDGE_ROW_4_Right_4.VNB 0.005753f
C1680 VSS.n162 PHY_EDGE_ROW_4_Right_4.VNB 0.007841f
C1681 VSS.n163 PHY_EDGE_ROW_4_Right_4.VNB 0.016123f
C1682 VSS.n164 PHY_EDGE_ROW_4_Right_4.VNB 0.007958f
C1683 VSS.n165 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1684 VSS.n166 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1685 VSS.n167 PHY_EDGE_ROW_4_Right_4.VNB 0.364181f
C1686 VSS.n168 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1687 VSS.n169 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1688 VSS.n170 PHY_EDGE_ROW_4_Right_4.VNB 0.011087f
C1689 VSS.n171 PHY_EDGE_ROW_4_Right_4.VNB 0.019492f
C1690 VSS.n172 PHY_EDGE_ROW_4_Right_4.VNB 0.020335f
C1691 VSS.n173 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1692 VSS.n174 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1693 VSS.n175 PHY_EDGE_ROW_4_Right_4.VNB 0.012875f
C1694 VSS.n176 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1695 VSS.n177 PHY_EDGE_ROW_4_Right_4.VNB 0.019974f
C1696 VSS.n178 PHY_EDGE_ROW_4_Right_4.VNB 0.005199f
C1697 VSS.n179 PHY_EDGE_ROW_4_Right_4.VNB 0.035874f
C1698 VSS.n180 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1699 VSS.n181 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1700 VSS.n182 PHY_EDGE_ROW_4_Right_4.VNB 0.020094f
C1701 VSS.n183 PHY_EDGE_ROW_4_Right_4.VNB 0.013115f
C1702 VSS.n184 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1703 VSS.n185 PHY_EDGE_ROW_4_Right_4.VNB 0.022556f
C1704 VSS.n186 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1705 VSS.n187 PHY_EDGE_ROW_4_Right_4.VNB 0.019974f
C1706 VSS.n188 PHY_EDGE_ROW_4_Right_4.VNB 0.009282f
C1707 VSS.n189 PHY_EDGE_ROW_4_Right_4.VNB 0.011484f
C1708 VSS.n190 PHY_EDGE_ROW_4_Right_4.VNB 0.012905f
C1709 VSS.n191 PHY_EDGE_ROW_4_Right_4.VNB 0.364181f
C1710 VSS.n192 PHY_EDGE_ROW_4_Right_4.VNB 1.73554f
C1711 VSS.n193 PHY_EDGE_ROW_4_Right_4.VNB 0.701419f
C1712 VSS.n194 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1713 VSS.n195 PHY_EDGE_ROW_4_Right_4.VNB 0.009041f
C1714 VSS.n196 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1715 VSS.t79 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1716 VSS.t49 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1717 VSS.n197 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1718 VSS.n198 PHY_EDGE_ROW_4_Right_4.VNB 0.022556f
C1719 VSS.n199 PHY_EDGE_ROW_4_Right_4.VNB 0.02108f
C1720 VSS.t92 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1721 VSS.t46 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1722 VSS.t47 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1723 VSS.n200 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1724 VSS.t71 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1725 VSS.t93 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1726 VSS.t72 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1727 VSS.n201 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1728 VSS.n202 PHY_EDGE_ROW_4_Right_4.VNB 0.060111f
C1729 VSS.n203 PHY_EDGE_ROW_4_Right_4.VNB 0.005199f
C1730 VSS.n204 PHY_EDGE_ROW_4_Right_4.VNB 0.026861f
C1731 VSS.n205 PHY_EDGE_ROW_4_Right_4.VNB 0.011912f
C1732 VSS.n206 PHY_EDGE_ROW_4_Right_4.VNB 0.009987f
C1733 VSS.n207 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1734 VSS.t85 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1735 VSS.t16 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1736 VSS.n208 PHY_EDGE_ROW_4_Right_4.VNB 0.008008f
C1737 VSS.n209 PHY_EDGE_ROW_4_Right_4.VNB 0.017836f
C1738 VSS.n210 PHY_EDGE_ROW_4_Right_4.VNB 0.007841f
C1739 VSS.n211 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1740 VSS.n212 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1741 VSS.n213 PHY_EDGE_ROW_4_Right_4.VNB 0.009867f
C1742 VSS.n214 PHY_EDGE_ROW_4_Right_4.VNB 0.008904f
C1743 VSS.n215 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1744 VSS.n216 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1745 VSS.n217 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1746 VSS.n218 PHY_EDGE_ROW_4_Right_4.VNB 0.527822f
C1747 VSS.n219 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1748 VSS.n220 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1749 VSS.n221 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1750 VSS.n222 PHY_EDGE_ROW_4_Right_4.VNB 0.01107f
C1751 VSS.n223 PHY_EDGE_ROW_4_Right_4.VNB 0.00758f
C1752 VSS.n224 PHY_EDGE_ROW_4_Right_4.VNB 0.00555f
C1753 VSS.n225 PHY_EDGE_ROW_4_Right_4.VNB 0.01671f
C1754 VSS.n226 PHY_EDGE_ROW_4_Right_4.VNB 0.019974f
C1755 VSS.n227 PHY_EDGE_ROW_4_Right_4.VNB 0.013115f
C1756 VSS.n228 PHY_EDGE_ROW_4_Right_4.VNB 0.035746f
C1757 VSS.n229 PHY_EDGE_ROW_4_Right_4.VNB 0.054365f
C1758 VSS.t18 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1759 VSS.n230 PHY_EDGE_ROW_4_Right_4.VNB 0.006301f
C1760 VSS.t86 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1761 VSS.t28 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1762 VSS.n231 PHY_EDGE_ROW_4_Right_4.VNB 0.007658f
C1763 VSS.n232 PHY_EDGE_ROW_4_Right_4.VNB 0.009418f
C1764 VSS.n233 PHY_EDGE_ROW_4_Right_4.VNB 0.004337f
C1765 VSS.n234 PHY_EDGE_ROW_4_Right_4.VNB 0.007149f
C1766 VSS.n235 PHY_EDGE_ROW_4_Right_4.VNB 0.01107f
C1767 VSS.n236 PHY_EDGE_ROW_4_Right_4.VNB 0.011311f
C1768 VSS.n237 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1769 VSS.t6 PHY_EDGE_ROW_4_Right_4.VNB 0.010265f
C1770 VSS.n238 PHY_EDGE_ROW_4_Right_4.VNB 0.021569f
C1771 VSS.n239 PHY_EDGE_ROW_4_Right_4.VNB 0.016302f
C1772 VSS.n240 PHY_EDGE_ROW_4_Right_4.VNB 0.010829f
C1773 VSS.n241 PHY_EDGE_ROW_4_Right_4.VNB 0.020094f
C1774 VSS.n242 PHY_EDGE_ROW_4_Right_4.VNB 0.013356f
C1775 VSS.n243 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1776 VSS.t1 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1777 VSS.t13 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1778 VSS.n244 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1779 VSS.n245 PHY_EDGE_ROW_4_Right_4.VNB 0.020681f
C1780 VSS.t32 PHY_EDGE_ROW_4_Right_4.VNB 0.004317f
C1781 VSS.t80 PHY_EDGE_ROW_4_Right_4.VNB 0.004649f
C1782 VSS.n246 PHY_EDGE_ROW_4_Right_4.VNB 0.012389f
C1783 VSS.n247 PHY_EDGE_ROW_4_Right_4.VNB 0.028367f
C1784 VSS.n248 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1785 VSS.n249 PHY_EDGE_ROW_4_Right_4.VNB 0.013356f
C1786 VSS.n250 PHY_EDGE_ROW_4_Right_4.VNB 0.017206f
C1787 VSS.n251 PHY_EDGE_ROW_4_Right_4.VNB 0.02132f
C1788 VSS.t38 PHY_EDGE_ROW_4_Right_4.VNB 0.002751f
C1789 VSS.t30 PHY_EDGE_ROW_4_Right_4.VNB 0.003895f
C1790 VSS.n252 PHY_EDGE_ROW_4_Right_4.VNB 0.014519f
C1791 VSS.n253 PHY_EDGE_ROW_4_Right_4.VNB 0.023112f
C1792 VSS.t29 PHY_EDGE_ROW_4_Right_4.VNB 0.0165f
C1793 VSS.t40 PHY_EDGE_ROW_4_Right_4.VNB 0.010377f
C1794 VSS.t7 PHY_EDGE_ROW_4_Right_4.VNB 0.010436f
C1795 VSS.n254 PHY_EDGE_ROW_4_Right_4.VNB 0.011558f
C1796 VSS.n255 PHY_EDGE_ROW_4_Right_4.VNB 0.038509f
C1797 VSS.n256 PHY_EDGE_ROW_4_Right_4.VNB 0.008904f
C1798 VSS.n257 PHY_EDGE_ROW_4_Right_4.VNB 0.012995f
C1799 VSS.t5 PHY_EDGE_ROW_4_Right_4.VNB 0.015862f
C1800 VSS.t62 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1801 VSS.t55 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1802 VSS.n258 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1803 VSS.n259 PHY_EDGE_ROW_4_Right_4.VNB 0.020214f
C1804 VSS.n260 PHY_EDGE_ROW_4_Right_4.VNB 0.013115f
C1805 VSS.t12 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1806 VSS.t58 PHY_EDGE_ROW_4_Right_4.VNB 0.00378f
C1807 VSS.n261 PHY_EDGE_ROW_4_Right_4.VNB 0.008232f
C1808 VSS.t98 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1809 VSS.t19 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1810 VSS.t20 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1811 VSS.n262 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1812 VSS.t25 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1813 VSS.t100 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1814 VSS.t26 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1815 VSS.n263 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1816 VSS.n264 PHY_EDGE_ROW_4_Right_4.VNB 0.060079f
C1817 VSS.n265 PHY_EDGE_ROW_4_Right_4.VNB 0.021946f
C1818 VSS.n266 PHY_EDGE_ROW_4_Right_4.VNB 0.010829f
C1819 VSS.n267 PHY_EDGE_ROW_4_Right_4.VNB 0.005199f
C1820 VSS.n268 PHY_EDGE_ROW_4_Right_4.VNB 0.02115f
C1821 VSS.n269 PHY_EDGE_ROW_4_Right_4.VNB 0.02115f
C1822 VSS.n270 PHY_EDGE_ROW_4_Right_4.VNB 0.006435f
C1823 VSS.n271 PHY_EDGE_ROW_4_Right_4.VNB 0.029192f
C1824 VSS.n272 PHY_EDGE_ROW_4_Right_4.VNB 0.016123f
C1825 VSS.n273 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1826 VSS.n274 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1827 VSS.n275 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1828 VSS.n276 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1829 VSS.n277 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1830 VSS.n278 PHY_EDGE_ROW_4_Right_4.VNB 0.011087f
C1831 VSS.n279 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1832 VSS.n280 PHY_EDGE_ROW_4_Right_4.VNB 0.004602f
C1833 VSS.n281 PHY_EDGE_ROW_4_Right_4.VNB 0.027822f
C1834 VSS.n282 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1835 VSS.n283 PHY_EDGE_ROW_4_Right_4.VNB 0.01107f
C1836 VSS.n284 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1837 VSS.n285 PHY_EDGE_ROW_4_Right_4.VNB 0.011592f
C1838 VSS.n286 PHY_EDGE_ROW_4_Right_4.VNB 0.012797f
C1839 VSS.n287 PHY_EDGE_ROW_4_Right_4.VNB 0.527822f
C1840 VSS.n288 PHY_EDGE_ROW_4_Right_4.VNB 0.910524f
C1841 VSS.n290 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1842 VSS.n291 PHY_EDGE_ROW_4_Right_4.VNB 0.01107f
C1843 VSS.n292 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1844 VSS.n293 PHY_EDGE_ROW_4_Right_4.VNB 0.007701f
C1845 VSS.n294 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1846 VSS.n295 PHY_EDGE_ROW_4_Right_4.VNB 0.032979f
C1847 VSS.n296 PHY_EDGE_ROW_4_Right_4.VNB 0.032979f
C1848 VSS.t60 PHY_EDGE_ROW_4_Right_4.VNB 0.004649f
C1849 VSS.t11 PHY_EDGE_ROW_4_Right_4.VNB 0.004317f
C1850 VSS.n297 PHY_EDGE_ROW_4_Right_4.VNB 0.012106f
C1851 VSS.t95 PHY_EDGE_ROW_4_Right_4.VNB 0.424091f
C1852 VSS.n298 PHY_EDGE_ROW_4_Right_4.VNB 0.031903f
C1853 VSS.t36 PHY_EDGE_ROW_4_Right_4.VNB 0.010265f
C1854 VSS.t68 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1855 VSS.n299 PHY_EDGE_ROW_4_Right_4.VNB 0.01705f
C1856 VSS.n300 PHY_EDGE_ROW_4_Right_4.VNB 0.018721f
C1857 VSS.t88 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1858 VSS.t73 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1859 VSS.t74 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1860 VSS.n301 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1861 VSS.t69 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1862 VSS.t89 PHY_EDGE_ROW_4_Right_4.VNB 0.058172f
C1863 VSS.t70 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1864 VSS.n302 PHY_EDGE_ROW_4_Right_4.VNB 0.108548f
C1865 VSS.n303 PHY_EDGE_ROW_4_Right_4.VNB 0.022993f
C1866 VSS.n304 PHY_EDGE_ROW_4_Right_4.VNB 0.059964f
C1867 VSS.n305 PHY_EDGE_ROW_4_Right_4.VNB 0.011616f
C1868 VSS.n306 PHY_EDGE_ROW_4_Right_4.VNB 0.013115f
C1869 VSS.n307 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1870 VSS.n308 PHY_EDGE_ROW_4_Right_4.VNB 0.02214f
C1871 VSS.n309 PHY_EDGE_ROW_4_Right_4.VNB 0.032979f
C1872 VSS.n310 PHY_EDGE_ROW_4_Right_4.VNB 0.024734f
C1873 VSS.n311 PHY_EDGE_ROW_4_Right_4.VNB 0.113638f
C1874 VSS.n312 PHY_EDGE_ROW_4_Right_4.VNB 0.027088f
C1875 VSS.n313 PHY_EDGE_ROW_4_Right_4.VNB 0.017384f
C1876 VSS.n314 PHY_EDGE_ROW_4_Right_4.VNB 0.016123f
C1877 VSS.n315 PHY_EDGE_ROW_4_Right_4.VNB 0.011087f
C1878 VSS.n316 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1879 VSS.n317 PHY_EDGE_ROW_4_Right_4.VNB 0.012905f
C1880 VSS.n318 PHY_EDGE_ROW_4_Right_4.VNB 0.011484f
C1881 VSS.n319 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1882 VSS.n320 PHY_EDGE_ROW_4_Right_4.VNB 0.009385f
C1883 VSS.n321 PHY_EDGE_ROW_4_Right_4.VNB 0.009385f
C1884 VSS.n322 PHY_EDGE_ROW_4_Right_4.VNB 0.00742f
C1885 VSS.n323 PHY_EDGE_ROW_4_Right_4.VNB 0.005936f
C1886 VSS.n324 PHY_EDGE_ROW_4_Right_4.VNB 0.013236f
C1887 VSS.n325 PHY_EDGE_ROW_4_Right_4.VNB 0.012905f
C1888 VSS.n326 PHY_EDGE_ROW_4_Right_4.VNB 0.011484f
C1889 VSS.n327 PHY_EDGE_ROW_4_Right_4.VNB 0.009041f
C1890 VSS.n328 PHY_EDGE_ROW_4_Right_4.VNB 0.01119f
C1891 VSS.n329 PHY_EDGE_ROW_4_Right_4.VNB 0.032979f
C1892 VSS.n330 PHY_EDGE_ROW_4_Right_4.VNB 0.029394f
C1893 VSS.n331 PHY_EDGE_ROW_4_Right_4.VNB 0.020384f
C1894 VSS.n332 PHY_EDGE_ROW_4_Right_4.VNB 0.027196f
C1895 VSS.n333 PHY_EDGE_ROW_4_Right_4.VNB 0.017468f
C1896 VSS.t66 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1897 VSS.n334 PHY_EDGE_ROW_4_Right_4.VNB 0.006762f
C1898 VSS.n335 PHY_EDGE_ROW_4_Right_4.VNB 0.05229f
C1899 VSS.n336 PHY_EDGE_ROW_4_Right_4.VNB 0.030653f
C1900 VSS.n337 PHY_EDGE_ROW_4_Right_4.VNB 0.021909f
C1901 VSS.t65 PHY_EDGE_ROW_4_Right_4.VNB 0.012881f
C1902 VSS.n338 PHY_EDGE_ROW_4_Right_4.VNB 0.022675f
C1903 VSS.n339 PHY_EDGE_ROW_4_Right_4.VNB 0.01671f
C1904 VSS.n340 PHY_EDGE_ROW_4_Right_4.VNB 0.019492f
.ends

