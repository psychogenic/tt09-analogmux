** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tb_anamux.sch
**.subckt tb_anamux
x1 net1 net2 net3 net4 VCC net5 net6 net7 VSS net8 net9 net10 net11 net12 net13 net14 net15 net16 net17 net18 net19 net20 net21
+ net22 net23 net24 net25 net26 net27 RSEL0 net28 net29 RSEL1 net30 RSEL2 net31 SEL0 net32 SEL1 net33 EN_COUNTER net34 EN_RING net35
+ net36 net37 net38 net39 VRES RINGOUT MUXOUT LADOUT tt_um_patdeegan_anamux_parax
R6 RINGOUT VSS 100k m=1
R1 MUXOUT VSS 100k m=1
R2 LADOUT VSS 100k m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sym # of pins=52
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sch
.subckt tt_um_patdeegan_anamux uo_out[0] uo_out[1] uo_out[2] uio_oe[0] VSS uo_out[3] uio_oe[1] uio_oe[2] VDD uo_out[4] uio_oe[3]
+ ena uo_out[5] uio_oe[4] clk uo_out[6] uio_oe[5] rst_n uo_out[7] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] ui_in[0] uio_out[6] uio_in[0] ui_in[1] uio_out[7] uio_in[1] ui_in[2] uio_in[2] ui_in[3] uio_in[3] ui_in[4] uio_in[4]
+ ui_in[5] uio_in[5] ui_in[6] uio_in[6] ui_in[7] uio_in[7] ua[4] ua[5] ua[6] ua[0] ua[1] ua[2] ua[3]
*.ipin ena
*.ipin clk
*.ipin rst_n
*.iopin ua[4]
*.iopin ua[5]
*.iopin ua[6]
*.ipin ui_in[7]
*.ipin uio_in[0]
*.ipin uio_in[1]
*.ipin uio_in[2]
*.ipin uio_in[3]
*.ipin uio_in[4]
*.ipin uio_in[5]
*.ipin uio_in[6]
*.ipin uio_in[7]
*.opin uio_oe[0]
*.opin uio_oe[1]
*.opin uio_oe[2]
*.opin uio_oe[3]
*.opin uio_oe[4]
*.opin uio_oe[5]
*.opin uio_oe[6]
*.opin uio_oe[7]
*.iopin uio_out[0]
*.iopin uio_out[1]
*.iopin uio_out[2]
*.iopin uio_out[3]
*.iopin uio_out[4]
*.iopin uio_out[5]
*.iopin uio_out[6]
*.iopin uio_out[7]
*.opin uo_out[0]
*.opin uo_out[1]
*.opin uo_out[2]
*.opin uo_out[3]
*.opin uo_out[4]
*.opin uo_out[5]
*.opin uo_out[6]
*.opin uo_out[7]
*.ipin ui_in[0]
*.ipin ui_in[1]
*.ipin ui_in[2]
*.ipin ui_in[3]
*.ipin ui_in[4]
*.ipin ui_in[5]
*.ipin ui_in[6]
*.iopin ua[0]
*.iopin ua[1]
*.iopin ua[2]
*.iopin ua[3]
*.ipin VSS
*.ipin VDD
x1 ua[0] ui_in[3] VDD ui_in[4] ua[1] VSS ui_in[0] ui_in[1] ua[2] ui_in[2] ua[3] ui_in[6] ui_in[5] fulltest_userarea
.ends


* expanding   symbol:  tt_um_patdeegan_anamux_parax.sym # of pins=52
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tt_um_patdeegan_anamux.sym
.include /home/ttuser/vmswap/tt09-analogmux/xschem/extracted/tt_um_patdeegan_anamux_parax.spice

* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sym # of pins=13
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/fulltest_userarea.sch
.subckt fulltest_userarea VRES select0 VDD select1 ring_out VSS rsel0 rsel1 muxtest_out rsel2 ladderout enable_ring
+ enable_counter
*.ipin VDD
*.ipin VSS
*.ipin select0
*.ipin select1
*.ipin rsel0
*.ipin rsel1
*.ipin rsel2
*.ipin enable_ring
*.ipin enable_counter
*.opin ring_out
*.opin muxtest_out
*.opin ladderout
*.ipin VRES
x1 VDD VSS VRES select0 select1 rsel0 rsel1 rsel2 muxtest_out ladderout muxtest
x2 select0 VDD select1 VSS ring_out enable_ring enable_counter ringtest
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sym # of pins=10
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/muxtest.sch
.subckt muxtest VDD VSS VRES SELECT0 SELECT1 RSEL0 RSEL1 RSEL2 OUT LADDEROUT
*.ipin VSS
*.ipin VDD
*.ipin SELECT0
*.ipin SELECT1
*.ipin VRES
*.ipin RSEL0
*.ipin RSEL1
*.ipin RSEL2
*.opin OUT
*.opin LADDEROUT
x1 VDD VSS RSEL0 RSEL1 A1 A5 A6 A2 A7 A3 RSEL2 VRES A4 LADDEROUT mux8onehot
x2 SELECT1 VDD VSS A5 VRES LADDEROUT OUT OUT OUT A1 OUT SELECT0 VDD net1 mux4onehot_b
XR1 A7 VRES VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR2 A6 A7 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR3 A5 A6 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR4 A4 A5 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR5 A3 A4 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR6 A2 A3 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR7 A1 A2 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
XR8 VSS A1 VSS sky130_fd_pr__res_high_po_1p41 L=1.75 mult=1 m=1
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sym # of pins=7
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/ringtest.sch
.subckt ringtest select0 VDD select1 VSS mux_out enable_ring enable_counter
*.ipin VDD
*.ipin VSS
*.ipin enable_ring
*.ipin select0
*.ipin select1
*.ipin enable_counter
*.opin mux_out
x3 select1 VDD VSS counter3 drv_out ring_out mux_out mux_out mux_out counter7 mux_out select0 VDD net1 mux4onehot_b
x4 enable_counter drv_out net2 net3 net4 counter3 net5 net6 net7 counter7 net8 net9 VDD VSS simplecounter
x1 VDD VSS enable_ring ring_out ring
x2 VDD VSS ring_out drv_out driver
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux8onehot.sch
.subckt mux8onehot VDD VSS select0 select1 A1 A5 A6 A2 A7 A3 select2 A8 A4 Z
*.ipin select0
*.ipin select1
*.ipin select2
*.ipin VDD
*.ipin VSS
*.iopin Z
*.iopin A1
*.iopin A2
*.iopin A3
*.iopin A4
*.iopin A5
*.iopin A6
*.iopin A7
*.iopin A8
x4 Z OUT_HIGH nSEL2 select2 VSS VDD passgate
x5 Z OUT_LOW select2 nSEL2 VSS VDD passgate
x2 gpo2 gpo1 gpo0 VDD gpo3 VSS A3 A2 A1 OUT_LOW OUT_LOW OUT_LOW A4 OUT_LOW gno2 gno1 gno0 gno3 passgatex4
x1 gpo0 gno0 gno1 gpo1 select0 select1 gno2 gpo2 nSEL2 select2 gno3 gpo3 VDD VSS passgatesCtrlManual
x3 gpo2 gpo1 gpo0 VDD gpo3 VSS A7 A6 A5 OUT_HIGH OUT_HIGH OUT_HIGH A8 OUT_HIGH gno2 gno1 gno0 gno3 passgatex4
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sch
.subckt mux4onehot_b select1 VDD VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 select0 select2 nselect2
*.ipin select0
*.ipin select1
*.ipin select2
*.iopin A1
*.iopin A2
*.iopin A3
*.iopin A4
*.iopin Z1
*.iopin Z2
*.iopin Z3
*.iopin Z4
*.opin nselect2
*.ipin VDD
*.ipin VSS
x2 gpo2 gpo1 gpo0 VDD gpo3 VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 gno2 gno1 gno0 gno3 passgatex4
x1 gpo0 gno0 gno1 gpo1 select0 select1 gno2 gpo2 nselect2 select2 gno3 gpo3 VDD VSS passgatesCtrlManual
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/ring.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/ring.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/ring.sch
.subckt ring VDD VSS enable out
*.iopin VDD
*.ipin enable
*.iopin VSS
*.opin out
x2 enable net18 VSS VSS VDD VDD out sky130_fd_sc_hd__nand2_2
x1 VDD VSS out net1 inverter
x3 VDD VSS net1 net2 inverter
x4 VDD VSS net2 net3 inverter
x5 VDD VSS net3 net4 inverter
x6 VDD VSS net4 net5 inverter
x7 VDD VSS net5 net6 inverter
x8 VDD VSS net6 net7 inverter
x9 VDD VSS net7 net8 inverter
x10 VDD VSS net8 net9 inverter
x11 VDD VSS net9 net10 inverter
x12 VDD VSS net10 net11 inverter
x13 VDD VSS net11 net12 inverter
x14 VDD VSS net12 net13 inverter
x15 VDD VSS net13 net14 inverter
x16 VDD VSS net14 net15 inverter
x17 VDD VSS net15 net16 inverter
x18 VDD VSS net16 net17 inverter
x19 VDD VSS net17 net18 inverter
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/driver.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/driver.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mattring/driver.sch
.subckt driver VDD VSS in out
*.iopin VDD
*.iopin VSS
*.opin out
*.ipin in
XM9 net1 in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net1 in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=72 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=24 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym # of pins=6
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgate.sch
.subckt passgate Z A GP GN VSSBPIN VCCBPIN
*.ipin GN
*.ipin VCCBPIN
*.ipin VSSBPIN
*.ipin GP
*.iopin A
*.iopin Z
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym # of pins=18
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sch
.subckt passgatex4 GP3 GP2 GP1 VDD GP4 VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 GN3 GN2 GN1 GN4
*.ipin VDD
*.ipin VSS
*.ipin GP1
*.ipin GN1
*.iopin A1
*.iopin Z1
*.ipin GP2
*.ipin GN2
*.iopin A2
*.iopin Z2
*.ipin GP3
*.ipin GN3
*.iopin A3
*.iopin Z3
*.ipin GP4
*.ipin GN4
*.iopin A4
*.iopin Z4
x1 Z1 A1 GP1 GN1 VSS VDD passgate
x2 Z2 A2 GP2 GN2 VSS VDD passgate
x3 Z3 A3 GP3 GN3 VSS VDD passgate
x4 Z4 A4 GP4 GN4 VSS VDD passgate
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sch
.subckt passgatesCtrlManual gpo0 gno0 gno1 gpo1 SEL0 SEL1 gno2 gpo2 nSEL2 SEL2 gno3 gpo3 VDD VSS
*.ipin SEL0
*.ipin SEL1
*.ipin SEL2
*.opin gno0
*.opin gpo0
*.opin gno1
*.opin gpo1
*.opin gno2
*.opin gpo2
*.opin gno3
*.opin gpo3
*.opin nSEL2
*.ipin VDD
*.ipin VSS
x1 SEL0 VSS VSS VDD VDD nSEL0 sky130_fd_sc_hd__inv_2
x2 SEL1 VSS VSS VDD VDD nSEL1 sky130_fd_sc_hd__inv_2
x7 nSEL0 nSEL1 VSS VSS VDD VDD gno0 sky130_fd_sc_hd__and2_1
x10 SEL1 SEL0 VSS VSS VDD VDD gno3 sky130_fd_sc_hd__and2_1
x11 gno0 VSS VSS VDD VDD gpo0 sky130_fd_sc_hd__inv_2
x12 gno1 VSS VSS VDD VDD gpo1 sky130_fd_sc_hd__inv_2
x13 gno2 VSS VSS VDD VDD gpo2 sky130_fd_sc_hd__inv_2
x14 gno3 VSS VSS VDD VDD gpo3 sky130_fd_sc_hd__inv_2
x15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x16 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x17 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x8 SEL1 SEL0 VSS VSS VDD VDD gno1 sky130_fd_sc_hd__and2b_1
x9 SEL0 SEL1 VSS VSS VDD VDD gno2 sky130_fd_sc_hd__and2b_1
x18 SEL2 VSS VSS VDD VDD nSEL2 sky130_fd_sc_hd__inv_2
x19 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/inverter.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/inverter.sch
.subckt inverter VDD VSS in out
*.opin out
*.iopin VDD
*.iopin VSS
*.ipin in
x1 in VSS VSS VDD VDD out sky130_fd_sc_hd__inv_2
.ends

**** begin user architecture code


* ngspice commands
* .options savecurrents
.param VCC = 1.8
.param SRCRES = 1k
.include stimuli_tb_anamux.cir
.control
save all
op
write tb_anamux.raw
set appendwrite
tran 0.3n 260n uic
write tb_anamux.raw
* quit 0
.endc



**** end user architecture code
.end
