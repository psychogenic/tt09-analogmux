** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/tb_passgatex4.sch
**.subckt tb_passgatex4
x1 nEN3 nEN2 nEN1 VCC nEN4 VSS IN3 IN2 IN1 OUT OUT OUT IN4 OUT EN3 EN2 EN1 EN4 passgatex4
x2 nEN1 EN1 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
V2 net1 VSS sin(0.9 0.9 250k)
x3 nEN2 EN2 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x4 nEN3 EN3 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
x5 nEN4 EN4 VCC VSS not W_N=1 L_N=0.15 W_P=2 L_P=0.15 m=1
V3 net2 VSS sin(0.9 0.9 8Meg)
V5 net3 VSS sin(0.9 0.9 500k)
V6 net4 VSS sin(0.9 0.9 1Meg)
R1 OUT VSS 10k m=1
R2 IN1 net1 1 m=1
R3 IN2 net3 1 m=1
R4 IN3 net4 1 m=1
R5 IN4 net2 1 m=1
x6 nEN3 nEN2 nEN1 VCC nEN4 VSS IN3 IN2 IN1 OUTPX OUTPX OUTPX IN4 OUTPX EN3 EN2 EN1 EN4 passgatex4_parax
R6 OUTPX VSS 10k m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  /home/ttuser/work/tt09-analogmux/xschem/passgatex4.sym # of pins=18
** sym_path: /home/ttuser/work/tt09-analogmux/xschem/passgatex4.sym
** sch_path: /home/ttuser/work/tt09-analogmux/xschem/passgatex4.sch
.subckt passgatex4 GP3 GP2 GP1 VDD GP4 VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 GN3 GN2 GN1 GN4
*.ipin VDD
*.ipin VSS
*.ipin GP1
*.ipin GN1
*.iopin A1
*.iopin Z1
*.ipin GP2
*.ipin GN2
*.iopin A2
*.iopin Z2
*.ipin GP3
*.ipin GN3
*.iopin A3
*.iopin Z3
*.ipin GP4
*.ipin GN4
*.iopin A4
*.iopin Z4
x1 Z1 A1 GP1 GN1 VSS VDD passgate
x2 Z2 A2 GP2 GN2 VSS VDD passgate
x3 Z3 A3 GP3 GN3 VSS VDD passgate
x4 Z4 A4 GP4 GN4 VSS VDD passgate
.ends


* expanding   symbol:  sky130_tests/not.sym # of pins=2
** sym_path: /home/ttuser/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sym
** sch_path: /home/ttuser/pdk/sky130A/libs.tech/xschem/sky130_tests/not.sch
.subckt not y a VCCPIN VSSPIN     W_N=1 L_N=0.15 W_P=2 L_P=0.15
*.opin y
*.ipin a
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8 L=L_N W=W_N nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8 L=L_P W=W_P nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  passgatex4_parax.sym # of pins=18
** sym_path: /home/ttuser/work/tt09-analogmux/xschem/passgatex4.sym
.include /home/ttuser/vmswap/tt09-analogmux/xschem/extracted/passgatex4_parax.spice

* expanding   symbol:  /home/ttuser/tt08-wowa2/xschem/passgate.sym # of pins=6
** sym_path: /home/ttuser/tt08-wowa2/xschem/passgate.sym
** sch_path: /home/ttuser/tt08-wowa2/xschem/passgate.sch
.subckt passgate Z A GP GN VSSBPIN VCCBPIN
*.ipin GN
*.ipin VCCBPIN
*.ipin VSSBPIN
*.ipin GP
*.iopin A
*.iopin Z
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends

**** begin user architecture code


* ngspice commands
* .options savecurrents
.param VCC = 1.8
.param SRCRES = 1k
.include stimuli_tb_passgatex4.cir
.control
save all
op
write tb_passgatex4.raw
set appendwrite
tran 10n 50u
write tb_passgatex4.raw
quit 0
.endc



**** end user architecture code
.end
