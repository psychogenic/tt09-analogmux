* NGSPICE file created from mux8onehot_parax.ext - technology: sky130A

.subckt mux8onehot_parax select1 select2 A1 A3 A2 A4 Z A8 select0 A7 A6 VDD A5 VSS
X0 a_5645_5909# a_5645_6085# a_5671_6037# VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1 VSS.t6 select1.t0 a_5645_6085# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 x5.A select2.t0 Z.t5 VDD.t31 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X3 x3.Z3 x1.gno0.t2 A5.t3 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X4 VSS.t50 a_5645_6461# x1.gno2 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X5 x1.gpo3.t3 x1.gno3.t2 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 x1.nSEL2 select2.t1 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VSS.t38 a_5645_5909# x1.gno1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VDD.t59 select0.t0 x1.nSEL0 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 x5.A select2.t2 Z.t4 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X10 A1.t1 x1.gpo0.t4 x5.A VDD.t60 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X11 x5.A x1.gno1 A2.t2 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X12 VDD.t74 VSS.t76 VDD.t73 VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X13 x3.Z3 x1.nSEL2 Z.t3 VDD.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X14 x1.nSEL0 select0.t1 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 x5.A x1.gno3.t3 A4.t1 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X16 VSS.t67 VDD.t79 VSS.t66 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X17 a_5671_6037# select0.t2 VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X18 A7.t3 x1.gpo2 x3.Z3 VDD.t77 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X19 x3.Z3 x1.nSEL2 Z.t2 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X20 Z.t1 x1.nSEL2 x5.A VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X21 A3.t3 x1.gpo2 x5.A VDD.t78 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X22 VSS.t75 select1.t1 x1.nSEL1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 x1.gpo3.t1 x1.gno3.t4 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 Z.t7 select2.t3 x3.Z3 VSS.t70 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X25 VSS.t3 a_5645_7149# x1.gno3.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X26 VDD.t57 a_5645_6637# a_5645_6461# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X27 x3.Z3 x1.gno1 A6.t3 VSS.t44 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X28 a_5645_7149# select1.t2 a_5699_7287# VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X29 x3.Z3 x1.gno0.t3 A5.t2 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X30 a_5645_6637# select0.t3 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X31 VSS.t24 x1.gno0.t4 x1.gpo0.t3 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 a_5699_7287# select0.t4 VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X33 VSS.t9 VDD.t80 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X34 x5.A x1.gno2 A3.t1 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X35 A8.t3 x1.gpo3.t4 x3.Z3 VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X36 A1.t0 x1.gpo0.t5 x5.A VDD.t60 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X37 a_5645_6461# a_5645_6637# a_5671_6589# VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X38 x5.A x1.gno3.t5 A4.t0 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X39 VSS.t32 x1.gno2 x1.gpo2 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 x1.gpo0.t2 x1.gno0.t5 VSS.t34 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X41 VSS.t64 select0.t5 a_5645_6637# VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X42 Z.t0 x1.nSEL2 x5.A VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X43 VDD.t19 select1.t3 x1.nSEL1 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X44 VDD.t17 select1.t4 a_5645_7149# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X45 A5.t1 x1.gpo0.t6 x3.Z3 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X46 VDD.t71 VSS.t77 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X47 Z.t6 select2.t4 x3.Z3 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X48 VDD.t41 a_5645_5493# x1.gno0.t0 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X49 a_5645_7149# select0.t6 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X50 VDD.t76 x1.gno0.t6 x1.gpo0.t1 VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X51 x3.Z3 x1.gno2 A7.t1 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X52 x3.Z3 x1.gno1 A6.t2 VSS.t44 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X53 A4.t3 x1.gpo3.t5 x5.A VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X54 VSS.t19 select2.t5 x1.nSEL2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 a_5645_5493# x1.nSEL0 a_5699_5631# VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X56 x1.nSEL1 select1.t5 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X57 x5.A x1.gno0.t7 A1.t3 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X58 VDD.t25 x1.gno2 x1.gpo2 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X59 x1.gpo0.t0 x1.gno0.t8 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 a_5645_5909# select0.t7 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X61 x5.A x1.gno2 A3.t0 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X62 A2.t3 x1.gpo1.t4 x5.A VDD.t5 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X63 x5.A x1.gno0.t9 A1.t2 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X64 A3.t2 x1.gpo2 x5.A VDD.t78 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X65 VDD.t68 VSS.t78 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X66 a_5699_5631# x1.nSEL1 VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X67 VSS.t73 VDD.t81 VSS.t72 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X68 x3.Z3 x1.gno3.t6 A8.t1 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X69 VDD.t45 a_5645_6461# x1.gno2 VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X70 VSS.t43 x1.gno1 x1.gpo1.t3 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X71 A6.t1 x1.gpo1.t5 x3.Z3 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X72 A5.t0 x1.gpo0.t7 x3.Z3 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X73 VDD.t51 x1.nSEL0 a_5645_5493# VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X74 x1.gpo1.t2 x1.gno1 VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X75 VSS.t69 x1.gno3.t7 x1.gpo3.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X76 VDD.t35 a_5645_5909# x1.gno1 VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X77 x1.gpo2 x1.gno2 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X78 A7.t2 x1.gpo2 x3.Z3 VDD.t77 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X79 x1.nSEL1 select1.t6 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X80 VDD.t27 select2.t6 x1.nSEL2 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X81 a_5671_6589# select1.t7 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X82 x3.Z3 x1.gno2 A7.t0 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X83 A8.t2 x1.gpo3.t6 x3.Z3 VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X84 A4.t2 x1.gpo3.t7 x5.A VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X85 a_5645_5493# x1.nSEL1 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X86 VSS.t46 a_5645_5493# x1.gno0.t1 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X87 VSS.t55 VDD.t82 VSS.t54 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X88 x5.A x1.gno1 A2.t1 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X89 VDD.t39 x1.gno1 x1.gpo1.t1 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X90 A2.t0 x1.gpo1.t6 x5.A VDD.t5 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X91 VDD.t3 a_5645_7149# x1.gno3.t0 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X92 x1.nSEL2 select2.t7 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X93 VSS.t48 select0.t8 x1.nSEL0 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X94 x1.gpo1.t0 x1.gno1 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X95 VDD.t49 x1.gno3.t8 x1.gpo3.t0 VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X96 x3.Z3 x1.gno3.t9 A8.t0 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X97 VDD.t55 a_5645_6085# a_5645_5909# VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X98 x1.gpo2 x1.gno2 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X99 VDD.t65 VSS.t79 VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X100 a_5645_6085# select1.t8 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X101 x1.nSEL0 select0.t9 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X102 a_5645_6461# select1.t9 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X103 A6.t0 x1.gpo1.t7 x3.Z3 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
R0 VSS.n237 VSS.n236 587674
R1 VSS.n171 VSS.n170 153375
R2 VSS.n193 VSS.n178 117542
R3 VSS.n249 VSS.n172 71206.2
R4 VSS.n249 VSS.n248 64736.2
R5 VSS.n238 VSS.n9 16580.8
R6 VSS.n242 VSS.n173 11744.7
R7 VSS.n247 VSS.n173 11744.7
R8 VSS.n242 VSS.n174 11744.7
R9 VSS.n247 VSS.n174 11744.7
R10 VSS.n253 VSS.n28 11744.7
R11 VSS.n253 VSS.n29 11744.7
R12 VSS.n257 VSS.n29 11744.7
R13 VSS.n257 VSS.n28 11744.7
R14 VSS.n264 VSS.n22 11744.7
R15 VSS.n260 VSS.n22 11744.7
R16 VSS.n264 VSS.n23 11744.7
R17 VSS.n260 VSS.n23 11744.7
R18 VSS.n271 VSS.n16 11744.7
R19 VSS.n267 VSS.n16 11744.7
R20 VSS.n271 VSS.n17 11744.7
R21 VSS.n267 VSS.n17 11744.7
R22 VSS.n278 VSS.n10 11744.7
R23 VSS.n274 VSS.n10 11744.7
R24 VSS.n278 VSS.n11 11744.7
R25 VSS.n274 VSS.n11 11744.7
R26 VSS.n190 VSS.n179 11744.7
R27 VSS.n185 VSS.n179 11744.7
R28 VSS.n190 VSS.n181 11744.7
R29 VSS.n185 VSS.n181 11744.7
R30 VSS.n205 VSS.n204 11744.7
R31 VSS.n201 VSS.n200 11744.7
R32 VSS.n204 VSS.n201 11744.7
R33 VSS.n234 VSS.n194 11744.7
R34 VSS.n230 VSS.n195 11744.7
R35 VSS.n234 VSS.n195 11744.7
R36 VSS.n218 VSS.n217 11744.7
R37 VSS.n214 VSS.n213 11744.7
R38 VSS.n217 VSS.n214 11744.7
R39 VSS.n281 VSS.n4 11744.7
R40 VSS.n281 VSS.n5 11744.7
R41 VSS.n7 VSS.n4 11744.7
R42 VSS.n237 VSS.n178 10428.2
R43 VSS.n238 VSS.n191 7573.12
R44 VSS.n191 VSS.t0 7065.1
R45 VSS.t1 VSS.n172 7065.1
R46 VSS.n180 VSS.t0 6710.74
R47 VSS.n180 VSS.t1 6710.74
R48 VSS.n241 VSS.n239 6647.5
R49 VSS.n273 VSS.n272 6049.9
R50 VSS.n241 VSS.t70 6006.85
R51 VSS.n248 VSS.t57 6006.85
R52 VSS.n259 VSS.n258 6004.3
R53 VSS.n280 VSS.n279 5972.7
R54 VSS.n266 VSS.n265 5963.12
R55 VSS.t70 VSS.n240 5705.56
R56 VSS.n240 VSS.t57 5705.56
R57 VSS.n239 VSS.n178 4796.58
R58 VSS.n238 VSS.n237 3666.67
R59 VSS.n192 VSS.n9 3385.09
R60 VSS.n15 VSS.n9 3361.58
R61 VSS.n27 VSS.n21 3305.56
R62 VSS.n235 VSS.n193 3279.94
R63 VSS.n21 VSS.n15 3275.35
R64 VSS.n62 VSS.n27 2366.85
R65 VSS.n250 VSS.n249 2235.82
R66 VSS.n236 VSS.n235 1652.78
R67 VSS.n236 VSS.n192 1652.78
R68 VSS.t2 VSS.n169 1550.96
R69 VSS VSS.t63 1289.66
R70 VSS.n137 VSS.n136 1198.25
R71 VSS.n159 VSS.n40 1198.25
R72 VSS.n169 VSS.n168 1194.5
R73 VSS.n140 VSS.n139 1171.32
R74 VSS.n251 VSS.n250 1006.48
R75 VSS.n169 VSS 918.774
R76 VSS.t45 VSS 918.774
R77 VSS.t61 VSS.t2 910.346
R78 VSS.t20 VSS.t49 826.054
R79 VSS.t35 VSS.t37 826.054
R80 VSS.t5 VSS.t74 792.337
R81 VSS.n256 VSS.n255 767.294
R82 VSS.n270 VSS.n269 767.294
R83 VSS.n232 VSS.n231 767.294
R84 VSS.n6 VSS.n3 767.294
R85 VSS.n263 VSS.n262 763.106
R86 VSS.n277 VSS.n276 763.106
R87 VSS.n202 VSS.n198 763.106
R88 VSS.n215 VSS.n211 763.106
R89 VSS.n243 VSS.n177 763.09
R90 VSS.n189 VSS.n182 763.09
R91 VSS.n177 VSS.n175 732.236
R92 VSS.n256 VSS.n30 732.236
R93 VSS.n270 VSS.n18 732.236
R94 VSS.n263 VSS.n24 732.236
R95 VSS.n277 VSS.n12 732.236
R96 VSS.n184 VSS.n182 732.236
R97 VSS.n207 VSS.n198 732.236
R98 VSS.n231 VSS.n228 732.236
R99 VSS.n220 VSS.n211 732.236
R100 VSS.n6 VSS.n1 732.236
R101 VSS.n250 VSS.n171 709.912
R102 VSS.t18 VSS.t25 708.047
R103 VSS.t74 VSS.t16 708.047
R104 VSS.t47 VSS.t10 708.047
R105 VSS.t58 VSS.t51 708.047
R106 VSS.n139 VSS.t65 606.351
R107 VSS.t56 VSS 564.751
R108 VSS.t25 VSS 564.751
R109 VSS.t10 VSS 564.751
R110 VSS VSS.t58 564.751
R111 VSS.n171 VSS 564.751
R112 VSS.n170 VSS.t56 522.606
R113 VSS.t51 VSS.t71 522.606
R114 VSS.t59 VSS 480.461
R115 VSS VSS.t53 408.628
R116 VSS.t71 VSS.t45 387.74
R117 VSS.n138 VSS 384.901
R118 VSS.t42 VSS.n137 374.356
R119 VSS.n40 VSS.t60 337.166
R120 VSS.n252 VSS.n251 332.642
R121 VSS.t68 VSS 329.539
R122 VSS.t31 VSS 329.539
R123 VSS.t23 VSS 329.539
R124 VSS.n255 VSS.n254 325.502
R125 VSS.n269 VSS.n268 325.502
R126 VSS.n233 VSS.n232 325.502
R127 VSS.n282 VSS.n3 325.502
R128 VSS.n40 VSS.t20 320.307
R129 VSS.n244 VSS.n243 304.553
R130 VSS.n189 VSS.n188 304.553
R131 VSS.n262 VSS.n261 304.204
R132 VSS.n276 VSS.n275 304.204
R133 VSS.n203 VSS.n202 304.204
R134 VSS.n216 VSS.n215 304.204
R135 VSS.t60 VSS 295.019
R136 VSS.n245 VSS.n244 266.349
R137 VSS.n188 VSS.n187 266.349
R138 VSS VSS.t5 261.303
R139 VSS.t7 VSS 244.445
R140 VSS.n254 VSS.n32 242.448
R141 VSS.n268 VSS.n20 242.448
R142 VSS.n261 VSS.n26 242.448
R143 VSS.n275 VSS.n14 242.448
R144 VSS.n203 VSS.n197 242.448
R145 VSS.n233 VSS.n196 242.448
R146 VSS.n216 VSS.n210 242.448
R147 VSS.n283 VSS.n282 242.448
R148 VSS.n152 VSS.t6 240.575
R149 VSS.n164 VSS.t64 237.327
R150 VSS.t12 VSS.t68 221.451
R151 VSS.t28 VSS.t31 221.451
R152 VSS.t40 VSS.t42 221.451
R153 VSS.t33 VSS.t23 221.451
R154 VSS.n106 VSS.t79 218.308
R155 VSS.n82 VSS.t78 218.308
R156 VSS.n50 VSS.t77 218.308
R157 VSS.n36 VSS.t76 218.308
R158 VSS.n103 VSS.t66 214.456
R159 VSS.n105 VSS.t67 214.456
R160 VSS.n80 VSS.t54 214.456
R161 VSS.n67 VSS.t55 214.456
R162 VSS.n45 VSS.t72 214.456
R163 VSS.n49 VSS.t73 214.456
R164 VSS.n34 VSS.t8 214.456
R165 VSS.n37 VSS.t9 214.456
R166 VSS.n74 VSS.n70 204.457
R167 VSS.n146 VSS.n44 200.231
R168 VSS.n39 VSS.n38 200.231
R169 VSS.n52 VSS.n47 200.105
R170 VSS.n137 VSS 197.724
R171 VSS.n139 VSS 197.724
R172 VSS.n276 VSS.n11 195
R173 VSS.n11 VSS.t22 195
R174 VSS.n13 VSS.n10 195
R175 VSS.n10 VSS.t22 195
R176 VSS.n269 VSS.n17 195
R177 VSS.n17 VSS.t30 195
R178 VSS.n19 VSS.n16 195
R179 VSS.n16 VSS.t30 195
R180 VSS.n262 VSS.n23 195
R181 VSS.n23 VSS.t39 195
R182 VSS.n25 VSS.n22 195
R183 VSS.n22 VSS.t39 195
R184 VSS.n31 VSS.n28 195
R185 VSS.n138 VSS.n28 195
R186 VSS.n255 VSS.n29 195
R187 VSS.n29 VSS.t4 195
R188 VSS.n186 VSS.n185 195
R189 VSS.n185 VSS.n172 195
R190 VSS.n190 VSS.n189 195
R191 VSS.n191 VSS.n190 195
R192 VSS.n247 VSS.n246 195
R193 VSS.n248 VSS.n247 195
R194 VSS.n243 VSS.n242 195
R195 VSS.n242 VSS.n241 195
R196 VSS.n202 VSS.n201 195
R197 VSS.n201 VSS.t14 195
R198 VSS.n206 VSS.n205 195
R199 VSS.n232 VSS.n195 195
R200 VSS.n195 VSS.t27 195
R201 VSS.n227 VSS.n194 195
R202 VSS.n215 VSS.n214 195
R203 VSS.n214 VSS.t44 195
R204 VSS.n219 VSS.n218 195
R205 VSS.n4 VSS.n2 195
R206 VSS.t15 VSS.n4 195
R207 VSS.n5 VSS.n3 195
R208 VSS.n8 VSS.n5 188.989
R209 VSS.n218 VSS.n212 188.988
R210 VSS.n229 VSS.n194 188.986
R211 VSS.n205 VSS.n199 188.984
R212 VSS.n170 VSS.t61 185.441
R213 VSS.n258 VSS.t4 183.936
R214 VSS VSS.t35 177.012
R215 VSS VSS.t28 176.633
R216 VSS VSS.t40 176.633
R217 VSS VSS.t33 176.633
R218 VSS.n251 VSS 176.633
R219 VSS.n200 VSS.n199 173.373
R220 VSS.n230 VSS.n229 173.304
R221 VSS.n213 VSS.n212 173.167
R222 VSS.n8 VSS.n7 173.097
R223 VSS.n115 VSS.t69 162.471
R224 VSS.n120 VSS.t32 162.471
R225 VSS.n64 VSS.t43 162.471
R226 VSS.n130 VSS.t24 162.471
R227 VSS.n41 VSS.t75 162.471
R228 VSS.n146 VSS.t48 160.046
R229 VSS.n39 VSS.t19 160.046
R230 VSS.n119 VSS.t13 160.017
R231 VSS.n63 VSS.t29 160.017
R232 VSS.n131 VSS.t41 160.017
R233 VSS.n126 VSS.t34 160.017
R234 VSS.n57 VSS.t11 160.017
R235 VSS.n147 VSS.t17 160.017
R236 VSS.n152 VSS.t26 158.534
R237 VSS.n279 VSS.t22 155.954
R238 VSS.n272 VSS.t30 155.954
R239 VSS.n265 VSS.t39 155.831
R240 VSS.n252 VSS.t4 139.648
R241 VSS.n204 VSS.n193 118.54
R242 VSS.n235 VSS.n234 111.895
R243 VSS.n217 VSS.n192 111.808
R244 VSS.n273 VSS.n15 99.881
R245 VSS.n266 VSS.n21 93.748
R246 VSS.n259 VSS.n27 93.6734
R247 VSS.n62 VSS.t12 89.635
R248 VSS.n9 VSS.t15 89.4314
R249 VSS VSS.n62 86.9987
R250 VSS.t16 VSS.t59 84.2917
R251 VSS.n239 VSS.n238 79.0175
R252 VSS.n47 VSS.t52 72.8576
R253 VSS.n70 VSS.t62 72.8576
R254 VSS.n280 VSS.n9 72.6343
R255 VSS.n235 VSS.t27 66.9242
R256 VSS.t44 VSS.n192 66.8669
R257 VSS.n21 VSS.t30 62.2068
R258 VSS.n27 VSS.t39 62.1573
R259 VSS.t14 VSS.n193 60.352
R260 VSS.n44 VSS.t36 58.5719
R261 VSS.n38 VSS.t21 58.5719
R262 VSS.n15 VSS.t22 56.0738
R263 VSS.n246 VSS.n245 54.2123
R264 VSS.n187 VSS.n186 54.2123
R265 VSS.t49 VSS.t18 50.5752
R266 VSS.t37 VSS.t47 50.5752
R267 VSS.n76 VSS 43.9579
R268 VSS.n253 VSS.n252 42.2329
R269 VSS.n76 VSS.n75 34.6358
R270 VSS.n73 VSS.n33 34.6358
R271 VSS.n246 VSS.n175 30.8711
R272 VSS.n31 VSS.n30 30.8711
R273 VSS.n19 VSS.n18 30.8711
R274 VSS.n25 VSS.n24 30.8711
R275 VSS.n13 VSS.n12 30.8711
R276 VSS.n186 VSS.n184 30.8711
R277 VSS.n207 VSS.n206 30.8711
R278 VSS.n228 VSS.n227 30.8711
R279 VSS.n220 VSS.n219 30.8711
R280 VSS.n2 VSS.n1 30.8711
R281 VSS.n140 VSS.n61 26.9246
R282 VSS.n168 VSS.n33 25.6926
R283 VSS.n44 VSS.t38 25.4291
R284 VSS.n38 VSS.t50 25.4291
R285 VSS.n115 VSS.n66 25.224
R286 VSS.n119 VSS.n66 25.224
R287 VSS.n121 VSS.n120 25.224
R288 VSS.n121 VSS.n63 25.224
R289 VSS.n132 VSS.n64 25.224
R290 VSS.n132 VSS.n131 25.224
R291 VSS.n130 VSS.n129 25.224
R292 VSS.n129 VSS.n126 25.224
R293 VSS.n57 VSS.n43 25.224
R294 VSS.n148 VSS.n41 25.224
R295 VSS.n148 VSS.n147 25.224
R296 VSS.n153 VSS.n152 24.0946
R297 VSS.t65 VSS.n138 23.7273
R298 VSS.n47 VSS.t46 22.3257
R299 VSS.n70 VSS.t3 22.3257
R300 VSS.n146 VSS.n43 21.4593
R301 VSS.n153 VSS.n39 21.4593
R302 VSS.n120 VSS.n119 20.3299
R303 VSS.n131 VSS.n130 20.3299
R304 VSS.n115 VSS.n114 19.2926
R305 VSS.n57 VSS.n56 17.7867
R306 VSS.n136 VSS.n64 17.3181
R307 VSS.t63 VSS.t7 16.8587
R308 VSS.n136 VSS.n63 15.8123
R309 VSS.n126 VSS.n61 15.8123
R310 VSS.n281 VSS.n280 15.1478
R311 VSS.n102 VSS.n61 14.775
R312 VSS.n160 VSS.n159 14.775
R313 VSS.n152 VSS.n41 13.5534
R314 VSS.n79 VSS.n78 11.2844
R315 VSS.n275 VSS.n274 11.0382
R316 VSS.n274 VSS.n273 11.0382
R317 VSS.n278 VSS.n277 11.0382
R318 VSS.n279 VSS.n278 11.0382
R319 VSS.n268 VSS.n267 11.0382
R320 VSS.n267 VSS.n266 11.0382
R321 VSS.n271 VSS.n270 11.0382
R322 VSS.n272 VSS.n271 11.0382
R323 VSS.n261 VSS.n260 11.0382
R324 VSS.n260 VSS.n259 11.0382
R325 VSS.n264 VSS.n263 11.0382
R326 VSS.n265 VSS.n264 11.0382
R327 VSS.n254 VSS.n253 11.0382
R328 VSS.n257 VSS.n256 11.0382
R329 VSS.n258 VSS.n257 11.0382
R330 VSS.n188 VSS.n181 11.0382
R331 VSS.n181 VSS.n180 11.0382
R332 VSS.n182 VSS.n179 11.0382
R333 VSS.n180 VSS.n179 11.0382
R334 VSS.n244 VSS.n174 11.0382
R335 VSS.n240 VSS.n174 11.0382
R336 VSS.n177 VSS.n173 11.0382
R337 VSS.n240 VSS.n173 11.0382
R338 VSS.n204 VSS.n203 11.0382
R339 VSS.n200 VSS.n198 11.0382
R340 VSS.n234 VSS.n233 11.0382
R341 VSS.n231 VSS.n230 11.0382
R342 VSS.n217 VSS.n216 11.0382
R343 VSS.n213 VSS.n211 11.0382
R344 VSS.n7 VSS.n6 11.0382
R345 VSS.n282 VSS.n281 11.0382
R346 VSS.n32 VSS.n31 10.9181
R347 VSS.n20 VSS.n19 10.9181
R348 VSS.n26 VSS.n25 10.9181
R349 VSS.n14 VSS.n13 10.9181
R350 VSS.n206 VSS.n197 10.9181
R351 VSS.n227 VSS.n196 10.9181
R352 VSS.n219 VSS.n210 10.9181
R353 VSS.n283 VSS.n2 10.9181
R354 VSS.n176 VSS.n175 10.4476
R355 VSS.n85 VSS.n30 10.4476
R356 VSS.n89 VSS.n18 10.4476
R357 VSS.n87 VSS.n24 10.4476
R358 VSS.n91 VSS.n12 10.4476
R359 VSS.n184 VSS.n183 10.4476
R360 VSS.n208 VSS.n207 10.4476
R361 VSS.n228 VSS.n226 10.4476
R362 VSS.n221 VSS.n220 10.4476
R363 VSS.n284 VSS.n1 10.4476
R364 VSS.n147 VSS.n146 10.1652
R365 VSS.n105 VSS.n100 9.70901
R366 VSS.n80 VSS.n79 9.70901
R367 VSS.n49 VSS.n48 9.70901
R368 VSS.n74 VSS.n73 9.41227
R369 VSS.n141 VSS.n140 9.3005
R370 VSS.n127 VSS.n126 9.3005
R371 VSS.n131 VSS.n124 9.3005
R372 VSS.n136 VSS.n135 9.3005
R373 VSS.n123 VSS.n63 9.3005
R374 VSS.n119 VSS.n118 9.3005
R375 VSS.n114 VSS.n113 9.3005
R376 VSS.n84 VSS.n83 9.3005
R377 VSS.n81 VSS.n68 9.3005
R378 VSS.n116 VSS.n115 9.3005
R379 VSS.n117 VSS.n66 9.3005
R380 VSS.n120 VSS.n65 9.3005
R381 VSS.n122 VSS.n121 9.3005
R382 VSS.n134 VSS.n64 9.3005
R383 VSS.n133 VSS.n132 9.3005
R384 VSS.n130 VSS.n125 9.3005
R385 VSS.n129 VSS.n128 9.3005
R386 VSS.n108 VSS.n107 9.3005
R387 VSS.n104 VSS.n99 9.3005
R388 VSS.n102 VSS.n101 9.3005
R389 VSS.n61 VSS.n59 9.3005
R390 VSS.n168 VSS.n167 9.3005
R391 VSS.n166 VSS.n165 9.3005
R392 VSS.n157 VSS.n39 9.3005
R393 VSS.n152 VSS.n151 9.3005
R394 VSS.n146 VSS.n145 9.3005
R395 VSS.n51 VSS.n46 9.3005
R396 VSS.n54 VSS.n53 9.3005
R397 VSS.n56 VSS.n55 9.3005
R398 VSS.n58 VSS.n57 9.3005
R399 VSS.n144 VSS.n43 9.3005
R400 VSS.n147 VSS.n42 9.3005
R401 VSS.n149 VSS.n148 9.3005
R402 VSS.n150 VSS.n41 9.3005
R403 VSS.n154 VSS.n153 9.3005
R404 VSS.n161 VSS.n160 9.3005
R405 VSS.n163 VSS.n162 9.3005
R406 VSS.n71 VSS.n33 9.3005
R407 VSS.n73 VSS.n72 9.3005
R408 VSS.n75 VSS.n69 9.3005
R409 VSS.n77 VSS.n76 9.3005
R410 VSS.n159 VSS.n158 9.3005
R411 VSS.n93 VSS.n92 8.45078
R412 VSS.n224 VSS.n209 8.45078
R413 VSS.n95 VSS.n86 8.30267
R414 VSS.n285 VSS.n0 8.30267
R415 VSS.n94 VSS.n88 7.97888
R416 VSS.n223 VSS.n222 7.97888
R417 VSS.n93 VSS.n90 7.97601
R418 VSS.n225 VSS.n224 7.97601
R419 VSS.n176 VSS 7.23036
R420 VSS.n183 VSS 7.23036
R421 VSS.n86 VSS.n85 7.16724
R422 VSS.n90 VSS.n89 7.16724
R423 VSS.n88 VSS.n87 7.16724
R424 VSS.n92 VSS.n91 7.16724
R425 VSS.n209 VSS.n208 7.16724
R426 VSS.n226 VSS.n225 7.16724
R427 VSS.n222 VSS.n221 7.16724
R428 VSS.n285 VSS.n284 7.16724
R429 VSS.n159 VSS.n39 7.15344
R430 VSS.n143 VSS.n142 6.50373
R431 VSS.n75 VSS.n74 6.4005
R432 VSS.n107 VSS.n104 6.26433
R433 VSS.n83 VSS.n81 6.26433
R434 VSS.n104 VSS.n103 5.85582
R435 VSS.n81 VSS.n80 5.85582
R436 VSS.n53 VSS.n45 5.85582
R437 VSS.n165 VSS.n34 5.85582
R438 VSS.n164 VSS.n163 5.85582
R439 VSS.n142 VSS.n59 4.788
R440 VSS.n85 VSS.n32 4.73093
R441 VSS.n89 VSS.n20 4.73093
R442 VSS.n87 VSS.n26 4.73093
R443 VSS.n91 VSS.n14 4.73093
R444 VSS.n208 VSS.n197 4.73093
R445 VSS.n226 VSS.n196 4.73093
R446 VSS.n221 VSS.n210 4.73093
R447 VSS.n284 VSS.n283 4.73093
R448 VSS.n142 VSS.n141 4.50726
R449 VSS.n97 VSS 4.01425
R450 VSS.n96 VSS 4.01425
R451 VSS.n245 VSS.n176 3.78485
R452 VSS.n187 VSS.n183 3.78485
R453 VSS.n52 VSS.n51 3.40476
R454 VSS.n107 VSS.n106 3.13241
R455 VSS.n83 VSS.n82 3.13241
R456 VSS.n51 VSS.n50 3.13241
R457 VSS.n163 VSS.n36 3.13241
R458 VSS.n155 VSS.n35 2.88636
R459 VSS.t14 VSS.n199 2.87953
R460 VSS.n229 VSS.t27 2.87839
R461 VSS.t44 VSS.n212 2.87611
R462 VSS.t15 VSS.n8 2.87497
R463 VSS.n53 VSS.n52 2.86007
R464 VSS.n106 VSS.n105 2.7239
R465 VSS.n82 VSS.n67 2.7239
R466 VSS.n50 VSS.n49 2.7239
R467 VSS.n37 VSS.n36 2.7239
R468 VSS.n112 VSS.n111 1.753
R469 VSS.n110 VSS.n109 1.753
R470 VSS VSS.n98 1.48125
R471 VSS.n156 VSS.n155 1.21169
R472 VSS.n98 VSS.n97 1.11894
R473 VSS.n111 VSS 0.95037
R474 VSS.n111 VSS.n110 0.761313
R475 VSS.n155 VSS 0.531208
R476 VSS.n94 VSS.n93 0.467019
R477 VSS.n224 VSS.n223 0.467019
R478 VSS.n103 VSS.n102 0.409011
R479 VSS.n114 VSS.n67 0.409011
R480 VSS.n56 VSS.n45 0.409011
R481 VSS.n168 VSS.n34 0.409011
R482 VSS.n165 VSS.n164 0.409011
R483 VSS.n160 VSS.n37 0.409011
R484 VSS.n97 VSS.n0 0.198729
R485 VSS.n96 VSS.n95 0.194976
R486 VSS.n141 VSS.n60 0.1255
R487 VSS.n79 VSS.n68 0.120292
R488 VSS.n84 VSS.n68 0.120292
R489 VSS.n117 VSS.n116 0.120292
R490 VSS.n118 VSS.n117 0.120292
R491 VSS.n122 VSS.n65 0.120292
R492 VSS.n123 VSS.n122 0.120292
R493 VSS.n134 VSS.n133 0.120292
R494 VSS.n133 VSS.n124 0.120292
R495 VSS.n128 VSS.n125 0.120292
R496 VSS.n128 VSS.n127 0.120292
R497 VSS.n101 VSS.n99 0.120292
R498 VSS.n108 VSS.n100 0.120292
R499 VSS.n77 VSS.n69 0.120292
R500 VSS.n72 VSS.n69 0.120292
R501 VSS.n72 VSS.n71 0.120292
R502 VSS.n162 VSS.n161 0.120292
R503 VSS.n150 VSS.n149 0.120292
R504 VSS.n149 VSS.n42 0.120292
R505 VSS.n145 VSS.n144 0.120292
R506 VSS.n55 VSS.n54 0.120292
R507 VSS.n54 VSS.n46 0.120292
R508 VSS.n48 VSS.n46 0.120292
R509 VSS.n162 VSS 0.0981562
R510 VSS.n78 VSS 0.09425
R511 VSS.n110 VSS 0.0881354
R512 VSS.n95 VSS.n94 0.0766574
R513 VSS.n223 VSS.n0 0.0766574
R514 VSS.n109 VSS.n108 0.0721146
R515 VSS.n156 VSS.n154 0.0708125
R516 VSS.n86 VSS 0.064875
R517 VSS.n90 VSS 0.064875
R518 VSS.n88 VSS 0.064875
R519 VSS.n225 VSS 0.064875
R520 VSS.n222 VSS 0.064875
R521 VSS VSS.n285 0.064875
R522 VSS.n92 VSS 0.063625
R523 VSS.n209 VSS 0.063625
R524 VSS.n112 VSS.n84 0.0616979
R525 VSS.n116 VSS 0.0603958
R526 VSS VSS.n65 0.0603958
R527 VSS.n135 VSS 0.0603958
R528 VSS VSS.n134 0.0603958
R529 VSS.n125 VSS 0.0603958
R530 VSS VSS.n59 0.0603958
R531 VSS.n101 VSS 0.0603958
R532 VSS.n71 VSS 0.0603958
R533 VSS VSS.n166 0.0603958
R534 VSS.n158 VSS 0.0603958
R535 VSS VSS.n157 0.0603958
R536 VSS.n154 VSS 0.0603958
R537 VSS.n151 VSS 0.0603958
R538 VSS VSS.n150 0.0603958
R539 VSS.n145 VSS 0.0603958
R540 VSS.n144 VSS 0.0603958
R541 VSS.n55 VSS 0.0603958
R542 VSS.n113 VSS.n112 0.0590938
R543 VSS VSS.n143 0.0590938
R544 VSS.n157 VSS.n156 0.0499792
R545 VSS.n109 VSS.n99 0.0486771
R546 VSS VSS.n35 0.0460729
R547 VSS.n98 VSS.n96 0.040297
R548 VSS.n167 VSS 0.0343542
R549 VSS.n135 VSS 0.0330521
R550 VSS.n158 VSS 0.0330521
R551 VSS VSS.n60 0.03175
R552 VSS.n113 VSS 0.0226354
R553 VSS.n118 VSS 0.0226354
R554 VSS VSS.n123 0.0226354
R555 VSS VSS.n124 0.0226354
R556 VSS.n127 VSS 0.0226354
R557 VSS.n100 VSS 0.0226354
R558 VSS.n166 VSS 0.0226354
R559 VSS.n161 VSS 0.0226354
R560 VSS.n151 VSS 0.0226354
R561 VSS VSS.n42 0.0226354
R562 VSS.n58 VSS 0.0226354
R563 VSS.n48 VSS 0.0226354
R564 VSS.n167 VSS.n35 0.0148229
R565 VSS.n78 VSS.n77 0.00440625
R566 VSS.n60 VSS.n59 0.00180208
R567 VSS.n143 VSS.n58 0.00180208
R568 select1.n10 select1.t8 327.99
R569 select1.n3 select1.t7 293.969
R570 select1.n6 select1.t4 256.07
R571 select1.n1 select1.t6 212.081
R572 select1.n0 select1.t3 212.081
R573 select1.n10 select1.t0 199.457
R574 select1.n2 select1.n1 182.929
R575 select1 select1.n3 154.065
R576 select1.n11 select1.n10 152
R577 select1.n7 select1.n6 152
R578 select1.n6 select1.t2 150.03
R579 select1.n1 select1.t5 139.78
R580 select1.n0 select1.t1 139.78
R581 select1.n3 select1.t9 138.338
R582 select1.n1 select1.n0 61.346
R583 select1.n5 select1 22.1096
R584 select1.n14 select1.n13 14.6836
R585 select1.n13 select1.n12 14.6704
R586 select1.n12 select1 13.8672
R587 select1.n4 select1 13.8328
R588 select1.n11 select1 12.1605
R589 select1.n14 select1.n2 10.6811
R590 select1.n7 select1.n5 10.4374
R591 select1.n9 select1.n8 8.15359
R592 select1.n2 select1 6.1445
R593 select1.n4 select1 5.16179
R594 select1.n9 select1.n4 4.65206
R595 select1.n8 select1 3.93896
R596 select1 select1.n11 2.34717
R597 select1.n5 select1 2.16665
R598 select1.n8 select1.n7 1.57588
R599 select1.n13 select1.n9 0.79438
R600 select1.n12 select1 0.6405
R601 select1 select1.n14 0.248606
R602 select2.n5 select2.t0 450.938
R603 select2.n5 select2.t2 445.666
R604 select2.n0 select2.t3 377.486
R605 select2.n0 select2.t4 374.202
R606 select2.n2 select2.t1 212.081
R607 select2.n1 select2.t6 212.081
R608 select2.n3 select2.n2 183.441
R609 select2.n2 select2.t7 139.78
R610 select2.n1 select2.t5 139.78
R611 select2.n2 select2.n1 61.346
R612 select2.n8 select2.n7 12.4093
R613 select2 select2.n3 11.4331
R614 select2.n7 select2.n6 9.10647
R615 select2.n7 select2.n4 8.98648
R616 select2.n3 select2 5.6325
R617 select2.n4 select2 5.02323
R618 select2.n6 select2.n5 3.1748
R619 select2.n8 select2.n0 2.10165
R620 select2.n9 select2 1.09425
R621 select2.n4 select2 0.941788
R622 select2.n6 select2 0.063625
R623 select2.n9 select2.n8 0.062375
R624 select2 select2.n9 0.003
R625 Z.n1 Z.t4 23.6581
R626 Z.n7 Z.t3 23.6581
R627 Z.n0 Z.t5 23.3739
R628 Z.n6 Z.t2 23.3739
R629 Z.n1 Z.t1 10.7528
R630 Z.n7 Z.t6 10.7528
R631 Z.n3 Z.t0 10.6417
R632 Z.n9 Z.t7 10.6417
R633 Z.n2 Z.n1 1.30064
R634 Z.n8 Z.n7 1.30064
R635 Z.n11 Z.n10 1.04212
R636 Z Z.n5 0.919875
R637 Z.n5 Z.n4 0.859481
R638 Z.n11 Z 0.754624
R639 Z.n2 Z.n0 0.726502
R640 Z.n8 Z.n6 0.726502
R641 Z.n3 Z.n2 0.512491
R642 Z.n9 Z.n8 0.512491
R643 Z.n4 Z.n3 0.359663
R644 Z.n10 Z.n9 0.359663
R645 Z.n4 Z.n0 0.216071
R646 Z.n10 Z.n6 0.216071
R647 Z Z.n11 0.0100278
R648 Z.n5 Z 0.001125
R649 VDD.n190 VDD.n188 8629.41
R650 VDD.n193 VDD.n187 8629.41
R651 VDD.n206 VDD.n205 8629.41
R652 VDD.n208 VDD.n203 8629.41
R653 VDD.n226 VDD.n220 8629.41
R654 VDD.n229 VDD.n219 8629.41
R655 VDD.n242 VDD.n241 8629.41
R656 VDD.n244 VDD.n238 8629.41
R657 VDD.n259 VDD.n252 8629.41
R658 VDD.n256 VDD.n253 8629.41
R659 VDD.n53 VDD.n52 8629.41
R660 VDD.n55 VDD.n50 8629.41
R661 VDD.n36 VDD.n35 8629.41
R662 VDD.n38 VDD.n33 8629.41
R663 VDD.n19 VDD.n17 8629.41
R664 VDD.n22 VDD.n16 8629.41
R665 VDD.n8 VDD.n2 8629.41
R666 VDD.n8 VDD.n3 8629.41
R667 VDD.n6 VDD.n2 8629.41
R668 VDD.n6 VDD.n3 8629.41
R669 VDD.n276 VDD.n270 8629.41
R670 VDD.n276 VDD.n271 8629.41
R671 VDD.n274 VDD.n270 8629.41
R672 VDD.n274 VDD.n271 8629.41
R673 VDD.n8 VDD.t0 2459.29
R674 VDD.t1 VDD.n6 2459.29
R675 VDD.n276 VDD.t31 2459.29
R676 VDD.t28 VDD.n274 2459.29
R677 VDD.t0 VDD.n7 2298.92
R678 VDD.n7 VDD.t1 2298.92
R679 VDD.t31 VDD.n275 2298.92
R680 VDD.n275 VDD.t28 2298.92
R681 VDD.n189 VDD.n186 920.471
R682 VDD.n209 VDD.n202 920.471
R683 VDD.n225 VDD.n221 920.471
R684 VDD.n245 VDD.n237 920.471
R685 VDD.n255 VDD.n254 920.471
R686 VDD.n56 VDD.n49 920.471
R687 VDD.n39 VDD.n32 920.471
R688 VDD.n18 VDD.n15 920.471
R689 VDD.n5 VDD.n4 920.471
R690 VDD.n273 VDD.n272 920.471
R691 VDD.n195 VDD.n186 914.447
R692 VDD.n210 VDD.n209 914.447
R693 VDD.n221 VDD.n217 914.447
R694 VDD.n246 VDD.n245 914.447
R695 VDD.n254 VDD.n251 914.447
R696 VDD.n58 VDD.n56 914.447
R697 VDD.n41 VDD.n39 914.447
R698 VDD.n24 VDD.n15 914.447
R699 VDD.n4 VDD.n0 914.447
R700 VDD.n272 VDD.n268 914.447
R701 VDD.t70 VDD.n124 804.731
R702 VDD.n126 VDD.t70 751.692
R703 VDD.n98 VDD.t17 671.408
R704 VDD.n87 VDD.t51 671.408
R705 VDD VDD.t69 630.375
R706 VDD.n157 VDD.n156 602.456
R707 VDD.n179 VDD.n67 602.456
R708 VDD.n71 VDD.n70 585
R709 VDD.n73 VDD.n72 585
R710 VDD.n5 VDD.n1 480.764
R711 VDD.n273 VDD.n269 480.764
R712 VDD.n189 VDD.n184 480.764
R713 VDD.n202 VDD.n200 480.764
R714 VDD.n225 VDD.n224 480.764
R715 VDD.n239 VDD.n237 480.764
R716 VDD.n255 VDD.n250 480.764
R717 VDD.n49 VDD.n47 480.764
R718 VDD.n32 VDD.n30 480.764
R719 VDD.n18 VDD.n14 480.764
R720 VDD VDD.t72 458.724
R721 VDD.t69 VDD 458.724
R722 VDD.n119 VDD.t26 420.25
R723 VDD.n115 VDD.t73 388.656
R724 VDD.n150 VDD.t74 388.656
R725 VDD.n128 VDD.t71 388.656
R726 VDD.n101 VDD.t67 388.656
R727 VDD.n110 VDD.t68 388.656
R728 VDD.n75 VDD.t64 388.656
R729 VDD.n80 VDD.t65 388.656
R730 VDD.n197 VDD.n184 379.2
R731 VDD.n212 VDD.n200 379.2
R732 VDD.n224 VDD.n223 379.2
R733 VDD.n239 VDD.n236 379.2
R734 VDD.n263 VDD.n250 379.2
R735 VDD.n60 VDD.n47 379.2
R736 VDD.n43 VDD.n30 379.2
R737 VDD.n26 VDD.n14 379.2
R738 VDD.n10 VDD.n1 379.2
R739 VDD.n278 VDD.n269 379.2
R740 VDD VDD.t18 369.938
R741 VDD VDD.t58 369.938
R742 VDD.n104 VDD.n97 322.329
R743 VDD.n82 VDD.n78 322.329
R744 VDD.n161 VDD.n159 259.697
R745 VDD.n137 VDD.t59 255.905
R746 VDD.n142 VDD.t19 255.905
R747 VDD.n118 VDD.t27 255.905
R748 VDD.n158 VDD.t25 255.905
R749 VDD.n108 VDD.t49 254.475
R750 VDD.n133 VDD.t53 252.95
R751 VDD.n138 VDD.t15 252.95
R752 VDD.n143 VDD.t30 252.95
R753 VDD.n178 VDD.t37 252.95
R754 VDD.n157 VDD.t33 251.516
R755 VDD.n68 VDD.t76 250.724
R756 VDD.n66 VDD.t39 250.724
R757 VDD.t26 VDD.t29 248.599
R758 VDD.t18 VDD.t14 248.599
R759 VDD.t58 VDD.t52 248.599
R760 VDD.n173 VDD.t9 248.219
R761 VDD.n160 VDD.t24 248.219
R762 VDD.n119 VDD 221.964
R763 VDD.n126 VDD.t81 215.827
R764 VDD.n108 VDD.n107 213.119
R765 VDD.n148 VDD.n119 213.119
R766 VDD.n116 VDD.t80 210.964
R767 VDD.n102 VDD.t82 210.964
R768 VDD.n77 VDD.t79 210.964
R769 VDD.n168 VDD.n167 209.368
R770 VDD.t29 VDD 198.287
R771 VDD.t14 VDD 198.287
R772 VDD.t52 VDD 198.287
R773 VDD.n170 VDD.n169 183.673
R774 VDD VDD.t2 182.952
R775 VDD VDD.n168 182.952
R776 VDD.t40 VDD 182.952
R777 VDD.n72 VDD.n71 159.476
R778 VDD.n159 VDD.t11 157.014
R779 VDD.t75 VDD.t42 154.417
R780 VDD.t56 VDD.t10 147.703
R781 VDD.t61 VDD.t16 140.989
R782 VDD.t10 VDD.t23 140.989
R783 VDD.t36 VDD.t38 140.989
R784 VDD.t8 VDD.t75 140.989
R785 VDD.t50 VDD.t46 140.989
R786 VDD.n159 VDD.t45 137.079
R787 VDD.n107 VDD 125.883
R788 VDD.n169 VDD 125.883
R789 VDD.n97 VDD.t62 116.341
R790 VDD.n78 VDD.t47 116.341
R791 VDD.t16 VDD 112.457
R792 VDD.t23 VDD 112.457
R793 VDD VDD.t50 112.457
R794 VDD VDD.t34 109.1
R795 VDD.n11 VDD.n0 105.788
R796 VDD.n279 VDD.n268 105.788
R797 VDD.t66 VDD.t61 104.064
R798 VDD.t46 VDD.t63 104.064
R799 VDD.t20 VDD 102.385
R800 VDD.t48 VDD 99.0288
R801 VDD.n156 VDD.t57 96.1553
R802 VDD.n67 VDD.t55 96.1553
R803 VDD VDD.t54 92.315
R804 VDD.n71 VDD.t43 86.7743
R805 VDD.n107 VDD.t48 83.9228
R806 VDD.n168 VDD.t44 80.5659
R807 VDD.t2 VDD.t66 77.209
R808 VDD.t63 VDD.t40 77.209
R809 VDD.n72 VDD.t35 66.8398
R810 VDD.n196 VDD.n195 66.6358
R811 VDD.n211 VDD.n210 66.6358
R812 VDD.n218 VDD.n217 66.6358
R813 VDD.n247 VDD.n246 66.6358
R814 VDD.n262 VDD.n251 66.6358
R815 VDD.n59 VDD.n58 66.6358
R816 VDD.n42 VDD.n41 66.6358
R817 VDD.n25 VDD.n24 66.6358
R818 VDD.n10 VDD.n9 63.3551
R819 VDD.n278 VDD.n277 63.3551
R820 VDD.n156 VDD.t21 63.3219
R821 VDD.n67 VDD.t13 63.3219
R822 VDD VDD.t56 62.103
R823 VDD.n190 VDD.n189 61.6672
R824 VDD.n194 VDD.n193 61.6672
R825 VDD.n206 VDD.n202 61.6672
R826 VDD.n203 VDD.n201 61.6672
R827 VDD.n226 VDD.n225 61.6672
R828 VDD.n230 VDD.n229 61.6672
R829 VDD.n242 VDD.n237 61.6672
R830 VDD.n238 VDD.n234 61.6672
R831 VDD.n260 VDD.n259 61.6672
R832 VDD.n256 VDD.n255 61.6672
R833 VDD.n53 VDD.n49 61.6672
R834 VDD.n50 VDD.n48 61.6672
R835 VDD.n36 VDD.n32 61.6672
R836 VDD.n33 VDD.n31 61.6672
R837 VDD.n19 VDD.n18 61.6672
R838 VDD.n23 VDD.n22 61.6672
R839 VDD.n6 VDD.n5 61.6672
R840 VDD.n9 VDD.n8 61.6672
R841 VDD.n274 VDD.n273 61.6672
R842 VDD.n277 VDD.n276 61.6672
R843 VDD.n191 VDD.n190 60.9564
R844 VDD.n193 VDD.n192 60.9564
R845 VDD.n207 VDD.n206 60.9564
R846 VDD.n204 VDD.n203 60.9564
R847 VDD.n227 VDD.n226 60.9564
R848 VDD.n229 VDD.n228 60.9564
R849 VDD.n243 VDD.n242 60.9564
R850 VDD.n240 VDD.n238 60.9564
R851 VDD.n259 VDD.n258 60.9564
R852 VDD.n257 VDD.n256 60.9564
R853 VDD.n54 VDD.n53 60.9564
R854 VDD.n51 VDD.n50 60.9564
R855 VDD.n37 VDD.n36 60.9564
R856 VDD.n34 VDD.n33 60.9564
R857 VDD.n20 VDD.n19 60.9564
R858 VDD.n22 VDD.n21 60.9564
R859 VDD.n211 VDD.n201 60.6123
R860 VDD.n230 VDD.n218 60.6123
R861 VDD.n59 VDD.n48 60.6123
R862 VDD.n42 VDD.n31 60.6123
R863 VDD.n196 VDD.n185 59.4829
R864 VDD.n262 VDD.n261 59.4829
R865 VDD.n248 VDD.n247 58.7299
R866 VDD.n25 VDD.n13 58.7299
R867 VDD.t42 VDD 55.3892
R868 VDD.t12 VDD 52.0323
R869 VDD VDD.t44 45.3185
R870 VDD VDD.t32 41.9616
R871 VDD.n191 VDD.n187 38.5759
R872 VDD.n192 VDD.n188 38.5759
R873 VDD.n208 VDD.n207 38.5759
R874 VDD.n205 VDD.n204 38.5759
R875 VDD.n227 VDD.n219 38.5759
R876 VDD.n228 VDD.n220 38.5759
R877 VDD.n244 VDD.n243 38.5759
R878 VDD.n241 VDD.n240 38.5759
R879 VDD.n257 VDD.n252 38.5759
R880 VDD.n258 VDD.n253 38.5759
R881 VDD.n55 VDD.n54 38.5759
R882 VDD.n52 VDD.n51 38.5759
R883 VDD.n38 VDD.n37 38.5759
R884 VDD.n35 VDD.n34 38.5759
R885 VDD.n20 VDD.n16 38.5759
R886 VDD.n21 VDD.n17 38.5759
R887 VDD.n167 VDD.n89 34.6358
R888 VDD.n167 VDD.n90 34.6358
R889 VDD.n172 VDD.n171 34.6358
R890 VDD.n169 VDD 28.5341
R891 VDD.n97 VDD.t3 28.4453
R892 VDD.n78 VDD.t41 28.4453
R893 VDD.n174 VDD.n173 28.3534
R894 VDD.n171 VDD.n170 25.6953
R895 VDD.n137 VDD.n122 25.224
R896 VDD.n133 VDD.n122 25.224
R897 VDD.n142 VDD.n121 25.224
R898 VDD.n138 VDD.n121 25.224
R899 VDD.n144 VDD.n118 25.224
R900 VDD.n144 VDD.n143 25.224
R901 VDD.n162 VDD.n158 25.224
R902 VDD.n108 VDD.n92 23.7181
R903 VDD VDD.n98 23.252
R904 VDD.n157 VDD.n92 21.4593
R905 VDD.n138 VDD.n137 20.3299
R906 VDD.n143 VDD.n142 20.3299
R907 VDD.t54 VDD.t36 20.1418
R908 VDD.n179 VDD.n66 19.9534
R909 VDD.n178 VDD.n177 19.8181
R910 VDD.n148 VDD.n118 17.3181
R911 VDD.n161 VDD.n160 17.3181
R912 VDD.n158 VDD.n157 16.5652
R913 VDD.n162 VDD.n161 16.5652
R914 VDD.n133 VDD.n132 15.8123
R915 VDD.n149 VDD.n148 14.2735
R916 VDD.n109 VDD.n108 14.2735
R917 VDD.n171 VDD.n87 13.9299
R918 VDD.n179 VDD.n178 13.5534
R919 VDD.n114 VDD.n113 11.4366
R920 VDD.n198 VDD.n197 11.3235
R921 VDD.n213 VDD.n212 11.3235
R922 VDD.n223 VDD.n222 11.3235
R923 VDD.n236 VDD.n235 11.3235
R924 VDD.n264 VDD.n263 11.3235
R925 VDD.n61 VDD.n60 11.3235
R926 VDD.n44 VDD.n43 11.3235
R927 VDD.n27 VDD.n26 11.3235
R928 VDD.n170 VDD.n88 11.2937
R929 VDD.n154 VDD.n153 11.2737
R930 VDD.t32 VDD.t20 10.0712
R931 VDD.n128 VDD.n125 9.60526
R932 VDD.n115 VDD.n114 9.60526
R933 VDD.n80 VDD.n79 9.60526
R934 VDD.n117 VDD.n93 9.3005
R935 VDD.n152 VDD.n151 9.3005
R936 VDD.n149 VDD.n94 9.3005
R937 VDD.n148 VDD.n147 9.3005
R938 VDD.n143 VDD.n120 9.3005
R939 VDD.n139 VDD.n138 9.3005
R940 VDD.n134 VDD.n133 9.3005
R941 VDD.n130 VDD.n129 9.3005
R942 VDD.n135 VDD.n122 9.3005
R943 VDD.n137 VDD.n136 9.3005
R944 VDD.n140 VDD.n121 9.3005
R945 VDD.n142 VDD.n141 9.3005
R946 VDD.n145 VDD.n144 9.3005
R947 VDD.n146 VDD.n118 9.3005
R948 VDD.n175 VDD.n174 9.3005
R949 VDD.n180 VDD.n179 9.3005
R950 VDD.n164 VDD.n89 9.3005
R951 VDD.n157 VDD.n155 9.3005
R952 VDD.n108 VDD.n106 9.3005
R953 VDD.n100 VDD.n99 9.3005
R954 VDD.n103 VDD.n95 9.3005
R955 VDD.n112 VDD.n111 9.3005
R956 VDD.n109 VDD.n96 9.3005
R957 VDD.n105 VDD.n92 9.3005
R958 VDD.n158 VDD.n91 9.3005
R959 VDD.n163 VDD.n162 9.3005
R960 VDD.n167 VDD.n166 9.3005
R961 VDD.n165 VDD.n90 9.3005
R962 VDD.n178 VDD.n65 9.3005
R963 VDD.n177 VDD.n176 9.3005
R964 VDD.n172 VDD.n69 9.3005
R965 VDD.n171 VDD.n74 9.3005
R966 VDD.n86 VDD.n85 9.3005
R967 VDD.n84 VDD.n83 9.3005
R968 VDD.n81 VDD.n76 9.3005
R969 VDD.n28 VDD.n13 8.23557
R970 VDD.n12 VDD.n11 7.54844
R971 VDD.n280 VDD.n279 7.54407
R972 VDD.n185 VDD.n183 6.88686
R973 VDD.n73 VDD.n70 6.8005
R974 VDD.n132 VDD.n124 6.48583
R975 VDD.n195 VDD.n194 6.02403
R976 VDD.n246 VDD.n234 6.02403
R977 VDD.n260 VDD.n251 6.02403
R978 VDD.n24 VDD.n23 6.02403
R979 VDD.n9 VDD.n0 6.02403
R980 VDD.n277 VDD.n268 6.02403
R981 VDD.n127 VDD.n126 5.8885
R982 VDD.n11 VDD.n10 5.18145
R983 VDD.n279 VDD.n278 5.18145
R984 VDD.n201 VDD.n64 4.89462
R985 VDD.n231 VDD.n217 4.89462
R986 VDD.n57 VDD.n48 4.89462
R987 VDD.n41 VDD.n40 4.89462
R988 VDD.n151 VDD.n117 4.67352
R989 VDD.n132 VDD.n131 4.62124
R990 VDD.n129 VDD.n128 4.36875
R991 VDD.n151 VDD.n150 4.36875
R992 VDD.n111 VDD.n110 4.36875
R993 VDD.n81 VDD.n80 4.36875
R994 VDD.t38 VDD.t12 3.35739
R995 VDD.t34 VDD.t8 3.35739
R996 VDD.n183 VDD 3.29986
R997 VDD.n215 VDD.n64 3.25464
R998 VDD.n249 VDD.n248 3.24308
R999 VDD.n57 VDD.n46 3.23917
R1000 VDD.n232 VDD.n231 3.23136
R1001 VDD.n40 VDD.n29 3.23136
R1002 VDD.n261 VDD.n63 3.22655
R1003 VDD.n129 VDD.n127 3.2005
R1004 VDD.n187 VDD.n186 2.84665
R1005 VDD.n188 VDD.n184 2.84665
R1006 VDD.n209 VDD.n208 2.84665
R1007 VDD.n205 VDD.n200 2.84665
R1008 VDD.n221 VDD.n219 2.84665
R1009 VDD.n224 VDD.n220 2.84665
R1010 VDD.n245 VDD.n244 2.84665
R1011 VDD.n241 VDD.n239 2.84665
R1012 VDD.n254 VDD.n252 2.84665
R1013 VDD.n253 VDD.n250 2.84665
R1014 VDD.n56 VDD.n55 2.84665
R1015 VDD.n52 VDD.n47 2.84665
R1016 VDD.n39 VDD.n38 2.84665
R1017 VDD.n35 VDD.n30 2.84665
R1018 VDD.n16 VDD.n15 2.84665
R1019 VDD.n17 VDD.n14 2.84665
R1020 VDD.n3 VDD.n1 2.84665
R1021 VDD.n7 VDD.n3 2.84665
R1022 VDD.n4 VDD.n2 2.84665
R1023 VDD.n7 VDD.n2 2.84665
R1024 VDD.n271 VDD.n269 2.84665
R1025 VDD.n275 VDD.n271 2.84665
R1026 VDD.n272 VDD.n270 2.84665
R1027 VDD.n275 VDD.n270 2.84665
R1028 VDD.n127 VDD.n124 2.8165
R1029 VDD.n104 VDD.n103 2.54018
R1030 VDD.n83 VDD.n82 2.54018
R1031 VDD.n117 VDD.n116 2.33701
R1032 VDD.n103 VDD.n102 2.33701
R1033 VDD.n83 VDD.n77 2.33701
R1034 VDD.n197 VDD.n196 2.28169
R1035 VDD.n212 VDD.n211 2.28169
R1036 VDD.n223 VDD.n218 2.28169
R1037 VDD.n247 VDD.n236 2.28169
R1038 VDD.n263 VDD.n262 2.28169
R1039 VDD.n60 VDD.n59 2.28169
R1040 VDD.n43 VDD.n42 2.28169
R1041 VDD.n26 VDD.n25 2.28169
R1042 VDD.n233 VDD.n232 2.13544
R1043 VDD.n111 VDD.n104 2.13383
R1044 VDD.n82 VDD.n81 2.13383
R1045 VDD.n267 VDD.n12 2.06883
R1046 VDD.n116 VDD.n115 2.03225
R1047 VDD.n102 VDD.n101 2.03225
R1048 VDD.n77 VDD.n75 2.03225
R1049 VDD.n249 VDD.n233 1.95379
R1050 VDD.n248 VDD.n234 1.88285
R1051 VDD.n23 VDD.n13 1.88285
R1052 VDD.n182 VDD.n181 1.753
R1053 VDD VDD.n182 1.64258
R1054 VDD.n90 VDD.n66 1.50638
R1055 VDD.n174 VDD.n73 1.4005
R1056 VDD.n100 VDD.n98 1.37193
R1057 VDD.n87 VDD.n86 1.37193
R1058 VDD.n280 VDD.n267 1.33758
R1059 VDD.n214 VDD.n213 1.143
R1060 VDD.n222 VDD.n216 1.143
R1061 VDD.n62 VDD.n61 1.143
R1062 VDD.n45 VDD.n44 1.143
R1063 VDD.n199 VDD.n198 1.13925
R1064 VDD.n265 VDD.n264 1.13925
R1065 VDD.n235 VDD.n233 1.13675
R1066 VDD.n28 VDD.n27 1.13675
R1067 VDD.n194 VDD.n185 1.12991
R1068 VDD.n210 VDD.n64 1.12991
R1069 VDD.n231 VDD.n230 1.12991
R1070 VDD.n261 VDD.n260 1.12991
R1071 VDD.n58 VDD.n57 1.12991
R1072 VDD.n40 VDD.n31 1.12991
R1073 VDD.n123 VDD 1.06099
R1074 VDD.n46 VDD.n45 0.862816
R1075 VDD.n214 VDD.n199 0.854667
R1076 VDD.n29 VDD.n28 0.770881
R1077 VDD.n160 VDD.n89 0.753441
R1078 VDD.n173 VDD.n172 0.753441
R1079 VDD.n63 VDD.n62 0.747859
R1080 VDD.n267 VDD.n266 0.704667
R1081 VDD.n70 VDD.n68 0.6005
R1082 VDD.n216 VDD.n215 0.588641
R1083 VDD.n265 VDD.n249 0.518882
R1084 VDD.n182 VDD 0.460219
R1085 VDD.n177 VDD.n68 0.4005
R1086 VDD.n45 VDD.n29 0.392323
R1087 VDD.n62 VDD.n46 0.360318
R1088 VDD.n150 VDD.n149 0.305262
R1089 VDD.n101 VDD.n100 0.305262
R1090 VDD.n110 VDD.n109 0.305262
R1091 VDD.n86 VDD.n75 0.305262
R1092 VDD.t60 VDD.n191 0.27666
R1093 VDD.n192 VDD.t60 0.27666
R1094 VDD.n207 VDD.t5 0.27666
R1095 VDD.n204 VDD.t5 0.27666
R1096 VDD.t78 VDD.n227 0.27666
R1097 VDD.n228 VDD.t78 0.27666
R1098 VDD.n243 VDD.t22 0.27666
R1099 VDD.n240 VDD.t22 0.27666
R1100 VDD.t4 VDD.n257 0.27666
R1101 VDD.n258 VDD.t4 0.27666
R1102 VDD.n54 VDD.t6 0.27666
R1103 VDD.n51 VDD.t6 0.27666
R1104 VDD.n37 VDD.t77 0.27666
R1105 VDD.n34 VDD.t77 0.27666
R1106 VDD.t7 VDD.n20 0.27666
R1107 VDD.n21 VDD.t7 0.27666
R1108 VDD.n215 VDD.n214 0.268128
R1109 VDD.n232 VDD.n216 0.223986
R1110 VDD.n199 VDD.n183 0.202423
R1111 VDD.n131 VDD.n130 0.180304
R1112 VDD.n131 VDD 0.120408
R1113 VDD.n114 VDD.n93 0.120292
R1114 VDD.n152 VDD.n94 0.120292
R1115 VDD.n146 VDD.n145 0.120292
R1116 VDD.n145 VDD.n120 0.120292
R1117 VDD.n141 VDD.n140 0.120292
R1118 VDD.n140 VDD.n139 0.120292
R1119 VDD.n136 VDD.n135 0.120292
R1120 VDD.n135 VDD.n134 0.120292
R1121 VDD.n130 VDD.n125 0.120292
R1122 VDD.n99 VDD.n95 0.120292
R1123 VDD.n112 VDD.n96 0.120292
R1124 VDD.n163 VDD.n91 0.120292
R1125 VDD.n164 VDD.n163 0.120292
R1126 VDD.n180 VDD.n65 0.120292
R1127 VDD.n176 VDD.n175 0.120292
R1128 VDD.n175 VDD.n69 0.120292
R1129 VDD.n85 VDD.n84 0.120292
R1130 VDD.n84 VDD.n76 0.120292
R1131 VDD.n79 VDD.n76 0.120292
R1132 VDD.n153 VDD.n93 0.11899
R1133 VDD.n266 VDD.n63 0.1125
R1134 VDD.n99 VDD 0.0981562
R1135 VDD.n154 VDD 0.0955521
R1136 VDD.n113 VDD.n95 0.0916458
R1137 VDD.n198 VDD 0.06425
R1138 VDD.n213 VDD 0.06425
R1139 VDD.n222 VDD 0.06425
R1140 VDD.n235 VDD 0.06425
R1141 VDD.n264 VDD 0.06425
R1142 VDD.n61 VDD 0.06425
R1143 VDD.n44 VDD 0.06425
R1144 VDD.n27 VDD 0.06425
R1145 VDD VDD.n280 0.06425
R1146 VDD.n147 VDD 0.0603958
R1147 VDD VDD.n146 0.0603958
R1148 VDD.n141 VDD 0.0603958
R1149 VDD.n136 VDD 0.0603958
R1150 VDD.n106 VDD 0.0603958
R1151 VDD VDD.n105 0.0603958
R1152 VDD VDD.n91 0.0603958
R1153 VDD.n166 VDD 0.0603958
R1154 VDD VDD.n165 0.0603958
R1155 VDD.n176 VDD 0.0603958
R1156 VDD.n85 VDD 0.0603958
R1157 VDD.n12 VDD 0.059875
R1158 VDD.n88 VDD 0.0590938
R1159 VDD.n266 VDD.n265 0.054
R1160 VDD.n181 VDD 0.0525833
R1161 VDD.n181 VDD.n180 0.0460729
R1162 VDD.n106 VDD 0.0382604
R1163 VDD VDD.n123 0.0369583
R1164 VDD.n147 VDD 0.03175
R1165 VDD.n166 VDD 0.03175
R1166 VDD.n113 VDD.n112 0.0291458
R1167 VDD VDD.n94 0.0226354
R1168 VDD VDD.n120 0.0226354
R1169 VDD.n139 VDD 0.0226354
R1170 VDD.n134 VDD 0.0226354
R1171 VDD.n125 VDD 0.0226354
R1172 VDD VDD.n96 0.0226354
R1173 VDD.n105 VDD 0.0226354
R1174 VDD.n155 VDD 0.0226354
R1175 VDD VDD.n164 0.0226354
R1176 VDD.n165 VDD 0.0226354
R1177 VDD VDD.n65 0.0226354
R1178 VDD VDD.n69 0.0226354
R1179 VDD VDD.n74 0.0226354
R1180 VDD.n79 VDD 0.0226354
R1181 VDD.n155 VDD.n154 0.00310417
R1182 VDD.n153 VDD.n152 0.00180208
R1183 VDD.n123 VDD 0.00180208
R1184 VDD.n88 VDD.n74 0.00180208
R1185 x1.gno0.n2 x1.gno0.t9 377.486
R1186 x1.gno0.n3 x1.gno0.t2 377.486
R1187 x1.gno0.n2 x1.gno0.t7 374.202
R1188 x1.gno0.n3 x1.gno0.t3 374.202
R1189 x1.gno0.n10 x1.gno0.t0 339.418
R1190 x1.gno0.n1 x1.gno0.t1 274.06
R1191 x1.gno0.n7 x1.gno0.t8 212.081
R1192 x1.gno0.n6 x1.gno0.t6 212.081
R1193 x1.gno0.n8 x1.gno0.n7 182.673
R1194 x1.gno0.n7 x1.gno0.t5 139.78
R1195 x1.gno0.n6 x1.gno0.t4 139.78
R1196 x1.gno0.n7 x1.gno0.n6 61.346
R1197 x1.gno0.n5 x1.gno0.n8 15.8606
R1198 x1.gno0 x1.gno0.n9 13.8044
R1199 x1.gno0.n0 x1.gno0.n4 13.4101
R1200 x1.gno0.n0 x1.gno0 11.5859
R1201 x1.gno0.n4 x1.gno0 11.5859
R1202 x1.gno0 x1.gno0.n1 11.0989
R1203 x1.gno0.n9 x1.gno0.n5 6.94768
R1204 x1.gno0 x1.gno0.n0 6.73859
R1205 x1.gno0.n11 x1.gno0 6.6565
R1206 x1.gno0.n8 x1.gno0 6.4005
R1207 x1.gno0.n1 x1.gno0 6.1445
R1208 x1.gno0.n0 x1.gno0 5.13959
R1209 x1.gno0.n4 x1.gno0 4.55738
R1210 x1.gno0.n11 x1.gno0.n10 4.0914
R1211 x1.gno0 x1.gno0.n11 3.61789
R1212 x1.gno0.n9 x1.gno0 3.26325
R1213 x1.gno0.n1 x1.gno0 2.86947
R1214 x1.gno0 x1.gno0.n2 2.04102
R1215 x1.gno0 x1.gno0.n3 2.04102
R1216 x1.gno0.n10 x1.gno0 1.74382
R1217 x1.gno0.n5 x1.gno0 1.47326
R1218 A5.n1 A5.t0 26.3998
R1219 A5.n1 A5.t1 23.5483
R1220 A5.n0 A5.t3 12.7127
R1221 A5.n0 A5.t2 10.8578
R1222 A5.n2 A5.n1 3.12177
R1223 A5.n2 A5.n0 1.81453
R1224 A5.n3 A5.n2 1.1255
R1225 A5.n3 A5 0.21549
R1226 A5 A5.n3 0.0655
R1227 x1.gno3.n3 x1.gno3.t3 377.486
R1228 x1.gno3.n1 x1.gno3.t6 377.486
R1229 x1.gno3.n3 x1.gno3.t5 374.202
R1230 x1.gno3.n1 x1.gno3.t9 374.202
R1231 x1.gno3.n9 x1.gno3.t0 339.418
R1232 x1.gno3.n0 x1.gno3.t1 274.06
R1233 x1.gno3.n6 x1.gno3.t4 212.081
R1234 x1.gno3.n5 x1.gno3.t8 212.081
R1235 x1.gno3.n7 x1.gno3.n6 184.977
R1236 x1.gno3.n6 x1.gno3.t2 139.78
R1237 x1.gno3.n5 x1.gno3.t7 139.78
R1238 x1.gno3.n6 x1.gno3.n5 61.346
R1239 x1.gno3.n8 x1.gno3 18.2601
R1240 x1.gno3 x1.gno3.n7 13.8193
R1241 x1.gno3 x1.gno3.n4 11.7568
R1242 x1.gno3.n4 x1.gno3.n2 11.6628
R1243 x1.gno3 x1.gno3.n0 11.2645
R1244 x1.gno3 x1.gno3.n8 8.9605
R1245 x1.gno3.n8 x1.gno3 8.4485
R1246 x1.gno3.n2 x1.gno3 8.16743
R1247 x1.gno3.n10 x1.gno3 6.6565
R1248 x1.gno3.n0 x1.gno3 6.1445
R1249 x1.gno3.n4 x1.gno3 5.8185
R1250 x1.gno3.n2 x1.gno3 4.58237
R1251 x1.gno3.n7 x1.gno3 4.0965
R1252 x1.gno3.n10 x1.gno3.n9 4.0914
R1253 x1.gno3 x1.gno3.n10 3.61789
R1254 x1.gno3.n0 x1.gno3 2.86947
R1255 x1.gno3 x1.gno3.n3 2.04102
R1256 x1.gno3 x1.gno3.n1 2.04102
R1257 x1.gno3.n9 x1.gno3 1.74382
R1258 x1.gpo3.n3 x1.gpo3.t7 450.938
R1259 x1.gpo3.n2 x1.gpo3.t4 450.938
R1260 x1.gpo3.n3 x1.gpo3.t5 445.666
R1261 x1.gpo3.n2 x1.gpo3.t6 445.666
R1262 x1.gpo3 x1.gpo3.n7 203.923
R1263 x1.gpo3.n1 x1.gpo3.n0 101.49
R1264 x1.gpo3.n7 x1.gpo3.t0 26.5955
R1265 x1.gpo3.n7 x1.gpo3.t1 26.5955
R1266 x1.gpo3.n0 x1.gpo3.t2 24.9236
R1267 x1.gpo3.n0 x1.gpo3.t3 24.9236
R1268 x1.gpo3.n4 x1.gpo3 11.0619
R1269 x1.gpo3.n6 x1.gpo3 10.7525
R1270 x1.gpo3 x1.gpo3.n4 9.34192
R1271 x1.gpo3.n5 x1.gpo3 7.73829
R1272 x1.gpo3.n6 x1.gpo3 6.6565
R1273 x1.gpo3.n4 x1.gpo3 5.84951
R1274 x1.gpo3 x1.gpo3.n6 5.04292
R1275 x1.gpo3 x1.gpo3.n3 2.95993
R1276 x1.gpo3 x1.gpo3.n2 2.95993
R1277 x1.gpo3.n1 x1.gpo3 1.93989
R1278 x1.gpo3 x1.gpo3.n5 1.5365
R1279 x1.gpo3.n5 x1.gpo3.n1 1.0245
R1280 select0.n5 select0.t3 327.99
R1281 select0.n9 select0.t2 293.969
R1282 select0.n3 select0.t6 261.887
R1283 select0.n1 select0.t1 212.081
R1284 select0.n0 select0.t0 212.081
R1285 select0.n5 select0.t5 199.457
R1286 select0.n2 select0.n1 183.185
R1287 select0.n3 select0.t4 155.847
R1288 select0 select0.n9 154.065
R1289 select0.n6 select0.n5 152
R1290 select0.n4 select0.n3 152
R1291 select0.n1 select0.t9 139.78
R1292 select0.n0 select0.t8 139.78
R1293 select0.n9 select0.t7 138.338
R1294 select0.n1 select0.n0 61.346
R1295 select0.n10 select0 13.4199
R1296 select0.n8 select0.n4 11.9062
R1297 select0.n11 select0.n8 11.7395
R1298 select0.n12 select0.n11 11.5949
R1299 select0.n12 select0.n2 9.68118
R1300 select0.n7 select0 9.17383
R1301 select0.n2 select0 5.8885
R1302 select0.n10 select0 5.57469
R1303 select0.n8 select0.n7 4.6505
R1304 select0.n11 select0.n10 4.6505
R1305 select0.n7 select0.n6 2.98717
R1306 select0.n6 select0 2.34717
R1307 select0.n4 select0 2.07109
R1308 select0 select0.n12 0.559212
R1309 x1.gpo0.n4 x1.gpo0.t5 450.938
R1310 x1.gpo0.n3 x1.gpo0.t7 450.938
R1311 x1.gpo0.n4 x1.gpo0.t4 445.666
R1312 x1.gpo0.n3 x1.gpo0.t6 445.666
R1313 x1.gpo0.n7 x1.gpo0.n6 195.832
R1314 x1.gpo0.n1 x1.gpo0.n0 101.49
R1315 x1.gpo0.n6 x1.gpo0.t1 26.5955
R1316 x1.gpo0.n6 x1.gpo0.t0 26.5955
R1317 x1.gpo0.n0 x1.gpo0.t3 24.9236
R1318 x1.gpo0.n0 x1.gpo0.t2 24.9236
R1319 x1.gpo0.n5 x1.gpo0 13.3282
R1320 x1.gpo0.n7 x1.gpo0 11.8923
R1321 x1.gpo0.n2 x1.gpo0 10.7525
R1322 x1.gpo0 x1.gpo0.n7 8.09215
R1323 x1.gpo0.n2 x1.gpo0 6.6565
R1324 x1.gpo0 x1.gpo0.n5 5.46644
R1325 x1.gpo0.n5 x1.gpo0 5.31412
R1326 x1.gpo0 x1.gpo0.n2 5.04292
R1327 x1.gpo0 x1.gpo0.n4 3.18415
R1328 x1.gpo0 x1.gpo0.n3 2.90754
R1329 x1.gpo0 x1.gpo0.n1 2.5605
R1330 x1.gpo0.n1 x1.gpo0 1.93989
R1331 A1.n1 A1.t0 26.3998
R1332 A1.n1 A1.t1 23.5483
R1333 A1.n0 A1.t2 12.7127
R1334 A1.n0 A1.t3 10.8578
R1335 A1.n2 A1.n1 3.12177
R1336 A1.n2 A1.n0 1.81453
R1337 A1.n3 A1.n2 1.1255
R1338 A1.n3 A1 0.21549
R1339 A1 A1.n3 0.0655
R1340 A2.n1 A2.t0 26.3998
R1341 A2.n1 A2.t3 23.5483
R1342 A2.n0 A2.t1 12.7127
R1343 A2.n0 A2.t2 10.8578
R1344 A2.n2 A2.n1 3.12177
R1345 A2.n2 A2.n0 1.81453
R1346 A2.n3 A2.n2 1.1255
R1347 A2.n3 A2 0.219402
R1348 A2 A2.n3 0.0655
R1349 A4.n1 A4.t2 26.3998
R1350 A4.n1 A4.t3 23.5483
R1351 A4.n0 A4.t1 12.7127
R1352 A4.n0 A4.t0 10.8578
R1353 A4.n2 A4.n1 3.12177
R1354 A4.n2 A4.n0 1.81453
R1355 A4.n3 A4.n2 1.1255
R1356 A4 A4.n3 0.203263
R1357 A4.n3 A4 0.0655
R1358 A7.n1 A7.t2 26.3998
R1359 A7.n1 A7.t3 23.5483
R1360 A7.n0 A7.t1 12.7127
R1361 A7.n0 A7.t0 10.8578
R1362 A7.n2 A7.n1 3.12177
R1363 A7.n2 A7.n0 1.81453
R1364 A7.n3 A7.n2 1.1255
R1365 A7.n3 A7 0.210543
R1366 A7 A7.n3 0.0655
R1367 A3.n1 A3.t3 26.3998
R1368 A3.n1 A3.t2 23.5483
R1369 A3.n0 A3.t1 12.7127
R1370 A3.n0 A3.t0 10.8578
R1371 A3.n2 A3.n1 3.12177
R1372 A3.n2 A3.n0 1.81453
R1373 A3.n3 A3.n2 1.1255
R1374 A3.n3 A3 0.210543
R1375 A3 A3.n3 0.0655
R1376 A6.n1 A6.t0 26.3998
R1377 A6.n1 A6.t1 23.5483
R1378 A6.n0 A6.t3 12.7127
R1379 A6.n0 A6.t2 10.8578
R1380 A6.n2 A6.n1 3.12177
R1381 A6.n2 A6.n0 1.81453
R1382 A6.n3 A6.n2 1.1255
R1383 A6.n3 A6 0.219402
R1384 A6 A6.n3 0.0655
R1385 A8.n1 A8.t3 26.3998
R1386 A8.n1 A8.t2 23.5483
R1387 A8.n0 A8.t1 12.7127
R1388 A8.n0 A8.t0 10.8578
R1389 A8.n2 A8.n1 3.12177
R1390 A8.n2 A8.n0 1.81453
R1391 A8.n3 A8.n2 1.1255
R1392 A8 A8.n3 0.203263
R1393 A8.n3 A8 0.0655
R1394 x1.gpo1.n4 x1.gpo1.t6 450.938
R1395 x1.gpo1.n3 x1.gpo1.t7 450.938
R1396 x1.gpo1.n4 x1.gpo1.t4 445.666
R1397 x1.gpo1.n3 x1.gpo1.t5 445.666
R1398 x1.gpo1.n7 x1.gpo1.n6 195.958
R1399 x1.gpo1.n1 x1.gpo1.n0 101.49
R1400 x1.gpo1.n6 x1.gpo1.t1 26.5955
R1401 x1.gpo1.n6 x1.gpo1.t0 26.5955
R1402 x1.gpo1.n0 x1.gpo1.t3 24.9236
R1403 x1.gpo1.n0 x1.gpo1.t2 24.9236
R1404 x1.gpo1.n5 x1.gpo1 14.964
R1405 x1.gpo1.n7 x1.gpo1 11.8408
R1406 x1.gpo1.n2 x1.gpo1 10.7525
R1407 x1.gpo1 x1.gpo1.n5 8.86265
R1408 x1.gpo1 x1.gpo1.n7 7.96524
R1409 x1.gpo1.n2 x1.gpo1 6.6565
R1410 x1.gpo1.n5 x1.gpo1 5.75481
R1411 x1.gpo1 x1.gpo1.n2 5.04292
R1412 x1.gpo1 x1.gpo1.n4 2.94361
R1413 x1.gpo1 x1.gpo1.n3 2.94361
R1414 x1.gpo1 x1.gpo1.n1 2.5605
R1415 x1.gpo1.n1 x1.gpo1 1.93989
C0 x1.nSEL0 x1.nSEL2 0.043717f
C1 x1.gno1 select2 0.001516f
C2 VDD a_5645_5493# 0.21052f
C3 x1.nSEL1 x1.nSEL2 0.10521f
C4 x5.A x1.gpo1 0.350703f
C5 x1.gno0 x1.gpo3 0.848624f
C6 x5.A x1.gno3 0.446599f
C7 x1.gpo2 x1.gpo0 0.062293f
C8 a_5671_6589# select0 0.001558f
C9 A3 x1.nSEL2 7.03e-21
C10 x1.gno1 A4 6.05e-19
C11 x1.gno3 a_5645_7149# 0.134079f
C12 x1.gno0 A6 3.66e-20
C13 x1.gpo3 A8 4.00906f
C14 select2 x1.nSEL2 4.00521f
C15 select0 x1.gno2 0.254198f
C16 a_5645_7149# a_5699_7287# 0.006584f
C17 x1.nSEL0 x1.gno0 0.002613f
C18 x1.gno0 x1.nSEL1 0.034871f
C19 A8 A6 2.39e-19
C20 select1 VDD 2.65613f
C21 x1.gpo2 x1.gpo3 0.109471f
C22 x1.gno1 a_5645_6461# 1.61e-19
C23 A7 x3.Z3 4.5214f
C24 x1.gpo3 a_5645_6637# 4.96e-19
C25 A3 x1.gno0 0.131584f
C26 Z select2 0.799881f
C27 a_5645_5909# x1.gno1 0.106139f
C28 m2_5776_5494# VDD 0.139797f
C29 select1 a_5645_5493# 0.02803f
C30 x3.Z3 x1.gno2 0.429865f
C31 x1.gpo1 x1.gno1 3.78638f
C32 A2 x1.gno2 0.137879f
C33 x1.gpo2 A6 0.001573f
C34 x1.gno3 x1.gno1 0.061048f
C35 m2_5776_5494# a_5645_5493# 0.01297f
C36 x1.gno0 select2 0.054258f
C37 A1 VDD 1.6325f
C38 a_5671_6589# x1.gno2 0.001073f
C39 a_5645_6085# x1.gno1 0.016995f
C40 x1.nSEL2 a_5645_6461# 3.51e-19
C41 x1.gno1 a_5699_7287# 8.14e-21
C42 A7 x1.gno2 3.80762f
C43 x1.nSEL0 a_5645_6637# 1.21e-20
C44 a_5645_5909# x1.nSEL2 3.56e-19
C45 x1.nSEL1 a_5645_6637# 1.59e-19
C46 x1.gno0 A4 0.218459f
C47 A5 x3.Z3 4.52088f
C48 x1.gpo1 x1.nSEL2 1.7e-20
C49 x1.gno3 x1.nSEL2 9.02e-19
C50 A3 x1.gpo2 3.96087f
C51 a_5645_7149# select0 0.220366f
C52 a_5699_5631# select0 9.55e-19
C53 a_5645_6085# x1.nSEL2 3.26e-19
C54 x1.gpo2 select2 1.6e-19
C55 select1 m2_5776_5494# 0.183786f
C56 x5.A x3.Z3 2.05508f
C57 Z x1.gpo1 2.41e-19
C58 A2 x5.A 4.52052f
C59 x1.gpo0 VDD 3.28453f
C60 x1.gno0 a_5645_6461# 7.95e-20
C61 A5 x1.gno2 2.86e-19
C62 Z x1.gno3 9.07e-20
C63 a_5645_5909# x1.gno0 0.012357f
C64 x1.gpo1 x1.gno0 0.069439f
C65 select1 A1 4.98e-22
C66 x1.gpo2 A4 0.162086f
C67 x1.gno3 x1.gno0 0.145529f
C68 a_5671_6037# x1.gno2 5.17e-20
C69 x1.gno0 a_5645_6085# 1.45e-19
C70 x1.gno1 select0 0.114399f
C71 x5.A x1.gno2 0.429924f
C72 x1.gpo1 A8 2.07e-19
C73 x1.gpo3 VDD 2.92994f
C74 x1.gno3 A8 3.84592f
C75 a_5645_7149# x1.gno2 1.07e-20
C76 x1.gpo2 a_5645_6461# 0.001353f
C77 a_5645_6637# a_5645_6461# 0.185422f
C78 x1.gno1 x3.Z3 0.429208f
C79 x1.gpo1 x1.gpo2 0.096269f
C80 VDD A6 1.60651f
C81 A2 x1.gno1 3.7791f
C82 select1 x1.gpo0 8.43e-19
C83 select0 x1.nSEL2 0.131913f
C84 x1.gpo1 a_5645_6637# 2.95e-20
C85 x5.A A5 4.07e-21
C86 x1.gno3 x1.gpo2 5.65242f
C87 x1.gno3 a_5645_6637# 0.003645f
C88 a_5671_6589# x1.gno1 3.11e-20
C89 x1.nSEL0 VDD 0.386805f
C90 x1.nSEL1 VDD 0.472688f
C91 A7 x1.gno1 0.006482f
C92 x1.nSEL0 a_5645_5493# 0.081627f
C93 A1 x1.gpo0 3.9665f
C94 x3.Z3 x1.nSEL2 4.15404f
C95 x1.nSEL1 a_5645_5493# 0.193944f
C96 A2 x1.nSEL2 0.011628f
C97 A3 VDD 1.61205f
C98 x1.gno1 x1.gno2 0.179257f
C99 select1 x1.gpo3 3.7e-19
C100 x1.gno0 select0 0.020289f
C101 a_5671_6589# x1.nSEL2 9.76e-20
C102 select2 VDD 3.46438f
C103 Z x3.Z3 5.48465f
C104 select2 a_5645_5493# 4.33e-19
C105 x1.gno1 A5 0.145599f
C106 x1.nSEL2 x1.gno2 1.63e-19
C107 A4 VDD 1.56602f
C108 A1 x1.gpo3 1.62e-19
C109 x1.gno0 x3.Z3 0.428132f
C110 A2 x1.gno0 0.135398f
C111 select1 x1.nSEL0 0.137595f
C112 select1 x1.nSEL1 0.275603f
C113 x1.gno1 a_5671_6037# 0.002395f
C114 m2_5776_5494# x1.nSEL0 3.43e-19
C115 x1.gpo2 select0 2.74e-19
C116 m2_5776_5494# x1.nSEL1 0.00815f
C117 select0 a_5645_6637# 0.279858f
C118 x5.A x1.gno1 0.429382f
C119 x3.Z3 A8 4.51511f
C120 VDD a_5645_6461# 0.171399f
C121 a_5645_7149# x1.gno1 7.58e-21
C122 x1.gno0 x1.gno2 0.089083f
C123 a_5699_5631# x1.gno1 8.86e-19
C124 select1 select2 0.289185f
C125 a_5645_5909# VDD 0.162117f
C126 x1.nSEL2 a_5671_6037# 1.08e-19
C127 x1.gpo1 VDD 3.26715f
C128 x1.gpo2 x3.Z3 0.358391f
C129 x1.gpo0 x1.gpo3 0.080341f
C130 x1.gno3 VDD 1.35568f
C131 A2 x1.gpo2 0.001569f
C132 m2_5776_5494# select2 4.4e-19
C133 a_5645_5909# a_5645_5493# 0.002207f
C134 A7 A8 2.08862f
C135 x5.A x1.nSEL2 4.05923f
C136 a_5645_6085# VDD 0.193284f
C137 A8 x1.gno2 0.006957f
C138 a_5671_6589# x1.gpo2 4.39e-19
C139 x1.gpo0 A6 0.12311f
C140 a_5699_7287# VDD 8.97e-19
C141 A1 select2 0.054741f
C142 a_5645_7149# x1.nSEL2 1.19e-19
C143 x1.gno0 A5 3.85224f
C144 a_5699_5631# x1.nSEL2 1.95e-19
C145 A7 x1.gpo2 4.00999f
C146 x1.nSEL0 x1.gpo0 6.21e-20
C147 Z x5.A 4.51604f
C148 x1.gno0 a_5671_6037# 1.22e-20
C149 x1.gpo2 x1.gno2 5.02054f
C150 x1.gpo0 x1.nSEL1 1.17e-19
C151 a_5645_6637# x1.gno2 0.004289f
C152 select1 a_5645_6461# 0.261734f
C153 x5.A x1.gno0 0.430802f
C154 A3 x1.gpo0 0.001407f
C155 select1 a_5645_5909# 0.03417f
C156 select1 x1.gpo1 3.1e-20
C157 x1.gpo3 A6 1.72e-19
C158 select1 x1.gno3 0.059776f
C159 x1.gno0 a_5699_5631# 0.001144f
C160 x1.gpo0 select2 5.94e-19
C161 x1.gpo2 A5 2.05e-19
C162 x1.gno1 x1.nSEL2 0.019435f
C163 select1 a_5645_6085# 0.254026f
C164 select1 a_5699_7287# 8.84e-19
C165 x1.gpo1 A1 0.002755f
C166 select0 VDD 1.13942f
C167 x1.gpo0 A4 0.002819f
C168 x1.gno3 A1 1.72e-19
C169 A3 x1.gpo3 0.00162f
C170 x5.A x1.gpo2 0.358718f
C171 Z x1.gno1 9.36e-20
C172 select0 a_5645_5493# 0.048888f
C173 x1.gpo3 select2 0.006992f
C174 x1.gno0 x1.gno1 0.146872f
C175 x1.nSEL0 x1.nSEL1 0.352716f
C176 x3.Z3 VDD 14.4075f
C177 A2 VDD 1.60691f
C178 x1.gpo0 a_5645_6461# 1.19e-20
C179 Z x1.nSEL2 0.833318f
C180 a_5645_5909# x1.gpo0 9.98e-19
C181 x1.gpo3 A4 3.96247f
C182 a_5671_6589# VDD 0.001496f
C183 x1.gpo1 x1.gpo0 0.101838f
C184 x1.gno3 x1.gpo0 0.066343f
C185 A7 VDD 1.61205f
C186 x1.gno0 x1.nSEL2 0.645006f
C187 x1.nSEL0 select2 0.131256f
C188 select2 x1.nSEL1 0.164995f
C189 A4 A6 7.47e-20
C190 select1 select0 1.85585f
C191 VDD x1.gno2 0.767412f
C192 x1.gpo2 x1.gno1 0.060968f
C193 m2_5776_5494# select0 0.130999f
C194 A3 select2 2.39e-19
C195 x1.gno1 a_5645_6637# 1.03e-19
C196 Z x1.gno0 4.27e-20
C197 x1.gpo1 x1.gpo3 0.069892f
C198 A1 select0 2.25e-21
C199 x1.gno3 x1.gpo3 5.58658f
C200 A3 A4 2.08862f
C201 A5 VDD 1.60179f
C202 x1.gpo2 x1.nSEL2 3.82e-20
C203 x1.gpo1 A6 4.01113f
C204 x1.nSEL2 a_5645_6637# 2.27e-19
C205 a_5699_7287# x1.gpo3 1e-19
C206 x1.nSEL0 a_5645_6461# 1.91e-20
C207 select2 A4 6.76e-20
C208 x1.gno3 A6 1.76e-19
C209 VDD a_5671_6037# 4.32e-19
C210 x1.nSEL1 a_5645_6461# 7.84e-19
C211 a_5645_5909# x1.nSEL0 0.03096f
C212 A2 A1 1.81909f
C213 a_5645_5909# x1.nSEL1 0.073392f
C214 x5.A VDD 14.1327f
C215 x1.nSEL0 x1.gno3 2.26e-20
C216 select1 x1.gno2 0.272271f
C217 Z x1.gpo2 2.44e-19
C218 a_5645_7149# VDD 0.217381f
C219 x1.nSEL0 a_5645_6085# 0.001174f
C220 x1.gpo0 select0 8.18e-19
C221 A3 x1.gpo1 0.1453f
C222 a_5699_5631# VDD 9.09e-19
C223 a_5645_6085# x1.nSEL1 0.041068f
C224 select2 a_5645_6461# 0.009143f
C225 A3 x1.gno3 0.16467f
C226 x1.gno0 x1.gpo2 0.076333f
C227 x1.gno0 a_5645_6637# 1.69e-20
C228 a_5645_5909# select2 8.66e-20
C229 a_5699_5631# a_5645_5493# 0.006584f
C230 A1 x1.gno2 2.84e-19
C231 x1.gpo1 select2 4.34e-19
C232 x1.gno3 select2 5.71e-20
C233 x1.gpo0 x3.Z3 0.354991f
C234 A2 x1.gpo0 0.124367f
C235 x1.gpo2 A8 0.161339f
C236 a_5645_6085# select2 1.67e-19
C237 x1.gpo1 A4 4.15e-19
C238 x1.gpo3 select0 0.001185f
C239 x1.gno3 A4 3.82666f
C240 x1.gno1 VDD 0.699246f
C241 A7 x1.gpo0 2.46e-21
C242 x1.gpo2 a_5645_6637# 4.69e-19
C243 x1.gno1 a_5645_5493# 0.039612f
C244 select1 a_5645_7149# 0.125445f
C245 x1.gpo0 x1.gno2 0.056456f
C246 x1.gpo3 x3.Z3 0.3315f
C247 x1.gpo1 a_5645_6461# 2.46e-19
C248 A2 x1.gpo3 1.55e-19
C249 x5.A A1 4.52065f
C250 x1.nSEL0 select0 0.325123f
C251 x1.gno3 a_5645_6461# 6.84e-19
C252 x1.nSEL1 select0 0.169954f
C253 VDD x1.nSEL2 3.6311f
C254 x3.Z3 A6 4.52053f
C255 a_5645_6085# a_5645_6461# 3.02e-19
C256 x1.gpo1 x1.gno3 0.062916f
C257 a_5645_5493# x1.nSEL2 0.001336f
C258 a_5645_5909# a_5645_6085# 0.185422f
C259 A7 x1.gpo3 0.00162f
C260 x1.gpo0 A5 4.0165f
C261 x1.gpo3 x1.gno2 0.072782f
C262 Z VDD 5.306779f
C263 select2 select0 0.446748f
C264 select1 x1.gno1 0.108644f
C265 x1.gno3 a_5699_7287# 0.001562f
C266 A7 A6 1.81997f
C267 A3 x3.Z3 1.64e-20
C268 x1.gno0 VDD 0.889132f
C269 x5.A x1.gpo0 0.35382f
C270 A6 x1.gno2 0.156179f
C271 a_5671_6589# x1.nSEL1 4.08e-19
C272 A3 A2 1.81997f
C273 x1.gno0 a_5645_5493# 0.128677f
C274 select2 x3.Z3 5.00334f
C275 A5 x1.gpo3 0.098584f
C276 A1 x1.gno1 0.13437f
C277 x1.nSEL0 x1.gno2 4.01e-20
C278 select1 x1.nSEL2 0.140519f
C279 x1.nSEL1 x1.gno2 0.012418f
C280 VDD A8 1.54289f
C281 m2_5776_5494# x1.nSEL2 4e-19
C282 A5 A6 1.81909f
C283 x3.Z3 A4 0.003925f
C284 A3 x1.gno2 3.78522f
C285 A2 A4 2.39e-19
C286 select0 a_5645_6461# 0.086353f
C287 x5.A x1.gpo3 0.278763f
C288 x1.gpo2 VDD 3.24607f
C289 A1 x1.nSEL2 0.566094f
C290 a_5645_5909# select0 0.246189f
C291 VDD a_5645_6637# 0.262163f
C292 select2 x1.gno2 0.00233f
C293 x1.gpo1 select0 4.71e-19
C294 a_5645_7149# x1.gpo3 2.98e-19
C295 x1.gno3 select0 0.218342f
C296 select1 x1.gno0 0.312176f
C297 x1.gpo0 x1.gno1 4.59887f
C298 x1.nSEL0 a_5671_6037# 2.51e-19
C299 x1.nSEL1 a_5671_6037# 9.57e-19
C300 a_5645_6085# select0 0.143958f
C301 A4 x1.gno2 0.007342f
C302 m2_5776_5494# x1.gno0 0.06935f
C303 a_5699_7287# select0 1.4e-19
C304 x1.gpo1 x3.Z3 0.350405f
C305 A5 select2 2.94e-19
C306 A2 x1.gpo1 3.95776f
C307 a_5671_6589# a_5645_6461# 0.004764f
C308 x1.gno3 x3.Z3 0.446539f
C309 A2 x1.gno3 1.76e-19
C310 A1 x1.gno0 4.31208f
C311 A3 x5.A 4.5214f
C312 x1.gpo0 x1.nSEL2 0.045168f
C313 a_5699_5631# x1.nSEL1 0.00175f
C314 x1.gno3 a_5671_6589# 3.22e-19
C315 A5 A4 1.27332f
C316 x1.gno1 x1.gpo3 0.068595f
C317 a_5645_6461# x1.gno2 0.104374f
C318 A7 x1.gpo1 0.145249f
C319 select1 x1.gpo2 0.003325f
C320 x5.A select2 5.67997f
C321 select1 a_5645_6637# 0.127717f
C322 A7 x1.gno3 0.180503f
C323 a_5645_5909# x1.gno2 6.68e-19
C324 x1.gpo1 x1.gno2 4.59188f
C325 x1.gno3 x1.gno2 0.195239f
C326 x1.gno1 A6 3.81297f
C327 Z x1.gpo0 2.38e-19
C328 x5.A A4 4.5151f
C329 a_5645_6085# x1.gno2 0.048646f
C330 A1 x1.gpo2 1.96e-19
C331 x1.gpo3 x1.nSEL2 1.12e-19
C332 x1.gno0 x1.gpo0 2.99937f
C333 a_5699_7287# x1.gno2 1.07e-20
C334 x1.nSEL0 x1.gno1 0.154394f
C335 x1.gno1 x1.nSEL1 0.209954f
C336 x1.gpo1 A5 0.001763f
C337 x1.gno3 A5 0.005885f
C338 A3 x1.gno1 0.007138f
C339 a_5645_5909# a_5671_6037# 0.004764f
C340 Z x1.gpo3 1.68e-19
C341 Z VSS 6.578722f
C342 A8 VSS 3.687544f
C343 A7 VSS 3.163578f
C344 A6 VSS 3.279698f
C345 A5 VSS 3.5005f
C346 A4 VSS 3.017403f
C347 A3 VSS 3.186499f
C348 A2 VSS 3.320398f
C349 A1 VSS 4.042872f
C350 select2 VSS 6.567346f
C351 select0 VSS 1.45124f
C352 select1 VSS 1.80202f
C353 VDD VSS 0.117673p
C354 m2_5776_5494# VSS 0.065655f $ **FLOATING
C355 x3.Z3 VSS 16.058199f
C356 x5.A VSS 12.524099f
C357 a_5699_5631# VSS 0.006505f
C358 a_5645_5493# VSS 0.266782f
C359 x1.nSEL0 VSS 0.650696f
C360 x1.gpo0 VSS 10.456742f
C361 x1.gno0 VSS 11.723553f
C362 a_5671_6037# VSS 0.004461f
C363 a_5645_5909# VSS 0.220868f
C364 x1.nSEL1 VSS 0.682637f
C365 x1.gpo1 VSS 10.05377f
C366 x1.gno1 VSS 7.03383f
C367 a_5645_6085# VSS 0.23458f
C368 x1.nSEL2 VSS 5.45531f
C369 x1.gpo2 VSS 3.19357f
C370 a_5671_6589# VSS 0.006801f
C371 x1.gno2 VSS 6.82653f
C372 a_5645_6461# VSS 0.232731f
C373 x1.gpo3 VSS 12.517524f
C374 a_5645_6637# VSS 0.249604f
C375 x1.gno3 VSS 13.497057f
C376 a_5699_7287# VSS 0.006583f
C377 a_5645_7149# VSS 0.307391f
C378 x1.gpo1.t3 VSS 0.018013f
C379 x1.gpo1.t2 VSS 0.018013f
C380 x1.gpo1.n0 VSS 0.042951f
C381 x1.gpo1.n1 VSS 0.084381f
C382 x1.gpo1.n2 VSS 0.026255f
C383 x1.gpo1.t5 VSS 0.911601f
C384 x1.gpo1.t7 VSS 0.937021f
C385 x1.gpo1.n3 VSS 3.3244f
C386 x1.gpo1.t4 VSS 0.911601f
C387 x1.gpo1.t6 VSS 0.937021f
C388 x1.gpo1.n4 VSS 3.3244f
C389 x1.gpo1.n5 VSS 1.96615f
C390 x1.gpo1.t1 VSS 0.027712f
C391 x1.gpo1.t0 VSS 0.027712f
C392 x1.gpo1.n6 VSS 0.057149f
C393 x1.gpo1.n7 VSS 0.119653f
C394 A8.t1 VSS 0.893325f
C395 A8.t0 VSS 0.512841f
C396 A8.n0 VSS 4.96695f
C397 A8.t3 VSS 0.924602f
C398 A8.t2 VSS 0.65407f
C399 A8.n1 VSS 5.0783f
C400 A8.n2 VSS 0.803255f
C401 A8.n3 VSS 0.258761f
C402 A6.t3 VSS 0.763965f
C403 A6.t2 VSS 0.438578f
C404 A6.n0 VSS 4.2477f
C405 A6.t0 VSS 0.790712f
C406 A6.t1 VSS 0.559356f
C407 A6.n1 VSS 4.34292f
C408 A6.n2 VSS 0.686937f
C409 A6.n3 VSS 0.222065f
C410 A3.t1 VSS 0.893857f
C411 A3.t0 VSS 0.513146f
C412 A3.n0 VSS 4.9699f
C413 A3.t3 VSS 0.925152f
C414 A3.t2 VSS 0.654459f
C415 A3.n1 VSS 5.08132f
C416 A3.n2 VSS 0.803733f
C417 A3.n3 VSS 0.264783f
C418 A7.t1 VSS 0.893857f
C419 A7.t0 VSS 0.513146f
C420 A7.n0 VSS 4.9699f
C421 A7.t2 VSS 0.925152f
C422 A7.t3 VSS 0.654459f
C423 A7.n1 VSS 5.08132f
C424 A7.n2 VSS 0.803733f
C425 A7.n3 VSS 0.264783f
C426 A4.t1 VSS 0.893325f
C427 A4.t0 VSS 0.512841f
C428 A4.n0 VSS 4.96695f
C429 A4.t2 VSS 0.924602f
C430 A4.t3 VSS 0.65407f
C431 A4.n1 VSS 5.0783f
C432 A4.n2 VSS 0.803255f
C433 A4.n3 VSS 0.258761f
C434 A2.t1 VSS 0.763965f
C435 A2.t2 VSS 0.438578f
C436 A2.n0 VSS 4.2477f
C437 A2.t0 VSS 0.790712f
C438 A2.t3 VSS 0.559356f
C439 A2.n1 VSS 4.34292f
C440 A2.n2 VSS 0.686937f
C441 A2.n3 VSS 0.222065f
C442 A1.t2 VSS 0.795131f
C443 A1.t3 VSS 0.45647f
C444 A1.n0 VSS 4.42098f
C445 A1.t0 VSS 0.82297f
C446 A1.t1 VSS 0.582175f
C447 A1.n1 VSS 4.52009f
C448 A1.n2 VSS 0.714961f
C449 A1.n3 VSS 0.223162f
C450 x1.gpo0.t3 VSS 0.01774f
C451 x1.gpo0.t2 VSS 0.01774f
C452 x1.gpo0.n0 VSS 0.0423f
C453 x1.gpo0.n1 VSS 0.083102f
C454 x1.gpo0.n2 VSS 0.025857f
C455 x1.gpo0.t6 VSS 0.897787f
C456 x1.gpo0.t7 VSS 0.922822f
C457 x1.gpo0.n3 VSS 3.26002f
C458 x1.gpo0.t4 VSS 0.897787f
C459 x1.gpo0.t5 VSS 0.922822f
C460 x1.gpo0.n4 VSS 3.29215f
C461 x1.gpo0.n5 VSS 1.7367f
C462 x1.gpo0.t1 VSS 0.027292f
C463 x1.gpo0.t0 VSS 0.027292f
C464 x1.gpo0.n6 VSS 0.056236f
C465 x1.gpo0.n7 VSS 0.120059f
C466 x1.gpo3.t2 VSS 0.01237f
C467 x1.gpo3.t3 VSS 0.01237f
C468 x1.gpo3.n0 VSS 0.029497f
C469 x1.gpo3.n1 VSS 0.056891f
C470 x1.gpo3.t6 VSS 0.626043f
C471 x1.gpo3.t4 VSS 0.643501f
C472 x1.gpo3.n2 VSS 2.2877f
C473 x1.gpo3.t5 VSS 0.626043f
C474 x1.gpo3.t7 VSS 0.643501f
C475 x1.gpo3.n3 VSS 2.2877f
C476 x1.gpo3.n4 VSS 2.68712f
C477 x1.gpo3.n5 VSS 0.0412f
C478 x1.gpo3.n6 VSS 0.01803f
C479 x1.gpo3.t0 VSS 0.019031f
C480 x1.gpo3.t1 VSS 0.019031f
C481 x1.gpo3.n7 VSS 0.041797f
C482 x1.gno3.t1 VSS 0.053338f
C483 x1.gno3.n0 VSS 0.061486f
C484 x1.gno3.t6 VSS 0.60277f
C485 x1.gno3.t9 VSS 0.588227f
C486 x1.gno3.n1 VSS 2.63915f
C487 x1.gno3.n2 VSS 1.63117f
C488 x1.gno3.t3 VSS 0.60277f
C489 x1.gno3.t5 VSS 0.588227f
C490 x1.gno3.n3 VSS 2.63915f
C491 x1.gno3.n4 VSS 2.31307f
C492 x1.gno3.t4 VSS 0.033483f
C493 x1.gno3.t2 VSS 0.019731f
C494 x1.gno3.t8 VSS 0.033483f
C495 x1.gno3.t7 VSS 0.019731f
C496 x1.gno3.n5 VSS 0.05618f
C497 x1.gno3.n6 VSS 0.083224f
C498 x1.gno3.n7 VSS 0.037258f
C499 x1.gno3.n8 VSS 0.301796f
C500 x1.gno3.t0 VSS 0.13622f
C501 x1.gno3.n9 VSS 0.024501f
C502 x1.gno3.n10 VSS 0.027448f
C503 A5.t3 VSS 0.770284f
C504 A5.t2 VSS 0.442205f
C505 A5.n0 VSS 4.28283f
C506 A5.t0 VSS 0.797252f
C507 A5.t1 VSS 0.563982f
C508 A5.n1 VSS 4.37884f
C509 A5.n2 VSS 0.692619f
C510 A5.n3 VSS 0.216188f
C511 x1.gno0.n0 VSS 1.21068f
C512 x1.gno0.t1 VSS 0.038064f
C513 x1.gno0.n1 VSS 0.043923f
C514 x1.gno0.t9 VSS 0.430161f
C515 x1.gno0.t7 VSS 0.419783f
C516 x1.gno0.n2 VSS 1.8834f
C517 x1.gno0.t2 VSS 0.430161f
C518 x1.gno0.t3 VSS 0.419783f
C519 x1.gno0.n3 VSS 1.8834f
C520 x1.gno0.n4 VSS 0.892351f
C521 x1.gno0.n5 VSS 0.304041f
C522 x1.gno0.t8 VSS 0.023895f
C523 x1.gno0.t5 VSS 0.014081f
C524 x1.gno0.t6 VSS 0.023895f
C525 x1.gno0.t4 VSS 0.014081f
C526 x1.gno0.n6 VSS 0.040092f
C527 x1.gno0.n7 VSS 0.059217f
C528 x1.gno0.n8 VSS 0.057595f
C529 x1.gno0.n9 VSS 0.1251f
C530 x1.gno0.t0 VSS 0.097212f
C531 x1.gno0.n10 VSS 0.017485f
C532 x1.gno0.n11 VSS 0.019588f
C533 VDD.n0 VSS 0.078152f
C534 VDD.n1 VSS 0.253693f
C535 VDD.n2 VSS 0.122926f
C536 VDD.n3 VSS 0.122926f
C537 VDD.n4 VSS 0.122525f
C538 VDD.n5 VSS 0.169863f
C539 VDD.n6 VSS 0.547624f
C540 VDD.t1 VSS 0.790353f
C541 VDD.n7 VSS 0.763087f
C542 VDD.t0 VSS 0.790353f
C543 VDD.n8 VSS 0.547624f
C544 VDD.n9 VSS 0.004814f
C545 VDD.n10 VSS 0.134493f
C546 VDD.n11 VSS 0.040318f
C547 VDD.n12 VSS 0.138067f
C548 VDD.n13 VSS 0.057005f
C549 VDD.n14 VSS 0.253704f
C550 VDD.n15 VSS 0.122531f
C551 VDD.n16 VSS 1.03197f
C552 VDD.n17 VSS 1.03197f
C553 VDD.n18 VSS 0.169845f
C554 VDD.n19 VSS 0.124397f
C555 VDD.t7 VSS 1.37216f
C556 VDD.n22 VSS 0.124397f
C557 VDD.n23 VSS 5.27e-19
C558 VDD.n24 VSS 0.07554f
C559 VDD.n25 VSS 0.013735f
C560 VDD.n26 VSS 0.149327f
C561 VDD.n27 VSS 0.079843f
C562 VDD.n28 VSS 0.162134f
C563 VDD.n29 VSS 0.188097f
C564 VDD.n30 VSS 0.253704f
C565 VDD.n31 VSS 0.004119f
C566 VDD.n32 VSS 0.169845f
C567 VDD.n33 VSS 0.124397f
C568 VDD.t77 VSS 1.37216f
C569 VDD.n35 VSS 1.03197f
C570 VDD.n36 VSS 0.124397f
C571 VDD.n38 VSS 1.03197f
C572 VDD.n39 VSS 0.122531f
C573 VDD.n40 VSS 0.009862f
C574 VDD.n41 VSS 0.075465f
C575 VDD.n42 VSS 0.013861f
C576 VDD.n43 VSS 0.149327f
C577 VDD.n44 VSS 0.079211f
C578 VDD.n45 VSS 0.128376f
C579 VDD.n46 VSS 0.184404f
C580 VDD.n47 VSS 0.253704f
C581 VDD.n48 VSS 0.00437f
C582 VDD.n49 VSS 0.169845f
C583 VDD.n50 VSS 0.124397f
C584 VDD.t6 VSS 1.37216f
C585 VDD.n52 VSS 1.03197f
C586 VDD.n53 VSS 0.124397f
C587 VDD.n55 VSS 1.03197f
C588 VDD.n56 VSS 0.122531f
C589 VDD.n57 VSS 0.009878f
C590 VDD.n58 VSS 0.075214f
C591 VDD.n59 VSS 0.013861f
C592 VDD.n60 VSS 0.149327f
C593 VDD.n61 VSS 0.079211f
C594 VDD.n62 VSS 0.125941f
C595 VDD.n63 VSS 0.167914f
C596 VDD.n64 VSS 0.010164f
C597 VDD.n65 VSS 0.00773f
C598 VDD.t39 VSS 0.015599f
C599 VDD.n66 VSS 0.015344f
C600 VDD.t13 VSS 0.001675f
C601 VDD.t55 VSS 0.002544f
C602 VDD.n67 VSS 0.004395f
C603 VDD.t37 VSS 0.015899f
C604 VDD.t76 VSS 0.015599f
C605 VDD.n68 VSS 0.014858f
C606 VDD.n69 VSS 0.00773f
C607 VDD.n70 VSS 0.006997f
C608 VDD.t43 VSS 0.002296f
C609 VDD.n71 VSS 0.006515f
C610 VDD.t35 VSS 0.009437f
C611 VDD.n72 VSS 0.008687f
C612 VDD.n73 VSS 0.007753f
C613 VDD.t9 VSS 0.015603f
C614 VDD.n74 VSS 0.001276f
C615 VDD.t51 VSS 0.00669f
C616 VDD.t64 VSS 0.011043f
C617 VDD.n75 VSS 0.010887f
C618 VDD.n76 VSS 0.013048f
C619 VDD.t79 VSS 0.046088f
C620 VDD.n77 VSS 0.041686f
C621 VDD.t41 VSS 0.00125f
C622 VDD.t47 VSS 0.003352f
C623 VDD.n78 VSS 0.0153f
C624 VDD.t65 VSS 0.011043f
C625 VDD.n79 VSS 0.008081f
C626 VDD.n80 VSS 0.030158f
C627 VDD.n81 VSS 0.023827f
C628 VDD.n82 VSS 0.030949f
C629 VDD.n83 VSS 0.01787f
C630 VDD.n84 VSS 0.013048f
C631 VDD.n85 VSS 0.009786f
C632 VDD.n86 VSS 0.006143f
C633 VDD.n87 VSS 0.019352f
C634 VDD.n88 VSS 0.030339f
C635 VDD.t44 VSS 0.031357f
C636 VDD.n89 VSS 0.002361f
C637 VDD.n90 VSS 0.002411f
C638 VDD.n91 VSS 0.009786f
C639 VDD.n92 VSS 0.003014f
C640 VDD.t33 VSS 0.015814f
C641 VDD.n93 VSS 0.012977f
C642 VDD.n94 VSS 0.00773f
C643 VDD.t80 VSS 0.046088f
C644 VDD.n95 VSS 0.011488f
C645 VDD.n96 VSS 0.00773f
C646 VDD.t3 VSS 0.00125f
C647 VDD.t62 VSS 0.003352f
C648 VDD.n97 VSS 0.0153f
C649 VDD.t82 VSS 0.046088f
C650 VDD.t17 VSS 0.00669f
C651 VDD.n98 VSS 0.020658f
C652 VDD.n99 VSS 0.011843f
C653 VDD.n100 VSS 0.006143f
C654 VDD.t67 VSS 0.011043f
C655 VDD.n101 VSS 0.010887f
C656 VDD.n102 VSS 0.041686f
C657 VDD.n103 VSS 0.01787f
C658 VDD.n104 VSS 0.030949f
C659 VDD.t68 VSS 0.011043f
C660 VDD.t49 VSS 0.015815f
C661 VDD.n105 VSS 0.004468f
C662 VDD.n106 VSS 0.005319f
C663 VDD.t16 VSS 0.063133f
C664 VDD.t61 VSS 0.061042f
C665 VDD.t66 VSS 0.045154f
C666 VDD.t2 VSS 0.064805f
C667 VDD.t23 VSS 0.063133f
C668 VDD.t10 VSS 0.071913f
C669 VDD.t56 VSS 0.052262f
C670 VDD.t20 VSS 0.028013f
C671 VDD.t32 VSS 0.012961f
C672 VDD.t48 VSS 0.045572f
C673 VDD.n107 VSS 0.059469f
C674 VDD.n108 VSS 0.041241f
C675 VDD.n109 VSS 0.012122f
C676 VDD.n110 VSS 0.01945f
C677 VDD.n111 VSS 0.023827f
C678 VDD.n112 VSS 0.008084f
C679 VDD.n113 VSS 0.064395f
C680 VDD.n114 VSS 0.087594f
C681 VDD.t73 VSS 0.011043f
C682 VDD.n115 VSS 0.021596f
C683 VDD.n116 VSS 0.041686f
C684 VDD.n117 VSS 0.025689f
C685 VDD.t74 VSS 0.011043f
C686 VDD.t27 VSS 0.015891f
C687 VDD.n118 VSS 0.018568f
C688 VDD.t72 VSS 0.142033f
C689 VDD.t69 VSS 0.087258f
C690 VDD.t52 VSS 0.035804f
C691 VDD.t58 VSS 0.049557f
C692 VDD.t14 VSS 0.035804f
C693 VDD.t18 VSS 0.049557f
C694 VDD.t29 VSS 0.035804f
C695 VDD.t26 VSS 0.053589f
C696 VDD.n119 VSS 0.058661f
C697 VDD.n120 VSS 0.00773f
C698 VDD.n121 VSS 0.003365f
C699 VDD.t19 VSS 0.015891f
C700 VDD.n122 VSS 0.003365f
C701 VDD.t59 VSS 0.015891f
C702 VDD.n123 VSS 0.227132f
C703 VDD.n124 VSS 0.013294f
C704 VDD.n125 VSS 0.008081f
C705 VDD.t81 VSS 0.046809f
C706 VDD.t70 VSS 0.011043f
C707 VDD.n126 VSS 0.04634f
C708 VDD.n127 VSS 0.023029f
C709 VDD.t71 VSS 0.011043f
C710 VDD.n128 VSS 0.030158f
C711 VDD.n129 VSS 0.027736f
C712 VDD.n130 VSS 0.017403f
C713 VDD.n131 VSS 0.013581f
C714 VDD.n132 VSS 0.013243f
C715 VDD.t53 VSS 0.015899f
C716 VDD.n133 VSS 0.020008f
C717 VDD.n134 VSS 0.00773f
C718 VDD.n135 VSS 0.013048f
C719 VDD.n136 VSS 0.009786f
C720 VDD.n137 VSS 0.018769f
C721 VDD.t15 VSS 0.015899f
C722 VDD.n138 VSS 0.02031f
C723 VDD.n139 VSS 0.00773f
C724 VDD.n140 VSS 0.013048f
C725 VDD.n141 VSS 0.009786f
C726 VDD.n142 VSS 0.018769f
C727 VDD.t30 VSS 0.015899f
C728 VDD.n143 VSS 0.02031f
C729 VDD.n144 VSS 0.003365f
C730 VDD.n145 VSS 0.013048f
C731 VDD.n146 VSS 0.009786f
C732 VDD.n147 VSS 0.004964f
C733 VDD.n148 VSS 0.027117f
C734 VDD.n149 VSS 0.012122f
C735 VDD.n150 VSS 0.01945f
C736 VDD.n151 VSS 0.033134f
C737 VDD.n152 VSS 0.006595f
C738 VDD.n153 VSS 0.059927f
C739 VDD.n154 VSS 0.058109f
C740 VDD.n155 VSS 0.001347f
C741 VDD.t21 VSS 0.001675f
C742 VDD.t57 VSS 0.002544f
C743 VDD.n156 VSS 0.004395f
C744 VDD.n157 VSS 0.029498f
C745 VDD.t25 VSS 0.015891f
C746 VDD.n158 VSS 0.018518f
C747 VDD.t11 VSS 0.005236f
C748 VDD.t45 VSS 0.013917f
C749 VDD.n159 VSS 0.007895f
C750 VDD.t24 VSS 0.015603f
C751 VDD.n160 VSS 0.016462f
C752 VDD.n161 VSS 0.021174f
C753 VDD.n162 VSS 0.002788f
C754 VDD.n163 VSS 0.013048f
C755 VDD.n164 VSS 0.00773f
C756 VDD.n165 VSS 0.004468f
C757 VDD.n166 VSS 0.004964f
C758 VDD.n167 VSS 0.026569f
C759 VDD.n168 VSS 0.072449f
C760 VDD.t12 VSS 0.013797f
C761 VDD.t38 VSS 0.035956f
C762 VDD.t36 VSS 0.040137f
C763 VDD.t54 VSS 0.028013f
C764 VDD.t42 VSS 0.052262f
C765 VDD.t75 VSS 0.073585f
C766 VDD.t8 VSS 0.035956f
C767 VDD.t34 VSS 0.028013f
C768 VDD.t40 VSS 0.064805f
C769 VDD.t63 VSS 0.045154f
C770 VDD.t46 VSS 0.061042f
C771 VDD.t50 VSS 0.063133f
C772 VDD.n169 VSS 0.042993f
C773 VDD.n170 VSS 0.01249f
C774 VDD.n171 VSS 0.008891f
C775 VDD.n172 VSS 0.002361f
C776 VDD.n173 VSS 0.017322f
C777 VDD.n174 VSS 0.006606f
C778 VDD.n175 VSS 0.013048f
C779 VDD.n176 VSS 0.009786f
C780 VDD.n177 VSS 0.005817f
C781 VDD.n178 VSS 0.019774f
C782 VDD.n179 VSS 0.014151f
C783 VDD.n180 VSS 0.009006f
C784 VDD.n181 VSS 0.025467f
C785 VDD.n182 VSS 0.279991f
C786 VDD.n183 VSS 0.651519f
C787 VDD.n184 VSS 0.253704f
C788 VDD.n185 VSS 0.051921f
C789 VDD.n186 VSS 0.122531f
C790 VDD.n187 VSS 1.03197f
C791 VDD.n188 VSS 1.03197f
C792 VDD.n189 VSS 0.169845f
C793 VDD.n190 VSS 0.124397f
C794 VDD.t60 VSS 1.37216f
C795 VDD.n193 VSS 0.124397f
C796 VDD.n194 VSS 4.77e-19
C797 VDD.n195 VSS 0.07554f
C798 VDD.n196 VSS 0.013785f
C799 VDD.n197 VSS 0.149327f
C800 VDD.n198 VSS 0.079793f
C801 VDD.n199 VSS 0.15219f
C802 VDD.n200 VSS 0.253704f
C803 VDD.n201 VSS 0.00437f
C804 VDD.n202 VSS 0.169845f
C805 VDD.n203 VSS 0.124397f
C806 VDD.t5 VSS 1.37216f
C807 VDD.n205 VSS 1.03197f
C808 VDD.n206 VSS 0.124397f
C809 VDD.n208 VSS 1.03197f
C810 VDD.n209 VSS 0.122531f
C811 VDD.n210 VSS 0.075214f
C812 VDD.n211 VSS 0.013861f
C813 VDD.n212 VSS 0.149327f
C814 VDD.n213 VSS 0.079211f
C815 VDD.n214 VSS 0.153404f
C816 VDD.n215 VSS 0.196603f
C817 VDD.n216 VSS 0.116414f
C818 VDD.n217 VSS 0.075465f
C819 VDD.n218 VSS 0.013861f
C820 VDD.n219 VSS 1.03197f
C821 VDD.n220 VSS 1.03197f
C822 VDD.n221 VSS 0.122531f
C823 VDD.n222 VSS 0.079211f
C824 VDD.n223 VSS 0.149327f
C825 VDD.n224 VSS 0.253704f
C826 VDD.n225 VSS 0.169845f
C827 VDD.n226 VSS 0.124397f
C828 VDD.t78 VSS 1.37216f
C829 VDD.n229 VSS 0.124397f
C830 VDD.n230 VSS 0.004119f
C831 VDD.n231 VSS 0.009862f
C832 VDD.n232 VSS 0.235683f
C833 VDD.n233 VSS 0.097082f
C834 VDD.n234 VSS 5.27e-19
C835 VDD.n235 VSS 0.079843f
C836 VDD.n236 VSS 0.149327f
C837 VDD.n237 VSS 0.169845f
C838 VDD.n238 VSS 0.124397f
C839 VDD.t22 VSS 1.37216f
C840 VDD.n239 VSS 0.253704f
C841 VDD.n241 VSS 1.03197f
C842 VDD.n242 VSS 0.124397f
C843 VDD.n244 VSS 1.03197f
C844 VDD.n245 VSS 0.122531f
C845 VDD.n246 VSS 0.07554f
C846 VDD.n247 VSS 0.013735f
C847 VDD.n248 VSS 0.013528f
C848 VDD.n249 VSS 0.191035f
C849 VDD.n250 VSS 0.253704f
C850 VDD.n251 VSS 0.07554f
C851 VDD.n252 VSS 1.03197f
C852 VDD.n253 VSS 1.03197f
C853 VDD.n254 VSS 0.122531f
C854 VDD.n255 VSS 0.169845f
C855 VDD.n256 VSS 0.124397f
C856 VDD.t4 VSS 1.37216f
C857 VDD.n259 VSS 0.124397f
C858 VDD.n260 VSS 4.77e-19
C859 VDD.n261 VSS 0.013492f
C860 VDD.n262 VSS 0.013785f
C861 VDD.n263 VSS 0.149327f
C862 VDD.n264 VSS 0.079793f
C863 VDD.n265 VSS 0.142932f
C864 VDD.n266 VSS 0.154755f
C865 VDD.n267 VSS 0.390936f
C866 VDD.n268 VSS 0.078152f
C867 VDD.n269 VSS 0.253693f
C868 VDD.n270 VSS 0.122926f
C869 VDD.n271 VSS 0.122926f
C870 VDD.n272 VSS 0.122525f
C871 VDD.n273 VSS 0.169863f
C872 VDD.n274 VSS 0.547624f
C873 VDD.t28 VSS 0.790353f
C874 VDD.n275 VSS 0.763087f
C875 VDD.t31 VSS 0.790353f
C876 VDD.n276 VSS 0.547624f
C877 VDD.n277 VSS 0.004814f
C878 VDD.n278 VSS 0.134493f
C879 VDD.n279 VSS 0.040288f
C880 VDD.n280 VSS 0.072753f
C881 Z.t5 VSS 0.434416f
C882 Z.n0 VSS 0.540283f
C883 Z.t4 VSS 0.446377f
C884 Z.t1 VSS 0.336375f
C885 Z.n1 VSS 2.25255f
C886 Z.n2 VSS 0.762169f
C887 Z.t0 VSS 0.329756f
C888 Z.n3 VSS 0.492384f
C889 Z.n4 VSS 0.648657f
C890 Z.n5 VSS 0.805956f
C891 Z.t2 VSS 0.434416f
C892 Z.n6 VSS 0.540283f
C893 Z.t3 VSS 0.446377f
C894 Z.t6 VSS 0.336375f
C895 Z.n7 VSS 2.25255f
C896 Z.n8 VSS 0.762169f
C897 Z.t7 VSS 0.329756f
C898 Z.n9 VSS 0.492384f
C899 Z.n10 VSS 0.664311f
C900 Z.n11 VSS 0.690962f
C901 select2.t3 VSS 0.587307f
C902 select2.t4 VSS 0.573137f
C903 select2.n0 VSS 2.59595f
C904 select2.t1 VSS 0.032624f
C905 select2.t7 VSS 0.019225f
C906 select2.t6 VSS 0.032624f
C907 select2.t5 VSS 0.019225f
C908 select2.n1 VSS 0.054739f
C909 select2.n2 VSS 0.080926f
C910 select2.n3 VSS 0.080283f
C911 select2.n4 VSS 1.30573f
C912 select2.t2 VSS 0.689904f
C913 select2.t0 VSS 0.709143f
C914 select2.n5 VSS 2.58376f
C915 select2.n6 VSS 1.7346f
C916 select2.n7 VSS 4.54427f
C917 select2.n8 VSS 1.56778f
C918 select2.n9 VSS 0.081638f
C919 select1.t6 VSS 0.031316f
C920 select1.t5 VSS 0.018454f
C921 select1.t3 VSS 0.031316f
C922 select1.t1 VSS 0.018454f
C923 select1.n0 VSS 0.052544f
C924 select1.n1 VSS 0.077632f
C925 select1.n2 VSS 0.047269f
C926 select1.t9 VSS 0.014491f
C927 select1.t7 VSS 0.03056f
C928 select1.n3 VSS 0.109737f
C929 select1.n4 VSS 0.021277f
C930 select1.n5 VSS 0.018327f
C931 select1.t4 VSS 0.022078f
C932 select1.t2 VSS 0.015172f
C933 select1.n6 VSS 0.064155f
C934 select1.n7 VSS 0.014778f
C935 select1.n8 VSS 0.105859f
C936 select1.n9 VSS 0.383423f
C937 select1.t8 VSS 0.026898f
C938 select1.t0 VSS 0.018264f
C939 select1.n10 VSS 0.063549f
C940 select1.n11 VSS 0.015211f
C941 select1.n12 VSS 0.098666f
C942 select1.n13 VSS 0.442567f
C943 select1.n14 VSS 0.578172f
.ends

