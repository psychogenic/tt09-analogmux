** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/mux4onehot_b.sch
.subckt mux4onehot_b select1 VDD VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 select0 select2 nselect2
*.PININFO select0:I select1:I select2:I A1:B A2:B A3:B A4:B Z1:B Z2:B Z3:B Z4:B nselect2:O VDD:I VSS:I
x2 gpo2 gpo1 gpo0 VDD gpo3 VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 gno2 gno1 gno0 gno3 passgatex4
x1 gpo0 gno0 gno1 gpo1 select0 select1 gno2 gpo2 nselect2 select2 gno3 gpo3 VDD VSS passgatesCtrlManual
.ends

* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym # of pins=18
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatex4.sch
.subckt passgatex4 GP3 GP2 GP1 VDD GP4 VSS A3 A2 A1 Z3 Z1 Z2 A4 Z4 GN3 GN2 GN1 GN4
*.PININFO VDD:I VSS:I GP1:I GN1:I A1:B Z1:B GP2:I GN2:I A2:B Z2:B GP3:I GN3:I A3:B Z3:B GP4:I GN4:I A4:B Z4:B
x1 Z1 A1 GP1 GN1 VSS VDD passgate
x2 Z2 A2 GP2 GN2 VSS VDD passgate
x3 Z3 A3 GP3 GN3 VSS VDD passgate
x4 Z4 A4 GP4 GN4 VSS VDD passgate
.ends


* expanding   symbol:  /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym # of pins=14
** sym_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sym
** sch_path: /home/ttuser/vmswap/tt09-analogmux/xschem/passgatesCtrlManual.sch
.subckt passgatesCtrlManual gpo0 gno0 gno1 gpo1 SEL0 SEL1 gno2 gpo2 nSEL2 SEL2 gno3 gpo3 VDD VSS
*.PININFO SEL0:I SEL1:I SEL2:I gno0:O gpo0:O gno1:O gpo1:O gno2:O gpo2:O gno3:O gpo3:O nSEL2:O VDD:I VSS:I
x1 SEL0 VSS VSS VDD VDD nSEL0 sky130_fd_sc_hd__inv_2
x2 SEL1 VSS VSS VDD VDD nSEL1 sky130_fd_sc_hd__inv_2
x7 nSEL0 nSEL1 VSS VSS VDD VDD gno0 sky130_fd_sc_hd__and2_1
x10 SEL1 SEL0 VSS VSS VDD VDD gno3 sky130_fd_sc_hd__and2_1
x11 gno0 VSS VSS VDD VDD gpo0 sky130_fd_sc_hd__inv_2
x12 gno1 VSS VSS VDD VDD gpo1 sky130_fd_sc_hd__inv_2
x13 gno2 VSS VSS VDD VDD gpo2 sky130_fd_sc_hd__inv_2
x14 gno3 VSS VSS VDD VDD gpo3 sky130_fd_sc_hd__inv_2
x15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x16 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x17 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
x8 SEL1 SEL0 VSS VSS VDD VDD gno1 sky130_fd_sc_hd__and2b_1
x9 SEL0 SEL1 VSS VSS VDD VDD gno2 sky130_fd_sc_hd__and2b_1
x18 SEL2 VSS VSS VDD VDD nSEL2 sky130_fd_sc_hd__inv_2
x19 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
.ends


* expanding   symbol:  /home/ttuser/tt08-wowa2/xschem/passgate.sym # of pins=6
** sym_path: /home/ttuser/tt08-wowa2/xschem/passgate.sym
** sch_path: /home/ttuser/tt08-wowa2/xschem/passgate.sch
.subckt passgate Z A GP GN VSSBPIN VCCBPIN
*.PININFO GN:I VCCBPIN:I VSSBPIN:I GP:I A:B Z:B
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 m=2
XM3 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 m=2
.ends

.end
