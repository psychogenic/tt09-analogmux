magic
tech sky130A
magscale 1 2
timestamp 1728254216
<< metal1 >>
rect 4142 774 4194 776
rect 4138 770 4198 774
rect 4138 718 4142 770
rect 4194 718 4198 770
rect 3898 643 3950 648
rect 3895 642 3953 643
rect 3895 586 3898 642
rect 3950 586 3953 642
rect 3088 502 3140 506
rect 3084 500 3144 502
rect 3084 444 3088 500
rect 3140 444 3144 500
rect 2858 367 2910 372
rect 2856 366 2913 367
rect 2856 310 2858 366
rect 2910 310 2913 366
rect 2040 238 2092 242
rect 2038 236 2094 238
rect 2038 184 2040 236
rect 2092 184 2094 236
rect 1804 116 1856 120
rect 1801 114 1860 116
rect 1801 58 1804 114
rect 1856 58 1860 114
rect 998 14 1050 20
rect 1050 -42 1051 13
rect 754 -88 806 -84
rect 752 -90 808 -88
rect 752 -142 754 -90
rect 806 -142 808 -90
rect 452 -422 652 -222
rect 752 -384 808 -142
rect 998 -344 1051 -42
rect 1508 -424 1708 -224
rect 1801 -387 1860 58
rect 2038 -358 2094 184
rect 2550 -428 2750 -228
rect 2856 -382 2913 310
rect 3084 -380 3144 444
rect 3584 -412 3778 -212
rect 3895 -369 3953 586
rect 4138 -324 4198 718
rect 426 -5154 622 -4796
rect 1492 -5154 1694 -4956
rect 2562 -5192 2764 -4994
rect 3622 -5194 3820 -4792
<< via1 >>
rect 4142 718 4194 770
rect 3898 586 3950 642
rect 3088 444 3140 500
rect 2858 310 2910 366
rect 2040 184 2092 236
rect 1804 58 1856 114
rect 998 -42 1050 14
rect 754 -142 806 -90
<< metal2 >>
rect -3508 772 -3075 773
rect -3562 770 -3075 772
rect -3562 718 4142 770
rect 4194 718 4200 770
rect -3562 714 -3075 718
rect -3562 -574 -3506 714
rect -2760 640 3898 642
rect -3264 586 3898 640
rect 3950 586 3956 642
rect -3264 584 -2564 586
rect -3264 -568 -3208 584
rect -2620 500 -2184 502
rect -2620 446 3088 500
rect -2620 -584 -2564 446
rect -2330 444 3088 446
rect 3140 444 3146 500
rect -1978 310 2858 366
rect 2910 310 2916 366
rect -1976 308 -1750 310
rect -1976 -492 -1920 308
rect -1332 238 -1276 240
rect -1332 236 2096 238
rect -1332 184 2040 236
rect 2092 184 2098 236
rect -1332 182 2096 184
rect -1332 -550 -1276 182
rect -686 58 1804 114
rect 1856 58 1862 114
rect -686 -574 -630 58
rect -40 -42 998 14
rect 1050 -42 1056 14
rect -40 -580 16 -42
rect 290 -90 806 -89
rect 290 -142 754 -90
rect 806 -142 812 -90
rect 290 -146 806 -142
rect 290 -586 347 -146
rect -112 -4896 74 -4894
rect 188 -4896 848 -4894
rect -112 -4904 848 -4896
rect 74 -5058 848 -4904
rect -112 -5068 848 -5058
rect -104 -5094 848 -5068
rect -104 -5096 630 -5094
rect -756 -5316 -584 -5158
rect -288 -5302 -116 -5144
<< via2 >>
rect -112 -5058 74 -4904
<< metal3 >>
rect -1145 -208 1434 -10
rect -1145 -783 -947 -208
rect 1236 -422 1434 -208
rect -2299 -808 -659 -783
rect -2299 -952 -2272 -808
rect -1992 -952 -974 -808
rect -694 -952 -659 -808
rect -2299 -981 -659 -952
rect -2992 -4628 110 -4574
rect -2992 -4634 -1642 -4628
rect -2992 -4842 -2968 -4634
rect -2662 -4836 -1642 -4634
rect -1336 -4634 110 -4628
rect -1336 -4836 -334 -4634
rect -2662 -4842 -334 -4836
rect -28 -4714 110 -4634
rect -28 -4842 114 -4714
rect -2992 -4896 114 -4842
rect -124 -4904 114 -4896
rect -124 -5058 -112 -4904
rect 74 -5058 114 -4904
rect -124 -5086 114 -5058
<< via3 >>
rect -2272 -952 -1992 -808
rect -974 -952 -694 -808
rect -2968 -4842 -2662 -4634
rect -1642 -4836 -1336 -4628
rect -334 -4842 -28 -4634
<< metal4 >>
rect -2304 -807 -1992 -792
rect -2304 -808 -1991 -807
rect -2304 -952 -2272 -808
rect -1992 -952 -1991 -808
rect -2304 -953 -1991 -952
rect -988 -808 -676 -806
rect -988 -952 -974 -808
rect -694 -952 -676 -808
rect -2304 -1176 -1992 -953
rect -988 -1190 -676 -952
rect -2968 -4633 -2648 -4145
rect -2969 -4634 -2648 -4633
rect -2969 -4842 -2968 -4634
rect -2662 -4842 -2648 -4634
rect -2969 -4843 -2648 -4842
rect -2968 -4858 -2648 -4843
rect -1648 -4628 -1328 -4145
rect -1648 -4836 -1642 -4628
rect -1336 -4836 -1328 -4628
rect -328 -4633 -8 -4145
rect -1648 -4844 -1328 -4836
rect -335 -4634 -8 -4633
rect -335 -4842 -334 -4634
rect -28 -4842 -8 -4634
rect -335 -4843 -8 -4842
rect -328 -4844 -8 -4843
use passgatesCtrl  passgatesCtrl_0
timestamp 1728249049
transform -1 0 1138 0 -1 1025
box 784 1432 4700 6262
use passgatex4  passgatex4_0
timestamp 1728165396
transform 1 0 -10990 0 1 -4896
box 11366 -356 15589 4682
<< labels >>
flabel metal1 452 -422 652 -222 0 FreeSans 1600 0 0 0 A1
port 3 nsew
flabel metal1 1508 -424 1708 -224 0 FreeSans 1600 0 0 0 A2
port 4 nsew
flabel metal1 2552 -428 2752 -228 0 FreeSans 1600 0 0 0 A3
port 5 nsew
flabel metal1 1492 -5154 1692 -4954 0 FreeSans 1600 0 0 0 Z2
port 8 nsew
flabel metal1 2562 -5190 2762 -4990 0 FreeSans 1600 0 0 0 Z3
port 9 nsew
flabel metal1 424 -5158 624 -4794 0 FreeSans 1600 0 0 0 Z1
port 7 nsew
flabel metal2 -288 -5302 -116 -5144 0 FreeSans 1600 0 0 0 select0
port 1 nsew
flabel metal2 -756 -5316 -584 -5158 0 FreeSans 1600 0 0 0 select1
port 2 nsew
flabel metal3 -336 -4848 -32 -4636 0 FreeSans 1600 0 0 0 VDD
port 11 nsew
flabel metal3 -1138 -202 -906 -20 0 FreeSans 1600 0 0 0 VSS
port 12 nsew
flabel metal1 3584 -412 3778 -212 0 FreeSans 1600 0 0 0 A4
port 6 nsew
flabel metal1 3622 -5186 3816 -4986 0 FreeSans 1600 0 0 0 Z4
port 10 nsew
<< end >>
