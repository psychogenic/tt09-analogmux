* NGSPICE file created from mux4onehot_parax.ext - technology: sky130A

.subckt mux4onehot_parax select0 select1 A1 Z4 Z3 Z2 A2 Z1 A4 A3 VSS VDD
X0 VSS.t97 passgatesCtrl_0.net2.t2 a_n597_n2040# VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VSS.t140 VDD.t176 VSS.t139 VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2 VDD.t66 VSS.t177 VDD.t65 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3 VSS.t142 VDD.t177 VSS.t141 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4 VDD.t64 VSS.t178 VDD.t63 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5 VSS.t41 a_n1361_n1429# passgatex4_0.GN3 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6 a_n1361_n1429# passgatesCtrl_0.net5 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7 VSS.t99 select1.t0 a_n2480_n4368# VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VSS.t157 VDD.t178 VSS.t156 VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X9 VSS.t53 a_n2189_n1429# passgatex4_0.GP3 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X10 a_n2189_n1429# passgatesCtrl_0.net9 VDD.t134 VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11 passgatesCtrl_0.net6 a_n2975_n2192# VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X12 a_n1084_n4216# a_n988_n4394# VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X13 VSS.t160 VDD.t179 VSS.t159 VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X14 VDD.t117 passgatesCtrl_0.net2.t3 a_n2161_n4368# VDD.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 VDD.t138 a_n715_n3850# passgatesCtrl_0._04_ VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X16 VDD.t62 VSS.t179 VDD.t61 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X17 a_n1913_n1429# passgatesCtrl_0.net10.t3 VSS.t68 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X18 a_n1173_n2218# a_n1003_n2040# a_n1045_n1942# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X19 passgatex4_0.GN2 a_n951_n2736# VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X20 a_n801_n4216# passgatesCtrl_0.net1.t2 VSS.t168 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X21 VDD.t98 a_n1085_n1429# passgatex4_0.GP2 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X22 Z3.t1 passgatex4_0.GN3 A3.t1 VSS.t154 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X23 VDD.t60 VSS.t180 VDD.t59 VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X24 Z3.t0 passgatex4_0.GN3 A3.t0 VSS.t154 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X25 VDD.t175 a_n1459_n3306# a_n1635_n3306# VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X26 passgatesCtrl_0.net10.t2 passgatesCtrl_0.net1.t3 a_n2429_n1328# VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VSS.t7 passgatesCtrl_0._01_ a_n1503_n2192# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X28 VSS.t137 passgatesCtrl_0.net3 a_n1227_n2736# VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X29 VDD.t4 a_n995_n3605# passgatesCtrl_0.net4 VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X30 passgatex4_0.GP1 a_n491_n3280# VSS.t145 VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X31 VSS.t105 passgatesCtrl_0.net7 a_n491_n3280# VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X32 VDD.t74 passgatesCtrl_0._00_ a_n2883_n1648# VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X33 VSS.t173 VDD.t180 VSS.t172 VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X34 a_n715_n3850# passgatesCtrl_0.net1.t4 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X35 VDD.t125 a_n1637_n1429# passgatex4_0.GN4 VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X36 passgatex4_0.GN1 a_n1227_n2736# VDD.t159 VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X37 passgatesCtrl_0.net7 a_n675_n1648# VDD.t121 VDD.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X38 VSS.t155 passgatesCtrl_0._02_ a_n675_n1648# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X39 A3.t2 passgatex4_0.GP3 Z3.t3 VDD.t172 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X40 VDD.t58 VSS.t181 VDD.t57 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X41 a_n482_n4216# select0.t0 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X42 VSS.t175 VDD.t181 VSS.t174 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X43 a_n2185_n2218# a_n2015_n2040# a_n2057_n1942# VDD.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X44 VDD.t56 VSS.t182 VDD.t55 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X45 VSS.t107 a_n1635_n3306# passgatesCtrl_0._03_ VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X46 VDD.t54 VSS.t183 VDD.t53 VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X47 VDD.t52 VSS.t184 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X48 VDD.t140 passgatesCtrl_0._05_ a_n2975_n2192# VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X49 VSS.t119 VDD.t182 VSS.t118 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X50 VDD.t128 a_n1635_n3306# passgatesCtrl_0._03_ VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X51 A2.t1 passgatex4_0.GP2 Z2.t0 VDD.t85 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X52 VSS.t122 VDD.t183 VSS.t121 VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X53 VSS.t55 a_n1984_n4368# a_n1878_n4368# VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X54 VDD.t49 VSS.t185 VDD.t48 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X55 a_n2189_n1429# passgatesCtrl_0.net9 VSS.t113 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X56 VDD.t146 a_n1173_n2218# passgatesCtrl_0._01_ VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X57 VSS.t76 VDD.t184 VSS.t75 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X58 VSS.t52 a_n1003_n2040# a_n1173_n2218# VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X59 a_n2429_n1328# passgatesCtrl_0.net2.t4 VSS.t95 VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 VSS.t131 a_n1173_n2218# passgatesCtrl_0._01_ VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1755 ps=1.84 w=0.65 l=0.15
X61 VSS.t5 a_n995_n3605# passgatesCtrl_0.net4 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X62 VSS.t79 VDD.t185 VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X63 a_n1003_n2040# passgatesCtrl_0.net1.t5 VSS.t135 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1575 ps=1.17 w=0.42 l=0.15
X64 VSS.t65 a_n1085_n1429# passgatex4_0.GP2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X65 passgatesCtrl_0.net2.t1 a_n2480_n4368# VSS.t134 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X66 a_n1459_n3306# passgatesCtrl_0.net1.t6 VDD.t155 VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X67 VDD.t47 VSS.t186 VDD.t46 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X68 a_n1085_n1429# passgatesCtrl_0.net8 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X69 a_n715_n3850# a_n539_n3518# a_n587_n3458# VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X70 a_n587_n3458# passgatesCtrl_0.net1.t7 VSS.t115 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X71 VSS.t21 VDD.t186 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X72 passgatesCtrl_0.net2.t0 a_n2480_n4368# VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X73 passgatesCtrl_0.net8 a_n1503_n2192# VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X74 passgatex4_0.GN1 a_n1227_n2736# VSS.t153 VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X75 A4.t3 passgatex4_0.GP4 Z4.t2 VDD.t163 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X76 Z4.t0 passgatex4_0.GN4 A4.t1 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X77 Z2.t2 passgatex4_0.GN2 A2.t3 VSS.t108 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X78 VDD.t2 passgatesCtrl_0._03_ a_n1963_n3280# VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X79 VSS.t38 a_n801_n4216# a_n988_n4394# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X80 passgatesCtrl_0.net9 a_n2883_n1648# VDD.t144 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X81 VSS.t24 VDD.t187 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X82 VDD.t153 a_n539_n3518# a_n715_n3850# VDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X83 VSS.t36 passgatesCtrl_0._00_ a_n2883_n1648# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X84 a_n1637_n1429# passgatesCtrl_0.net6 VDD.t148 VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X85 VDD.t76 a_n801_n4216# a_n988_n4394# VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X86 VSS.t103 a_n1637_n1429# passgatex4_0.GN4 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X87 VDD.t45 VSS.t187 VDD.t44 VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X88 VDD.t119 a_n2185_n2218# passgatesCtrl_0._00_ VDD.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X89 Z2.t3 passgatex4_0.GN2 A2.t2 VSS.t108 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X90 VSS.t149 a_n1084_n4216# a_n1135_n4368# VSS.t148 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X91 passgatesCtrl_0.net7 a_n675_n1648# VSS.t102 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X92 VDD.t123 passgatesCtrl_0.net1.t8 passgatesCtrl_0.net10.t1 VDD.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X93 VDD.t157 a_n1084_n4216# a_n1135_n4368# VDD.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X94 VSS.t101 a_n2185_n2218# passgatesCtrl_0._00_ VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1755 ps=1.84 w=0.65 l=0.15
X95 VSS.t93 passgatesCtrl_0.net2.t5 a_n539_n3518# VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X96 a_n1173_n2218# passgatesCtrl_0.net2.t6 VSS.t91 VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X97 VSS.t89 passgatesCtrl_0.net2.t7 a_n2161_n4368# VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X98 VSS.t14 VDD.t188 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X99 passgatesCtrl_0.net6 a_n2975_n2192# VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X100 VDD.t43 VSS.t188 VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X101 VSS.t17 VDD.t189 VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X102 VDD.t82 a_n2639_n2040# passgatesCtrl_0._05_ VDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X103 VSS.t61 VDD.t190 VSS.t60 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X104 VSS.t64 VDD.t191 VSS.t63 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X105 a_n2465_n2164# passgatesCtrl_0.net2.t8 VSS.t87 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X106 VSS.t49 a_n2639_n2040# passgatesCtrl_0._05_ VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X107 VDD.t158 passgatesCtrl_0.net4 a_n951_n2736# VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X108 a_n2015_n2040# passgatesCtrl_0.net2.t9 VSS.t85 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1575 ps=1.17 w=0.42 l=0.15
X109 VDD.t40 VSS.t189 VDD.t39 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X110 VDD.t68 a_n1913_n1429# passgatex4_0.GP4 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X111 VDD.t6 passgatesCtrl_0._01_ a_n1503_n2192# VDD.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X112 VDD.t38 VSS.t190 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X113 VSS.t83 passgatesCtrl_0.net2.t10 passgatesCtrl_0.net3 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X114 A1.t3 passgatex4_0.GP1 Z1.t2 VDD.t171 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X115 VSS.t128 a_n482_n4216# passgatesCtrl_0.net1.t0 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X116 VDD.t136 select1.t1 a_n2480_n4368# VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X117 a_n2185_n2218# passgatesCtrl_0.net1.t9 VSS.t126 VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X118 a_n1701_n4368# a_n1878_n4368# VSS.t162 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X119 VDD.t142 a_n482_n4216# passgatesCtrl_0.net1.t1 VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X120 a_n1085_n1429# passgatesCtrl_0.net8 VSS.t50 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X121 VDD.t35 VSS.t191 VDD.t34 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X122 VSS.t44 VDD.t192 VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X123 Z4.t1 passgatex4_0.GN4 A4.t0 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X124 a_n1701_n4368# a_n1878_n4368# VDD.t169 VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X125 passgatesCtrl_0.net10.t0 passgatesCtrl_0.net2.t11 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X126 a_n2639_n2040# passgatesCtrl_0.net2.t12 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X127 VDD.t102 passgatesCtrl_0.net1.t10 a_n1003_n2040# VDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1176 ps=1.4 w=0.42 l=0.15
X128 VSS.t3 passgatesCtrl_0._03_ a_n1963_n3280# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X129 passgatesCtrl_0.net5 a_n1963_n3280# VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X130 a_n1084_n4216# a_n988_n4394# VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X131 a_n539_n3518# passgatesCtrl_0.net2.t13 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X132 passgatesCtrl_0.net9 a_n2883_n1648# VSS.t129 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X133 a_n1637_n1429# passgatesCtrl_0.net6 VSS.t132 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X134 a_n801_n4216# passgatesCtrl_0.net1.t11 VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X135 a_n2639_n2040# passgatesCtrl_0.net1.t12 a_n2465_n2164# VSS.t144 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X136 A3.t3 passgatex4_0.GP3 Z3.t2 VDD.t172 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X137 VDD.t12 a_n597_n2040# passgatesCtrl_0._02_ VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X138 VDD.t33 VSS.t192 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X139 VSS.t47 VDD.t193 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X140 a_n995_n3605# passgatesCtrl_0._04_ VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X141 a_n1507_n3280# passgatesCtrl_0.net2.t14 VSS.t81 VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X142 a_n1635_n3306# a_n1459_n3306# a_n1507_n3280# VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X143 VSS.t11 a_n597_n2040# passgatesCtrl_0._02_ VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X144 VSS.t32 VDD.t194 VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X145 A2.t0 passgatex4_0.GP2 Z2.t1 VDD.t85 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X146 VDD.t30 VSS.t193 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X147 VSS.t151 passgatesCtrl_0.net4 a_n951_n2736# VSS.t150 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X148 VSS.t117 a_n715_n3850# passgatesCtrl_0._04_ VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X149 VDD.t80 a_n1361_n1429# passgatex4_0.GN3 VDD.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X150 a_n1361_n1429# passgatesCtrl_0.net5 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X151 VSS.t164 a_n2015_n2040# a_n2185_n2218# VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X152 VSS.t35 VDD.t195 VSS.t34 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X153 VDD.t27 VSS.t194 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X154 VSS.t71 VDD.t196 VSS.t70 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X155 VDD.t90 passgatesCtrl_0.net1.t13 a_n2639_n2040# VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X156 a_n1045_n1942# passgatesCtrl_0.net2.t15 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14825 ps=1.34 w=0.42 l=0.15
X157 VDD.t92 a_n2189_n1429# passgatex4_0.GP3 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X158 VSS.t124 passgatesCtrl_0._05_ a_n2975_n2192# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X159 a_n482_n4216# select0.t1 VDD.t162 VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X160 passgatesCtrl_0.net3 passgatesCtrl_0.net1.t14 VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X161 A1.t2 passgatex4_0.GP1 Z1.t3 VDD.t171 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X162 VDD.t24 VSS.t195 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X163 VSS.t74 VDD.t197 VSS.t73 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X164 VSS.t147 passgatesCtrl_0.net1.t15 a_n1459_n3306# VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X165 a_n1984_n4368# a_n2161_n4368# VSS.t110 VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X166 VSS.t18 a_n1913_n1429# passgatex4_0.GP4 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X167 a_n1913_n1429# passgatesCtrl_0.net10.t4 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X168 a_n1984_n4368# a_n2161_n4368# VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X169 passgatesCtrl_0.net8 a_n1503_n2192# VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X170 a_n597_n2040# passgatesCtrl_0.net2.t16 a_n434_n1942# VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X171 VDD.t106 passgatesCtrl_0.net2.t17 a_n2015_n2040# VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1176 ps=1.4 w=0.42 l=0.15
X172 VDD.t94 a_n1984_n4368# a_n1878_n4368# VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X173 a_n1635_n3306# passgatesCtrl_0.net2.t18 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X174 passgatex4_0.GN2 a_n951_n2736# VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X175 VDD.t21 VSS.t196 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X176 passgatesCtrl_0.net5 a_n1963_n3280# VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X177 a_n434_n1942# passgatesCtrl_0.net1.t16 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X178 passgatex4_0.GP1 a_n491_n3280# VDD.t154 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X179 A4.t2 passgatex4_0.GP4 Z4.t3 VDD.t163 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X180 VDD.t126 passgatesCtrl_0.net7 a_n491_n3280# VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X181 a_n2057_n1942# passgatesCtrl_0.net1.t17 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14825 ps=1.34 w=0.42 l=0.15
X182 Z1.t0 passgatex4_0.GN1 A1.t1 VSS.t166 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X183 a_n995_n3605# passgatesCtrl_0._04_ VSS.t57 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X184 VDD.t18 VSS.t197 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X185 a_n597_n2040# passgatesCtrl_0.net1.t18 VSS.t170 VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X186 passgatesCtrl_0.net3 passgatesCtrl_0.net2.t19 a_n485_n2736# VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X187 VDD.t151 passgatesCtrl_0.net3 a_n1227_n2736# VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X188 Z1.t1 passgatex4_0.GN1 A1.t0 VSS.t165 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X189 VDD.t165 passgatesCtrl_0._02_ a_n675_n1648# VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X190 VDD.t15 VSS.t198 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X191 a_n485_n2736# passgatesCtrl_0.net1.t19 VDD.t160 VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
R0 passgatesCtrl_0.net2.n5 passgatesCtrl_0.net2.t15 562.236
R1 passgatesCtrl_0.net2.t15 passgatesCtrl_0.net2.t6 392.027
R2 passgatesCtrl_0.net2.n21 passgatesCtrl_0.net2.t13 327.99
R3 passgatesCtrl_0.net2.n2 passgatesCtrl_0.net2.t3 323.55
R4 passgatesCtrl_0.net2.n1 passgatesCtrl_0.net2.t0 319.171
R5 passgatesCtrl_0.net2.n18 passgatesCtrl_0.net2.t14 293.969
R6 passgatesCtrl_0.net2.n13 passgatesCtrl_0.net2.t12 261.887
R7 passgatesCtrl_0.net2.n6 passgatesCtrl_0.net2.t19 230.363
R8 passgatesCtrl_0.net2.n15 passgatesCtrl_0.net2.t11 229.369
R9 passgatesCtrl_0.net2 passgatesCtrl_0.net2.t1 209.923
R10 passgatesCtrl_0.net2.n21 passgatesCtrl_0.net2.t5 199.457
R11 passgatesCtrl_0.net2.n2 passgatesCtrl_0.net2.t7 195.017
R12 passgatesCtrl_0.net2.n8 passgatesCtrl_0.net2.t2 192.639
R13 passgatesCtrl_0.net2.n11 passgatesCtrl_0.net2.t9 185.376
R14 passgatesCtrl_0.net2.n6 passgatesCtrl_0.net2.t10 158.064
R15 passgatesCtrl_0.net2.n15 passgatesCtrl_0.net2.t4 157.07
R16 passgatesCtrl_0.net2.n13 passgatesCtrl_0.net2.t8 155.847
R17 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n8 154.286
R18 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n18 154.065
R19 passgatesCtrl_0.net2.n16 passgatesCtrl_0.net2.n15 153.66
R20 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n2 153.409
R21 passgatesCtrl_0.net2.n7 passgatesCtrl_0.net2.n6 153.097
R22 passgatesCtrl_0.net2.n22 passgatesCtrl_0.net2.n21 152
R23 passgatesCtrl_0.net2.n14 passgatesCtrl_0.net2.n13 152
R24 passgatesCtrl_0.net2.n12 passgatesCtrl_0.net2.n11 152
R25 passgatesCtrl_0.net2.n18 passgatesCtrl_0.net2.t18 138.338
R26 passgatesCtrl_0.net2.n11 passgatesCtrl_0.net2.t17 137.177
R27 passgatesCtrl_0.net2.n8 passgatesCtrl_0.net2.t16 134.799
R28 passgatesCtrl_0.net2.n10 passgatesCtrl_0.net2.n5 26.6879
R29 passgatesCtrl_0.net2.n23 passgatesCtrl_0.net2 24.7034
R30 passgatesCtrl_0.net2.n17 passgatesCtrl_0.net2.n16 21.1865
R31 passgatesCtrl_0.net2.n9 passgatesCtrl_0.net2.n7 21.1676
R32 passgatesCtrl_0.net2.n24 passgatesCtrl_0.net2.n23 17.5163
R33 passgatesCtrl_0.net2.n4 passgatesCtrl_0.net2 16.0005
R34 passgatesCtrl_0.net2.n19 passgatesCtrl_0.net2 15.4844
R35 passgatesCtrl_0.net2.n9 passgatesCtrl_0.net2 11.2434
R36 passgatesCtrl_0.net2.n0 passgatesCtrl_0.net2.n12 10.8365
R37 passgatesCtrl_0.net2.n17 passgatesCtrl_0.net2.n14 10.1066
R38 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n19 10.0713
R39 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n22 9.6005
R40 passgatesCtrl_0.net2.n0 passgatesCtrl_0.net2.n10 9.15538
R41 passgatesCtrl_0.net2.n5 passgatesCtrl_0.net2 8.92171
R42 passgatesCtrl_0.net2.n24 passgatesCtrl_0.net2.n4 8.88939
R43 passgatesCtrl_0.net2.n20 passgatesCtrl_0.net2.n0 8.61863
R44 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n24 7.82272
R45 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n1 7.73474
R46 passgatesCtrl_0.net2.n10 passgatesCtrl_0.net2.n9 7.03724
R47 passgatesCtrl_0.net2 passgatesCtrl_0.net2.n3 6.34564
R48 passgatesCtrl_0.net2.n4 passgatesCtrl_0.net2 6.0165
R49 passgatesCtrl_0.net2.n4 passgatesCtrl_0.net2 5.7605
R50 passgatesCtrl_0.net2.n20 passgatesCtrl_0.net2 5.25599
R51 passgatesCtrl_0.net2.n22 passgatesCtrl_0.net2 4.90717
R52 passgatesCtrl_0.net2.n16 passgatesCtrl_0.net2 4.26717
R53 passgatesCtrl_0.net2.n14 passgatesCtrl_0.net2 3.8405
R54 passgatesCtrl_0.net2.n19 passgatesCtrl_0.net2 3.51018
R55 passgatesCtrl_0.net2.n7 passgatesCtrl_0.net2 3.10907
R56 passgatesCtrl_0.net2.n12 passgatesCtrl_0.net2 3.0725
R57 passgatesCtrl_0.net2.n0 passgatesCtrl_0.net2.n17 2.62704
R58 passgatesCtrl_0.net2.n1 passgatesCtrl_0.net2 2.48634
R59 passgatesCtrl_0.net2.n23 passgatesCtrl_0.net2.n20 2.2972
R60 passgatesCtrl_0.net2.n3 passgatesCtrl_0.net2 2.19479
R61 passgatesCtrl_0.net2.n3 passgatesCtrl_0.net2 1.80756
R62 VSS.t165 VSS.n7 13018.9
R63 VSS.n115 VSS.n114 12462.1
R64 VSS.n108 VSS.n92 12047.7
R65 VSS.n135 VSS.n94 11744.7
R66 VSS.n135 VSS.n95 11744.7
R67 VSS.n94 VSS.n93 11744.7
R68 VSS.n95 VSS.n93 11744.7
R69 VSS.n121 VSS.n100 11744.7
R70 VSS.n121 VSS.n101 11744.7
R71 VSS.n120 VSS.n100 11744.7
R72 VSS.n120 VSS.n101 11744.7
R73 VSS.n113 VSS.n102 11744.7
R74 VSS.n109 VSS.n102 11744.7
R75 VSS.n113 VSS.n103 11744.7
R76 VSS.n109 VSS.n103 11744.7
R77 VSS.n562 VSS.n4 11744.7
R78 VSS.n562 VSS.n5 11744.7
R79 VSS.n560 VSS.n5 11744.7
R80 VSS.n560 VSS.n4 11744.7
R81 VSS.n387 VSS 10843
R82 VSS.n387 VSS.n386 10123.6
R83 VSS.n386 VSS.n385 10123.6
R84 VSS.n137 VSS.n136 3869.02
R85 VSS.n136 VSS.n91 3771.63
R86 VSS.n116 VSS.n91 3735.78
R87 VSS.n561 VSS.n6 3570.22
R88 VSS.n558 VSS.t165 2593.05
R89 VSS.t165 VSS 2390.62
R90 VSS.n561 VSS.n558 2369.23
R91 VSS.t69 VSS.t138 2326.44
R92 VSS.n388 VSS.t19 1938.7
R93 VSS VSS.t12 1694.25
R94 VSS VSS.t15 1601.53
R95 VSS.n386 VSS 1601.53
R96 VSS VSS.n387 1601.53
R97 VSS.t176 VSS.t146 1584.67
R98 VSS.t0 VSS.t77 1567.82
R99 VSS.t163 VSS.t84 1517.24
R100 VSS VSS.t30 1407.66
R101 VSS.t166 VSS.n6 1392.06
R102 VSS VSS.t100 1340.23
R103 VSS VSS.t4 1230.65
R104 VSS.t120 VSS.t158 1219.28
R105 VSS.n384 VSS.n383 1194.5
R106 VSS.n254 VSS.t48 1194.5
R107 VSS.n557 VSS.n556 1194.5
R108 VSS.n389 VSS.n388 1194.5
R109 VSS VSS.t62 1019.92
R110 VSS.t19 VSS 1019.92
R111 VSS VSS.t10 977.779
R112 VSS.t48 VSS 918.774
R113 VSS.t30 VSS 918.774
R114 VSS.n388 VSS 918.774
R115 VSS.t138 VSS 918.774
R116 VSS.t48 VSS.t86 910.346
R117 VSS.t22 VSS 893.633
R118 VSS VSS.n6 851.341
R119 VSS.n558 VSS 851.341
R120 VSS.t127 VSS.t167 848.193
R121 VSS.t88 VSS.t133 848.193
R122 VSS.t100 VSS.t125 826.054
R123 VSS.t116 VSS.t114 826.054
R124 VSS.t106 VSS.t80 826.054
R125 VSS.t42 VSS.t116 792.337
R126 VSS.n112 VSS.n111 767.294
R127 VSS.n559 VSS.n3 767.294
R128 VSS.n131 VSS.n130 763.106
R129 VSS.n119 VSS.n99 763.106
R130 VSS.t33 VSS 742.169
R131 VSS.t150 VSS.t66 741.763
R132 VSS.t6 VSS.t25 741.763
R133 VSS.t39 VSS.t123 741.763
R134 VSS.t104 VSS.t92 741.763
R135 VSS.t4 VSS.t56 741.763
R136 VSS.t2 VSS.t0 741.763
R137 VSS.n130 VSS.n96 732.236
R138 VSS.n123 VSS.n99 732.236
R139 VSS.n112 VSS.n104 732.236
R140 VSS.n559 VSS.n1 732.236
R141 VSS.t130 VSS.t152 724.904
R142 VSS.t37 VSS.t111 711.876
R143 VSS.t54 VSS.t109 711.876
R144 VSS.t90 VSS.t51 708.047
R145 VSS.t125 VSS.t163 708.047
R146 VSS.t80 VSS.t176 657.471
R147 VSS.t15 VSS 632.184
R148 VSS.t12 VSS 632.184
R149 VSS.t148 VSS 594.492
R150 VSS.t144 VSS 564.751
R151 VSS VSS.t6 547.894
R152 VSS.t123 VSS 547.894
R153 VSS VSS.t2 547.894
R154 VSS.t58 VSS.t169 531.034
R155 VSS VSS.t150 531.034
R156 VSS VSS.t136 531.034
R157 VSS VSS.t104 531.034
R158 VSS VSS.t42 531.034
R159 VSS VSS.t161 507.401
R160 VSS.t96 VSS 505.748
R161 VSS.t86 VSS 497.318
R162 VSS VSS.t143 480.461
R163 VSS.n385 VSS.t166 479.757
R164 VSS VSS.t22 458.176
R165 VSS.t158 VSS 458.176
R166 VSS.n557 VSS 412.738
R167 VSS VSS.t120 412.738
R168 VSS.t98 VSS 397.591
R169 VSS.t72 VSS.t69 387.74
R170 VSS.t28 VSS.t127 359.726
R171 VSS.t167 VSS.t37 359.726
R172 VSS.t111 VSS.t148 359.726
R173 VSS.t161 VSS.t54 359.726
R174 VSS.t109 VSS.t88 359.726
R175 VSS.t133 VSS.t98 359.726
R176 VSS.n111 VSS.n110 325.502
R177 VSS.n563 VSS.n3 325.502
R178 VSS.t143 VSS 311.877
R179 VSS.n132 VSS.n131 304.204
R180 VSS.n119 VSS.n118 304.204
R181 VSS.t10 VSS.t58 286.591
R182 VSS VSS.t33 283.993
R183 VSS VSS.t96 278.161
R184 VSS.n226 VSS.t173 273.171
R185 VSS.n431 VSS.t79 273.171
R186 VSS VSS.t28 268.848
R187 VSS VSS.n557 265.06
R188 VSS.n158 VSS.t191 262.719
R189 VSS.n70 VSS.t195 262.719
R190 VSS.t25 VSS 261.303
R191 VSS.t92 VSS 261.303
R192 VSS.t56 VSS 261.303
R193 VSS.t146 VSS 261.303
R194 VSS.n393 VSS.t186 259.082
R195 VSS.n49 VSS.t179 259.082
R196 VSS.n48 VSS.t177 259.082
R197 VSS.n395 VSS.t189 259.082
R198 VSS.n394 VSS.t188 259.082
R199 VSS.n372 VSS.t197 259.082
R200 VSS.n304 VSS.t187 259.082
R201 VSS.n175 VSS.t193 259.082
R202 VSS.n174 VSS.t192 259.082
R203 VSS.n243 VSS.t183 259.082
R204 VSS.n242 VSS.t181 259.082
R205 VSS.n468 VSS.t190 259.082
R206 VSS.n544 VSS.t180 259.082
R207 VSS.t82 VSS 252.875
R208 VSS.t66 VSS 252.875
R209 VSS.n158 VSS.t172 251.564
R210 VSS.n70 VSS.t78 251.564
R211 VSS.t51 VSS 244.445
R212 VSS VSS.t72 244.445
R213 VSS.n133 VSS.n132 242.448
R214 VSS.n118 VSS.n98 242.448
R215 VSS.n110 VSS.n107 242.448
R216 VSS.n564 VSS.n563 242.448
R217 VSS.n179 VSS.t97 241.971
R218 VSS.n411 VSS.t21 240.72
R219 VSS.n439 VSS.t147 237.327
R220 VSS.n53 VSS.t93 237.327
R221 VSS.t171 VSS 236.016
R222 VSS.n64 VSS.t44 233.073
R223 VSS.n241 VSS.t64 225.427
R224 VSS.n504 VSS.t24 225.427
R225 VSS.n551 VSS.t160 225.427
R226 VSS.n411 VSS.t76 225.427
R227 VSS.n391 VSS.t74 225.427
R228 VSS.n89 VSS.t20 225.261
R229 VSS.n401 VSS.t71 221.793
R230 VSS.n51 VSS.t14 221.793
R231 VSS.n51 VSS.t61 221.793
R232 VSS.n396 VSS.t139 221.793
R233 VSS.n396 VSS.t156 221.793
R234 VSS.n373 VSS.t174 221.793
R235 VSS.n305 VSS.t47 221.793
R236 VSS.n177 VSS.t17 221.793
R237 VSS.n177 VSS.t119 221.793
R238 VSS.n244 VSS.t141 221.793
R239 VSS.n244 VSS.t31 221.793
R240 VSS.n469 VSS.t35 221.793
R241 VSS.n545 VSS.t121 221.793
R242 VSS.n42 VSS.t43 221.603
R243 VSS.n240 VSS.t178 218.308
R244 VSS.n24 VSS.t184 218.308
R245 VSS.n542 VSS.t196 218.308
R246 VSS.n90 VSS.t194 218.308
R247 VSS.n390 VSS.t185 218.308
R248 VSS.n240 VSS.t63 217.78
R249 VSS.n24 VSS.t23 217.78
R250 VSS.n542 VSS.t159 217.78
R251 VSS.n90 VSS.t75 217.78
R252 VSS.n390 VSS.t73 217.78
R253 VSS.n393 VSS.t70 215.905
R254 VSS.n49 VSS.t13 215.905
R255 VSS.n48 VSS.t60 215.905
R256 VSS.n395 VSS.t140 215.905
R257 VSS.n394 VSS.t157 215.905
R258 VSS.n372 VSS.t175 215.905
R259 VSS.n304 VSS.t46 215.905
R260 VSS.n175 VSS.t16 215.905
R261 VSS.n174 VSS.t118 215.905
R262 VSS.n243 VSS.t142 215.905
R263 VSS.n242 VSS.t32 215.905
R264 VSS.n468 VSS.t34 215.905
R265 VSS.n544 VSS.t122 215.905
R266 VSS VSS.t144 210.728
R267 VSS.n185 VSS.n184 205.541
R268 VSS.n236 VSS.n235 200.105
R269 VSS.n433 VSS.n69 197.476
R270 VSS.n44 VSS.n43 197.476
R271 VSS.n426 VSS.n73 196.442
R272 VSS.n445 VSS.n41 196.442
R273 VSS.n46 VSS.n45 196.442
R274 VSS.n379 VSS.n370 196.442
R275 VSS.n142 VSS.n141 196.442
R276 VSS.n281 VSS.n280 196.442
R277 VSS.n341 VSS.n283 196.442
R278 VSS.n336 VSS.n286 196.442
R279 VSS.n331 VSS.n289 196.442
R280 VSS.n301 VSS.n300 196.442
R281 VSS.n249 VSS.n239 196.442
R282 VSS.n161 VSS.n160 196.442
R283 VSS.n163 VSS.n162 196.442
R284 VSS.n192 VSS.n191 196.442
R285 VSS.n210 VSS.n209 195.612
R286 VSS.n232 VSS.n155 195.612
R287 VSS.n111 VSS.n103 195
R288 VSS.n103 VSS.t154 195
R289 VSS.n106 VSS.n102 195
R290 VSS.n102 VSS.t154 195
R291 VSS.n120 VSS.n119 195
R292 VSS.t27 VSS.n120 195
R293 VSS.n122 VSS.n121 195
R294 VSS.n121 VSS.t27 195
R295 VSS.n131 VSS.n93 195
R296 VSS.t108 VSS.n93 195
R297 VSS.n135 VSS.n134 195
R298 VSS.t108 VSS.n135 195
R299 VSS.n4 VSS.n2 195
R300 VSS.n137 VSS.n4 195
R301 VSS.n5 VSS.n3 195
R302 VSS.t165 VSS.n5 195
R303 VSS.n475 VSS.n466 194.809
R304 VSS.n481 VSS.n463 194.809
R305 VSS.n497 VSS.n27 194.809
R306 VSS.n512 VSS.n511 194.809
R307 VSS.n519 VSS.n518 194.809
R308 VSS.n537 VSS.n11 194.809
R309 VSS.t169 VSS.t82 177.012
R310 VSS.t114 VSS 177.012
R311 VSS.n117 VSS.n100 172.754
R312 VSS.n114 VSS.t154 161.819
R313 VSS.t108 VSS.n92 161.685
R314 VSS.n172 VSS.t83 152.381
R315 VSS.n171 VSS.t59 150.101
R316 VSS.n365 VSS.t95 147.411
R317 VSS VSS.n137 133.785
R318 VSS.n385 VSS.n384 131.803
R319 VSS.n42 VSS.t182 116.734
R320 VSS.n116 VSS.n115 103.636
R321 VSS.t152 VSS.t90 101.15
R322 VSS.n89 VSS.t198 99.7822
R323 VSS.n108 VSS.n91 97.2732
R324 VSS.n136 VSS.n7 97.1929
R325 VSS.n165 VSS.t135 89.3384
R326 VSS.n156 VSS.t85 89.3384
R327 VSS.n165 VSS.t52 88.7758
R328 VSS.n156 VSS.t164 88.7758
R329 VSS.t8 VSS 81.2618
R330 VSS.n235 VSS.t87 72.8576
R331 VSS.n166 VSS.n165 70.4565
R332 VSS.n157 VSS.n156 70.4565
R333 VSS.t154 VSS.n91 64.546
R334 VSS.n136 VSS.t108 64.4927
R335 VSS.n69 VSS.t81 58.5719
R336 VSS.n43 VSS.t115 58.5719
R337 VSS.n117 VSS.n116 58.1458
R338 VSS.n184 VSS.t170 55.7148
R339 VSS.n209 VSS.t91 52.8576
R340 VSS.n155 VSS.t126 52.8576
R341 VSS.n466 VSS.t29 45.7148
R342 VSS.n463 VSS.t168 45.7148
R343 VSS.n27 VSS.t112 45.7148
R344 VSS.n511 VSS.t55 45.7148
R345 VSS.n518 VSS.t89 45.7148
R346 VSS.n11 VSS.t99 45.7148
R347 VSS.n305 VSS.n303 34.6358
R348 VSS.n309 VSS.n303 34.6358
R349 VSS.n310 VSS.n309 34.6358
R350 VSS.n311 VSS.n310 34.6358
R351 VSS.n311 VSS.n301 34.6358
R352 VSS.n315 VSS.n301 34.6358
R353 VSS.n316 VSS.n315 34.6358
R354 VSS.n316 VSS.n290 34.6358
R355 VSS.n330 VSS.n290 34.6358
R356 VSS.n331 VSS.n330 34.6358
R357 VSS.n331 VSS.n287 34.6358
R358 VSS.n335 VSS.n287 34.6358
R359 VSS.n336 VSS.n335 34.6358
R360 VSS.n337 VSS.n336 34.6358
R361 VSS.n337 VSS.n284 34.6358
R362 VSS.n341 VSS.n284 34.6358
R363 VSS.n342 VSS.n341 34.6358
R364 VSS.n343 VSS.n342 34.6358
R365 VSS.n343 VSS.n281 34.6358
R366 VSS.n347 VSS.n281 34.6358
R367 VSS.n348 VSS.n347 34.6358
R368 VSS.n348 VSS.n142 34.6358
R369 VSS.n363 VSS.n142 34.6358
R370 VSS.n364 VSS.n363 34.6358
R371 VSS.n366 VSS.n364 34.6358
R372 VSS.n383 VSS.n138 34.6358
R373 VSS.n383 VSS.n139 34.6358
R374 VSS.n379 VSS.n139 34.6358
R375 VSS.n379 VSS.n378 34.6358
R376 VSS.n378 VSS.n377 34.6358
R377 VSS.n377 VSS.n371 34.6358
R378 VSS.n373 VSS.n371 34.6358
R379 VSS.n178 VSS.n177 34.6358
R380 VSS.n180 VSS.n178 34.6358
R381 VSS.n186 VSS.n183 34.6358
R382 VSS.n190 VSS.n171 34.6358
R383 VSS.n193 VSS.n190 34.6358
R384 VSS.n193 VSS.n192 34.6358
R385 VSS.n211 VSS.n208 34.6358
R386 VSS.n215 VSS.n163 34.6358
R387 VSS.n216 VSS.n215 34.6358
R388 VSS.n216 VSS.n161 34.6358
R389 VSS.n220 VSS.n161 34.6358
R390 VSS.n221 VSS.n220 34.6358
R391 VSS.n221 VSS.n159 34.6358
R392 VSS.n225 VSS.n159 34.6358
R393 VSS.n231 VSS.n230 34.6358
R394 VSS.n269 VSS.n268 34.6358
R395 VSS.n268 VSS.n233 34.6358
R396 VSS.n258 VSS.n233 34.6358
R397 VSS.n258 VSS.n257 34.6358
R398 VSS.n254 VSS.n253 34.6358
R399 VSS.n253 VSS.n237 34.6358
R400 VSS.n249 VSS.n248 34.6358
R401 VSS.n248 VSS.n247 34.6358
R402 VSS.n247 VSS.n244 34.6358
R403 VSS.n469 VSS.n467 34.6358
R404 VSS.n473 VSS.n467 34.6358
R405 VSS.n474 VSS.n473 34.6358
R406 VSS.n476 VSS.n464 34.6358
R407 VSS.n480 VSS.n464 34.6358
R408 VSS.n482 VSS.n28 34.6358
R409 VSS.n496 VSS.n28 34.6358
R410 VSS.n498 VSS.n25 34.6358
R411 VSS.n502 VSS.n25 34.6358
R412 VSS.n503 VSS.n502 34.6358
R413 VSS.n505 VSS.n22 34.6358
R414 VSS.n509 VSS.n22 34.6358
R415 VSS.n510 VSS.n509 34.6358
R416 VSS.n513 VSS.n510 34.6358
R417 VSS.n517 VSS.n20 34.6358
R418 VSS.n520 VSS.n517 34.6358
R419 VSS.n535 VSS.n12 34.6358
R420 VSS.n536 VSS.n535 34.6358
R421 VSS.n538 VSS.n8 34.6358
R422 VSS.n556 VSS.n8 34.6358
R423 VSS.n556 VSS.n9 34.6358
R424 VSS.n552 VSS.n9 34.6358
R425 VSS.n550 VSS.n549 34.6358
R426 VSS.n549 VSS.n543 34.6358
R427 VSS.n545 VSS.n543 34.6358
R428 VSS.n52 VSS.n51 34.6358
R429 VSS.n54 VSS.n52 34.6358
R430 VSS.n58 VSS.n46 34.6358
R431 VSS.n59 VSS.n58 34.6358
R432 VSS.n63 VSS.n62 34.6358
R433 VSS.n445 VSS.n65 34.6358
R434 VSS.n445 VSS.n444 34.6358
R435 VSS.n444 VSS.n66 34.6358
R436 VSS.n440 VSS.n66 34.6358
R437 VSS.n438 VSS.n67 34.6358
R438 VSS.n434 VSS.n67 34.6358
R439 VSS.n430 VSS.n71 34.6358
R440 VSS.n426 VSS.n71 34.6358
R441 VSS.n426 VSS.n425 34.6358
R442 VSS.n425 VSS.n424 34.6358
R443 VSS.n424 VSS.n74 34.6358
R444 VSS.n88 VSS.n74 34.6358
R445 VSS.n412 VSS.n88 34.6358
R446 VSS.n410 VSS.n409 34.6358
R447 VSS.n409 VSS.n389 34.6358
R448 VSS.n405 VSS.n389 34.6358
R449 VSS.n405 VSS.n404 34.6358
R450 VSS.n401 VSS.n400 34.6358
R451 VSS.n400 VSS.n399 34.6358
R452 VSS.n399 VSS.n396 34.6358
R453 VSS.n466 VSS.t128 34.506
R454 VSS.n463 VSS.t38 34.506
R455 VSS.n27 VSS.t149 34.506
R456 VSS.n511 VSS.t162 34.506
R457 VSS.n518 VSS.t110 34.506
R458 VSS.n11 VSS.t134 34.506
R459 VSS.n366 VSS.n365 33.8829
R460 VSS.n497 VSS.n496 33.5064
R461 VSS.n73 VSS.t1 33.462
R462 VSS.n73 VSS.t3 33.462
R463 VSS.n41 VSS.t57 33.462
R464 VSS.n41 VSS.t5 33.462
R465 VSS.n45 VSS.t145 33.462
R466 VSS.n45 VSS.t105 33.462
R467 VSS.n370 VSS.t129 33.462
R468 VSS.n370 VSS.t36 33.462
R469 VSS.n141 VSS.t113 33.462
R470 VSS.n141 VSS.t53 33.462
R471 VSS.n280 VSS.t68 33.462
R472 VSS.n280 VSS.t18 33.462
R473 VSS.n283 VSS.t132 33.462
R474 VSS.n283 VSS.t103 33.462
R475 VSS.n286 VSS.t9 33.462
R476 VSS.n286 VSS.t41 33.462
R477 VSS.n289 VSS.t50 33.462
R478 VSS.n289 VSS.t65 33.462
R479 VSS.n300 VSS.t102 33.462
R480 VSS.n300 VSS.t155 33.462
R481 VSS.n239 VSS.t40 33.462
R482 VSS.n239 VSS.t124 33.462
R483 VSS.n160 VSS.t26 33.462
R484 VSS.n160 VSS.t7 33.462
R485 VSS.n162 VSS.t153 33.462
R486 VSS.n162 VSS.t137 33.462
R487 VSS.n191 VSS.t67 33.462
R488 VSS.n191 VSS.t151 33.462
R489 VSS.n512 VSS.n20 33.1299
R490 VSS.n59 VSS.n44 33.1299
R491 VSS.n434 VSS.n433 33.1299
R492 VSS.n53 VSS.n46 32.377
R493 VSS.n439 VSS.n438 32.377
R494 VSS.n211 VSS.n210 31.2476
R495 VSS.n232 VSS.n231 31.2476
R496 VSS.n134 VSS.n96 30.8711
R497 VSS.n123 VSS.n122 30.8711
R498 VSS.n106 VSS.n104 30.8711
R499 VSS.n481 VSS.n480 30.8711
R500 VSS.n2 VSS.n1 30.8711
R501 VSS.n519 VSS.n12 30.4946
R502 VSS.n209 VSS.t131 28.3166
R503 VSS.n155 VSS.t101 28.3166
R504 VSS.n184 VSS.t11 26.8576
R505 VSS.n69 VSS.t107 25.4291
R506 VSS.n43 VSS.t117 25.4291
R507 VSS.n185 VSS.n171 24.0946
R508 VSS.n179 VSS.n172 23.7181
R509 VSS.n235 VSS.t49 22.3257
R510 VSS.n226 VSS.n158 21.6078
R511 VSS.n431 VSS.n70 21.6078
R512 VSS.n192 VSS.n166 20.3299
R513 VSS.n227 VSS.n157 20.3299
R514 VSS.n537 VSS.n536 20.3299
R515 VSS.n476 VSS.n475 19.9534
R516 VSS.n254 VSS.n236 18.824
R517 VSS.n226 VSS.n225 17.3181
R518 VSS.n227 VSS.n226 17.3181
R519 VSS.n241 VSS.n237 17.3181
R520 VSS.n249 VSS.n241 17.3181
R521 VSS.n504 VSS.n503 17.3181
R522 VSS.n505 VSS.n504 17.3181
R523 VSS.n552 VSS.n551 17.3181
R524 VSS.n551 VSS.n550 17.3181
R525 VSS.n64 VSS.n63 17.3181
R526 VSS.n65 VSS.n64 17.3181
R527 VSS.n432 VSS.n431 17.3181
R528 VSS.n431 VSS.n430 17.3181
R529 VSS.n412 VSS.n411 17.3181
R530 VSS.n411 VSS.n410 17.3181
R531 VSS.n404 VSS.n391 17.3181
R532 VSS.n401 VSS.n391 17.3181
R533 VSS.t136 VSS.t130 16.8587
R534 VSS.t84 VSS.t171 16.8587
R535 VSS.t62 VSS.t39 16.8587
R536 VSS.t77 VSS.t106 16.8587
R537 VSS.n384 VSS.t94 15.8564
R538 VSS.n257 VSS.n236 15.8123
R539 VSS.n411 VSS.n89 15.4602
R540 VSS.n475 VSS.n474 14.6829
R541 VSS.n208 VSS.n166 14.3064
R542 VSS.n230 VSS.n157 14.3064
R543 VSS.n538 VSS.n537 14.3064
R544 VSS.n81 VSS 13.1605
R545 VSS.n64 VSS.n42 11.4706
R546 VSS.n110 VSS.n109 11.0382
R547 VSS.n109 VSS.n108 11.0382
R548 VSS.n113 VSS.n112 11.0382
R549 VSS.n114 VSS.n113 11.0382
R550 VSS.n118 VSS.n101 11.0382
R551 VSS.n115 VSS.n101 11.0382
R552 VSS.n100 VSS.n99 11.0382
R553 VSS.n132 VSS.n95 11.0382
R554 VSS.n95 VSS.n7 11.0382
R555 VSS.n130 VSS.n94 11.0382
R556 VSS.n94 VSS.n92 11.0382
R557 VSS.n560 VSS.n559 11.0382
R558 VSS.n561 VSS.n560 11.0382
R559 VSS.n563 VSS.n562 11.0382
R560 VSS.n562 VSS.n561 11.0382
R561 VSS.n134 VSS.n133 10.9181
R562 VSS.n122 VSS.n98 10.9181
R563 VSS.n107 VSS.n106 10.9181
R564 VSS.n564 VSS.n2 10.9181
R565 VSS.n180 VSS.n179 10.5417
R566 VSS.n186 VSS.n185 10.5417
R567 VSS.n129 VSS.n96 10.4476
R568 VSS.n124 VSS.n123 10.4476
R569 VSS.n105 VSS.n104 10.4476
R570 VSS.n565 VSS.n1 10.4476
R571 VSS.t94 VSS.t45 9.91041
R572 VSS.n307 VSS.n303 9.3005
R573 VSS.n309 VSS.n308 9.3005
R574 VSS.n310 VSS.n302 9.3005
R575 VSS.n312 VSS.n311 9.3005
R576 VSS.n313 VSS.n301 9.3005
R577 VSS.n315 VSS.n314 9.3005
R578 VSS.n317 VSS.n316 9.3005
R579 VSS.n291 VSS.n290 9.3005
R580 VSS.n330 VSS.n329 9.3005
R581 VSS.n332 VSS.n331 9.3005
R582 VSS.n333 VSS.n287 9.3005
R583 VSS.n335 VSS.n334 9.3005
R584 VSS.n336 VSS.n285 9.3005
R585 VSS.n338 VSS.n337 9.3005
R586 VSS.n339 VSS.n284 9.3005
R587 VSS.n341 VSS.n340 9.3005
R588 VSS.n342 VSS.n282 9.3005
R589 VSS.n344 VSS.n343 9.3005
R590 VSS.n345 VSS.n281 9.3005
R591 VSS.n347 VSS.n346 9.3005
R592 VSS.n349 VSS.n348 9.3005
R593 VSS.n353 VSS.n142 9.3005
R594 VSS.n363 VSS.n362 9.3005
R595 VSS.n364 VSS.n140 9.3005
R596 VSS.n367 VSS.n366 9.3005
R597 VSS.n368 VSS.n138 9.3005
R598 VSS.n383 VSS.n382 9.3005
R599 VSS.n381 VSS.n139 9.3005
R600 VSS.n380 VSS.n379 9.3005
R601 VSS.n378 VSS.n369 9.3005
R602 VSS.n377 VSS.n376 9.3005
R603 VSS.n375 VSS.n371 9.3005
R604 VSS.n247 VSS.n246 9.3005
R605 VSS.n178 VSS.n173 9.3005
R606 VSS.n181 VSS.n180 9.3005
R607 VSS.n183 VSS.n182 9.3005
R608 VSS.n187 VSS.n186 9.3005
R609 VSS.n188 VSS.n171 9.3005
R610 VSS.n190 VSS.n189 9.3005
R611 VSS.n194 VSS.n193 9.3005
R612 VSS.n192 VSS.n167 9.3005
R613 VSS.n208 VSS.n207 9.3005
R614 VSS.n212 VSS.n211 9.3005
R615 VSS.n213 VSS.n163 9.3005
R616 VSS.n215 VSS.n214 9.3005
R617 VSS.n217 VSS.n216 9.3005
R618 VSS.n218 VSS.n161 9.3005
R619 VSS.n220 VSS.n219 9.3005
R620 VSS.n222 VSS.n221 9.3005
R621 VSS.n223 VSS.n159 9.3005
R622 VSS.n225 VSS.n224 9.3005
R623 VSS.n228 VSS.n227 9.3005
R624 VSS.n230 VSS.n229 9.3005
R625 VSS.n231 VSS.n153 9.3005
R626 VSS.n270 VSS.n269 9.3005
R627 VSS.n268 VSS.n267 9.3005
R628 VSS.n260 VSS.n233 9.3005
R629 VSS.n259 VSS.n258 9.3005
R630 VSS.n257 VSS.n256 9.3005
R631 VSS.n255 VSS.n254 9.3005
R632 VSS.n253 VSS.n252 9.3005
R633 VSS.n251 VSS.n237 9.3005
R634 VSS.n250 VSS.n249 9.3005
R635 VSS.n248 VSS.n238 9.3005
R636 VSS.n547 VSS.n543 9.3005
R637 VSS.n471 VSS.n467 9.3005
R638 VSS.n473 VSS.n472 9.3005
R639 VSS.n474 VSS.n465 9.3005
R640 VSS.n477 VSS.n476 9.3005
R641 VSS.n478 VSS.n464 9.3005
R642 VSS.n480 VSS.n479 9.3005
R643 VSS.n483 VSS.n482 9.3005
R644 VSS.n29 VSS.n28 9.3005
R645 VSS.n496 VSS.n495 9.3005
R646 VSS.n499 VSS.n498 9.3005
R647 VSS.n500 VSS.n25 9.3005
R648 VSS.n502 VSS.n501 9.3005
R649 VSS.n503 VSS.n23 9.3005
R650 VSS.n506 VSS.n505 9.3005
R651 VSS.n507 VSS.n22 9.3005
R652 VSS.n509 VSS.n508 9.3005
R653 VSS.n510 VSS.n21 9.3005
R654 VSS.n514 VSS.n513 9.3005
R655 VSS.n515 VSS.n20 9.3005
R656 VSS.n517 VSS.n516 9.3005
R657 VSS.n521 VSS.n520 9.3005
R658 VSS.n525 VSS.n12 9.3005
R659 VSS.n535 VSS.n534 9.3005
R660 VSS.n536 VSS.n10 9.3005
R661 VSS.n539 VSS.n538 9.3005
R662 VSS.n540 VSS.n8 9.3005
R663 VSS.n556 VSS.n555 9.3005
R664 VSS.n554 VSS.n9 9.3005
R665 VSS.n553 VSS.n552 9.3005
R666 VSS.n550 VSS.n541 9.3005
R667 VSS.n549 VSS.n548 9.3005
R668 VSS.n399 VSS.n398 9.3005
R669 VSS.n52 VSS.n47 9.3005
R670 VSS.n55 VSS.n54 9.3005
R671 VSS.n56 VSS.n46 9.3005
R672 VSS.n58 VSS.n57 9.3005
R673 VSS.n60 VSS.n59 9.3005
R674 VSS.n62 VSS.n61 9.3005
R675 VSS.n63 VSS.n37 9.3005
R676 VSS.n65 VSS.n38 9.3005
R677 VSS.n446 VSS.n445 9.3005
R678 VSS.n444 VSS.n443 9.3005
R679 VSS.n442 VSS.n66 9.3005
R680 VSS.n441 VSS.n440 9.3005
R681 VSS.n438 VSS.n437 9.3005
R682 VSS.n436 VSS.n67 9.3005
R683 VSS.n435 VSS.n434 9.3005
R684 VSS.n432 VSS.n68 9.3005
R685 VSS.n430 VSS.n429 9.3005
R686 VSS.n428 VSS.n71 9.3005
R687 VSS.n427 VSS.n426 9.3005
R688 VSS.n425 VSS.n72 9.3005
R689 VSS.n424 VSS.n423 9.3005
R690 VSS.n76 VSS.n74 9.3005
R691 VSS.n88 VSS.n87 9.3005
R692 VSS.n413 VSS.n412 9.3005
R693 VSS.n410 VSS.n84 9.3005
R694 VSS.n409 VSS.n408 9.3005
R695 VSS.n407 VSS.n389 9.3005
R696 VSS.n406 VSS.n405 9.3005
R697 VSS.n404 VSS.n403 9.3005
R698 VSS.n402 VSS.n401 9.3005
R699 VSS.n400 VSS.n392 9.3005
R700 VSS.n126 VSS.n125 8.45078
R701 VSS.n566 VSS.n0 8.30267
R702 VSS.n128 VSS.n127 7.97888
R703 VSS.n126 VSS.n97 7.97601
R704 VSS.n306 VSS.n305 7.66295
R705 VSS.n177 VSS.n176 7.66295
R706 VSS.n470 VSS.n469 7.66295
R707 VSS.n51 VSS.n50 7.66295
R708 VSS.n374 VSS.n373 7.65909
R709 VSS.n245 VSS.n244 7.65909
R710 VSS.n546 VSS.n545 7.65909
R711 VSS.n397 VSS.n396 7.65909
R712 VSS.n241 VSS.n240 7.64725
R713 VSS.n504 VSS.n24 7.64725
R714 VSS.n551 VSS.n542 7.64725
R715 VSS.n411 VSS.n90 7.64725
R716 VSS.n391 VSS.n390 7.64725
R717 VSS.n129 VSS.n128 7.16724
R718 VSS.n125 VSS.n124 7.16724
R719 VSS.n105 VSS.n97 7.16724
R720 VSS.n566 VSS.n565 7.16724
R721 VSS.n401 VSS.n393 5.8885
R722 VSS.n51 VSS.n48 5.8885
R723 VSS.n51 VSS.n49 5.8885
R724 VSS.n396 VSS.n394 5.8885
R725 VSS.n396 VSS.n395 5.8885
R726 VSS.n373 VSS.n372 5.8885
R727 VSS.n305 VSS.n304 5.8885
R728 VSS.n177 VSS.n174 5.8885
R729 VSS.n177 VSS.n175 5.8885
R730 VSS.n244 VSS.n242 5.8885
R731 VSS.n244 VSS.n243 5.8885
R732 VSS.n469 VSS.n468 5.8885
R733 VSS.n545 VSS.n544 5.8885
R734 VSS.n133 VSS.n129 4.73093
R735 VSS.n124 VSS.n98 4.73093
R736 VSS.n107 VSS.n105 4.73093
R737 VSS.n565 VSS.n564 4.73093
R738 VSS.n356 VSS.n278 4.51401
R739 VSS.n361 VSS.n360 4.51401
R740 VSS.n322 VSS.n298 4.51401
R741 VSS.n326 VSS.n288 4.51401
R742 VSS.n273 VSS.n151 4.51401
R743 VSS.n266 VSS.n265 4.51401
R744 VSS.n199 VSS.n170 4.51401
R745 VSS.n204 VSS.n164 4.51401
R746 VSS.n455 VSS.n35 4.51401
R747 VSS.n40 VSS.n39 4.51401
R748 VSS.n528 VSS.n18 4.51401
R749 VSS.n533 VSS.n532 4.51401
R750 VSS.n488 VSS.n461 4.51401
R751 VSS.n492 VSS.n26 4.51401
R752 VSS.n77 VSS.n75 4.51401
R753 VSS.n415 VSS.n414 4.51401
R754 VSS.n144 VSS.n143 4.5005
R755 VSS.n355 VSS.n354 4.5005
R756 VSS.n352 VSS.n351 4.5005
R757 VSS.n321 VSS.n320 4.5005
R758 VSS.n319 VSS.n318 4.5005
R759 VSS.n328 VSS.n327 4.5005
R760 VSS.n264 VSS.n234 4.5005
R761 VSS.n272 VSS.n271 4.5005
R762 VSS.n261 VSS.n154 4.5005
R763 VSS.n198 VSS.n197 4.5005
R764 VSS.n196 VSS.n195 4.5005
R765 VSS.n206 VSS.n205 4.5005
R766 VSS.n14 VSS.n13 4.5005
R767 VSS.n527 VSS.n526 4.5005
R768 VSS.n524 VSS.n523 4.5005
R769 VSS.n487 VSS.n486 4.5005
R770 VSS.n485 VSS.n484 4.5005
R771 VSS.n494 VSS.n493 4.5005
R772 VSS.n86 VSS.n83 4.5005
R773 VSS.n454 VSS.n453 4.5005
R774 VSS.n452 VSS.n451 4.5005
R775 VSS.n448 VSS.n447 4.5005
R776 VSS.n422 VSS.n421 4.5005
R777 VSS.n85 VSS.n78 4.5005
R778 VSS.n520 VSS.n519 4.14168
R779 VSS.n146 VSS 4.01425
R780 VSS.n482 VSS.n481 3.76521
R781 VSS.n360 VSS.n359 3.43925
R782 VSS.n357 VSS.n356 3.43925
R783 VSS.n326 VSS.n325 3.43925
R784 VSS.n323 VSS.n322 3.43925
R785 VSS.n265 VSS.n149 3.43925
R786 VSS.n274 VSS.n273 3.43925
R787 VSS.n204 VSS.n203 3.43925
R788 VSS.n200 VSS.n199 3.43925
R789 VSS.n39 VSS.n33 3.43925
R790 VSS.n456 VSS.n455 3.43925
R791 VSS.n532 VSS.n531 3.43925
R792 VSS.n529 VSS.n528 3.43925
R793 VSS.n492 VSS.n491 3.43925
R794 VSS.n489 VSS.n488 3.43925
R795 VSS.n279 VSS.n277 3.4105
R796 VSS.n350 VSS.n145 3.4105
R797 VSS.n299 VSS.n297 3.4105
R798 VSS.n293 VSS.n292 3.4105
R799 VSS.n152 VSS.n150 3.4105
R800 VSS.n263 VSS.n262 3.4105
R801 VSS.n201 VSS.n169 3.4105
R802 VSS.n202 VSS.n168 3.4105
R803 VSS.n36 VSS.n34 3.4105
R804 VSS.n450 VSS.n449 3.4105
R805 VSS.n19 VSS.n17 3.4105
R806 VSS.n522 VSS.n15 3.4105
R807 VSS.n462 VSS.n460 3.4105
R808 VSS.n31 VSS.n30 3.4105
R809 VSS.n417 VSS.n416 3.4105
R810 VSS.n417 VSS.n79 3.4105
R811 VSS.n416 VSS.n415 3.4105
R812 VSS.n79 VSS.n77 3.4105
R813 VSS.n420 VSS.n419 3.4105
R814 VSS.n82 VSS.n80 3.4105
R815 VSS.n210 VSS.n163 3.38874
R816 VSS.n269 VSS.n232 3.38874
R817 VSS.t45 VSS.t8 2.97347
R818 VSS.n54 VSS.n53 2.25932
R819 VSS.n440 VSS.n439 2.25932
R820 VSS.n491 VSS.n490 1.69188
R821 VSS.n490 VSS.n489 1.69188
R822 VSS.n457 VSS.n33 1.69188
R823 VSS.n457 VSS.n456 1.69188
R824 VSS.n203 VSS.n32 1.69188
R825 VSS.n200 VSS.n32 1.69188
R826 VSS.n325 VSS.n324 1.69188
R827 VSS.n324 VSS.n323 1.69188
R828 VSS.n531 VSS.n530 1.69188
R829 VSS.n530 VSS.n529 1.69188
R830 VSS.n275 VSS.n149 1.69188
R831 VSS.n275 VSS.n274 1.69188
R832 VSS.n359 VSS.n358 1.69188
R833 VSS.n358 VSS.n357 1.69188
R834 VSS.n418 VSS.n417 1.69188
R835 VSS.n513 VSS.n512 1.50638
R836 VSS.n62 VSS.n44 1.50638
R837 VSS.n433 VSS.n432 1.50638
R838 VSS.n498 VSS.n497 1.12991
R839 VSS.n358 VSS.n148 0.867399
R840 VSS.n365 VSS.n138 0.753441
R841 VSS.n324 VSS.n148 0.659756
R842 VSS.n147 VSS.n146 0.595833
R843 VSS.n459 VSS.n458 0.500125
R844 VSS.n295 VSS.n294 0.500125
R845 VSS.n296 VSS 0.478236
R846 VSS.n127 VSS.n126 0.467019
R847 VSS.n294 VSS.n276 0.3805
R848 VSS.n458 VSS.n16 0.3805
R849 VSS.n183 VSS.n172 0.376971
R850 VSS.n146 VSS.n0 0.195328
R851 VSS.n530 VSS.n16 0.162755
R852 VSS.n457 VSS.n32 0.1603
R853 VSS.n490 VSS.n459 0.159712
R854 VSS.n375 VSS.n374 0.141672
R855 VSS.n246 VSS.n245 0.141672
R856 VSS.n547 VSS.n546 0.141672
R857 VSS.n398 VSS.n397 0.141672
R858 VSS.n307 VSS.n306 0.137814
R859 VSS.n176 VSS.n173 0.137814
R860 VSS.n471 VSS.n470 0.137814
R861 VSS.n50 VSS.n47 0.137814
R862 VSS.n148 VSS.n147 0.13699
R863 VSS.n358 VSS.n276 0.129226
R864 VSS.n374 VSS 0.121778
R865 VSS.n245 VSS 0.121778
R866 VSS.n546 VSS 0.121778
R867 VSS.n397 VSS 0.121778
R868 VSS.n296 VSS.n295 0.121084
R869 VSS.n308 VSS.n307 0.120292
R870 VSS.n312 VSS.n302 0.120292
R871 VSS.n313 VSS.n312 0.120292
R872 VSS.n314 VSS.n313 0.120292
R873 VSS.n333 VSS.n332 0.120292
R874 VSS.n334 VSS.n333 0.120292
R875 VSS.n338 VSS.n285 0.120292
R876 VSS.n339 VSS.n338 0.120292
R877 VSS.n340 VSS.n282 0.120292
R878 VSS.n344 VSS.n282 0.120292
R879 VSS.n346 VSS.n345 0.120292
R880 VSS.n367 VSS.n140 0.120292
R881 VSS.n368 VSS.n367 0.120292
R882 VSS.n381 VSS.n380 0.120292
R883 VSS.n380 VSS.n369 0.120292
R884 VSS.n181 VSS.n173 0.120292
R885 VSS.n188 VSS.n187 0.120292
R886 VSS.n189 VSS.n188 0.120292
R887 VSS.n213 VSS.n212 0.120292
R888 VSS.n214 VSS.n213 0.120292
R889 VSS.n219 VSS.n218 0.120292
R890 VSS.n224 VSS.n223 0.120292
R891 VSS.n229 VSS.n228 0.120292
R892 VSS.n256 VSS.n255 0.120292
R893 VSS.n251 VSS.n250 0.120292
R894 VSS.n250 VSS.n238 0.120292
R895 VSS.n472 VSS.n471 0.120292
R896 VSS.n477 VSS.n465 0.120292
R897 VSS.n478 VSS.n477 0.120292
R898 VSS.n479 VSS.n478 0.120292
R899 VSS.n500 VSS.n499 0.120292
R900 VSS.n501 VSS.n500 0.120292
R901 VSS.n506 VSS.n23 0.120292
R902 VSS.n507 VSS.n506 0.120292
R903 VSS.n508 VSS.n507 0.120292
R904 VSS.n514 VSS.n21 0.120292
R905 VSS.n515 VSS.n514 0.120292
R906 VSS.n516 VSS.n515 0.120292
R907 VSS.n539 VSS.n10 0.120292
R908 VSS.n540 VSS.n539 0.120292
R909 VSS.n553 VSS.n541 0.120292
R910 VSS.n548 VSS.n541 0.120292
R911 VSS.n548 VSS.n547 0.120292
R912 VSS.n55 VSS.n47 0.120292
R913 VSS.n57 VSS.n56 0.120292
R914 VSS.n443 VSS.n442 0.120292
R915 VSS.n437 VSS.n436 0.120292
R916 VSS.n436 VSS.n435 0.120292
R917 VSS.n435 VSS.n68 0.120292
R918 VSS.n429 VSS.n68 0.120292
R919 VSS.n429 VSS.n428 0.120292
R920 VSS.n428 VSS.n427 0.120292
R921 VSS.n427 VSS.n72 0.120292
R922 VSS.n413 VSS.n84 0.120292
R923 VSS.n408 VSS.n84 0.120292
R924 VSS.n408 VSS.n407 0.120292
R925 VSS.n402 VSS.n392 0.120292
R926 VSS.n398 VSS.n392 0.120292
R927 VSS.n458 VSS 0.107437
R928 VSS.n294 VSS 0.107437
R929 VSS VSS.n375 0.104667
R930 VSS VSS.n465 0.104667
R931 VSS.n217 VSS 0.10076
R932 VSS.n60 VSS 0.10076
R933 VSS.n376 VSS 0.0981562
R934 VSS.n182 VSS 0.0981562
R935 VSS.n218 VSS 0.0981562
R936 VSS.n222 VSS 0.0981562
R937 VSS VSS.n259 0.0981562
R938 VSS VSS.n251 0.0981562
R939 VSS.n246 VSS 0.0981562
R940 VSS VSS.n23 0.0981562
R941 VSS VSS.n553 0.0981562
R942 VSS.n56 VSS 0.0981562
R943 VSS.n61 VSS 0.0981562
R944 VSS VSS.n441 0.0981562
R945 VSS.n437 VSS 0.0981562
R946 VSS.n403 VSS 0.0981562
R947 VSS VSS.n402 0.0981562
R948 VSS.n346 VSS.n278 0.0968542
R949 VSS.n382 VSS 0.0968542
R950 VSS.n187 VSS 0.0968542
R951 VSS.n228 VSS 0.0968542
R952 VSS.n229 VSS.n151 0.0968542
R953 VSS.n516 VSS.n18 0.0968542
R954 VSS VSS.n285 0.0955521
R955 VSS.n340 VSS 0.0955521
R956 VSS.n345 VSS 0.0955521
R957 VSS.n356 VSS.n355 0.0950946
R958 VSS.n360 VSS.n144 0.0950946
R959 VSS.n322 VSS.n321 0.0950946
R960 VSS.n327 VSS.n326 0.0950946
R961 VSS.n273 VSS.n272 0.0950946
R962 VSS.n265 VSS.n264 0.0950946
R963 VSS.n199 VSS.n198 0.0950946
R964 VSS.n205 VSS.n204 0.0950946
R965 VSS.n455 VSS.n454 0.0950946
R966 VSS.n448 VSS.n39 0.0950946
R967 VSS.n528 VSS.n527 0.0950946
R968 VSS.n532 VSS.n14 0.0950946
R969 VSS.n488 VSS.n487 0.0950946
R970 VSS.n493 VSS.n492 0.0950946
R971 VSS.n421 VSS.n77 0.0950946
R972 VSS.n415 VSS.n83 0.0950946
R973 VSS.n332 VSS.n288 0.0916458
R974 VSS.n212 VSS.n164 0.0916458
R975 VSS.n499 VSS.n26 0.0916458
R976 VSS.n555 VSS 0.0916458
R977 VSS.n443 VSS.n40 0.0916458
R978 VSS VSS.n381 0.0864375
R979 VSS.n252 VSS 0.0864375
R980 VSS VSS.n554 0.0864375
R981 VSS VSS.n406 0.0864375
R982 VSS VSS.n302 0.0851354
R983 VSS.n223 VSS 0.0851354
R984 VSS.n256 VSS 0.0851354
R985 VSS.n352 VSS.n143 0.0838333
R986 VSS.n234 VSS.n154 0.0838333
R987 VSS.n486 VSS.n485 0.0838333
R988 VSS.n524 VSS.n13 0.0838333
R989 VSS.n453 VSS.n452 0.0838333
R990 VSS.n86 VSS.n85 0.0838333
R991 VSS.n275 VSS.n81 0.0819267
R992 VSS.n417 VSS.n81 0.0819267
R993 VSS.n306 VSS 0.0814556
R994 VSS.n176 VSS 0.0814556
R995 VSS.n470 VSS 0.0814556
R996 VSS.n50 VSS 0.0814556
R997 VSS VSS.n196 0.078625
R998 VSS.n127 VSS.n0 0.0766574
R999 VSS.n75 VSS 0.0747188
R1000 VSS.n362 VSS.n361 0.0708125
R1001 VSS.n267 VSS.n266 0.0708125
R1002 VSS.n534 VSS.n533 0.0708125
R1003 VSS.n351 VSS.n279 0.0680676
R1004 VSS.n351 VSS.n350 0.0680676
R1005 VSS.n318 VSS.n299 0.0680676
R1006 VSS.n318 VSS.n292 0.0680676
R1007 VSS.n261 VSS.n152 0.0680676
R1008 VSS.n263 VSS.n261 0.0680676
R1009 VSS.n195 VSS.n169 0.0680676
R1010 VSS.n195 VSS.n168 0.0680676
R1011 VSS.n451 VSS.n36 0.0680676
R1012 VSS.n451 VSS.n450 0.0680676
R1013 VSS.n523 VSS.n19 0.0680676
R1014 VSS.n523 VSS.n522 0.0680676
R1015 VSS.n484 VSS.n462 0.0680676
R1016 VSS.n484 VSS.n30 0.0680676
R1017 VSS.n420 VSS.n78 0.0680676
R1018 VSS.n82 VSS.n78 0.0680676
R1019 VSS VSS.n319 0.0669062
R1020 VSS.n317 VSS.n298 0.0656042
R1021 VSS.n328 VSS.n291 0.0656042
R1022 VSS.n194 VSS.n170 0.0656042
R1023 VSS.n206 VSS.n167 0.0656042
R1024 VSS.n483 VSS.n461 0.0656042
R1025 VSS.n494 VSS.n29 0.0656042
R1026 VSS.n37 VSS.n35 0.0656042
R1027 VSS.n128 VSS 0.064875
R1028 VSS.n97 VSS 0.064875
R1029 VSS VSS.n566 0.064875
R1030 VSS.n125 VSS 0.063625
R1031 VSS.n354 VSS.n353 0.0603958
R1032 VSS.n271 VSS.n153 0.0603958
R1033 VSS.n271 VSS.n270 0.0603958
R1034 VSS VSS.n21 0.0603958
R1035 VSS.n526 VSS.n521 0.0603958
R1036 VSS.n526 VSS.n525 0.0603958
R1037 VSS.n422 VSS.n76 0.0603958
R1038 VSS.n277 VSS.n145 0.0574697
R1039 VSS.n297 VSS.n293 0.0574697
R1040 VSS.n262 VSS.n150 0.0574697
R1041 VSS.n202 VSS.n201 0.0574697
R1042 VSS.n449 VSS.n34 0.0574697
R1043 VSS.n17 VSS.n15 0.0574697
R1044 VSS.n460 VSS.n31 0.0574697
R1045 VSS.n419 VSS.n79 0.0574697
R1046 VSS.n416 VSS.n80 0.0574697
R1047 VSS.n329 VSS.n328 0.0551875
R1048 VSS.n207 VSS.n206 0.0551875
R1049 VSS.n479 VSS.n461 0.0551875
R1050 VSS.n495 VSS.n494 0.0551875
R1051 VSS.n61 VSS.n35 0.0551875
R1052 VSS.n447 VSS.n446 0.0551875
R1053 VSS.n361 VSS.n140 0.0499792
R1054 VSS.n266 VSS.n260 0.0499792
R1055 VSS.n533 VSS.n10 0.0499792
R1056 VSS.n414 VSS.n413 0.0499792
R1057 VSS.n414 VSS 0.0486771
R1058 VSS.n447 VSS 0.0434688
R1059 VSS.n355 VSS.n279 0.0410405
R1060 VSS.n350 VSS.n144 0.0410405
R1061 VSS.n321 VSS.n299 0.0410405
R1062 VSS.n327 VSS.n292 0.0410405
R1063 VSS.n272 VSS.n152 0.0410405
R1064 VSS.n264 VSS.n263 0.0410405
R1065 VSS.n198 VSS.n169 0.0410405
R1066 VSS.n205 VSS.n168 0.0410405
R1067 VSS.n454 VSS.n36 0.0410405
R1068 VSS.n450 VSS.n448 0.0410405
R1069 VSS.n527 VSS.n19 0.0410405
R1070 VSS.n522 VSS.n14 0.0410405
R1071 VSS.n487 VSS.n462 0.0410405
R1072 VSS.n493 VSS.n30 0.0410405
R1073 VSS.n421 VSS.n420 0.0410405
R1074 VSS.n83 VSS.n82 0.0410405
R1075 VSS VSS.n170 0.0395625
R1076 VSS VSS.n422 0.0382604
R1077 VSS.n308 VSS 0.0356562
R1078 VSS.n354 VSS 0.0356562
R1079 VSS VSS.n222 0.0356562
R1080 VSS.n259 VSS 0.0356562
R1081 VSS.n276 VSS.n275 0.0346274
R1082 VSS.n382 VSS 0.0343542
R1083 VSS.n255 VSS 0.0343542
R1084 VSS.n555 VSS 0.0343542
R1085 VSS.n407 VSS 0.0343542
R1086 VSS.n295 VSS.n32 0.0339875
R1087 VSS VSS.n298 0.0330521
R1088 VSS.n489 VSS.n460 0.0292489
R1089 VSS.n491 VSS.n31 0.0292489
R1090 VSS.n456 VSS.n34 0.0292489
R1091 VSS.n449 VSS.n33 0.0292489
R1092 VSS.n201 VSS.n200 0.0292489
R1093 VSS.n203 VSS.n202 0.0292489
R1094 VSS.n323 VSS.n297 0.0292489
R1095 VSS.n325 VSS.n293 0.0292489
R1096 VSS.n529 VSS.n17 0.0292489
R1097 VSS.n531 VSS.n15 0.0292489
R1098 VSS.n274 VSS.n150 0.0292489
R1099 VSS.n262 VSS.n149 0.0292489
R1100 VSS.n357 VSS.n277 0.0292489
R1101 VSS.n359 VSS.n145 0.0292489
R1102 VSS.n418 VSS.n80 0.0292489
R1103 VSS.n419 VSS.n418 0.0292489
R1104 VSS.n495 VSS.n26 0.0291458
R1105 VSS VSS.n540 0.0291458
R1106 VSS.n446 VSS.n40 0.0291458
R1107 VSS.t27 VSS.n117 0.0282554
R1108 VSS.n329 VSS 0.0252396
R1109 VSS.n334 VSS 0.0252396
R1110 VSS VSS.n339 0.0252396
R1111 VSS VSS.n344 0.0252396
R1112 VSS VSS.n349 0.0252396
R1113 VSS.n349 VSS.n278 0.0239375
R1114 VSS.n353 VSS.n352 0.0239375
R1115 VSS VSS.n368 0.0239375
R1116 VSS.n182 VSS 0.0239375
R1117 VSS.n224 VSS 0.0239375
R1118 VSS.n153 VSS.n151 0.0239375
R1119 VSS.n270 VSS.n154 0.0239375
R1120 VSS.n521 VSS.n18 0.0239375
R1121 VSS.n525 VSS.n524 0.0239375
R1122 VSS.n423 VSS.n75 0.0239375
R1123 VSS.n85 VSS.n76 0.0239375
R1124 VSS.n314 VSS 0.0226354
R1125 VSS VSS.n369 0.0226354
R1126 VSS VSS.n217 0.0226354
R1127 VSS.n219 VSS 0.0226354
R1128 VSS.n260 VSS 0.0226354
R1129 VSS.n252 VSS 0.0226354
R1130 VSS VSS.n238 0.0226354
R1131 VSS.n501 VSS 0.0226354
R1132 VSS.n554 VSS 0.0226354
R1133 VSS VSS.n55 0.0226354
R1134 VSS VSS.n60 0.0226354
R1135 VSS VSS.n38 0.0226354
R1136 VSS.n441 VSS 0.0226354
R1137 VSS VSS.n72 0.0226354
R1138 VSS.n423 VSS 0.0226354
R1139 VSS.n87 VSS 0.0226354
R1140 VSS.n406 VSS 0.0226354
R1141 VSS.n403 VSS 0.0226354
R1142 VSS.n147 VSS 0.0223384
R1143 VSS.n207 VSS 0.0200312
R1144 VSS.n214 VSS 0.0200312
R1145 VSS.n57 VSS 0.0200312
R1146 VSS.n320 VSS.n317 0.0187292
R1147 VSS.n319 VSS.n291 0.0187292
R1148 VSS.n197 VSS.n194 0.0187292
R1149 VSS.n196 VSS.n167 0.0187292
R1150 VSS.n486 VSS.n483 0.0187292
R1151 VSS.n485 VSS.n29 0.0187292
R1152 VSS.n453 VSS.n37 0.0187292
R1153 VSS.n452 VSS.n38 0.0187292
R1154 VSS.n320 VSS 0.0174271
R1155 VSS.n376 VSS 0.016125
R1156 VSS VSS.n181 0.016125
R1157 VSS.n189 VSS 0.016125
R1158 VSS.n472 VSS 0.016125
R1159 VSS.n508 VSS 0.016125
R1160 VSS.n442 VSS 0.016125
R1161 VSS.n362 VSS.n143 0.0135208
R1162 VSS.n267 VSS.n234 0.0135208
R1163 VSS.n534 VSS.n13 0.0135208
R1164 VSS.n87 VSS.n86 0.0135208
R1165 VSS VSS.n164 0.00961458
R1166 VSS.n530 VSS 0.00768471
R1167 VSS.n490 VSS 0.00755
R1168 VSS.n324 VSS.n296 0.00619255
R1169 VSS.n197 VSS 0.00570833
R1170 VSS VSS.n288 0.00440625
R1171 VSS.n417 VSS.n16 0.00109873
R1172 VSS.n459 VSS.n457 0.0010875
R1173 VDD.n488 VDD.n487 8629.41
R1174 VDD.n490 VDD.n484 8629.41
R1175 VDD.n506 VDD.n500 8629.41
R1176 VDD.n509 VDD.n499 8629.41
R1177 VDD.n523 VDD.n517 8629.41
R1178 VDD.n526 VDD.n516 8629.41
R1179 VDD.n537 VDD.n535 8629.41
R1180 VDD.n540 VDD.n534 8629.41
R1181 VDD.n491 VDD.n483 920.471
R1182 VDD.n505 VDD.n501 920.471
R1183 VDD.n522 VDD.n518 920.471
R1184 VDD.n536 VDD.n533 920.471
R1185 VDD.n492 VDD.n491 914.447
R1186 VDD.n501 VDD.n497 914.447
R1187 VDD.n518 VDD.n514 914.447
R1188 VDD.n542 VDD.n533 914.447
R1189 VDD.n53 VDD.t45 804.731
R1190 VDD.n57 VDD.t30 804.731
R1191 VDD.n120 VDD.t18 804.731
R1192 VDD.n123 VDD.t54 804.731
R1193 VDD.n280 VDD.t47 804.731
R1194 VDD.n276 VDD.t15 804.731
R1195 VDD.n14 VDD.t35 804.731
R1196 VDD.n243 VDD.t34 804.731
R1197 VDD.n204 VDD.t33 804.731
R1198 VDD.n209 VDD.t62 804.731
R1199 VDD.n287 VDD.t58 804.731
R1200 VDD.n290 VDD.t40 804.731
R1201 VDD.n431 VDD.t24 804.731
R1202 VDD.n395 VDD.t23 804.731
R1203 VDD.n345 VDD.t66 804.731
R1204 VDD.n348 VDD.t38 804.731
R1205 VDD.n320 VDD.t49 804.731
R1206 VDD.n456 VDD.t21 804.731
R1207 VDD.n459 VDD.t43 804.731
R1208 VDD.n462 VDD.t60 804.731
R1209 VDD.t15 VDD.n275 751.692
R1210 VDD.t49 VDD.n319 751.692
R1211 VDD.t21 VDD.n455 751.692
R1212 VDD.t45 VDD.n52 725.173
R1213 VDD.t30 VDD.n56 725.173
R1214 VDD.t18 VDD.n119 725.173
R1215 VDD.t54 VDD.n122 725.173
R1216 VDD.t47 VDD.n279 725.173
R1217 VDD.t33 VDD.n203 725.173
R1218 VDD.t62 VDD.n208 725.173
R1219 VDD.t58 VDD.n286 725.173
R1220 VDD.t40 VDD.n289 725.173
R1221 VDD.t66 VDD.n344 725.173
R1222 VDD.t38 VDD.n347 725.173
R1223 VDD.t43 VDD.n458 725.173
R1224 VDD.t60 VDD.n461 725.173
R1225 VDD.n63 VDD.t102 701.529
R1226 VDD VDD.t106 697.264
R1227 VDD.n96 VDD.t90 671.408
R1228 VDD.n370 VDD.n342 599.159
R1229 VDD.n341 VDD.n340 594.144
R1230 VDD.n430 VDD.n327 594.144
R1231 VDD.n423 VDD.n330 594.144
R1232 VDD.n437 VDD.n324 594.144
R1233 VDD.n33 VDD.n32 590.973
R1234 VDD.n247 VDD.n246 585
R1235 VDD.n249 VDD.n248 585
R1236 VDD.n379 VDD.n378 585
R1237 VDD.n377 VDD.n376 585
R1238 VDD.n381 VDD.n380 585
R1239 VDD.n389 VDD.n388 585
R1240 VDD.t19 VDD.t41 540.46
R1241 VDD.n485 VDD.n483 480.764
R1242 VDD.n505 VDD.n504 480.764
R1243 VDD.n522 VDD.n521 480.764
R1244 VDD.n536 VDD.n531 480.764
R1245 VDD VDD.t50 394.435
R1246 VDD.n10 VDD.t63 393.002
R1247 VDD.n284 VDD.t64 388.656
R1248 VDD.n325 VDD.t26 388.656
R1249 VDD.n440 VDD.t27 388.656
R1250 VDD.n225 VDD.t55 388.656
R1251 VDD.n232 VDD.t56 388.656
R1252 VDD.n268 VDD.t14 388.656
R1253 VDD.n396 VDD.t51 388.656
R1254 VDD.n407 VDD.t52 388.656
R1255 VDD.n318 VDD.t48 387.682
R1256 VDD.n454 VDD.t20 387.682
R1257 VDD.n51 VDD.t44 380.193
R1258 VDD.n55 VDD.t29 380.193
R1259 VDD.n118 VDD.t17 380.193
R1260 VDD.n121 VDD.t53 380.193
R1261 VDD.n278 VDD.t46 380.193
R1262 VDD.n202 VDD.t32 380.193
R1263 VDD.n207 VDD.t61 380.193
R1264 VDD.n285 VDD.t57 380.193
R1265 VDD.n288 VDD.t39 380.193
R1266 VDD.n343 VDD.t65 380.193
R1267 VDD.n346 VDD.t37 380.193
R1268 VDD.n457 VDD.t42 380.193
R1269 VDD.n460 VDD.t59 380.193
R1270 VDD.n485 VDD.n482 379.2
R1271 VDD.n504 VDD.n503 379.2
R1272 VDD.n521 VDD.n520 379.2
R1273 VDD.n544 VDD.n531 379.2
R1274 VDD VDD.t28 335.69
R1275 VDD VDD.t36 328.976
R1276 VDD.n137 VDD.n98 322.329
R1277 VDD.n165 VDD.n68 317.104
R1278 VDD.n146 VDD.n95 316.515
R1279 VDD.t129 VDD.t93 315.548
R1280 VDD.n78 VDD.n77 312.053
R1281 VDD.n117 VDD.n116 312.053
R1282 VDD.n41 VDD.n40 312.053
R1283 VDD.n166 VDD.n65 312.051
R1284 VDD.n70 VDD.n69 312.051
R1285 VDD.n89 VDD.n80 312.051
R1286 VDD.n151 VDD.n90 312.051
R1287 VDD.n146 VDD.n94 312.051
R1288 VDD.n107 VDD.n106 312.051
R1289 VDD.n237 VDD.n36 312.051
R1290 VDD.n390 VDD.n387 312.051
R1291 VDD.n174 VDD.n61 312.005
R1292 VDD.n16 VDD.t180 310.853
R1293 VDD.n263 VDD.n18 308.755
R1294 VDD.n173 VDD.n62 308.755
R1295 VDD.n231 VDD.n38 308.755
R1296 VDD.n424 VDD.t185 306.735
R1297 VDD.n9 VDD.t103 293.159
R1298 VDD.t173 VDD.t7 281.979
R1299 VDD VDD.t16 280.3
R1300 VDD.n9 VDD.n8 269.485
R1301 VDD VDD.t124 263.517
R1302 VDD VDD.t91 263.517
R1303 VDD VDD.t101 256.803
R1304 VDD.n52 VDD.t193 245.667
R1305 VDD.n56 VDD.t189 245.667
R1306 VDD.n119 VDD.t181 245.667
R1307 VDD.n122 VDD.t177 245.667
R1308 VDD.n279 VDD.t196 245.667
R1309 VDD.n203 VDD.t182 245.667
R1310 VDD.n208 VDD.t188 245.667
R1311 VDD.n286 VDD.t194 245.667
R1312 VDD.n289 VDD.t176 245.667
R1313 VDD.n344 VDD.t190 245.667
R1314 VDD.n347 VDD.t195 245.667
R1315 VDD.n458 VDD.t178 245.667
R1316 VDD.n461 VDD.t183 245.667
R1317 VDD.n144 VDD.t123 245.178
R1318 VDD.n138 VDD.t115 243.508
R1319 VDD.n224 VDD.t160 240.939
R1320 VDD VDD.t116 240.018
R1321 VDD.t81 VDD.t143 234.982
R1322 VDD.n319 VDD.t197 213.148
R1323 VDD.n455 VDD.t179 213.148
R1324 VDD.n281 VDD.t191 210.964
R1325 VDD.n406 VDD.t187 210.964
R1326 VDD.n439 VDD.t184 210.964
R1327 VDD.n136 VDD.t81 209.368
R1328 VDD.t50 VDD 203.093
R1329 VDD VDD.t19 203.093
R1330 VDD.t16 VDD 182.952
R1331 VDD.n316 VDD 182.952
R1332 VDD.t41 VDD 182.952
R1333 VDD VDD.t135 176.238
R1334 VDD.t170 VDD.t67 174.559
R1335 VDD.n248 VDD.n247 159.476
R1336 VDD.n378 VDD.n377 159.476
R1337 VDD.t93 VDD.t168 159.452
R1338 VDD.t116 VDD.t129 159.452
R1339 VDD.t168 VDD.t22 157.774
R1340 VDD.t156 VDD.t3 154.417
R1341 VDD.t145 VDD.t97 151.06
R1342 VDD.t79 VDD.t9 147.703
R1343 VDD.t5 VDD.t69 147.703
R1344 VDD.t67 VDD.t71 147.703
R1345 VDD.t143 VDD.t73 147.703
R1346 VDD.t118 VDD.t133 144.346
R1347 VDD.t75 VDD.t137 142.668
R1348 VDD.t131 VDD.t95 142.668
R1349 VDD.t149 VDD 135.954
R1350 VDD.n34 VDD.n33 132.268
R1351 VDD.n233 VDD.t192 129.344
R1352 VDD.t28 VDD 125.883
R1353 VDD.t36 VDD 125.883
R1354 VDD.t81 VDD 124.206
R1355 VDD.t107 VDD 120.849
R1356 VDD.t166 VDD.t107 120.849
R1357 VDD.t108 VDD.t86 120.849
R1358 VDD VDD.t75 120.849
R1359 VDD.t120 VDD.t166 119.171
R1360 VDD.n275 VDD.t186 118.853
R1361 VDD.n316 VDD 117.492
R1362 VDD.n98 VDD.t113 116.341
R1363 VDD VDD.t145 112.457
R1364 VDD VDD.t164 109.1
R1365 VDD VDD.t5 109.1
R1366 VDD VDD.t156 109.1
R1367 VDD.n317 VDD.n316 106.561
R1368 VDD.t152 VDD.t161 105.743
R1369 VDD.t164 VDD.t11 104.064
R1370 VDD.t77 VDD 102.385
R1371 VDD VDD.t147 100.707
R1372 VDD.n68 VDD.t109 98.5005
R1373 VDD.n95 VDD.t88 98.5005
R1374 VDD.n61 VDD.t167 96.1553
R1375 VDD.n32 VDD.t175 96.1553
R1376 VDD.n342 VDD.t153 96.1553
R1377 VDD.t7 VDD.t141 93.9934
R1378 VDD.t135 VDD.t25 92.315
R1379 VDD VDD.t170 88.9581
R1380 VDD.t139 VDD 88.9581
R1381 VDD.n248 VDD.t105 86.7743
R1382 VDD.n377 VDD.t8 86.7743
R1383 VDD.t114 VDD.t89 80.5659
R1384 VDD.n388 VDD.t132 77.3934
R1385 VDD.n380 VDD.t174 77.3934
R1386 VDD.n340 VDD.t162 77.3934
R1387 VDD.n327 VDD.t117 77.3934
R1388 VDD.n330 VDD.t94 77.3934
R1389 VDD.n324 VDD.t136 77.3934
R1390 VDD.n10 VDD.n9 72.8099
R1391 VDD.t22 VDD 68.8168
R1392 VDD.t25 VDD.t149 67.1383
R1393 VDD.n247 VDD.t128 66.8398
R1394 VDD.n378 VDD.t138 66.8398
R1395 VDD.n493 VDD.n492 66.6358
R1396 VDD.n498 VDD.n497 66.6358
R1397 VDD.n515 VDD.n514 66.6358
R1398 VDD.n543 VDD.n542 66.6358
R1399 VDD.n32 VDD.t155 63.3219
R1400 VDD.n342 VDD.t111 63.3219
R1401 VDD.n488 VDD.n483 61.6672
R1402 VDD.n484 VDD.n480 61.6672
R1403 VDD.n506 VDD.n505 61.6672
R1404 VDD.n510 VDD.n509 61.6672
R1405 VDD.n523 VDD.n522 61.6672
R1406 VDD.n527 VDD.n526 61.6672
R1407 VDD.n537 VDD.n536 61.6672
R1408 VDD.n541 VDD.n540 61.6672
R1409 VDD.n489 VDD.n488 60.9564
R1410 VDD.n486 VDD.n484 60.9564
R1411 VDD.n507 VDD.n506 60.9564
R1412 VDD.n509 VDD.n508 60.9564
R1413 VDD.n524 VDD.n523 60.9564
R1414 VDD.n526 VDD.n525 60.9564
R1415 VDD.n538 VDD.n537 60.9564
R1416 VDD.n540 VDD.n539 60.9564
R1417 VDD.n510 VDD.n498 60.6123
R1418 VDD.n527 VDD.n515 60.6123
R1419 VDD.t89 VDD.t122 60.4245
R1420 VDD.t112 VDD.t114 60.4245
R1421 VDD.n494 VDD.n493 59.4829
R1422 VDD.t161 VDD.t110 58.7461
R1423 VDD.n543 VDD.n532 58.7299
R1424 VDD VDD.t112 57.0676
R1425 VDD.t141 VDD.t152 53.7107
R1426 VDD.t83 VDD 52.0323
R1427 VDD.t9 VDD 52.0323
R1428 VDD.t147 VDD 52.0323
R1429 VDD.t122 VDD 52.0323
R1430 VDD.t110 VDD 52.0323
R1431 VDD.t95 VDD 52.0323
R1432 VDD.t101 VDD 50.3539
R1433 VDD.t71 VDD 50.3539
R1434 VDD.t124 VDD 46.997
R1435 VDD VDD.t139 45.3185
R1436 VDD.t11 VDD.t120 43.6401
R1437 VDD.n388 VDD.t157 41.0422
R1438 VDD.n380 VDD.t76 41.0422
R1439 VDD.n340 VDD.t142 41.0422
R1440 VDD.n327 VDD.t130 41.0422
R1441 VDD.n330 VDD.t169 41.0422
R1442 VDD.n324 VDD.t150 41.0422
R1443 VDD.n490 VDD.n489 38.5759
R1444 VDD.n487 VDD.n486 38.5759
R1445 VDD.n507 VDD.n499 38.5759
R1446 VDD.n508 VDD.n500 38.5759
R1447 VDD.n524 VDD.n516 38.5759
R1448 VDD.n525 VDD.n517 38.5759
R1449 VDD.n538 VDD.n534 38.5759
R1450 VDD.n539 VDD.n535 38.5759
R1451 VDD.n62 VDD.t121 36.1587
R1452 VDD.n62 VDD.t165 36.1587
R1453 VDD.n65 VDD.t84 36.1587
R1454 VDD.n65 VDD.t98 36.1587
R1455 VDD.n69 VDD.t10 36.1587
R1456 VDD.n69 VDD.t80 36.1587
R1457 VDD.n77 VDD.t70 36.1587
R1458 VDD.n77 VDD.t6 36.1587
R1459 VDD.n80 VDD.t148 36.1587
R1460 VDD.n80 VDD.t125 36.1587
R1461 VDD.n90 VDD.t72 36.1587
R1462 VDD.n90 VDD.t68 36.1587
R1463 VDD.n94 VDD.t134 36.1587
R1464 VDD.n94 VDD.t92 36.1587
R1465 VDD.n106 VDD.t144 36.1587
R1466 VDD.n106 VDD.t74 36.1587
R1467 VDD.n116 VDD.t78 36.1587
R1468 VDD.n116 VDD.t140 36.1587
R1469 VDD.n18 VDD.t1 36.1587
R1470 VDD.n18 VDD.t2 36.1587
R1471 VDD.n38 VDD.t100 36.1587
R1472 VDD.n38 VDD.t158 36.1587
R1473 VDD.n40 VDD.t154 36.1587
R1474 VDD.n40 VDD.t126 36.1587
R1475 VDD.n36 VDD.t159 36.1587
R1476 VDD.n36 VDD.t151 36.1587
R1477 VDD.n387 VDD.t96 36.1587
R1478 VDD.n387 VDD.t4 36.1587
R1479 VDD.n173 VDD.n172 34.6358
R1480 VDD.n185 VDD.n58 34.6358
R1481 VDD.n175 VDD.n58 34.6358
R1482 VDD.n168 VDD.n167 34.6358
R1483 VDD.n150 VDD.n92 34.6358
R1484 VDD.n140 VDD.n139 34.6358
R1485 VDD.n136 VDD.n99 34.6358
R1486 VDD.n370 VDD.n369 33.8829
R1487 VDD.n145 VDD.n144 33.5064
R1488 VDD.t87 VDD 31.891
R1489 VDD.n8 VDD 31.4055
R1490 VDD.n98 VDD.t82 28.4453
R1491 VDD.n375 VDD.n374 27.724
R1492 VDD.n386 VDD.n338 27.1064
R1493 VDD.n168 VDD.n63 25.977
R1494 VDD.n61 VDD.t12 25.6105
R1495 VDD.n68 VDD.t146 25.6105
R1496 VDD.n95 VDD.t119 25.6105
R1497 VDD.n165 VDD.n164 25.224
R1498 VDD.n172 VDD.n63 24.0946
R1499 VDD.n153 VDD.n152 24.0946
R1500 VDD.n186 VDD.n185 23.7181
R1501 VDD.n126 VDD.n125 23.7181
R1502 VDD.n211 VDD.n210 23.7181
R1503 VDD.n369 VDD.n349 23.7181
R1504 VDD.n174 VDD.n173 22.5887
R1505 VDD.n167 VDD.n166 22.2123
R1506 VDD.n164 VDD.n70 22.2123
R1507 VDD.n79 VDD.n78 22.2123
R1508 VDD.n89 VDD.n79 22.2123
R1509 VDD.n153 VDD.n89 22.2123
R1510 VDD.n151 VDD.n150 22.2123
R1511 VDD.n146 VDD.n92 22.2123
R1512 VDD.n146 VDD.n145 22.2123
R1513 VDD.n107 VDD.n99 22.2123
R1514 VDD.n126 VDD.n117 22.2123
R1515 VDD.n210 VDD.n41 22.2123
R1516 VDD.n223 VDD.n41 22.2123
R1517 VDD.n238 VDD.n237 22.2123
R1518 VDD.n390 VDD.n386 22.2123
R1519 VDD.n238 VDD.n34 21.4593
R1520 VDD.n224 VDD.n223 21.2076
R1521 VDD VDD.t104 20.1894
R1522 VDD.t133 VDD.t87 20.1418
R1523 VDD.n140 VDD.n96 19.9534
R1524 VDD.n374 VDD.n341 19.9534
R1525 VDD.n138 VDD.n137 18.4476
R1526 VDD.n433 VDD.n432 17.612
R1527 VDD.n394 VDD.n337 17.3741
R1528 VDD.t137 VDD.t173 16.785
R1529 VDD.n137 VDD.n136 15.8123
R1530 VDD.n382 VDD.n381 14.8543
R1531 VDD.n143 VDD.n96 14.6829
R1532 VDD.n371 VDD.n341 14.6829
R1533 VDD.n292 VDD.n291 14.2735
R1534 VDD.n441 VDD.n317 14.2735
R1535 VDD.n152 VDD.n151 13.5534
R1536 VDD.t86 VDD.t83 13.4281
R1537 VDD.t97 VDD.t108 13.4281
R1538 VDD.n464 VDD.n317 12.8005
R1539 VDD.n464 VDD.n463 12.8005
R1540 VDD.n237 VDD.n35 12.7676
R1541 VDD.n175 VDD.n174 12.0476
R1542 VDD.n482 VDD.n481 11.3235
R1543 VDD.n503 VDD.n502 11.3235
R1544 VDD.n520 VDD.n519 11.3235
R1545 VDD.n545 VDD.n544 11.3235
R1546 VDD.n390 VDD.n389 10.5955
R1547 VDD.n166 VDD.n165 10.5417
R1548 VDD.t104 VDD.t0 10.3754
R1549 VDD.n78 VDD.n70 9.78874
R1550 VDD.n117 VDD.n107 9.78874
R1551 VDD.n262 VDD.n19 9.73273
R1552 VDD.n263 VDD.n262 9.73273
R1553 VDD.n264 VDD.n263 9.73273
R1554 VDD.n421 VDD.n331 9.73273
R1555 VDD.n422 VDD.n421 9.73273
R1556 VDD.n425 VDD.n328 9.73273
R1557 VDD.n429 VDD.n328 9.73273
R1558 VDD.n242 VDD.n33 9.6005
R1559 VDD.n186 VDD 9.32264
R1560 VDD.n211 VDD 9.32264
R1561 VDD VDD.n349 9.32264
R1562 VDD.n187 VDD.n186 9.3005
R1563 VDD.n186 VDD.n54 9.3005
R1564 VDD.n185 VDD.n184 9.3005
R1565 VDD.n177 VDD.n58 9.3005
R1566 VDD.n176 VDD.n175 9.3005
R1567 VDD.n173 VDD.n60 9.3005
R1568 VDD.n172 VDD.n171 9.3005
R1569 VDD.n170 VDD.n63 9.3005
R1570 VDD.n169 VDD.n168 9.3005
R1571 VDD.n167 VDD.n64 9.3005
R1572 VDD.n166 VDD.n66 9.3005
R1573 VDD.n165 VDD.n67 9.3005
R1574 VDD.n164 VDD.n163 9.3005
R1575 VDD.n162 VDD.n70 9.3005
R1576 VDD.n78 VDD.n71 9.3005
R1577 VDD.n82 VDD.n79 9.3005
R1578 VDD.n89 VDD.n88 9.3005
R1579 VDD.n154 VDD.n153 9.3005
R1580 VDD.n152 VDD.n76 9.3005
R1581 VDD.n151 VDD.n91 9.3005
R1582 VDD.n150 VDD.n149 9.3005
R1583 VDD.n148 VDD.n92 9.3005
R1584 VDD.n147 VDD.n146 9.3005
R1585 VDD.n145 VDD.n93 9.3005
R1586 VDD.n143 VDD.n142 9.3005
R1587 VDD.n141 VDD.n140 9.3005
R1588 VDD.n139 VDD.n97 9.3005
R1589 VDD.n136 VDD.n135 9.3005
R1590 VDD.n100 VDD.n99 9.3005
R1591 VDD.n109 VDD.n107 9.3005
R1592 VDD.n117 VDD.n115 9.3005
R1593 VDD.n127 VDD.n126 9.3005
R1594 VDD.n212 VDD.n211 9.3005
R1595 VDD.n211 VDD.n206 9.3005
R1596 VDD.n210 VDD.n42 9.3005
R1597 VDD.n221 VDD.n41 9.3005
R1598 VDD.n223 VDD.n222 9.3005
R1599 VDD.n227 VDD.n226 9.3005
R1600 VDD.n228 VDD.n39 9.3005
R1601 VDD.n230 VDD.n229 9.3005
R1602 VDD.n231 VDD.n37 9.3005
R1603 VDD.n234 VDD.n233 9.3005
R1604 VDD.n235 VDD.n35 9.3005
R1605 VDD.n237 VDD.n236 9.3005
R1606 VDD.n239 VDD.n238 9.3005
R1607 VDD.n241 VDD.n240 9.3005
R1608 VDD.n244 VDD.n27 9.3005
R1609 VDD.n251 VDD.n250 9.3005
R1610 VDD.n245 VDD.n20 9.3005
R1611 VDD.n260 VDD.n19 9.3005
R1612 VDD.n262 VDD.n261 9.3005
R1613 VDD.n263 VDD.n17 9.3005
R1614 VDD.n265 VDD.n264 9.3005
R1615 VDD.n267 VDD.n266 9.3005
R1616 VDD.n269 VDD.n15 9.3005
R1617 VDD.n271 VDD.n270 9.3005
R1618 VDD.n273 VDD.n272 9.3005
R1619 VDD.n277 VDD.n13 9.3005
R1620 VDD.n277 VDD.n11 9.3005
R1621 VDD.n304 VDD.n303 9.3005
R1622 VDD.n302 VDD.n301 9.3005
R1623 VDD.n293 VDD.n292 9.3005
R1624 VDD.n359 VDD.n349 9.3005
R1625 VDD.n360 VDD.n349 9.3005
R1626 VDD.n369 VDD.n368 9.3005
R1627 VDD.n372 VDD.n371 9.3005
R1628 VDD.n374 VDD.n373 9.3005
R1629 VDD.n375 VDD.n339 9.3005
R1630 VDD.n383 VDD.n382 9.3005
R1631 VDD.n384 VDD.n338 9.3005
R1632 VDD.n386 VDD.n385 9.3005
R1633 VDD.n391 VDD.n390 9.3005
R1634 VDD.n392 VDD.n337 9.3005
R1635 VDD.n394 VDD.n393 9.3005
R1636 VDD.n398 VDD.n397 9.3005
R1637 VDD.n399 VDD.n336 9.3005
R1638 VDD.n405 VDD.n404 9.3005
R1639 VDD.n409 VDD.n408 9.3005
R1640 VDD.n410 VDD.n331 9.3005
R1641 VDD.n421 VDD.n420 9.3005
R1642 VDD.n422 VDD.n329 9.3005
R1643 VDD.n426 VDD.n425 9.3005
R1644 VDD.n427 VDD.n328 9.3005
R1645 VDD.n429 VDD.n428 9.3005
R1646 VDD.n432 VDD.n326 9.3005
R1647 VDD.n434 VDD.n433 9.3005
R1648 VDD.n436 VDD.n435 9.3005
R1649 VDD.n438 VDD.n323 9.3005
R1650 VDD.n442 VDD.n441 9.3005
R1651 VDD.n443 VDD.n317 9.3005
R1652 VDD.n464 VDD.n453 9.3005
R1653 VDD.n464 VDD.n322 9.3005
R1654 VDD.n464 VDD.n321 9.3005
R1655 VDD.n465 VDD.n464 9.3005
R1656 VDD.n244 VDD.n243 9.09802
R1657 VDD.n245 VDD.n19 8.80773
R1658 VDD.n250 VDD.n244 8.57648
R1659 VDD.n532 VDD.n530 8.23557
R1660 VDD.n431 VDD.n430 7.93438
R1661 VDD.n408 VDD.n331 7.75995
R1662 VDD.n397 VDD.n395 7.12524
R1663 VDD.n379 VDD.n376 6.8005
R1664 VDD.t69 VDD.t79 6.71428
R1665 VDD.t73 VDD.t77 6.71428
R1666 VDD.n492 VDD.n480 6.02403
R1667 VDD.n542 VDD.n541 6.02403
R1668 VDD.n8 VDD.t99 5.88893
R1669 VDD.n425 VDD.n424 5.18397
R1670 VDD.t3 VDD.t131 5.03584
R1671 VDD.n511 VDD.n510 4.89462
R1672 VDD.n528 VDD.n514 4.89462
R1673 VDD.n230 VDD.n39 4.67352
R1674 VDD.n231 VDD.n230 4.67352
R1675 VDD.n233 VDD.n231 4.67352
R1676 VDD.n303 VDD.n302 4.67352
R1677 VDD.n277 VDD.n12 4.62124
R1678 VDD.n161 VDD.n160 4.51401
R1679 VDD.n156 VDD.n155 4.51401
R1680 VDD.n134 VDD.n133 4.51401
R1681 VDD.n129 VDD.n128 4.51401
R1682 VDD.n190 VDD.n48 4.51401
R1683 VDD.n183 VDD.n182 4.51401
R1684 VDD.n254 VDD.n25 4.51401
R1685 VDD.n259 VDD.n258 4.51401
R1686 VDD.n307 VDD.n6 4.51401
R1687 VDD.n298 VDD.n294 4.51401
R1688 VDD.n215 VDD.n197 4.51401
R1689 VDD.n220 VDD.n219 4.51401
R1690 VDD.n356 VDD.n354 4.51401
R1691 VDD.n367 VDD.n366 4.51401
R1692 VDD.n445 VDD.n444 4.51401
R1693 VDD.n467 VDD.n466 4.51401
R1694 VDD.n403 VDD.n402 4.51401
R1695 VDD.n81 VDD.n72 4.5005
R1696 VDD.n86 VDD.n85 4.5005
R1697 VDD.n87 VDD.n75 4.5005
R1698 VDD.n108 VDD.n101 4.5005
R1699 VDD.n113 VDD.n112 4.5005
R1700 VDD.n114 VDD.n105 4.5005
R1701 VDD.n189 VDD.n188 4.5005
R1702 VDD.n178 VDD.n50 4.5005
R1703 VDD.n181 VDD.n59 4.5005
R1704 VDD.n253 VDD.n252 4.5005
R1705 VDD.n31 VDD.n30 4.5005
R1706 VDD.n28 VDD.n21 4.5005
R1707 VDD.n306 VDD.n305 4.5005
R1708 VDD.n295 VDD.n282 4.5005
R1709 VDD.n300 VDD.n299 4.5005
R1710 VDD.n214 VDD.n213 4.5005
R1711 VDD.n201 VDD.n200 4.5005
R1712 VDD.n205 VDD.n43 4.5005
R1713 VDD.n358 VDD.n357 4.5005
R1714 VDD.n362 VDD.n361 4.5005
R1715 VDD.n351 VDD.n350 4.5005
R1716 VDD.n452 VDD.n451 4.5005
R1717 VDD.n448 VDD.n447 4.5005
R1718 VDD.n314 VDD.n313 4.5005
R1719 VDD.n400 VDD.n335 4.5005
R1720 VDD.n413 VDD.n412 4.5005
R1721 VDD.n411 VDD.n332 4.5005
R1722 VDD.n419 VDD.n418 4.5005
R1723 VDD.n264 VDD.n16 4.47065
R1724 VDD.n225 VDD.n39 4.36875
R1725 VDD.n233 VDD.n232 4.36875
R1726 VDD.n436 VDD.n325 4.36875
R1727 VDD.n152 VDD 4.26717
R1728 VDD.n424 VDD.n423 4.12612
R1729 VDD.n249 VDD.n246 4.04887
R1730 VDD.n186 VDD.n53 4.02033
R1731 VDD.n186 VDD.n57 4.02033
R1732 VDD.n125 VDD.n120 4.02033
R1733 VDD.n125 VDD.n123 4.02033
R1734 VDD.n211 VDD.n204 4.02033
R1735 VDD.n211 VDD.n209 4.02033
R1736 VDD.n291 VDD.n287 4.02033
R1737 VDD.n291 VDD.n290 4.02033
R1738 VDD.n349 VDD.n345 4.02033
R1739 VDD.n349 VDD.n348 4.02033
R1740 VDD.n463 VDD.n459 4.02033
R1741 VDD.n463 VDD.n462 4.02033
R1742 VDD.t31 VDD.t103 3.64572
R1743 VDD.t13 VDD.t127 3.64572
R1744 VDD.n270 VDD.n269 3.47425
R1745 VDD.n405 VDD.n336 3.47425
R1746 VDD.n157 VDD.n156 3.43925
R1747 VDD.n160 VDD.n159 3.43925
R1748 VDD.n130 VDD.n129 3.43925
R1749 VDD.n133 VDD.n132 3.43925
R1750 VDD.n182 VDD.n46 3.43925
R1751 VDD.n191 VDD.n190 3.43925
R1752 VDD.n258 VDD.n257 3.43925
R1753 VDD.n255 VDD.n254 3.43925
R1754 VDD.n298 VDD.n4 3.43925
R1755 VDD.n308 VDD.n307 3.43925
R1756 VDD.n219 VDD.n218 3.43925
R1757 VDD.n216 VDD.n215 3.43925
R1758 VDD.n366 VDD.n365 3.43925
R1759 VDD.n356 VDD.n355 3.43925
R1760 VDD.n417 VDD.n416 3.43925
R1761 VDD.n402 VDD.n401 3.43925
R1762 VDD.n83 VDD.n73 3.4105
R1763 VDD.n84 VDD.n74 3.4105
R1764 VDD.n110 VDD.n102 3.4105
R1765 VDD.n111 VDD.n104 3.4105
R1766 VDD.n49 VDD.n47 3.4105
R1767 VDD.n180 VDD.n179 3.4105
R1768 VDD.n26 VDD.n24 3.4105
R1769 VDD.n29 VDD.n22 3.4105
R1770 VDD.n7 VDD.n5 3.4105
R1771 VDD.n297 VDD.n296 3.4105
R1772 VDD.n198 VDD.n196 3.4105
R1773 VDD.n199 VDD.n44 3.4105
R1774 VDD.n353 VDD.n352 3.4105
R1775 VDD.n364 VDD.n363 3.4105
R1776 VDD.n469 VDD.n468 3.4105
R1777 VDD.n469 VDD.n311 3.4105
R1778 VDD.n468 VDD.n467 3.4105
R1779 VDD.n445 VDD.n311 3.4105
R1780 VDD.n450 VDD.n449 3.4105
R1781 VDD.n446 VDD.n312 3.4105
R1782 VDD.n334 VDD.n333 3.4105
R1783 VDD.n415 VDD.n414 3.4105
R1784 VDD.t91 VDD.t118 3.35739
R1785 VDD.n269 VDD.n268 3.2477
R1786 VDD.n270 VDD.n14 3.2477
R1787 VDD.n396 VDD.n336 3.2477
R1788 VDD.n512 VDD.n511 3.23917
R1789 VDD.n529 VDD.n528 3.23136
R1790 VDD.n495 VDD.n494 3.22655
R1791 VDD.n267 VDD.n16 3.219
R1792 VDD.n303 VDD.n277 3.2005
R1793 VDD.n302 VDD.n280 3.12116
R1794 VDD.n241 VDD.n34 3.06827
R1795 VDD.n125 VDD.n124 3.04861
R1796 VDD.n291 VDD.n283 3.04861
R1797 VDD.n463 VDD.n315 3.04861
R1798 VDD.n464 VDD.n320 2.91308
R1799 VDD.n464 VDD.n456 2.91308
R1800 VDD.n277 VDD.n276 2.87861
R1801 VDD.n491 VDD.n490 2.84665
R1802 VDD.n487 VDD.n485 2.84665
R1803 VDD.n501 VDD.n499 2.84665
R1804 VDD.n504 VDD.n500 2.84665
R1805 VDD.n518 VDD.n516 2.84665
R1806 VDD.n521 VDD.n517 2.84665
R1807 VDD.n534 VDD.n533 2.84665
R1808 VDD.n535 VDD.n531 2.84665
R1809 VDD.n437 VDD.n436 2.74336
R1810 VDD.n53 VDD.n51 2.63539
R1811 VDD.n57 VDD.n55 2.63539
R1812 VDD.n120 VDD.n118 2.63539
R1813 VDD.n123 VDD.n121 2.63539
R1814 VDD.n280 VDD.n278 2.63539
R1815 VDD.n204 VDD.n202 2.63539
R1816 VDD.n209 VDD.n207 2.63539
R1817 VDD.n287 VDD.n285 2.63539
R1818 VDD.n290 VDD.n288 2.63539
R1819 VDD.n345 VDD.n343 2.63539
R1820 VDD.n348 VDD.n346 2.63539
R1821 VDD.n459 VDD.n457 2.63539
R1822 VDD.n462 VDD.n460 2.63539
R1823 VDD.n274 VDD.n273 2.63233
R1824 VDD.n275 VDD.n274 2.61352
R1825 VDD.n56 VDD.n55 2.37495
R1826 VDD.n52 VDD.n51 2.37495
R1827 VDD.n122 VDD.n121 2.37495
R1828 VDD.n119 VDD.n118 2.37495
R1829 VDD.n279 VDD.n278 2.37495
R1830 VDD.n208 VDD.n207 2.37495
R1831 VDD.n203 VDD.n202 2.37495
R1832 VDD.n289 VDD.n288 2.37495
R1833 VDD.n286 VDD.n285 2.37495
R1834 VDD.n347 VDD.n346 2.37495
R1835 VDD.n344 VDD.n343 2.37495
R1836 VDD.n461 VDD.n460 2.37495
R1837 VDD.n458 VDD.n457 2.37495
R1838 VDD.n302 VDD.n281 2.33701
R1839 VDD.n439 VDD.n438 2.33701
R1840 VDD.n493 VDD.n482 2.28169
R1841 VDD.n503 VDD.n498 2.28169
R1842 VDD.n520 VDD.n515 2.28169
R1843 VDD.n544 VDD.n543 2.28169
R1844 VDD.t99 VDD.t31 2.24371
R1845 VDD.t0 VDD.t13 2.24371
R1846 VDD.n284 VDD.n281 2.03225
R1847 VDD.n440 VDD.n439 2.03225
R1848 VDD.n320 VDD.n318 2.01703
R1849 VDD.n456 VDD.n454 2.01703
R1850 VDD.n438 VDD.n437 1.93066
R1851 VDD.n455 VDD.n454 1.88416
R1852 VDD.n319 VDD.n318 1.88416
R1853 VDD.n541 VDD.n532 1.88285
R1854 VDD.n406 VDD.n405 1.73737
R1855 VDD.n365 VDD.n0 1.69188
R1856 VDD.n355 VDD.n0 1.69188
R1857 VDD.n218 VDD.n217 1.69188
R1858 VDD.n217 VDD.n216 1.69188
R1859 VDD.n192 VDD.n46 1.69188
R1860 VDD.n192 VDD.n191 1.69188
R1861 VDD.n309 VDD.n4 1.69188
R1862 VDD.n309 VDD.n308 1.69188
R1863 VDD.n131 VDD.n130 1.69188
R1864 VDD.n132 VDD.n131 1.69188
R1865 VDD.n469 VDD.n310 1.69188
R1866 VDD.n416 VDD.n2 1.69188
R1867 VDD.n401 VDD.n2 1.69188
R1868 VDD.n257 VDD.n256 1.69188
R1869 VDD.n256 VDD.n255 1.69188
R1870 VDD.n158 VDD.n157 1.69188
R1871 VDD.n159 VDD.n158 1.69188
R1872 VDD.n407 VDD.n406 1.51082
R1873 VDD.n382 VDD.n379 1.4005
R1874 VDD.n479 VDD.n478 1.38219
R1875 VDD.n276 VDD.n274 1.2502
R1876 VDD.n430 VDD.n429 1.16414
R1877 VDD.n502 VDD.n496 1.143
R1878 VDD.n519 VDD.n513 1.143
R1879 VDD.n481 VDD.n479 1.13977
R1880 VDD.n545 VDD.n530 1.13675
R1881 VDD.n144 VDD.n143 1.12991
R1882 VDD.n494 VDD.n480 1.12991
R1883 VDD.n511 VDD.n497 1.12991
R1884 VDD.n528 VDD.n527 1.12991
R1885 VDD.n381 VDD.n338 1.07613
R1886 VDD.n376 VDD.n375 1.0005
R1887 VDD.n513 VDD.n512 0.862816
R1888 VDD.n246 VDD.n245 0.833988
R1889 VDD.n495 VDD.n479 0.823939
R1890 VDD.n530 VDD.n529 0.770881
R1891 VDD.n371 VDD.n370 0.753441
R1892 VDD.n496 VDD.n495 0.729231
R1893 VDD.n472 VDD 0.660687
R1894 VDD.n395 VDD.n394 0.635211
R1895 VDD.n432 VDD.n431 0.635211
R1896 VDD.n250 VDD.n249 0.595849
R1897 VDD.n192 VDD.n45 0.55065
R1898 VDD.n243 VDD.n242 0.529426
R1899 VDD.n476 VDD.n475 0.500125
R1900 VDD.n195 VDD.n194 0.500125
R1901 VDD.n478 VDD 0.467141
R1902 VDD VDD.n472 0.466259
R1903 VDD.n131 VDD.n103 0.431025
R1904 VDD.n158 VDD.n45 0.431025
R1905 VDD.n423 VDD.n422 0.42364
R1906 VDD.n529 VDD.n513 0.392323
R1907 VDD.n193 VDD.n3 0.3805
R1908 VDD.n470 VDD.n1 0.3805
R1909 VDD.n194 VDD.n23 0.3805
R1910 VDD.n475 VDD.n474 0.3805
R1911 VDD.n139 VDD.n138 0.376971
R1912 VDD.n512 VDD.n496 0.360318
R1913 VDD.n389 VDD.n337 0.323189
R1914 VDD.n226 VDD.n225 0.305262
R1915 VDD.n232 VDD.n35 0.305262
R1916 VDD.n292 VDD.n284 0.305262
R1917 VDD.n433 VDD.n325 0.305262
R1918 VDD.n441 VDD.n440 0.305262
R1919 VDD.n489 VDD.t171 0.27666
R1920 VDD.n486 VDD.t171 0.27666
R1921 VDD.t85 VDD.n507 0.27666
R1922 VDD.n508 VDD.t85 0.27666
R1923 VDD.t172 VDD.n524 0.27666
R1924 VDD.n525 VDD.t172 0.27666
R1925 VDD.t163 VDD.n538 0.27666
R1926 VDD.n539 VDD.t163 0.27666
R1927 VDD.n293 VDD.n283 0.239726
R1928 VDD.n465 VDD.n315 0.239726
R1929 VDD.n268 VDD.n267 0.227049
R1930 VDD.n273 VDD.n14 0.227049
R1931 VDD.n397 VDD.n396 0.227049
R1932 VDD.n408 VDD.n407 0.227049
R1933 VDD.n124 VDD 0.217591
R1934 VDD.n226 VDD.n224 0.209973
R1935 VDD.n472 VDD 0.168795
R1936 VDD.n217 VDD.n0 0.1603
R1937 VDD.n469 VDD.n309 0.1603
R1938 VDD.n256 VDD.n2 0.1603
R1939 VDD VDD.n12 0.145148
R1940 VDD.n195 VDD.n192 0.14385
R1941 VDD.n131 VDD.n3 0.14385
R1942 VDD.n158 VDD.n23 0.14385
R1943 VDD.n124 VDD 0.141725
R1944 VDD.n283 VDD 0.141725
R1945 VDD.n315 VDD 0.141725
R1946 VDD.n277 VDD.n10 0.140696
R1947 VDD.n177 VDD.n176 0.120292
R1948 VDD.n176 VDD.n60 0.120292
R1949 VDD.n171 VDD.n60 0.120292
R1950 VDD.n169 VDD.n64 0.120292
R1951 VDD.n67 VDD.n66 0.120292
R1952 VDD.n163 VDD.n67 0.120292
R1953 VDD.n154 VDD.n76 0.120292
R1954 VDD.n149 VDD.n91 0.120292
R1955 VDD.n149 VDD.n148 0.120292
R1956 VDD.n147 VDD.n93 0.120292
R1957 VDD.n142 VDD.n93 0.120292
R1958 VDD.n141 VDD.n97 0.120292
R1959 VDD.n229 VDD.n37 0.120292
R1960 VDD.n234 VDD.n37 0.120292
R1961 VDD.n236 VDD.n235 0.120292
R1962 VDD.n261 VDD.n260 0.120292
R1963 VDD.n261 VDD.n17 0.120292
R1964 VDD.n265 VDD.n17 0.120292
R1965 VDD.n271 VDD.n15 0.120292
R1966 VDD.n272 VDD.n271 0.120292
R1967 VDD.n272 VDD.n13 0.120292
R1968 VDD.n373 VDD.n372 0.120292
R1969 VDD.n373 VDD.n339 0.120292
R1970 VDD.n383 VDD.n339 0.120292
R1971 VDD.n384 VDD.n383 0.120292
R1972 VDD.n385 VDD.n384 0.120292
R1973 VDD.n392 VDD.n391 0.120292
R1974 VDD.n393 VDD.n392 0.120292
R1975 VDD.n420 VDD.n329 0.120292
R1976 VDD.n426 VDD.n329 0.120292
R1977 VDD.n427 VDD.n426 0.120292
R1978 VDD.n428 VDD.n427 0.120292
R1979 VDD.n428 VDD.n326 0.120292
R1980 VDD.n434 VDD.n326 0.120292
R1981 VDD.n435 VDD.n323 0.120292
R1982 VDD.n442 VDD.n323 0.120292
R1983 VDD.n475 VDD.n1 0.120125
R1984 VDD.n194 VDD.n193 0.120125
R1985 VDD.n103 VDD.n45 0.120125
R1986 VDD.n242 VDD.n241 0.106285
R1987 VDD.n221 VDD 0.104667
R1988 VDD.n229 VDD 0.104667
R1989 VDD.n239 VDD 0.104667
R1990 VDD.n12 VDD 0.098273
R1991 VDD VDD.n170 0.0981562
R1992 VDD.n66 VDD 0.0981562
R1993 VDD VDD.n162 0.0981562
R1994 VDD VDD.n147 0.0981562
R1995 VDD VDD.n141 0.0981562
R1996 VDD.n227 VDD 0.0981562
R1997 VDD.n228 VDD 0.0981562
R1998 VDD.n235 VDD 0.0981562
R1999 VDD.n240 VDD 0.0981562
R2000 VDD.n266 VDD 0.0981562
R2001 VDD VDD.n15 0.0981562
R2002 VDD.n372 VDD 0.0981562
R2003 VDD.n391 VDD 0.0981562
R2004 VDD.n398 VDD 0.0981562
R2005 VDD.n399 VDD 0.0981562
R2006 VDD.n435 VDD 0.0981562
R2007 VDD.n91 VDD 0.0968542
R2008 VDD.n135 VDD 0.0968542
R2009 VDD.n222 VDD 0.0968542
R2010 VDD.n160 VDD.n72 0.0950946
R2011 VDD.n156 VDD.n75 0.0950946
R2012 VDD.n133 VDD.n101 0.0950946
R2013 VDD.n129 VDD.n105 0.0950946
R2014 VDD.n190 VDD.n189 0.0950946
R2015 VDD.n182 VDD.n181 0.0950946
R2016 VDD.n254 VDD.n253 0.0950946
R2017 VDD.n258 VDD.n21 0.0950946
R2018 VDD.n307 VDD.n306 0.0950946
R2019 VDD.n299 VDD.n298 0.0950946
R2020 VDD.n215 VDD.n214 0.0950946
R2021 VDD.n219 VDD.n43 0.0950946
R2022 VDD.n357 VDD.n356 0.0950946
R2023 VDD.n366 VDD.n351 0.0950946
R2024 VDD.n451 VDD.n445 0.0950946
R2025 VDD.n467 VDD.n313 0.0950946
R2026 VDD.n402 VDD.n400 0.0950946
R2027 VDD.n417 VDD.n332 0.0950946
R2028 VDD.n443 VDD 0.0916458
R2029 VDD VDD.n177 0.0851354
R2030 VDD VDD.n169 0.0851354
R2031 VDD.n188 VDD.n48 0.0838333
R2032 VDD.n213 VDD.n197 0.0838333
R2033 VDD.n31 VDD.n28 0.0838333
R2034 VDD.n300 VDD.n294 0.0838333
R2035 VDD.n358 VDD.n354 0.0838333
R2036 VDD.n412 VDD.n411 0.0838333
R2037 VDD.n466 VDD.n314 0.0838333
R2038 VDD.n187 VDD.n50 0.0812292
R2039 VDD.n82 VDD.n81 0.0812292
R2040 VDD.n108 VDD.n100 0.0812292
R2041 VDD.n212 VDD.n201 0.0812292
R2042 VDD.n252 VDD.n251 0.0812292
R2043 VDD.n361 VDD.n359 0.0812292
R2044 VDD.n409 VDD.n335 0.0812292
R2045 VDD VDD.n134 0.0799271
R2046 VDD VDD.n6 0.0799271
R2047 VDD.n444 VDD 0.0799271
R2048 VDD.n184 VDD.n59 0.0760208
R2049 VDD.n162 VDD.n161 0.0760208
R2050 VDD.n115 VDD.n113 0.0760208
R2051 VDD.n205 VDD.n42 0.0760208
R2052 VDD.n301 VDD.n282 0.0760208
R2053 VDD.n368 VDD.n350 0.0760208
R2054 VDD.n403 VDD.n399 0.0760208
R2055 VDD.n447 VDD.n321 0.0760208
R2056 VDD.n155 VDD.n154 0.0708125
R2057 VDD.n260 VDD.n259 0.0708125
R2058 VDD.n420 VDD.n419 0.0708125
R2059 VDD.n128 VDD 0.0695104
R2060 VDD.n85 VDD.n83 0.0680676
R2061 VDD.n85 VDD.n84 0.0680676
R2062 VDD.n112 VDD.n110 0.0680676
R2063 VDD.n112 VDD.n111 0.0680676
R2064 VDD.n178 VDD.n49 0.0680676
R2065 VDD.n180 VDD.n178 0.0680676
R2066 VDD.n30 VDD.n26 0.0680676
R2067 VDD.n30 VDD.n29 0.0680676
R2068 VDD.n295 VDD.n7 0.0680676
R2069 VDD.n297 VDD.n295 0.0680676
R2070 VDD.n200 VDD.n198 0.0680676
R2071 VDD.n200 VDD.n199 0.0680676
R2072 VDD.n362 VDD.n353 0.0680676
R2073 VDD.n363 VDD.n362 0.0680676
R2074 VDD.n450 VDD.n448 0.0680676
R2075 VDD.n448 VDD.n446 0.0680676
R2076 VDD.n413 VDD.n334 0.0680676
R2077 VDD.n414 VDD.n413 0.0680676
R2078 VDD.n87 VDD 0.0643021
R2079 VDD.n481 VDD 0.06425
R2080 VDD.n502 VDD 0.06425
R2081 VDD.n519 VDD 0.06425
R2082 VDD VDD.n545 0.06425
R2083 VDD.n305 VDD 0.0590938
R2084 VDD VDD.n452 0.0590938
R2085 VDD.n74 VDD.n73 0.0574697
R2086 VDD.n104 VDD.n102 0.0574697
R2087 VDD.n179 VDD.n47 0.0574697
R2088 VDD.n24 VDD.n22 0.0574697
R2089 VDD.n296 VDD.n5 0.0574697
R2090 VDD.n196 VDD.n44 0.0574697
R2091 VDD.n364 VDD.n352 0.0574697
R2092 VDD.n449 VDD.n311 0.0574697
R2093 VDD.n468 VDD.n312 0.0574697
R2094 VDD.n415 VDD.n333 0.0574697
R2095 VDD VDD.n25 0.0538854
R2096 VDD.n259 VDD.n20 0.0499792
R2097 VDD.n1 VDD 0.047625
R2098 VDD.n193 VDD 0.047625
R2099 VDD.n103 VDD 0.047625
R2100 VDD.n477 VDD 0.0472062
R2101 VDD.n471 VDD 0.0472062
R2102 VDD.n473 VDD 0.0472062
R2103 VDD VDD.n477 0.0469161
R2104 VDD VDD.n471 0.0469161
R2105 VDD.n473 VDD 0.0469161
R2106 VDD.n59 VDD.n54 0.0447708
R2107 VDD.n161 VDD.n71 0.0447708
R2108 VDD.n113 VDD.n109 0.0447708
R2109 VDD.n206 VDD.n205 0.0447708
R2110 VDD.n27 VDD.n25 0.0447708
R2111 VDD.n360 VDD.n350 0.0447708
R2112 VDD.n404 VDD.n403 0.0447708
R2113 VDD.n447 VDD.n322 0.0447708
R2114 VDD.n83 VDD.n72 0.0410405
R2115 VDD.n84 VDD.n75 0.0410405
R2116 VDD.n110 VDD.n101 0.0410405
R2117 VDD.n111 VDD.n105 0.0410405
R2118 VDD.n189 VDD.n49 0.0410405
R2119 VDD.n181 VDD.n180 0.0410405
R2120 VDD.n253 VDD.n26 0.0410405
R2121 VDD.n29 VDD.n21 0.0410405
R2122 VDD.n306 VDD.n7 0.0410405
R2123 VDD.n299 VDD.n297 0.0410405
R2124 VDD.n214 VDD.n198 0.0410405
R2125 VDD.n199 VDD.n43 0.0410405
R2126 VDD.n357 VDD.n353 0.0410405
R2127 VDD.n363 VDD.n351 0.0410405
R2128 VDD.n451 VDD.n450 0.0410405
R2129 VDD.n446 VDD.n313 0.0410405
R2130 VDD.n400 VDD.n334 0.0410405
R2131 VDD.n414 VDD.n332 0.0410405
R2132 VDD.n54 VDD.n50 0.0395625
R2133 VDD.n81 VDD.n71 0.0395625
R2134 VDD.n109 VDD.n108 0.0395625
R2135 VDD.n206 VDD.n201 0.0395625
R2136 VDD.n252 VDD.n27 0.0395625
R2137 VDD.n305 VDD.n304 0.0395625
R2138 VDD.n361 VDD.n360 0.0395625
R2139 VDD.n404 VDD.n335 0.0395625
R2140 VDD.n452 VDD.n322 0.0395625
R2141 VDD.n135 VDD 0.0382604
R2142 VDD VDD.n443 0.0382604
R2143 VDD.n88 VDD 0.0356562
R2144 VDD.n13 VDD 0.0356562
R2145 VDD.n88 VDD.n87 0.0343542
R2146 VDD.n28 VDD.n20 0.0343542
R2147 VDD.n411 VDD.n410 0.0343542
R2148 VDD.n419 VDD 0.0343542
R2149 VDD.n355 VDD.n352 0.0292489
R2150 VDD.n365 VDD.n364 0.0292489
R2151 VDD.n216 VDD.n196 0.0292489
R2152 VDD.n218 VDD.n44 0.0292489
R2153 VDD.n191 VDD.n47 0.0292489
R2154 VDD.n179 VDD.n46 0.0292489
R2155 VDD.n308 VDD.n5 0.0292489
R2156 VDD.n296 VDD.n4 0.0292489
R2157 VDD.n132 VDD.n102 0.0292489
R2158 VDD.n130 VDD.n104 0.0292489
R2159 VDD.n312 VDD.n310 0.0292489
R2160 VDD.n449 VDD.n310 0.0292489
R2161 VDD.n401 VDD.n333 0.0292489
R2162 VDD.n416 VDD.n415 0.0292489
R2163 VDD.n255 VDD.n24 0.0292489
R2164 VDD.n257 VDD.n22 0.0292489
R2165 VDD.n159 VDD.n73 0.0292489
R2166 VDD.n157 VDD.n74 0.0292489
R2167 VDD.n128 VDD.n127 0.0291458
R2168 VDD.n294 VDD.n293 0.0291458
R2169 VDD VDD.n442 0.0291458
R2170 VDD.n466 VDD.n465 0.0291458
R2171 VDD.n170 VDD 0.0239375
R2172 VDD VDD.n76 0.0239375
R2173 VDD VDD.n97 0.0239375
R2174 VDD VDD.n221 0.0239375
R2175 VDD.n478 VDD 0.0231242
R2176 VDD.n477 VDD.n476 0.0231188
R2177 VDD.n471 VDD.n470 0.0231188
R2178 VDD.n474 VDD.n473 0.0231188
R2179 VDD.n171 VDD 0.0226354
R2180 VDD VDD.n64 0.0226354
R2181 VDD.n163 VDD 0.0226354
R2182 VDD.n148 VDD 0.0226354
R2183 VDD.n142 VDD 0.0226354
R2184 VDD.n222 VDD 0.0226354
R2185 VDD VDD.n227 0.0226354
R2186 VDD VDD.n234 0.0226354
R2187 VDD VDD.n239 0.0226354
R2188 VDD.n240 VDD 0.0226354
R2189 VDD VDD.n265 0.0226354
R2190 VDD.n266 VDD 0.0226354
R2191 VDD.n11 VDD 0.0226354
R2192 VDD.n304 VDD 0.0226354
R2193 VDD.n282 VDD 0.0226354
R2194 VDD.n385 VDD 0.0226354
R2195 VDD.n393 VDD 0.0226354
R2196 VDD VDD.n398 0.0226354
R2197 VDD VDD.n434 0.0226354
R2198 VDD.n453 VDD 0.0226354
R2199 VDD VDD.n86 0.0200312
R2200 VDD.n476 VDD.n0 0.018125
R2201 VDD.n470 VDD.n469 0.018125
R2202 VDD.n474 VDD.n2 0.018125
R2203 VDD.n217 VDD.n195 0.01695
R2204 VDD.n309 VDD.n3 0.01695
R2205 VDD.n256 VDD.n23 0.01695
R2206 VDD.n127 VDD 0.016125
R2207 VDD VDD.n228 0.016125
R2208 VDD.n236 VDD 0.016125
R2209 VDD.n410 VDD 0.016125
R2210 VDD.n183 VDD 0.0148229
R2211 VDD.n155 VDD 0.0148229
R2212 VDD.n114 VDD 0.0148229
R2213 VDD.n418 VDD.n417 0.0140135
R2214 VDD.n418 VDD 0.0140135
R2215 VDD VDD.n48 0.0122188
R2216 VDD VDD.n197 0.0122188
R2217 VDD.n354 VDD 0.0122188
R2218 VDD.n184 VDD.n183 0.0083125
R2219 VDD.n115 VDD.n114 0.0083125
R2220 VDD.n220 VDD.n42 0.0083125
R2221 VDD VDD.n220 0.0083125
R2222 VDD.n301 VDD.n300 0.0083125
R2223 VDD.n368 VDD.n367 0.0083125
R2224 VDD.n367 VDD 0.0083125
R2225 VDD.n321 VDD.n314 0.0083125
R2226 VDD.n188 VDD.n187 0.00310417
R2227 VDD.n86 VDD.n82 0.00310417
R2228 VDD.n134 VDD.n100 0.00310417
R2229 VDD.n213 VDD.n212 0.00310417
R2230 VDD.n251 VDD.n31 0.00310417
R2231 VDD.n11 VDD.n6 0.00310417
R2232 VDD.n359 VDD.n358 0.00310417
R2233 VDD.n412 VDD.n409 0.00310417
R2234 VDD.n453 VDD.n444 0.00310417
R2235 select1.n0 select1.t1 323.55
R2236 select1.n0 select1.t0 195.017
R2237 select1.n1 select1.n0 152
R2238 select1.n3 select1 18.8151
R2239 select1 select1.n2 10.2766
R2240 select1.n2 select1 6.7304
R2241 select1.n1 select1 1.45205
R2242 select1.n2 select1.n1 0.792253
R2243 select1.n3 select1 0.0384464
R2244 select1 select1.n3 0.0128547
R2245 passgatesCtrl_0.net10.n1 passgatesCtrl_0.net10.t4 260.322
R2246 passgatesCtrl_0.net10.n3 passgatesCtrl_0.net10.n0 207.22
R2247 passgatesCtrl_0.net10.n1 passgatesCtrl_0.net10.t3 175.169
R2248 passgatesCtrl_0.net10.n2 passgatesCtrl_0.net10.n1 153.13
R2249 passgatesCtrl_0.net10 passgatesCtrl_0.net10.t2 132.067
R2250 passgatesCtrl_0.net10.n0 passgatesCtrl_0.net10.t1 26.5955
R2251 passgatesCtrl_0.net10.n0 passgatesCtrl_0.net10.t0 26.5955
R2252 passgatesCtrl_0.net10 passgatesCtrl_0.net10.n3 17.4717
R2253 passgatesCtrl_0.net10.n3 passgatesCtrl_0.net10 12.2141
R2254 passgatesCtrl_0.net10 passgatesCtrl_0.net10.n2 9.39918
R2255 passgatesCtrl_0.net10.n2 passgatesCtrl_0.net10 3.2005
R2256 passgatesCtrl_0.net1.n12 passgatesCtrl_0.net1.t17 562.236
R2257 passgatesCtrl_0.net1.t17 passgatesCtrl_0.net1.t9 392.027
R2258 passgatesCtrl_0.net1.n20 passgatesCtrl_0.net1.t6 327.99
R2259 passgatesCtrl_0.net1.n3 passgatesCtrl_0.net1.t11 323.55
R2260 passgatesCtrl_0.net1.n1 passgatesCtrl_0.net1.t1 319.171
R2261 passgatesCtrl_0.net1.n24 passgatesCtrl_0.net1.t7 293.969
R2262 passgatesCtrl_0.net1.n8 passgatesCtrl_0.net1.t13 256.07
R2263 passgatesCtrl_0.net1.n17 passgatesCtrl_0.net1.t19 231.835
R2264 passgatesCtrl_0.net1.n6 passgatesCtrl_0.net1.t8 230.155
R2265 passgatesCtrl_0.net1 passgatesCtrl_0.net1.t0 209.923
R2266 passgatesCtrl_0.net1.n16 passgatesCtrl_0.net1.t18 206.19
R2267 passgatesCtrl_0.net1.n20 passgatesCtrl_0.net1.t15 199.457
R2268 passgatesCtrl_0.net1.n3 passgatesCtrl_0.net1.t2 195.017
R2269 passgatesCtrl_0.net1.n14 passgatesCtrl_0.net1.t5 185.376
R2270 passgatesCtrl_0.net1.n6 passgatesCtrl_0.net1.t3 157.856
R2271 passgatesCtrl_0.net1.n17 passgatesCtrl_0.net1.t14 157.07
R2272 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n16 154.657
R2273 passgatesCtrl_0.net1.n18 passgatesCtrl_0.net1.n17 154.048
R2274 passgatesCtrl_0.net1.n7 passgatesCtrl_0.net1.n6 153.147
R2275 passgatesCtrl_0.net1.n25 passgatesCtrl_0.net1.n24 152
R2276 passgatesCtrl_0.net1.n21 passgatesCtrl_0.net1.n20 152
R2277 passgatesCtrl_0.net1.n15 passgatesCtrl_0.net1.n14 152
R2278 passgatesCtrl_0.net1.n9 passgatesCtrl_0.net1.n8 152
R2279 passgatesCtrl_0.net1.n4 passgatesCtrl_0.net1.n3 152
R2280 passgatesCtrl_0.net1.n8 passgatesCtrl_0.net1.t12 150.03
R2281 passgatesCtrl_0.net1.n16 passgatesCtrl_0.net1.t16 148.35
R2282 passgatesCtrl_0.net1.n24 passgatesCtrl_0.net1.t4 138.338
R2283 passgatesCtrl_0.net1.n14 passgatesCtrl_0.net1.t10 137.177
R2284 passgatesCtrl_0.net1.n5 passgatesCtrl_0.net1 28.0894
R2285 passgatesCtrl_0.net1.n11 passgatesCtrl_0.net1.n10 25.2401
R2286 passgatesCtrl_0.net1.n13 passgatesCtrl_0.net1.n12 22.4834
R2287 passgatesCtrl_0.net1.n0 passgatesCtrl_0.net1 21.6175
R2288 passgatesCtrl_0.net1.n11 passgatesCtrl_0.net1.n7 20.5972
R2289 passgatesCtrl_0.net1.n23 passgatesCtrl_0.net1.n22 16.5589
R2290 passgatesCtrl_0.net1.n9 passgatesCtrl_0.net1 16.3845
R2291 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n25 15.2457
R2292 passgatesCtrl_0.net1.n26 passgatesCtrl_0.net1 14.6453
R2293 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n26 13.9801
R2294 passgatesCtrl_0.net1.n21 passgatesCtrl_0.net1 12.1605
R2295 passgatesCtrl_0.net1.n19 passgatesCtrl_0.net1.n0 11.55
R2296 passgatesCtrl_0.net1.n22 passgatesCtrl_0.net1 10.8805
R2297 passgatesCtrl_0.net1.n0 passgatesCtrl_0.net1.n15 10.8365
R2298 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n2 10.6976
R2299 passgatesCtrl_0.net1.n19 passgatesCtrl_0.net1.n18 9.3005
R2300 passgatesCtrl_0.net1.n12 passgatesCtrl_0.net1 8.92171
R2301 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n1 7.73474
R2302 passgatesCtrl_0.net1.n23 passgatesCtrl_0.net1.n19 7.40435
R2303 passgatesCtrl_0.net1.n5 passgatesCtrl_0.net1.n4 7.1685
R2304 passgatesCtrl_0.net1.n0 passgatesCtrl_0.net1.n13 6.03757
R2305 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n5 4.62272
R2306 passgatesCtrl_0.net1.n10 passgatesCtrl_0.net1.n9 4.6085
R2307 passgatesCtrl_0.net1.n10 passgatesCtrl_0.net1 4.58918
R2308 passgatesCtrl_0.net1.n18 passgatesCtrl_0.net1 4.3525
R2309 passgatesCtrl_0.net1.n26 passgatesCtrl_0.net1 4.26717
R2310 passgatesCtrl_0.net1.n22 passgatesCtrl_0.net1 3.62717
R2311 passgatesCtrl_0.net1.n13 passgatesCtrl_0.net1.n11 3.29171
R2312 passgatesCtrl_0.net1.n7 passgatesCtrl_0.net1 3.24826
R2313 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n23 3.14198
R2314 passgatesCtrl_0.net1.n15 passgatesCtrl_0.net1 3.0725
R2315 passgatesCtrl_0.net1.n4 passgatesCtrl_0.net1 2.9445
R2316 passgatesCtrl_0.net1.n1 passgatesCtrl_0.net1 2.48634
R2317 passgatesCtrl_0.net1 passgatesCtrl_0.net1.n21 2.34717
R2318 passgatesCtrl_0.net1.n2 passgatesCtrl_0.net1 2.19479
R2319 passgatesCtrl_0.net1.n25 passgatesCtrl_0.net1 2.06502
R2320 passgatesCtrl_0.net1.n2 passgatesCtrl_0.net1 1.80756
R2321 passgatesCtrl_0.net1.n5 passgatesCtrl_0.net1 1.6645
R2322 A3.n1 A3.t3 26.3998
R2323 A3.n1 A3.t2 23.5483
R2324 A3.n0 A3.t0 12.7127
R2325 A3.n0 A3.t1 10.8578
R2326 A3.n2 A3.n1 3.12177
R2327 A3.n2 A3.n0 1.81453
R2328 A3.n3 A3.n2 1.1255
R2329 A3.n3 A3 0.210543
R2330 A3 A3.n3 0.0655
R2331 Z3.n1 Z3.t3 23.6581
R2332 Z3.n3 Z3.t2 23.3739
R2333 Z3.n1 Z3.t1 10.7528
R2334 Z3.n0 Z3.t0 10.6417
R2335 Z3.n2 Z3.n1 1.30064
R2336 Z3.n5 Z3.n4 0.924585
R2337 Z3.n3 Z3.n2 0.726502
R2338 Z3.n2 Z3.n0 0.512491
R2339 Z3.n4 Z3.n0 0.359663
R2340 Z3.n4 Z3.n3 0.216071
R2341 Z3.n5 Z3 0.0656042
R2342 Z3 Z3.n5 0.0376287
R2343 select0.n0 select0.t1 323.55
R2344 select0.n0 select0.t0 195.017
R2345 select0.n1 select0.n0 152
R2346 select0 select0.n2 14.4176
R2347 select0.n2 select0 6.7304
R2348 select0.n3 select0 2.87104
R2349 select0.n1 select0 1.45205
R2350 select0.n2 select0.n1 0.792253
R2351 select0.n3 select0 0.0696964
R2352 select0 select0.n3 0.0230291
R2353 Z2.n1 Z2.t0 23.6581
R2354 Z2.n3 Z2.t1 23.3739
R2355 Z2.n1 Z2.t3 10.7528
R2356 Z2.n0 Z2.t2 10.6417
R2357 Z2.n2 Z2.n1 1.30064
R2358 Z2.n5 Z2.n4 0.936641
R2359 Z2.n3 Z2.n2 0.726502
R2360 Z2.n2 Z2.n0 0.512491
R2361 Z2.n4 Z2.n0 0.359663
R2362 Z2.n4 Z2.n3 0.216071
R2363 Z2.n5 Z2 0.0776605
R2364 Z2 Z2.n5 0.0561931
R2365 A2.n1 A2.t0 26.3998
R2366 A2.n1 A2.t1 23.5483
R2367 A2.n0 A2.t3 12.7127
R2368 A2.n0 A2.t2 10.8578
R2369 A2.n2 A2.n1 3.12177
R2370 A2.n2 A2.n0 1.81453
R2371 A2.n3 A2.n2 1.1255
R2372 A2.n3 A2 0.219402
R2373 A2 A2.n3 0.0655
R2374 Z4.n1 Z4.t3 23.6581
R2375 Z4.n3 Z4.t2 23.3739
R2376 Z4.n1 Z4.t0 10.7528
R2377 Z4.n0 Z4.t1 10.6417
R2378 Z4.n2 Z4.n1 1.30064
R2379 Z4 Z4.n4 0.983856
R2380 Z4.n3 Z4.n2 0.726502
R2381 Z4.n2 Z4.n0 0.512491
R2382 Z4.n4 Z4.n0 0.359663
R2383 Z4.n4 Z4.n3 0.216071
R2384 A4.n1 A4.t3 26.3998
R2385 A4.n1 A4.t2 23.5483
R2386 A4.n0 A4.t0 12.7127
R2387 A4.n0 A4.t1 10.8578
R2388 A4.n2 A4.n1 3.12177
R2389 A4.n2 A4.n0 1.81453
R2390 A4.n3 A4.n2 1.1255
R2391 A4 A4.n3 0.134513
R2392 A4.n3 A4 0.0655
R2393 Z1.n1 Z1.t2 23.6581
R2394 Z1.n3 Z1.t3 23.3739
R2395 Z1.n1 Z1.t0 10.7528
R2396 Z1.n0 Z1.t1 10.6417
R2397 Z1.n2 Z1.n1 1.30064
R2398 Z1 Z1.n4 0.983856
R2399 Z1.n3 Z1.n2 0.726502
R2400 Z1.n2 Z1.n0 0.512491
R2401 Z1.n4 Z1.n0 0.359663
R2402 Z1.n4 Z1.n3 0.216071
R2403 A1.n1 A1.t2 26.3998
R2404 A1.n1 A1.t3 23.5483
R2405 A1.n0 A1.t0 12.7127
R2406 A1.n0 A1.t1 10.8578
R2407 A1.n2 A1.n1 3.12177
R2408 A1.n2 A1.n0 1.81453
R2409 A1.n3 A1.n2 1.1255
R2410 A1.n3 A1 0.21549
R2411 A1 A1.n3 0.0655
C0 passgatesCtrl_0.net6 a_n2057_n1942# 0.001427f
C1 passgatex4_0.GN1 passgatesCtrl_0.net1 0.055547f
C2 passgatesCtrl_0.net7 a_n1459_n3306# 1.39e-19
C3 passgatex4_0.GP4 a_n2883_n1648# 0.033357f
C4 A1 passgatesCtrl_0._02_ 2.53e-20
C5 passgatex4_0.GN4 Z4 0.443709f
C6 passgatex4_0.GN3 passgatex4_0.GN1 5.26e-19
C7 a_n491_n3280# a_n539_n3518# 5.96e-19
C8 passgatesCtrl_0.net3 passgatesCtrl_0._02_ 6.01e-20
C9 a_n1878_n4368# a_n1984_n4368# 0.313533f
C10 a_n801_n4216# passgatesCtrl_0._04_ 5.33e-19
C11 passgatesCtrl_0.net8 passgatesCtrl_0.net3 8.71e-21
C12 a_n1503_n2192# a_n1459_n3306# 6.43e-21
C13 passgatesCtrl_0.net6 a_n2639_n2040# 0.046149f
C14 passgatesCtrl_0._05_ passgatesCtrl_0.net2 0.019534f
C15 passgatesCtrl_0._03_ passgatex4_0.GP1 4.32e-20
C16 passgatesCtrl_0.net1 a_n2015_n2040# 0.134894f
C17 passgatesCtrl_0.net9 a_n1913_n1429# 0.031948f
C18 passgatex4_0.GP4 passgatesCtrl_0.net7 3.05e-20
C19 a_n2429_n1328# passgatesCtrl_0.net9 2.52e-19
C20 passgatesCtrl_0.net4 passgatesCtrl_0.net5 0.024789f
C21 passgatesCtrl_0.net5 a_n1003_n2040# 6.98e-19
C22 passgatex4_0.GN1 a_n995_n3605# 3.14e-19
C23 passgatex4_0.GN1 a_n1173_n2218# 1.7e-19
C24 passgatex4_0.GN3 a_n2015_n2040# 7.19e-21
C25 passgatesCtrl_0.net1 passgatex4_0.GN2 0.117828f
C26 passgatesCtrl_0.net2 a_n2975_n2192# 0.006018f
C27 passgatex4_0.GP2 A1 0.002086f
C28 passgatesCtrl_0.net4 a_n715_n3850# 8.15e-19
C29 select0 a_n1878_n4368# 3.96e-19
C30 VDD a_n1637_n1429# 0.221714f
C31 passgatex4_0.GN3 passgatex4_0.GN2 0.051202f
C32 passgatex4_0.GP2 passgatesCtrl_0.net3 3.9e-21
C33 a_n1361_n1429# passgatesCtrl_0.net10 5.14e-19
C34 passgatesCtrl_0.net5 a_n1913_n1429# 0.038008f
C35 passgatesCtrl_0.net1 a_n2883_n1648# -6.59e-36
C36 passgatex4_0.GP4 passgatex4_0.GN4 3.44232f
C37 a_n1085_n1429# passgatesCtrl_0._00_ 4.99e-20
C38 a_n2429_n1328# passgatesCtrl_0.net5 8.98e-21
C39 select1 a_n1084_n4216# 0.005547f
C40 a_n1963_n3280# passgatesCtrl_0.net1 2.5e-19
C41 VDD a_n491_n3280# 0.291441f
C42 a_n1635_n3306# a_n1459_n3306# 0.185422f
C43 a_n1173_n2218# passgatex4_0.GN2 0.001025f
C44 select0 a_n1984_n4368# 1.65e-19
C45 passgatesCtrl_0.net7 passgatesCtrl_0.net1 0.492308f
C46 passgatesCtrl_0.net2 passgatesCtrl_0._00_ 0.181488f
C47 a_n482_n4216# a_n715_n3850# 0.001428f
C48 passgatesCtrl_0._01_ a_n1045_n1942# 3.51e-19
C49 a_n597_n2040# a_n675_n1648# 0.003066f
C50 passgatex4_0.GN1 passgatesCtrl_0.net5 0.002166f
C51 passgatex4_0.GN3 passgatesCtrl_0.net7 1.52e-19
C52 passgatesCtrl_0.net1 a_n587_n3458# 0.002306f
C53 Z3 passgatex4_0.GN2 2.12e-20
C54 passgatesCtrl_0.net6 a_n1003_n2040# 2.87e-20
C55 passgatesCtrl_0._01_ a_n2185_n2218# 0.001002f
C56 passgatex4_0.GN4 passgatesCtrl_0.net1 5.43e-19
C57 passgatex4_0.GN1 a_n715_n3850# 0.001005f
C58 a_n1503_n2192# passgatesCtrl_0.net1 0.040031f
C59 a_n1459_n3306# passgatesCtrl_0.net2 0.096716f
C60 select1 passgatesCtrl_0.net2 0.026514f
C61 passgatex4_0.GN3 passgatex4_0.GN4 0.155269f
C62 passgatesCtrl_0.net6 a_n1913_n1429# 0.008072f
C63 a_n1503_n2192# passgatex4_0.GN3 1.78e-19
C64 a_n2015_n2040# passgatesCtrl_0.net5 0.012287f
C65 passgatesCtrl_0.net9 a_n2883_n1648# 0.123724f
C66 passgatesCtrl_0.net10 a_n675_n1648# 7.12e-20
C67 a_n597_n2040# passgatex4_0.GP1 9.87e-19
C68 passgatex4_0.GN1 A2 3.14e-19
C69 a_n539_n3518# passgatesCtrl_0._04_ 0.001297f
C70 passgatesCtrl_0.net5 passgatex4_0.GN2 0.011028f
C71 a_n2015_n2040# a_n2057_n1942# 3.5e-20
C72 a_n1503_n2192# a_n1173_n2218# 0.018393f
C73 passgatex4_0.GN3 Z2 0.00126f
C74 VDD a_n1361_n1429# 0.211763f
C75 passgatesCtrl_0.net5 a_n2883_n1648# 4.81e-20
C76 passgatex4_0.GP4 passgatesCtrl_0.net2 0.005696f
C77 passgatesCtrl_0.net1 a_n1084_n4216# 0.004309f
C78 passgatesCtrl_0.net4 a_n1003_n2040# 0.001809f
C79 a_n1635_n3306# passgatesCtrl_0.net1 0.001693f
C80 passgatesCtrl_0.net7 passgatesCtrl_0.net9 1.77e-20
C81 VDD a_n951_n2736# 0.193152f
C82 a_n1963_n3280# passgatesCtrl_0.net5 0.115837f
C83 a_n1637_n1429# passgatesCtrl_0.net8 0.001796f
C84 passgatex4_0.GP3 passgatex4_0.GP1 5.06e-19
C85 passgatex4_0.GN4 Z3 0.00128f
C86 A2 passgatex4_0.GN2 3.8137f
C87 passgatesCtrl_0.net1 a_n1085_n1429# 1.87e-20
C88 a_n1459_n3306# passgatesCtrl_0.net3 2.01e-19
C89 VDD Z1 2.98463f
C90 a_n482_n4216# select0 0.266581f
C91 passgatex4_0.GN4 passgatesCtrl_0.net9 4.06e-19
C92 passgatesCtrl_0.net7 passgatesCtrl_0.net5 0.002751f
C93 passgatex4_0.GN3 a_n1085_n1429# 6.29e-19
C94 a_n1135_n4368# VDD 0.162421f
C95 a_n1084_n4216# a_n995_n3605# 1.65e-19
C96 passgatesCtrl_0.net6 a_n2015_n2040# 0.013011f
C97 VDD passgatesCtrl_0._04_ 0.211525f
C98 passgatesCtrl_0.net7 a_n715_n3850# 0.00214f
C99 passgatex4_0.GP2 a_n1637_n1429# 0.002575f
C100 Z3 Z2 7.67e-19
C101 passgatex4_0.GN1 select0 0.005832f
C102 passgatex4_0.GP4 A1 1.34e-19
C103 passgatesCtrl_0.net6 passgatex4_0.GN2 5.41e-20
C104 passgatesCtrl_0.net1 passgatesCtrl_0.net2 1.72543f
C105 passgatex4_0.GN4 passgatesCtrl_0.net5 0.05537f
C106 a_n1503_n2192# passgatesCtrl_0.net5 0.003576f
C107 a_n715_n3850# a_n587_n3458# 0.004764f
C108 a_n1173_n2218# a_n1085_n1429# 4.77e-20
C109 passgatex4_0.GN3 passgatesCtrl_0.net2 0.006039f
C110 passgatesCtrl_0.net6 a_n2883_n1648# 4.16e-19
C111 VDD a_n2161_n4368# 0.173581f
C112 passgatex4_0.GN1 passgatesCtrl_0.net4 0.083575f
C113 passgatex4_0.GN1 a_n1003_n2040# 4.06e-19
C114 VDD a_n675_n1648# 0.230164f
C115 passgatesCtrl_0.net2 a_n995_n3605# 0.043831f
C116 passgatesCtrl_0.net2 a_n1173_n2218# 0.177825f
C117 passgatex4_0.GN4 A2 1.95e-19
C118 a_n1085_n1429# passgatesCtrl_0.net9 4.15e-21
C119 passgatesCtrl_0.net6 passgatesCtrl_0.net7 5.12e-20
C120 passgatex4_0.GN4 a_n2639_n2040# 3.33e-20
C121 passgatesCtrl_0.net1 A1 0.049065f
C122 a_n1635_n3306# passgatesCtrl_0.net5 0.0036f
C123 VDD passgatesCtrl_0._03_ 0.196287f
C124 passgatesCtrl_0.net4 passgatex4_0.GN2 0.005352f
C125 a_n1003_n2040# passgatex4_0.GN2 0.003895f
C126 VDD passgatex4_0.GP1 2.34735f
C127 passgatesCtrl_0.net1 passgatesCtrl_0.net3 0.178768f
C128 passgatex4_0.GN3 A1 4.37e-19
C129 passgatesCtrl_0.net2 a_n2480_n4368# 0.162398f
C130 a_n2015_n2040# a_n1913_n1429# 1.05e-19
C131 passgatex4_0.GN1 a_n482_n4216# 0.00164f
C132 A2 Z2 4.51569f
C133 passgatesCtrl_0.net5 a_n1085_n1429# 0.032876f
C134 a_n1361_n1429# passgatesCtrl_0.net8 0.004727f
C135 passgatex4_0.GN4 passgatesCtrl_0.net6 0.043823f
C136 VDD a_n1227_n2736# 0.241578f
C137 a_n1503_n2192# passgatesCtrl_0.net6 0.001672f
C138 VDD a_n2465_n2164# 3.98e-19
C139 a_n1913_n1429# passgatex4_0.GN2 5.52e-20
C140 passgatesCtrl_0.net2 passgatesCtrl_0.net9 0.086587f
C141 a_n1135_n4368# a_n988_n4394# 0.003683f
C142 passgatesCtrl_0.net4 a_n1963_n3280# 0.001365f
C143 a_n1637_n1429# passgatesCtrl_0._00_ 1.44e-19
C144 VDD a_n1045_n1942# 6.29e-19
C145 a_n988_n4394# passgatesCtrl_0._04_ 0.001033f
C146 VDD passgatesCtrl_0._01_ 0.225859f
C147 passgatesCtrl_0._03_ a_n1507_n3280# 8.17e-20
C148 a_n995_n3605# passgatesCtrl_0.net3 1.28e-21
C149 a_n1173_n2218# passgatesCtrl_0.net3 0.010683f
C150 passgatesCtrl_0.net2 passgatesCtrl_0.net5 0.544042f
C151 passgatex4_0.GP2 a_n1361_n1429# 0.134077f
C152 VDD a_n2185_n2218# 0.130016f
C153 passgatex4_0.GP3 passgatesCtrl_0.net10 0.234131f
C154 passgatesCtrl_0.net4 passgatesCtrl_0.net7 3.73e-19
C155 passgatesCtrl_0.net2 a_n715_n3850# 0.067356f
C156 Z3 A1 4.74e-21
C157 VDD a_n801_n4216# 0.191329f
C158 a_n1084_n4216# a_n1984_n4368# 1.1e-19
C159 passgatesCtrl_0.net4 a_n587_n3458# 4.09e-19
C160 passgatex4_0.GN1 passgatex4_0.GN2 0.033541f
C161 passgatesCtrl_0.net7 a_n1913_n1429# 6.2e-20
C162 passgatex4_0.GP2 Z1 3.73e-21
C163 a_n1503_n2192# a_n1003_n2040# 4.74e-20
C164 passgatesCtrl_0.net2 a_n1878_n4368# 0.010759f
C165 passgatesCtrl_0.net6 a_n1085_n1429# 0.001258f
C166 passgatesCtrl_0._02_ a_n675_n1648# 0.194553f
C167 passgatex4_0.GN4 a_n1913_n1429# 0.112321f
C168 passgatesCtrl_0.net8 a_n675_n1648# 6.36e-19
C169 passgatesCtrl_0.net2 a_n2639_n2040# 0.180659f
C170 a_n2015_n2040# passgatex4_0.GN2 1.39e-19
C171 passgatesCtrl_0.net5 A1 5.61e-21
C172 select0 a_n1084_n4216# 0.001575f
C173 a_n482_n4216# passgatesCtrl_0.net7 6.47e-19
C174 passgatex4_0.GN4 a_n2429_n1328# 2.79e-21
C175 a_n715_n3850# A1 0.001233f
C176 passgatesCtrl_0.net5 passgatesCtrl_0.net3 0.001999f
C177 VDD a_n597_n2040# 0.179575f
C178 a_n434_n1942# passgatex4_0.GP1 2.65e-19
C179 passgatesCtrl_0.net6 passgatesCtrl_0.net2 0.0936f
C180 passgatex4_0.GN1 passgatesCtrl_0.net7 0.028089f
C181 passgatesCtrl_0.net2 a_n1984_n4368# 0.051248f
C182 passgatesCtrl_0.net4 a_n1084_n4216# 0.00141f
C183 passgatex4_0.GP1 passgatesCtrl_0._02_ 6.66e-20
C184 passgatex4_0.GP2 a_n675_n1648# 5.94e-19
C185 passgatesCtrl_0.net4 a_n1635_n3306# 0.007618f
C186 A4 passgatex4_0.GP3 0.16204f
C187 passgatex4_0.GN1 a_n587_n3458# 1.58e-19
C188 A1 A2 1.81909f
C189 passgatex4_0.GN1 passgatex4_0.GN4 2.04e-19
C190 a_n1227_n2736# passgatesCtrl_0.net8 1.26e-20
C191 passgatesCtrl_0.net4 a_n1085_n1429# 2.63e-19
C192 a_n1361_n1429# passgatesCtrl_0._00_ 8.1e-20
C193 VDD passgatesCtrl_0.net10 0.395163f
C194 A3 passgatex4_0.GP1 2.46e-21
C195 VDD passgatex4_0.GP3 1.84344f
C196 select0 passgatesCtrl_0.net2 0.002824f
C197 passgatesCtrl_0.net7 passgatex4_0.GN2 0.34798f
C198 a_n1637_n1429# passgatesCtrl_0.net1 1.96e-19
C199 passgatex4_0.GP2 passgatex4_0.GP1 0.008406f
C200 passgatesCtrl_0.net8 a_n1045_n1942# 9.1e-19
C201 passgatesCtrl_0._01_ passgatesCtrl_0.net8 0.208131f
C202 a_n801_n4216# a_n988_n4394# 0.159555f
C203 passgatex4_0.GN1 Z2 4.77e-21
C204 passgatex4_0.GN3 a_n1637_n1429# 0.14217f
C205 a_n1503_n2192# a_n2015_n2040# 0.014264f
C206 passgatesCtrl_0.net8 a_n2185_n2218# 1.99e-21
C207 VDD a_n1701_n4368# 0.143966f
C208 passgatex4_0.GP2 a_n1227_n2736# 4.59e-20
C209 passgatesCtrl_0.net4 passgatesCtrl_0.net2 0.097522f
C210 a_n1459_n3306# a_n1361_n1429# 8.17e-21
C211 passgatesCtrl_0.net2 a_n1003_n2040# 0.166925f
C212 passgatex4_0.GN4 passgatex4_0.GN2 5.8e-19
C213 a_n1503_n2192# passgatex4_0.GN2 4.62e-19
C214 a_n2189_n1429# a_n2185_n2218# 0.011493f
C215 a_n491_n3280# passgatesCtrl_0.net1 0.007927f
C216 VDD a_n539_n3518# 0.259999f
C217 passgatex4_0.GN1 a_n1084_n4216# 4.22e-19
C218 passgatesCtrl_0.net7 a_n1963_n3280# 3.8e-20
C219 passgatesCtrl_0.net2 a_n1913_n1429# 3.2e-19
C220 passgatex4_0.GN4 a_n2883_n1648# 2.19e-19
C221 passgatesCtrl_0.net2 a_n2429_n1328# 1.42e-19
C222 passgatesCtrl_0._01_ passgatex4_0.GP2 4.67e-20
C223 select1 Z1 2.26e-19
C224 select0 A1 0.040389f
C225 passgatex4_0.GN1 a_n1085_n1429# 3.8e-19
C226 passgatesCtrl_0._05_ a_n2465_n2164# 5.76e-19
C227 Z2 passgatex4_0.GN2 0.427031f
C228 select0 passgatesCtrl_0.net3 1.33e-20
C229 a_n1135_n4368# select1 0.004485f
C230 a_n597_n2040# a_n434_n1942# 0.004767f
C231 a_n482_n4216# passgatesCtrl_0.net2 0.001264f
C232 select1 passgatesCtrl_0._04_ 3.6e-20
C233 passgatesCtrl_0.net4 A1 6.83e-21
C234 a_n597_n2040# passgatesCtrl_0._02_ 0.106303f
C235 VDD A4 1.54289f
C236 passgatex4_0.GN4 passgatesCtrl_0.net7 4.64e-20
C237 a_n1503_n2192# passgatesCtrl_0.net7 2.69e-21
C238 passgatesCtrl_0._01_ passgatesCtrl_0._05_ 6.19e-21
C239 a_n1637_n1429# passgatesCtrl_0.net9 1.63e-19
C240 passgatesCtrl_0.net4 passgatesCtrl_0.net3 0.130377f
C241 a_n1003_n2040# passgatesCtrl_0.net3 7.73e-20
C242 passgatex4_0.GN1 passgatesCtrl_0.net2 0.068323f
C243 a_n1085_n1429# passgatex4_0.GN2 0.002397f
C244 select1 a_n2161_n4368# 0.002569f
C245 passgatesCtrl_0._01_ a_n2975_n2192# 3.25e-21
C246 a_n2975_n2192# a_n2185_n2218# 1.06e-20
C247 a_n1637_n1429# passgatesCtrl_0.net5 0.033814f
C248 passgatesCtrl_0.net10 passgatesCtrl_0._02_ 5.35e-20
C249 a_n1963_n3280# a_n1635_n3306# 0.017591f
C250 passgatesCtrl_0.net1 a_n1361_n1429# 2.44e-20
C251 passgatesCtrl_0.net2 a_n2015_n2040# 0.185322f
C252 passgatesCtrl_0.net8 passgatesCtrl_0.net10 1.06e-19
C253 a_n482_n4216# A1 0.001912f
C254 passgatex4_0.GN3 a_n1361_n1429# 0.109673f
C255 a_n1701_n4368# a_n988_n4394# 1.09e-19
C256 passgatesCtrl_0.net2 passgatex4_0.GN2 0.06846f
C257 a_n2189_n1429# passgatesCtrl_0.net10 0.041816f
C258 passgatesCtrl_0.net7 a_n1635_n3306# 1.83e-19
C259 a_n951_n2736# passgatesCtrl_0.net1 0.02864f
C260 a_n491_n3280# passgatesCtrl_0.net5 6.09e-20
C261 passgatex4_0.GP3 a_n2189_n1429# 0.110988f
C262 passgatesCtrl_0._03_ a_n1459_n3306# 9.63e-19
C263 select1 passgatesCtrl_0._03_ 4.71e-19
C264 passgatex4_0.GN1 A1 4.96968f
C265 a_n1459_n3306# passgatex4_0.GP1 1.14e-19
C266 VDD a_n1507_n3280# 0.003544f
C267 passgatesCtrl_0.net1 Z1 3.3e-21
C268 passgatesCtrl_0.net2 a_n2883_n1648# 0.012477f
C269 A3 passgatex4_0.GP3 3.97267f
C270 passgatesCtrl_0.net7 a_n1085_n1429# 4.02e-19
C271 passgatesCtrl_0._01_ passgatesCtrl_0._00_ 5.18e-20
C272 passgatex4_0.GN1 passgatesCtrl_0.net3 0.357097f
C273 a_n2185_n2218# passgatesCtrl_0._00_ 0.0957f
C274 passgatex4_0.GP2 passgatesCtrl_0.net10 9.63e-20
C275 a_n1135_n4368# passgatesCtrl_0.net1 0.001335f
C276 passgatex4_0.GP2 passgatex4_0.GP3 0.007549f
C277 passgatesCtrl_0.net1 passgatesCtrl_0._04_ 0.050056f
C278 a_n1963_n3280# passgatesCtrl_0.net2 0.04096f
C279 passgatex4_0.GP4 passgatex4_0.GP1 2.41e-19
C280 a_n1637_n1429# passgatesCtrl_0.net6 0.218518f
C281 passgatesCtrl_0.net7 passgatesCtrl_0.net2 0.090257f
C282 A1 passgatex4_0.GN2 0.151745f
C283 passgatesCtrl_0._05_ passgatex4_0.GP3 6.13e-19
C284 passgatesCtrl_0.net3 passgatex4_0.GN2 0.069726f
C285 passgatesCtrl_0.net2 a_n587_n3458# 0.001719f
C286 a_n1361_n1429# passgatesCtrl_0.net9 7.62e-20
C287 passgatesCtrl_0.net1 a_n675_n1648# 8.22e-19
C288 a_n995_n3605# passgatesCtrl_0._04_ 0.294104f
C289 VDD a_n988_n4394# 0.211037f
C290 a_n801_n4216# select1 0.001678f
C291 passgatex4_0.GN4 passgatesCtrl_0.net2 7.43e-19
C292 a_n1503_n2192# passgatesCtrl_0.net2 0.03779f
C293 passgatex4_0.GN1 a_n485_n2736# 0.003892f
C294 VDD a_n434_n1942# 0.002344f
C295 passgatex4_0.GN3 a_n675_n1648# 1.89e-19
C296 VDD passgatesCtrl_0._02_ 0.450634f
C297 a_n1361_n1429# passgatesCtrl_0.net5 0.230704f
C298 passgatex4_0.GP4 a_n2185_n2218# 2.89e-21
C299 VDD passgatesCtrl_0.net8 0.561328f
C300 A3 A4 2.08862f
C301 passgatesCtrl_0._03_ passgatesCtrl_0.net1 9.6e-19
C302 passgatesCtrl_0.net7 A1 0.012018f
C303 passgatesCtrl_0.net1 passgatex4_0.GP1 0.003098f
C304 VDD a_n2189_n1429# 0.195044f
C305 a_n951_n2736# passgatesCtrl_0.net5 6.35e-19
C306 passgatex4_0.GP2 A4 2.48e-20
C307 select0 a_n491_n3280# 4.9e-19
C308 passgatesCtrl_0.net7 passgatesCtrl_0.net3 0.034004f
C309 VDD A3 1.61205f
C310 a_n1227_n2736# passgatesCtrl_0.net1 8.11e-19
C311 passgatex4_0.GN3 passgatex4_0.GP1 8.28e-19
C312 a_n587_n3458# A1 4.82e-20
C313 passgatesCtrl_0.net2 a_n1084_n4216# 0.001027f
C314 passgatesCtrl_0.net10 passgatesCtrl_0._00_ 0.005756f
C315 passgatex4_0.GN4 A1 1.92e-19
C316 a_n1635_n3306# passgatesCtrl_0.net2 0.200956f
C317 VDD passgatex4_0.GP2 1.61055f
C318 passgatex4_0.GP3 passgatesCtrl_0._00_ 0.098299f
C319 a_n1637_n1429# a_n1913_n1429# 5.3e-19
C320 passgatesCtrl_0.net1 a_n1045_n1942# 0.001768f
C321 passgatesCtrl_0.net2 a_n1085_n1429# 0.006979f
C322 passgatesCtrl_0._01_ passgatesCtrl_0.net1 0.173572f
C323 a_n715_n3850# passgatesCtrl_0._04_ 0.099459f
C324 passgatesCtrl_0.net1 a_n2185_n2218# 0.184986f
C325 Z4 passgatex4_0.GP3 0.071646f
C326 a_n1227_n2736# a_n1173_n2218# 3.06e-19
C327 passgatesCtrl_0._01_ passgatex4_0.GN3 1.44e-19
C328 A1 Z2 0.004942f
C329 passgatex4_0.GN3 a_n2185_n2218# 4.42e-19
C330 passgatesCtrl_0.net6 a_n1361_n1429# 0.033794f
C331 VDD passgatesCtrl_0._05_ 0.358831f
C332 a_n801_n4216# passgatesCtrl_0.net1 0.329151f
C333 passgatesCtrl_0.net7 a_n485_n2736# 0.002755f
C334 Z3 passgatex4_0.GP1 1.86e-21
C335 passgatesCtrl_0.net5 a_n675_n1648# 2.48e-19
C336 a_n1173_n2218# a_n1045_n1942# 0.005162f
C337 a_n1084_n4216# A1 7.64e-21
C338 VDD a_n2975_n2192# 0.310075f
C339 passgatesCtrl_0._01_ a_n1173_n2218# 0.101852f
C340 a_n482_n4216# a_n491_n3280# 1.73e-21
C341 a_n1084_n4216# passgatesCtrl_0.net3 9.59e-22
C342 a_n1701_n4368# select1 0.004749f
C343 passgatex4_0.GP4 passgatesCtrl_0.net10 0.076097f
C344 a_n434_n1942# passgatesCtrl_0._02_ 4.96e-19
C345 passgatex4_0.GP4 passgatex4_0.GP3 0.057096f
C346 passgatex4_0.GN1 a_n491_n3280# 0.001658f
C347 a_n1135_n4368# a_n1984_n4368# 1.09e-19
C348 passgatesCtrl_0._03_ passgatesCtrl_0.net5 0.19429f
C349 passgatesCtrl_0.net5 passgatex4_0.GP1 0.0014f
C350 passgatesCtrl_0.net1 a_n597_n2040# 0.215616f
C351 passgatesCtrl_0.net8 passgatesCtrl_0._02_ 0.096563f
C352 a_n1637_n1429# passgatex4_0.GN2 2.05e-19
C353 a_n1227_n2736# passgatesCtrl_0.net5 0.002913f
C354 passgatesCtrl_0.net9 a_n2185_n2218# 6.62e-20
C355 select0 Z1 0.003513f
C356 VDD passgatesCtrl_0._00_ 0.89146f
C357 passgatesCtrl_0.net2 A1 0.002113f
C358 A4 Z4 4.51497f
C359 a_n2161_n4368# a_n1984_n4368# 0.159555f
C360 a_n951_n2736# passgatesCtrl_0.net4 0.194653f
C361 passgatesCtrl_0.net2 passgatesCtrl_0.net3 0.095367f
C362 a_n951_n2736# a_n1003_n2040# 3.63e-19
C363 a_n1135_n4368# select0 5.8e-19
C364 passgatesCtrl_0.net5 a_n1045_n1942# 3.13e-20
C365 passgatex4_0.GP1 A2 0.122954f
C366 passgatesCtrl_0._01_ passgatesCtrl_0.net5 0.003676f
C367 passgatex4_0.GP2 passgatesCtrl_0._02_ 2.58e-19
C368 passgatesCtrl_0.net1 passgatesCtrl_0.net10 0.160369f
C369 a_n1173_n2218# a_n597_n2040# 8.8e-19
C370 passgatesCtrl_0.net5 a_n2185_n2218# 0.00379f
C371 VDD Z4 2.81307f
C372 passgatesCtrl_0.net1 passgatex4_0.GP3 0.058232f
C373 passgatex4_0.GP2 passgatesCtrl_0.net8 0.008913f
C374 VDD a_n1459_n3306# 0.260783f
C375 VDD select1 1.30675f
C376 passgatex4_0.GN3 passgatesCtrl_0.net10 0.152678f
C377 passgatex4_0.GN3 passgatex4_0.GP3 2.37902f
C378 passgatesCtrl_0.net4 passgatesCtrl_0._04_ 0.00489f
C379 a_n1637_n1429# passgatesCtrl_0.net7 9.8e-20
C380 a_n2465_n2164# a_n2639_n2040# 0.006584f
C381 a_n2057_n1942# a_n2185_n2218# 0.005162f
C382 passgatesCtrl_0.net6 passgatesCtrl_0._03_ 2.14e-19
C383 passgatex4_0.GP2 A3 0.145029f
C384 passgatex4_0.GP4 A4 3.97306f
C385 a_n1701_n4368# passgatesCtrl_0.net1 3.89e-19
C386 a_n801_n4216# a_n715_n3850# 3.21e-19
C387 passgatex4_0.GN1 a_n1361_n1429# 2e-20
C388 passgatesCtrl_0.net1 a_n539_n3518# 0.107968f
C389 A1 passgatesCtrl_0.net3 1.84e-20
C390 passgatex4_0.GN4 a_n1637_n1429# 0.111188f
C391 passgatesCtrl_0._01_ a_n2639_n2040# 5.79e-21
C392 VDD passgatex4_0.GP4 1.50532f
C393 passgatesCtrl_0.net7 a_n491_n3280# 0.200958f
C394 a_n2639_n2040# a_n2185_n2218# 0.002367f
C395 a_n951_n2736# passgatex4_0.GN1 0.135217f
C396 passgatesCtrl_0.net6 a_n1045_n1942# 2.07e-20
C397 passgatex4_0.GN1 Z1 0.428012f
C398 passgatesCtrl_0._01_ passgatesCtrl_0.net6 0.002059f
C399 select0 passgatex4_0.GP1 7.71e-19
C400 passgatesCtrl_0.net6 a_n2185_n2218# 0.029048f
C401 Z3 passgatex4_0.GP3 0.278332f
C402 a_n1135_n4368# passgatex4_0.GN1 1.78e-19
C403 passgatesCtrl_0.net9 passgatesCtrl_0.net10 0.181065f
C404 a_n1361_n1429# passgatex4_0.GN2 6.44e-19
C405 passgatex4_0.GP3 passgatesCtrl_0.net9 0.117574f
C406 passgatesCtrl_0.net4 passgatesCtrl_0._03_ 0.002493f
C407 passgatex4_0.GN1 passgatesCtrl_0._04_ 0.004444f
C408 passgatesCtrl_0.net4 passgatex4_0.GP1 3.09e-20
C409 passgatex4_0.GN3 A4 0.007063f
C410 a_n951_n2736# passgatex4_0.GN2 0.110403f
C411 a_n1227_n2736# passgatesCtrl_0.net4 0.041847f
C412 passgatesCtrl_0.net5 passgatesCtrl_0.net10 0.099696f
C413 VDD passgatesCtrl_0.net1 2.63744f
C414 passgatesCtrl_0.net8 passgatesCtrl_0._00_ 1.17e-19
C415 Z1 passgatex4_0.GN2 6.82e-19
C416 passgatesCtrl_0.net3 a_n485_n2736# 0.011812f
C417 passgatex4_0.GP3 passgatesCtrl_0.net5 0.001185f
C418 VDD passgatex4_0.GN3 0.518775f
C419 a_n2189_n1429# passgatesCtrl_0._00_ 6.88e-19
C420 passgatex4_0.GN1 a_n675_n1648# 8.62e-19
C421 select1 a_n988_n4394# 5.9e-19
C422 passgatesCtrl_0.net4 a_n1045_n1942# 2.33e-19
C423 a_n1003_n2040# a_n1045_n1942# 3.5e-20
C424 passgatesCtrl_0._05_ a_n2975_n2192# 0.225698f
C425 a_n801_n4216# select0 0.004124f
C426 passgatesCtrl_0._01_ a_n1003_n2040# 2.42e-19
C427 passgatesCtrl_0.net7 a_n1361_n1429# 1.77e-19
C428 passgatex4_0.GP2 passgatesCtrl_0._00_ 3.42e-20
C429 VDD a_n995_n3605# 0.218874f
C430 VDD a_n1173_n2218# 0.118575f
C431 a_n1637_n1429# passgatesCtrl_0.net2 6.58e-20
C432 passgatex4_0.GP3 A2 0.001646f
C433 a_n951_n2736# passgatesCtrl_0.net7 0.001413f
C434 A3 Z4 0.005563f
C435 passgatex4_0.GN4 a_n1361_n1429# 5.36e-19
C436 a_n1503_n2192# a_n1361_n1429# 0.010239f
C437 passgatex4_0.GN1 passgatex4_0.GP1 1.11922f
C438 a_n715_n3850# a_n539_n3518# 0.185422f
C439 passgatex4_0.GP3 a_n2639_n2040# 0.002737f
C440 passgatex4_0.GN2 a_n675_n1648# 0.021336f
C441 passgatex4_0.GP2 Z4 6e-21
C442 a_n1701_n4368# a_n1878_n4368# 0.134298f
C443 VDD a_n2480_n4368# 0.27871f
C444 passgatex4_0.GN1 a_n1227_n2736# 0.109645f
C445 VDD Z3 2.85844f
C446 passgatesCtrl_0._05_ passgatesCtrl_0._00_ 0.005299f
C447 a_n491_n3280# passgatesCtrl_0.net2 0.013113f
C448 passgatesCtrl_0.net6 passgatesCtrl_0.net10 0.043833f
C449 passgatesCtrl_0.net6 passgatex4_0.GP3 2.34e-19
C450 VDD passgatesCtrl_0.net9 0.312028f
C451 passgatex4_0.GP4 a_n2189_n1429# 0.130626f
C452 passgatex4_0.GN1 a_n1045_n1942# 3.88e-20
C453 a_n587_n3458# passgatesCtrl_0._04_ 8.17e-20
C454 a_n2975_n2192# passgatesCtrl_0._00_ 0.012253f
C455 passgatesCtrl_0._01_ passgatex4_0.GN1 4.4e-20
C456 passgatex4_0.GP4 A3 0.001593f
C457 passgatex4_0.GP1 passgatex4_0.GN2 1.62948f
C458 a_n597_n2040# a_n1003_n2040# 4.09e-20
C459 a_n1701_n4368# a_n1984_n4368# 0.003683f
C460 VDD passgatesCtrl_0.net5 0.609808f
C461 passgatex4_0.GP2 passgatex4_0.GP4 3.49e-19
C462 passgatesCtrl_0.net1 a_n988_n4394# 0.019707f
C463 passgatesCtrl_0.net7 a_n675_n1648# 0.109167f
C464 a_n1227_n2736# passgatex4_0.GN2 9.69e-19
C465 passgatesCtrl_0.net1 a_n434_n1942# 3.05e-19
C466 passgatex4_0.GN1 a_n801_n4216# 6.45e-19
C467 VDD a_n715_n3850# 0.182247f
C468 passgatesCtrl_0._01_ a_n2015_n2040# 0.002311f
C469 passgatesCtrl_0.net1 passgatesCtrl_0._02_ 0.079473f
C470 a_n1361_n1429# a_n1085_n1429# 5.3e-19
C471 a_n491_n3280# A1 0.001919f
C472 passgatesCtrl_0._03_ a_n1963_n3280# 0.225915f
C473 A4 A2 2.39e-19
C474 VDD a_n2057_n1942# 4.1e-19
C475 a_n2015_n2040# a_n2185_n2218# 0.101254f
C476 passgatesCtrl_0.net1 passgatesCtrl_0.net8 0.194974f
C477 a_n491_n3280# passgatesCtrl_0.net3 1.85e-19
C478 passgatesCtrl_0._01_ passgatex4_0.GN2 6.19e-19
C479 passgatex4_0.GN3 passgatesCtrl_0._02_ 1.13e-19
C480 VDD a_n1878_n4368# 0.211692f
C481 a_n1701_n4368# select0 2.23e-19
C482 a_n1135_n4368# a_n1084_n4216# 0.134298f
C483 passgatex4_0.GP4 passgatesCtrl_0._05_ 6.86e-20
C484 passgatesCtrl_0.net1 a_n2189_n1429# 0.030465f
C485 passgatesCtrl_0.net7 passgatesCtrl_0._03_ 0.001559f
C486 passgatex4_0.GN3 passgatesCtrl_0.net8 0.002415f
C487 VDD A2 1.62685f
C488 a_n988_n4394# a_n995_n3605# 0.011149f
C489 a_n1084_n4216# passgatesCtrl_0._04_ 2.48e-19
C490 passgatesCtrl_0.net7 passgatex4_0.GP1 0.068983f
C491 a_n1913_n1429# passgatesCtrl_0.net10 0.219762f
C492 passgatex4_0.GN3 a_n2189_n1429# 0.011181f
C493 select0 a_n539_n3518# 8.27e-19
C494 passgatesCtrl_0.net2 a_n1361_n1429# 1.59e-20
C495 VDD a_n2639_n2040# 0.20743f
C496 a_n2429_n1328# passgatesCtrl_0.net10 0.009374f
C497 a_n1227_n2736# passgatesCtrl_0.net7 6.38e-19
C498 passgatex4_0.GP2 passgatesCtrl_0.net1 7.04e-20
C499 passgatex4_0.GN1 a_n597_n2040# 6.11e-19
C500 passgatex4_0.GN3 A3 3.80702f
C501 a_n2429_n1328# passgatex4_0.GP3 1.66e-19
C502 a_n1173_n2218# passgatesCtrl_0.net8 0.015061f
C503 passgatex4_0.GN4 passgatex4_0.GP1 3.45e-19
C504 a_n1503_n2192# passgatex4_0.GP1 3.01e-21
C505 a_n951_n2736# passgatesCtrl_0.net2 1.46e-19
C506 passgatesCtrl_0.net4 a_n539_n3518# 1.79e-19
C507 VDD passgatesCtrl_0.net6 0.615644f
C508 passgatex4_0.GN3 passgatex4_0.GP2 2.40528f
C509 VDD a_n1984_n4368# 0.222008f
C510 passgatesCtrl_0.net2 Z1 2.55e-19
C511 a_n1135_n4368# passgatesCtrl_0.net2 6.62e-19
C512 passgatesCtrl_0._05_ passgatesCtrl_0.net1 0.001365f
C513 passgatex4_0.GP1 Z2 0.065749f
C514 passgatex4_0.GP2 a_n1173_n2218# 5.22e-19
C515 passgatesCtrl_0.net2 passgatesCtrl_0._04_ 0.096582f
C516 select1 a_n1459_n3306# 3.4e-19
C517 a_n1085_n1429# a_n675_n1648# 0.031466f
C518 passgatex4_0.GN1 passgatex4_0.GP3 3.37e-19
C519 a_n597_n2040# passgatex4_0.GN2 0.009622f
C520 passgatex4_0.GP4 passgatesCtrl_0._00_ 0.039155f
C521 passgatesCtrl_0._01_ a_n1503_n2192# 0.213841f
C522 VDD select0 0.625418f
C523 passgatesCtrl_0.net1 a_n2975_n2192# 7.01e-19
C524 passgatex4_0.GN4 a_n2185_n2218# 2.2e-21
C525 a_n1361_n1429# passgatesCtrl_0.net3 6.41e-20
C526 A3 Z3 4.51555f
C527 passgatesCtrl_0._03_ a_n1635_n3306# 0.074703f
C528 a_n2189_n1429# passgatesCtrl_0.net9 0.219432f
C529 a_n482_n4216# a_n539_n3518# 0.003312f
C530 a_n1635_n3306# passgatex4_0.GP1 6.97e-20
C531 a_n951_n2736# A1 1.79e-20
C532 passgatesCtrl_0.net5 passgatesCtrl_0._02_ 4.38e-19
C533 passgatesCtrl_0.net2 a_n2161_n4368# 0.383661f
C534 passgatex4_0.GP2 Z3 0.063817f
C535 a_n1227_n2736# a_n1084_n4216# 4.03e-19
C536 passgatex4_0.GP4 Z4 0.278468f
C537 passgatesCtrl_0.net5 passgatesCtrl_0.net8 0.012208f
C538 passgatesCtrl_0.net2 a_n675_n1648# 1.87e-20
C539 A1 Z1 4.51541f
C540 a_n951_n2736# passgatesCtrl_0.net3 0.037807f
C541 VDD passgatesCtrl_0.net4 0.442407f
C542 VDD a_n1003_n2040# 0.076471f
C543 passgatex4_0.GN1 a_n539_n3518# 0.001234f
C544 passgatesCtrl_0.net10 passgatex4_0.GN2 4.61e-20
C545 passgatex4_0.GP2 passgatesCtrl_0.net9 8.22e-21
C546 passgatesCtrl_0.net5 a_n2189_n1429# 0.002712f
C547 a_n1135_n4368# A1 2.48e-21
C548 passgatex4_0.GP3 passgatex4_0.GN2 0.001327f
C549 a_n1878_n4368# a_n988_n4394# 1.1e-19
C550 passgatesCtrl_0._04_ A1 2.11e-20
C551 a_n1227_n2736# a_n1085_n1429# 2.57e-19
C552 passgatesCtrl_0.net7 a_n597_n2040# 0.010689f
C553 VDD a_n1913_n1429# 0.196943f
C554 passgatesCtrl_0.net10 a_n2883_n1648# 5.56e-19
C555 VDD a_n2429_n1328# 1.96e-19
C556 passgatex4_0.GP3 a_n2883_n1648# 0.008642f
C557 passgatesCtrl_0.net1 passgatesCtrl_0._00_ 0.110008f
C558 passgatex4_0.GP2 passgatesCtrl_0.net5 0.125101f
C559 passgatesCtrl_0._03_ passgatesCtrl_0.net2 0.265291f
C560 passgatesCtrl_0.net2 passgatex4_0.GP1 0.078988f
C561 passgatex4_0.GN3 passgatesCtrl_0._00_ 6.68e-20
C562 passgatesCtrl_0.net4 a_n1507_n3280# 5.55e-19
C563 a_n1503_n2192# a_n597_n2040# 1.1e-19
C564 VDD a_n482_n4216# 0.290651f
C565 a_n1227_n2736# passgatesCtrl_0.net2 0.006314f
C566 passgatesCtrl_0.net2 a_n2465_n2164# 0.001995f
C567 a_n988_n4394# a_n1984_n4368# 0.002297f
C568 A1 a_n675_n1648# 2.71e-20
C569 passgatesCtrl_0.net7 passgatesCtrl_0.net10 4.64e-20
C570 A3 A2 1.81997f
C571 a_n1459_n3306# passgatesCtrl_0.net1 0.20481f
C572 passgatex4_0.GN3 Z4 1.95e-20
C573 select1 passgatesCtrl_0.net1 0.002895f
C574 a_n1173_n2218# passgatesCtrl_0._00_ 1.7e-21
C575 VDD passgatex4_0.GN1 0.938241f
C576 passgatesCtrl_0.net6 passgatesCtrl_0.net8 0.02671f
C577 passgatesCtrl_0.net2 a_n1045_n1942# 0.001911f
C578 passgatex4_0.GP2 A2 3.97567f
C579 passgatesCtrl_0._01_ passgatesCtrl_0.net2 0.218705f
C580 passgatesCtrl_0.net6 a_n2189_n1429# 1.92e-20
C581 passgatex4_0.GN4 passgatesCtrl_0.net10 0.039325f
C582 passgatesCtrl_0.net2 a_n2185_n2218# 0.042928f
C583 select0 a_n988_n4394# 0.001977f
C584 passgatex4_0.GN4 passgatex4_0.GP3 3.23503f
C585 A1 passgatex4_0.GP1 4.03203f
C586 VDD a_n2015_n2040# 0.097823f
C587 passgatex4_0.GP4 passgatesCtrl_0.net1 0.00512f
C588 passgatesCtrl_0.net7 a_n539_n3518# 0.004605f
C589 a_n801_n4216# passgatesCtrl_0.net2 6.52e-19
C590 select1 a_n995_n3605# 2.55e-19
C591 passgatesCtrl_0.net3 passgatex4_0.GP1 0.001814f
C592 passgatex4_0.GP2 passgatesCtrl_0.net6 0.001965f
C593 passgatesCtrl_0.net9 passgatesCtrl_0._00_ 0.099215f
C594 VDD passgatex4_0.GN2 0.389408f
C595 passgatex4_0.GN3 passgatex4_0.GP4 0.048689f
C596 a_n1227_n2736# passgatesCtrl_0.net3 0.23425f
C597 passgatex4_0.GP3 Z2 1.03e-20
C598 passgatesCtrl_0._05_ a_n2639_n2040# 0.114102f
C599 Z3 Z4 0.002331f
C600 a_n1003_n2040# passgatesCtrl_0._02_ 0.054258f
C601 VDD a_n2883_n1648# 0.258847f
C602 select1 a_n2480_n4368# 0.270124f
C603 passgatesCtrl_0.net4 passgatesCtrl_0.net8 5.72e-20
C604 passgatesCtrl_0.net5 passgatesCtrl_0._00_ 0.002004f
C605 a_n1003_n2040# passgatesCtrl_0.net8 0.002587f
C606 a_n2975_n2192# a_n2639_n2040# 0.015664f
C607 passgatesCtrl_0.net6 passgatesCtrl_0._05_ 0.289483f
C608 a_n1637_n1429# a_n1361_n1429# 5.3e-19
C609 passgatesCtrl_0._01_ passgatesCtrl_0.net3 6.43e-19
C610 VDD a_n1963_n3280# 0.266692f
C611 passgatesCtrl_0.net2 a_n597_n2040# 0.154638f
C612 a_n801_n4216# A1 1.16e-20
C613 passgatesCtrl_0.net8 a_n1913_n1429# 3.98e-20
C614 a_n1085_n1429# passgatesCtrl_0.net10 2.12e-19
C615 a_n2057_n1942# passgatesCtrl_0._00_ 3.51e-19
C616 passgatesCtrl_0.net6 a_n2975_n2192# 0.108594f
C617 passgatex4_0.GP1 a_n485_n2736# 2.46e-19
C618 a_n2189_n1429# a_n1913_n1429# 5.3e-19
C619 VDD passgatesCtrl_0.net7 0.589224f
C620 passgatex4_0.GN4 A4 3.8425f
C621 passgatex4_0.GP4 Z3 1.58e-20
C622 a_n1459_n3306# passgatesCtrl_0.net5 7.33e-19
C623 passgatex4_0.GN3 passgatesCtrl_0.net1 0.027691f
C624 select1 passgatesCtrl_0.net5 2.72e-19
C625 passgatex4_0.GN1 a_n988_n4394# 4.16e-19
C626 VDD a_n587_n3458# 2.56e-19
C627 passgatex4_0.GP4 passgatesCtrl_0.net9 0.376983f
C628 select1 a_n715_n3850# 1.42e-19
C629 passgatex4_0.GN1 a_n434_n1942# 1.09e-19
C630 a_n2639_n2040# passgatesCtrl_0._00_ 0.054291f
C631 VDD passgatex4_0.GN4 0.255383f
C632 passgatesCtrl_0.net2 passgatesCtrl_0.net10 0.082322f
C633 VDD a_n1503_n2192# 0.26412f
C634 passgatesCtrl_0.net2 passgatex4_0.GP3 0.137787f
C635 passgatex4_0.GN1 passgatesCtrl_0._02_ 0.005251f
C636 passgatesCtrl_0.net1 a_n995_n3605# 0.008453f
C637 passgatesCtrl_0.net1 a_n1173_n2218# 0.059436f
C638 a_n491_n3280# Z1 1.26e-20
C639 passgatex4_0.GN1 passgatesCtrl_0.net8 1.87e-19
C640 passgatex4_0.GP4 passgatesCtrl_0.net5 0.005756f
C641 select1 a_n1878_n4368# 0.009355f
C642 passgatesCtrl_0.net6 passgatesCtrl_0._00_ 0.194746f
C643 a_n597_n2040# passgatesCtrl_0.net3 7.1e-21
C644 a_n1701_n4368# passgatesCtrl_0.net2 0.003464f
C645 VDD Z2 2.84785f
C646 passgatesCtrl_0.net2 a_n539_n3518# 0.242957f
C647 passgatex4_0.GP2 passgatex4_0.GN1 0.002408f
C648 passgatex4_0.GN2 passgatesCtrl_0._02_ 0.237149f
C649 VDD a_n1084_n4216# 0.201932f
C650 passgatex4_0.GN3 Z3 0.427101f
C651 passgatesCtrl_0.net1 passgatesCtrl_0.net9 0.061468f
C652 VDD a_n1635_n3306# 0.225849f
C653 select1 a_n1984_n4368# 0.00809f
C654 passgatex4_0.GP4 A2 1.28e-19
C655 passgatesCtrl_0.net8 passgatex4_0.GN2 0.00108f
C656 passgatex4_0.GP3 A1 2.76e-19
C657 passgatex4_0.GN3 passgatesCtrl_0.net9 0.015603f
C658 passgatex4_0.GP4 a_n2639_n2040# 1.28e-20
C659 VDD a_n1085_n1429# 0.219592f
C660 passgatesCtrl_0.net1 passgatesCtrl_0.net5 0.088832f
C661 A3 passgatex4_0.GN2 0.00661f
C662 a_n2189_n1429# a_n2883_n1648# 0.002068f
C663 passgatesCtrl_0.net1 a_n715_n3850# 0.224224f
C664 passgatex4_0.GN3 passgatesCtrl_0.net5 0.188564f
C665 passgatex4_0.GP4 passgatesCtrl_0.net6 2.47e-20
C666 passgatex4_0.GP2 passgatex4_0.GN2 1.51461f
C667 passgatesCtrl_0.net7 a_n434_n1942# 5.23e-19
C668 select1 select0 0.083731f
C669 a_n539_n3518# A1 0.002355f
C670 passgatesCtrl_0.net1 a_n2057_n1942# 0.00235f
C671 passgatesCtrl_0._03_ a_n491_n3280# 7.41e-20
C672 a_n491_n3280# passgatex4_0.GP1 0.109714f
C673 a_n1635_n3306# a_n1507_n3280# 0.004764f
C674 passgatesCtrl_0.net7 passgatesCtrl_0._02_ 0.003983f
C675 a_n1913_n1429# passgatesCtrl_0._00_ 2.75e-19
C676 a_n539_n3518# passgatesCtrl_0.net3 6.41e-21
C677 VDD passgatesCtrl_0.net2 3.00507f
C678 passgatesCtrl_0.net7 passgatesCtrl_0.net8 2.52e-19
C679 passgatesCtrl_0.net1 a_n1878_n4368# 6.03e-19
C680 a_n1173_n2218# passgatesCtrl_0.net5 0.001684f
C681 a_n951_n2736# Z1 1e-20
C682 passgatesCtrl_0.net4 a_n1459_n3306# 0.010474f
C683 passgatesCtrl_0._01_ a_n1637_n1429# 2.78e-19
C684 passgatesCtrl_0.net4 select1 0.003108f
C685 passgatesCtrl_0.net7 a_n2189_n1429# 2.69e-20
C686 a_n715_n3850# a_n995_n3605# 3.02e-19
C687 passgatesCtrl_0.net1 a_n2639_n2040# 0.084866f
C688 a_n1503_n2192# passgatesCtrl_0._02_ 4.67e-20
C689 passgatex4_0.GN3 A2 0.161523f
C690 passgatex4_0.GN4 passgatesCtrl_0.net8 5.26e-19
C691 a_n1503_n2192# passgatesCtrl_0.net8 0.107924f
C692 passgatesCtrl_0._05_ a_n2883_n1648# 6.71e-20
C693 passgatex4_0.GN4 a_n2189_n1429# 2.84e-19
C694 passgatex4_0.GP2 passgatesCtrl_0.net7 3.18e-19
C695 passgatesCtrl_0.net6 passgatesCtrl_0.net1 0.502444f
C696 passgatesCtrl_0.net2 a_n1507_n3280# 5.53e-19
C697 passgatesCtrl_0.net1 a_n1984_n4368# 2.27e-19
C698 passgatex4_0.GN4 A3 0.183073f
C699 passgatesCtrl_0.net5 passgatesCtrl_0.net9 0.011574f
C700 a_n1084_n4216# a_n988_n4394# 0.313533f
C701 VDD A1 1.84639f
C702 a_n2975_n2192# a_n2883_n1648# 1.44e-19
C703 passgatex4_0.GN3 passgatesCtrl_0.net6 0.151115f
C704 passgatex4_0.GP2 passgatex4_0.GN4 0.041571f
C705 a_n1503_n2192# passgatex4_0.GP2 3.34e-21
C706 VDD passgatesCtrl_0.net3 0.348944f
C707 passgatex4_0.GP4 a_n1913_n1429# 0.109546f
C708 Z1 a_n675_n1648# 3.24e-20
C709 passgatex4_0.GP4 a_n2429_n1328# 5.08e-19
C710 a_n2015_n2040# passgatesCtrl_0._00_ 1.34e-19
C711 passgatex4_0.GN1 a_n1459_n3306# 4.47e-21
C712 Z3 A2 0.004565f
C713 passgatex4_0.GN1 select1 1.61e-19
C714 A3 Z2 1.49e-20
C715 passgatesCtrl_0.net6 a_n1173_n2218# 2.62e-19
C716 select0 passgatesCtrl_0.net1 0.025769f
C717 a_n1085_n1429# passgatesCtrl_0._02_ 7.02e-19
C718 passgatex4_0.GP2 Z2 0.278333f
C719 passgatex4_0.GN4 passgatesCtrl_0._05_ 3.95e-20
C720 passgatesCtrl_0.net5 a_n2057_n1942# 2.64e-19
C721 a_n1085_n1429# passgatesCtrl_0.net8 0.201804f
C722 passgatesCtrl_0.net9 a_n2639_n2040# 2.03e-19
C723 a_n951_n2736# passgatex4_0.GP1 9.85e-21
C724 passgatesCtrl_0.net4 passgatesCtrl_0.net1 0.142351f
C725 passgatesCtrl_0._00_ a_n2883_n1648# 0.229802f
C726 passgatesCtrl_0.net1 a_n1003_n2040# 0.158092f
C727 passgatesCtrl_0.net2 a_n988_n4394# 7.27e-19
C728 Z1 passgatex4_0.GP1 0.278495f
C729 passgatesCtrl_0.net5 a_n1878_n4368# 3.52e-19
C730 passgatesCtrl_0.net2 a_n434_n1942# 9.54e-19
C731 a_n951_n2736# a_n1227_n2736# 5.3e-19
C732 passgatex4_0.GN1 passgatex4_0.GP4 1.4e-19
C733 a_n1637_n1429# passgatesCtrl_0.net10 0.030972f
C734 VDD a_n485_n2736# 0.00616f
C735 passgatesCtrl_0._01_ a_n1361_n1429# 1.94e-20
C736 passgatesCtrl_0.net6 passgatesCtrl_0.net9 5.48e-19
C737 passgatesCtrl_0.net2 passgatesCtrl_0._02_ 0.092244f
C738 passgatesCtrl_0.net1 a_n1913_n1429# 0.006122f
C739 passgatex4_0.GP2 a_n1085_n1429# 0.11066f
C740 passgatesCtrl_0.net2 passgatesCtrl_0.net8 0.129f
C741 passgatex4_0.GN3 a_n1913_n1429# 0.034066f
C742 a_n1135_n4368# a_n1227_n2736# 1.17e-20
C743 passgatesCtrl_0.net2 a_n2189_n1429# 3.62e-20
C744 passgatesCtrl_0.net4 a_n995_n3605# 0.110271f
C745 passgatesCtrl_0.net4 a_n1173_n2218# 0.001325f
C746 passgatex4_0.GN3 a_n2429_n1328# 9.54e-20
C747 a_n1003_n2040# a_n995_n3605# 4.27e-20
C748 a_n1173_n2218# a_n1003_n2040# 0.101254f
C749 passgatesCtrl_0.net6 passgatesCtrl_0.net5 0.372649f
C750 passgatesCtrl_0.net5 a_n1984_n4368# 1.71e-19
C751 select1 a_n1963_n3280# 3.96e-19
C752 a_n482_n4216# passgatesCtrl_0.net1 0.167305f
C753 passgatex4_0.GP4 passgatex4_0.GN2 3.27e-19
C754 passgatex4_0.GN4 passgatesCtrl_0._00_ 3.91e-19
C755 a_n988_n4394# A1 1.54e-20
C756 passgatex4_0.GP1 a_n675_n1648# 0.001422f
C757 passgatex4_0.GP2 passgatesCtrl_0.net2 3.91e-20
C758 a_n1503_n2192# passgatesCtrl_0._00_ 5.79e-21
C759 Z4 VSS 2.706298f
C760 A4 VSS 3.775201f
C761 Z3 VSS 2.493104f
C762 A3 VSS 3.16981f
C763 Z2 VSS 2.453408f
C764 A2 VSS 3.285328f
C765 Z1 VSS 2.856037f
C766 A1 VSS 3.713512f
C767 select0 VSS 0.611662f
C768 select1 VSS 1.92417f
C769 VDD VSS 0.101815p
C770 a_n1135_n4368# VSS 0.171495f
C771 a_n1701_n4368# VSS 0.108493f
C772 a_n482_n4216# VSS 0.309602f
C773 a_n801_n4216# VSS 0.268985f
C774 a_n988_n4394# VSS 0.277513f
C775 a_n1084_n4216# VSS 0.27241f
C776 a_n1878_n4368# VSS 0.260674f
C777 a_n1984_n4368# VSS 0.250918f
C778 a_n2161_n4368# VSS 0.286148f
C779 a_n2480_n4368# VSS 0.328097f
C780 a_n587_n3458# VSS 0.005492f
C781 a_n539_n3518# VSS 0.241098f
C782 a_n715_n3850# VSS 0.229487f
C783 passgatesCtrl_0._04_ VSS 0.264876f
C784 a_n995_n3605# VSS 0.260858f
C785 a_n1507_n3280# VSS 0.005035f
C786 passgatex4_0.GP1 VSS 2.27865f
C787 a_n491_n3280# VSS 0.274026f
C788 a_n1459_n3306# VSS 0.254131f
C789 a_n1635_n3306# VSS 0.235093f
C790 a_n1963_n3280# VSS 0.277418f
C791 passgatesCtrl_0._03_ VSS 0.368268f
C792 a_n485_n2736# VSS 2.19e-19
C793 passgatex4_0.GN2 VSS 4.32804f
C794 passgatex4_0.GN1 VSS 3.99205f
C795 a_n951_n2736# VSS 0.268527f
C796 passgatesCtrl_0.net4 VSS 0.647109f
C797 a_n1227_n2736# VSS 0.2678f
C798 passgatesCtrl_0.net3 VSS 0.42716f
C799 a_n434_n1942# VSS 5.62e-19
C800 a_n1045_n1942# VSS 7.49e-19
C801 a_n1003_n2040# VSS 0.298899f
C802 a_n2465_n2164# VSS 0.005723f
C803 a_n2057_n1942# VSS 8.59e-19
C804 a_n2015_n2040# VSS 0.295323f
C805 a_n597_n2040# VSS 0.234177f
C806 a_n1173_n2218# VSS 0.254047f
C807 a_n1503_n2192# VSS 0.224474f
C808 passgatesCtrl_0._01_ VSS 0.199048f
C809 a_n2185_n2218# VSS 0.267196f
C810 a_n2639_n2040# VSS 0.257089f
C811 a_n2975_n2192# VSS 0.252788f
C812 passgatesCtrl_0._05_ VSS 0.341727f
C813 passgatesCtrl_0.net7 VSS 0.453064f
C814 passgatex4_0.GP2 VSS 2.23556f
C815 passgatex4_0.GN3 VSS 3.82555f
C816 passgatex4_0.GN4 VSS 5.2369f
C817 passgatex4_0.GP4 VSS 5.2081f
C818 passgatex4_0.GP3 VSS 2.17467f
C819 a_n2429_n1328# VSS 0.001779f
C820 a_n675_n1648# VSS 0.258431f
C821 passgatesCtrl_0._02_ VSS 0.366887f
C822 passgatesCtrl_0.net8 VSS 0.333624f
C823 a_n1085_n1429# VSS 0.250109f
C824 passgatesCtrl_0.net5 VSS 0.6309f
C825 a_n1361_n1429# VSS 0.21514f
C826 passgatesCtrl_0.net6 VSS 0.300978f
C827 a_n1637_n1429# VSS 0.2182f
C828 passgatesCtrl_0.net10 VSS -0.162684f
C829 a_n1913_n1429# VSS 0.220816f
C830 passgatesCtrl_0.net9 VSS 0.33083f
C831 a_n2189_n1429# VSS 0.238577f
C832 passgatesCtrl_0.net1 VSS 3.170257f
C833 passgatesCtrl_0.net2 VSS 4.630451f
C834 a_n2883_n1648# VSS 0.241645f
C835 passgatesCtrl_0._00_ VSS 0.297612f
C836 A1.t0 VSS 0.838615f
C837 A1.t1 VSS 0.481433f
C838 A1.n0 VSS 4.66276f
C839 A1.t2 VSS 0.867976f
C840 A1.t3 VSS 0.614013f
C841 A1.n1 VSS 4.76729f
C842 A1.n2 VSS 0.754061f
C843 A1.n3 VSS 0.235366f
C844 Z1.t1 VSS 0.368287f
C845 Z1.n0 VSS 0.549919f
C846 Z1.t0 VSS 0.37568f
C847 Z1.t2 VSS 0.498536f
C848 Z1.n1 VSS 2.51576f
C849 Z1.n2 VSS 0.851227f
C850 Z1.t3 VSS 0.485176f
C851 Z1.n3 VSS 0.603414f
C852 Z1.n4 VSS 0.766774f
C853 A4.t0 VSS 0.893471f
C854 A4.t1 VSS 0.512925f
C855 A4.n0 VSS 4.96776f
C856 A4.t3 VSS 0.924752f
C857 A4.t2 VSS 0.654177f
C858 A4.n1 VSS 5.07912f
C859 A4.n2 VSS 0.803386f
C860 A4.n3 VSS 0.175929f
C861 Z4.t1 VSS 0.356732f
C862 Z4.n0 VSS 0.532664f
C863 Z4.t0 VSS 0.363892f
C864 Z4.t3 VSS 0.482893f
C865 Z4.n1 VSS 2.43682f
C866 Z4.n2 VSS 0.824519f
C867 Z4.t2 VSS 0.469953f
C868 Z4.n3 VSS 0.584481f
C869 Z4.n4 VSS 0.742715f
C870 A2.t3 VSS 0.763965f
C871 A2.t2 VSS 0.438578f
C872 A2.n0 VSS 4.2477f
C873 A2.t0 VSS 0.790712f
C874 A2.t1 VSS 0.559356f
C875 A2.n1 VSS 4.34292f
C876 A2.n2 VSS 0.686937f
C877 A2.n3 VSS 0.222065f
C878 Z2.t2 VSS 0.358466f
C879 Z2.n0 VSS 0.535254f
C880 Z2.t3 VSS 0.365662f
C881 Z2.t0 VSS 0.485241f
C882 Z2.n1 VSS 2.44867f
C883 Z2.n2 VSS 0.828528f
C884 Z2.t1 VSS 0.472238f
C885 Z2.n3 VSS 0.587323f
C886 Z2.n4 VSS 0.723782f
C887 Z2.n5 VSS 0.319875f
C888 Z3.t0 VSS 0.361967f
C889 Z3.n0 VSS 0.540482f
C890 Z3.t1 VSS 0.369233f
C891 Z3.t3 VSS 0.48998f
C892 Z3.n1 VSS 2.47259f
C893 Z3.n2 VSS 0.83662f
C894 Z3.t2 VSS 0.47685f
C895 Z3.n3 VSS 0.593059f
C896 Z3.n4 VSS 0.728589f
C897 Z3.n5 VSS 0.33185f
C898 A3.t0 VSS 0.893706f
C899 A3.t1 VSS 0.51306f
C900 A3.n0 VSS 4.969069f
C901 A3.t3 VSS 0.924996f
C902 A3.t2 VSS 0.654349f
C903 A3.n1 VSS 5.08046f
C904 A3.n2 VSS 0.803598f
C905 A3.n3 VSS 0.264739f
C906 passgatesCtrl_0.net1.n0 VSS 0.226539f
C907 passgatesCtrl_0.net1.t1 VSS 0.053408f
C908 passgatesCtrl_0.net1.n1 VSS 0.014253f
C909 passgatesCtrl_0.net1.t0 VSS 0.033625f
C910 passgatesCtrl_0.net1.n2 VSS 0.02627f
C911 passgatesCtrl_0.net1.t11 VSS 0.01948f
C912 passgatesCtrl_0.net1.t2 VSS 0.013193f
C913 passgatesCtrl_0.net1.n3 VSS 0.052945f
C914 passgatesCtrl_0.net1.n4 VSS 0.021541f
C915 passgatesCtrl_0.net1.n5 VSS 0.027845f
C916 passgatesCtrl_0.net1.t3 VSS 0.015219f
C917 passgatesCtrl_0.net1.t8 VSS 0.024374f
C918 passgatesCtrl_0.net1.n6 VSS 0.046451f
C919 passgatesCtrl_0.net1.n7 VSS 0.05146f
C920 passgatesCtrl_0.net1.t13 VSS 0.016147f
C921 passgatesCtrl_0.net1.t12 VSS 0.011096f
C922 passgatesCtrl_0.net1.n8 VSS 0.046923f
C923 passgatesCtrl_0.net1.n9 VSS 0.01118f
C924 passgatesCtrl_0.net1.n10 VSS 0.021551f
C925 passgatesCtrl_0.net1.n11 VSS 0.171457f
C926 passgatesCtrl_0.net1.t9 VSS 0.022577f
C927 passgatesCtrl_0.net1.t17 VSS 0.052767f
C928 passgatesCtrl_0.net1.n12 VSS 0.058498f
C929 passgatesCtrl_0.net1.n13 VSS 0.193324f
C930 passgatesCtrl_0.net1.t10 VSS 0.010521f
C931 passgatesCtrl_0.net1.t5 VSS 0.012736f
C932 passgatesCtrl_0.net1.n14 VSS 0.042403f
C933 passgatesCtrl_0.net1.n15 VSS 0.009709f
C934 passgatesCtrl_0.net1.t16 VSS 0.010838f
C935 passgatesCtrl_0.net1.t18 VSS 0.013595f
C936 passgatesCtrl_0.net1.n16 VSS 0.030532f
C937 passgatesCtrl_0.net1.t14 VSS 0.015192f
C938 passgatesCtrl_0.net1.t19 VSS 0.024522f
C939 passgatesCtrl_0.net1.n17 VSS 0.049813f
C940 passgatesCtrl_0.net1.n18 VSS 0.013363f
C941 passgatesCtrl_0.net1.n19 VSS 0.13082f
C942 passgatesCtrl_0.net1.t6 VSS 0.019673f
C943 passgatesCtrl_0.net1.t15 VSS 0.013358f
C944 passgatesCtrl_0.net1.n20 VSS 0.046479f
C945 passgatesCtrl_0.net1.n21 VSS 0.011125f
C946 passgatesCtrl_0.net1.n22 VSS 0.054042f
C947 passgatesCtrl_0.net1.n23 VSS 0.220245f
C948 passgatesCtrl_0.net1.t7 VSS 0.022351f
C949 passgatesCtrl_0.net1.t4 VSS 0.010599f
C950 passgatesCtrl_0.net1.n24 VSS 0.080089f
C951 passgatesCtrl_0.net1.n25 VSS 0.01726f
C952 passgatesCtrl_0.net1.n26 VSS 0.016365f
C953 passgatesCtrl_0.net10.t2 VSS -0.055929f
C954 passgatesCtrl_0.net10.t1 VSS -0.028065f
C955 passgatesCtrl_0.net10.t0 VSS -0.028065f
C956 passgatesCtrl_0.net10.n0 VSS -0.063496f
C957 passgatesCtrl_0.net10.t3 VSS -0.027227f
C958 passgatesCtrl_0.net10.t4 VSS -0.043656f
C959 passgatesCtrl_0.net10.n1 VSS -0.087973f
C960 passgatesCtrl_0.net10.n2 VSS -0.035052f
C961 passgatesCtrl_0.net10.n3 VSS -0.16161f
C962 VDD.n0 VSS 0.115638f
C963 VDD.n1 VSS 0.176137f
C964 VDD.n2 VSS 0.115638f
C965 VDD.n3 VSS 0.104151f
C966 VDD.n4 VSS 0.003054f
C967 VDD.n5 VSS 0.003159f
C968 VDD.n6 VSS 0.001813f
C969 VDD.n7 VSS 0.001417f
C970 VDD.t103 VSS 0.278603f
C971 VDD.t31 VSS 0.021284f
C972 VDD.t99 VSS 0.029392f
C973 VDD.t127 VSS 0.28885f
C974 VDD.t13 VSS 0.021284f
C975 VDD.t0 VSS 0.045608f
C976 VDD.t104 VSS 0.110472f
C977 VDD.n8 VSS 0.135354f
C978 VDD.n9 VSS 0.015324f
C979 VDD.t63 VSS 0.004539f
C980 VDD.n10 VSS 0.01112f
C981 VDD.n11 VSS 5.46e-19
C982 VDD.n12 VSS 0.00398f
C983 VDD.n13 VSS 0.003417f
C984 VDD.t35 VSS 0.004921f
C985 VDD.n14 VSS 0.009822f
C986 VDD.n15 VSS 0.004796f
C987 VDD.t180 VSS 0.065381f
C988 VDD.n16 VSS 0.029387f
C989 VDD.n17 VSS 0.005284f
C990 VDD.t1 VSS 0.001371f
C991 VDD.t2 VSS 0.001371f
C992 VDD.n18 VSS 0.002981f
C993 VDD.n19 VSS 0.006462f
C994 VDD.n20 VSS 0.001838f
C995 VDD.n21 VSS 0.001771f
C996 VDD.n22 VSS 0.003159f
C997 VDD.n23 VSS 0.104151f
C998 VDD.n24 VSS 0.003159f
C999 VDD.n25 VSS 0.002158f
C1000 VDD.n26 VSS 0.001417f
C1001 VDD.n27 VSS 0.001838f
C1002 VDD.n28 VSS 0.002585f
C1003 VDD.n29 VSS 0.001417f
C1004 VDD.n30 VSS 0.001771f
C1005 VDD.n31 VSS 0.001895f
C1006 VDD.t155 VSS 6.78e-19
C1007 VDD.t175 VSS 0.00103f
C1008 VDD.n32 VSS 0.00172f
C1009 VDD.n33 VSS 0.002685f
C1010 VDD.n34 VSS 0.001801f
C1011 VDD.n35 VSS 0.004842f
C1012 VDD.t159 VSS 0.001371f
C1013 VDD.t151 VSS 0.001371f
C1014 VDD.n36 VSS 0.003045f
C1015 VDD.n37 VSS 0.005284f
C1016 VDD.t192 VSS 0.026295f
C1017 VDD.t100 VSS 0.001371f
C1018 VDD.t158 VSS 0.001371f
C1019 VDD.n38 VSS 0.002981f
C1020 VDD.n39 VSS 0.013419f
C1021 VDD.t154 VSS 0.001371f
C1022 VDD.t126 VSS 0.001371f
C1023 VDD.n40 VSS 0.003045f
C1024 VDD.n41 VSS 0.008241f
C1025 VDD.n42 VSS 0.001838f
C1026 VDD.n43 VSS 0.001771f
C1027 VDD.n44 VSS 0.003159f
C1028 VDD.n45 VSS 0.40558f
C1029 VDD.n46 VSS 0.003054f
C1030 VDD.n47 VSS 0.003159f
C1031 VDD.n48 VSS 0.0021f
C1032 VDD.n49 VSS 0.001417f
C1033 VDD.n50 VSS 0.002642f
C1034 VDD.t44 VSS 0.004509f
C1035 VDD.t193 VSS 0.009569f
C1036 VDD.n52 VSS 0.024536f
C1037 VDD.t45 VSS 0.004509f
C1038 VDD.n53 VSS 0.013365f
C1039 VDD.n54 VSS 0.001838f
C1040 VDD.t29 VSS 0.004509f
C1041 VDD.t189 VSS 0.009569f
C1042 VDD.n56 VSS 0.024536f
C1043 VDD.t30 VSS 0.004509f
C1044 VDD.n57 VSS 0.013365f
C1045 VDD.n58 VSS 0.001871f
C1046 VDD.n59 VSS 0.002642f
C1047 VDD.n60 VSS 0.005284f
C1048 VDD.t167 VSS 0.00103f
C1049 VDD.t12 VSS 0.001556f
C1050 VDD.n61 VSS 0.004648f
C1051 VDD.t121 VSS 0.001371f
C1052 VDD.t165 VSS 0.001371f
C1053 VDD.n62 VSS 0.002981f
C1054 VDD.t102 VSS 0.00276f
C1055 VDD.n63 VSS 0.0092f
C1056 VDD.n64 VSS 0.00313f
C1057 VDD.t84 VSS 0.001371f
C1058 VDD.t98 VSS 0.001371f
C1059 VDD.n65 VSS 0.003045f
C1060 VDD.n66 VSS 0.004796f
C1061 VDD.n67 VSS 0.005284f
C1062 VDD.t109 VSS 0.001055f
C1063 VDD.t146 VSS 0.001556f
C1064 VDD.n68 VSS 0.004775f
C1065 VDD.t10 VSS 0.001371f
C1066 VDD.t80 VSS 0.001371f
C1067 VDD.n69 VSS 0.003045f
C1068 VDD.n70 VSS 0.007905f
C1069 VDD.n71 VSS 0.001838f
C1070 VDD.n72 VSS 0.001771f
C1071 VDD.n73 VSS 0.003159f
C1072 VDD.n74 VSS 0.003159f
C1073 VDD.n75 VSS 0.001771f
C1074 VDD.n76 VSS 0.003159f
C1075 VDD.t70 VSS 0.001371f
C1076 VDD.t6 VSS 0.001371f
C1077 VDD.n77 VSS 0.003045f
C1078 VDD.n78 VSS 0.007905f
C1079 VDD.n79 VSS 0.0012f
C1080 VDD.t148 VSS 0.001371f
C1081 VDD.t125 VSS 0.001371f
C1082 VDD.n80 VSS 0.003045f
C1083 VDD.n81 VSS 0.002642f
C1084 VDD.n82 VSS 0.001838f
C1085 VDD.n83 VSS 0.001417f
C1086 VDD.n84 VSS 0.001417f
C1087 VDD.n85 VSS 0.001771f
C1088 VDD.n86 VSS 4.88e-19
C1089 VDD.n87 VSS 0.002154f
C1090 VDD.n88 VSS 0.001522f
C1091 VDD.n89 VSS 0.008241f
C1092 VDD.t106 VSS 0.002717f
C1093 VDD.t72 VSS 0.001371f
C1094 VDD.t68 VSS 0.001371f
C1095 VDD.n90 VSS 0.003045f
C1096 VDD.n91 VSS 0.004767f
C1097 VDD.n92 VSS 0.001536f
C1098 VDD.n93 VSS 0.005284f
C1099 VDD.t134 VSS 0.001371f
C1100 VDD.t92 VSS 0.001371f
C1101 VDD.n94 VSS 0.003045f
C1102 VDD.t88 VSS 0.001055f
C1103 VDD.t119 VSS 0.001556f
C1104 VDD.n95 VSS 0.004765f
C1105 VDD.t123 VSS 0.006321f
C1106 VDD.t90 VSS 0.002709f
C1107 VDD.n96 VSS 0.005531f
C1108 VDD.n97 VSS 0.003159f
C1109 VDD.t115 VSS 0.006322f
C1110 VDD.t82 VSS 5.06e-19
C1111 VDD.t113 VSS 0.001358f
C1112 VDD.n98 VSS 0.006196f
C1113 VDD.t28 VSS 0.046562f
C1114 VDD.t107 VSS 0.024382f
C1115 VDD.t166 VSS 0.024212f
C1116 VDD.t120 VSS 0.016424f
C1117 VDD.t11 VSS 0.0149f
C1118 VDD.t164 VSS 0.021503f
C1119 VDD.t101 VSS 0.030985f
C1120 VDD.t83 VSS 0.006603f
C1121 VDD.t86 VSS 0.013545f
C1122 VDD.t108 VSS 0.013545f
C1123 VDD.t97 VSS 0.016593f
C1124 VDD.t145 VSS 0.026583f
C1125 VDD.t9 VSS 0.020149f
C1126 VDD.t79 VSS 0.015577f
C1127 VDD.t69 VSS 0.015577f
C1128 VDD.t5 VSS 0.025905f
C1129 VDD.t147 VSS 0.015408f
C1130 VDD.t124 VSS 0.031324f
C1131 VDD.t71 VSS 0.019979f
C1132 VDD.t67 VSS 0.032509f
C1133 VDD.t170 VSS 0.026583f
C1134 VDD.t87 VSS 0.005249f
C1135 VDD.t133 VSS 0.016593f
C1136 VDD.t118 VSS 0.0149f
C1137 VDD.t91 VSS 0.026921f
C1138 VDD.t122 VSS 0.011344f
C1139 VDD.t89 VSS 0.014223f
C1140 VDD.t114 VSS 0.014223f
C1141 VDD.t112 VSS 0.011852f
C1142 VDD.t16 VSS 0.046731f
C1143 VDD.t139 VSS 0.013545f
C1144 VDD.t77 VSS 0.011006f
C1145 VDD.t73 VSS 0.015577f
C1146 VDD.t143 VSS 0.038604f
C1147 VDD.t81 VSS 0.038991f
C1148 VDD.n99 VSS 0.001536f
C1149 VDD.n100 VSS 0.001838f
C1150 VDD.n101 VSS 0.001771f
C1151 VDD.n102 VSS 0.003159f
C1152 VDD.n103 VSS 0.185574f
C1153 VDD.n104 VSS 0.003159f
C1154 VDD.n105 VSS 0.001771f
C1155 VDD.t144 VSS 0.001371f
C1156 VDD.t74 VSS 0.001371f
C1157 VDD.n106 VSS 0.003045f
C1158 VDD.n107 VSS 0.007905f
C1159 VDD.n108 VSS 0.002642f
C1160 VDD.n109 VSS 0.001838f
C1161 VDD.n110 VSS 0.001417f
C1162 VDD.n111 VSS 0.001417f
C1163 VDD.n112 VSS 0.001771f
C1164 VDD.n113 VSS 0.002642f
C1165 VDD.n114 VSS 4.88e-19
C1166 VDD.n115 VSS 0.001838f
C1167 VDD.t78 VSS 0.001371f
C1168 VDD.t140 VSS 0.001371f
C1169 VDD.n116 VSS 0.003045f
C1170 VDD.n117 VSS 0.007905f
C1171 VDD.t17 VSS 0.004509f
C1172 VDD.t181 VSS 0.009569f
C1173 VDD.n119 VSS 0.024536f
C1174 VDD.t18 VSS 0.004509f
C1175 VDD.n120 VSS 0.013365f
C1176 VDD.t53 VSS 0.004509f
C1177 VDD.t177 VSS 0.009569f
C1178 VDD.n122 VSS 0.024536f
C1179 VDD.t54 VSS 0.004509f
C1180 VDD.n123 VSS 0.013365f
C1181 VDD.n124 VSS 0.005481f
C1182 VDD.n125 VSS 0.011299f
C1183 VDD.n126 VSS 0.001241f
C1184 VDD.n127 VSS 9.76e-19
C1185 VDD.n128 VSS 0.002158f
C1186 VDD.n129 VSS 0.002767f
C1187 VDD.n130 VSS 0.003054f
C1188 VDD.n131 VSS 0.197333f
C1189 VDD.n132 VSS 0.003054f
C1190 VDD.n133 VSS 0.002767f
C1191 VDD.n134 VSS 0.001813f
C1192 VDD.n135 VSS 0.002958f
C1193 VDD.n136 VSS 0.010251f
C1194 VDD.n137 VSS 0.006524f
C1195 VDD.n138 VSS 0.008048f
C1196 VDD.n139 VSS 9.46e-19
C1197 VDD.n140 VSS 0.001475f
C1198 VDD.n141 VSS 0.004796f
C1199 VDD.n142 VSS 0.00313f
C1200 VDD.n143 VSS 4.27e-19
C1201 VDD.n144 VSS 0.007931f
C1202 VDD.n145 VSS 0.001505f
C1203 VDD.n146 VSS 0.013321f
C1204 VDD.n147 VSS 0.004796f
C1205 VDD.n148 VSS 0.00313f
C1206 VDD.n149 VSS 0.005284f
C1207 VDD.n150 VSS 0.001536f
C1208 VDD.n151 VSS 0.008007f
C1209 VDD.n152 VSS 0.001795f
C1210 VDD.n153 VSS 0.001251f
C1211 VDD.n154 VSS 0.004193f
C1212 VDD.n155 VSS 0.001871f
C1213 VDD.n156 VSS 0.002767f
C1214 VDD.n157 VSS 0.003054f
C1215 VDD.n158 VSS 0.197333f
C1216 VDD.n159 VSS 0.003054f
C1217 VDD.n160 VSS 0.002767f
C1218 VDD.n161 VSS 0.002646f
C1219 VDD.n162 VSS 0.003819f
C1220 VDD.n163 VSS 0.00313f
C1221 VDD.n164 VSS 0.001282f
C1222 VDD.n165 VSS 0.007176f
C1223 VDD.n166 VSS 0.007926f
C1224 VDD.n167 VSS 0.001536f
C1225 VDD.n168 VSS 0.001638f
C1226 VDD.n169 VSS 0.004509f
C1227 VDD.n170 VSS 0.002671f
C1228 VDD.n171 VSS 0.00313f
C1229 VDD.n172 VSS 0.001587f
C1230 VDD.n173 VSS 0.007309f
C1231 VDD.n174 VSS 0.006996f
C1232 VDD.n175 VSS 0.001261f
C1233 VDD.n176 VSS 0.005284f
C1234 VDD.n177 VSS 0.004509f
C1235 VDD.n178 VSS 0.001771f
C1236 VDD.n179 VSS 0.003159f
C1237 VDD.n180 VSS 0.001417f
C1238 VDD.n181 VSS 0.001771f
C1239 VDD.n182 VSS 0.002767f
C1240 VDD.n183 VSS 4.92e-19
C1241 VDD.n184 VSS 0.001838f
C1242 VDD.n185 VSS 0.001577f
C1243 VDD.n186 VSS 0.011306f
C1244 VDD.n187 VSS 0.001838f
C1245 VDD.n188 VSS 0.001895f
C1246 VDD.n189 VSS 0.001771f
C1247 VDD.n190 VSS 0.002767f
C1248 VDD.n191 VSS 0.003054f
C1249 VDD.n192 VSS 0.237185f
C1250 VDD.n193 VSS 0.176137f
C1251 VDD.n194 VSS 0.384936f
C1252 VDD.n195 VSS 0.145773f
C1253 VDD.n196 VSS 0.003159f
C1254 VDD.n197 VSS 0.0021f
C1255 VDD.n198 VSS 0.001417f
C1256 VDD.n199 VSS 0.001417f
C1257 VDD.n200 VSS 0.001771f
C1258 VDD.n201 VSS 0.002642f
C1259 VDD.t32 VSS 0.004509f
C1260 VDD.t182 VSS 0.009569f
C1261 VDD.n203 VSS 0.024536f
C1262 VDD.t33 VSS 0.004509f
C1263 VDD.n204 VSS 0.013365f
C1264 VDD.n205 VSS 0.002642f
C1265 VDD.n206 VSS 0.001838f
C1266 VDD.t61 VSS 0.004509f
C1267 VDD.t188 VSS 0.009569f
C1268 VDD.n208 VSS 0.024536f
C1269 VDD.t62 VSS 0.004509f
C1270 VDD.n209 VSS 0.013365f
C1271 VDD.n210 VSS 0.001241f
C1272 VDD.n211 VSS 0.011306f
C1273 VDD.n212 VSS 0.001838f
C1274 VDD.n213 VSS 0.001895f
C1275 VDD.n214 VSS 0.001771f
C1276 VDD.n215 VSS 0.002767f
C1277 VDD.n216 VSS 0.003054f
C1278 VDD.n217 VSS 0.114872f
C1279 VDD.n218 VSS 0.003054f
C1280 VDD.n219 VSS 0.002767f
C1281 VDD.n220 VSS 3.49e-19
C1282 VDD.n221 VSS 0.002814f
C1283 VDD.n222 VSS 0.002613f
C1284 VDD.n223 VSS 0.001333f
C1285 VDD.t160 VSS 0.006334f
C1286 VDD.n224 VSS 0.010785f
C1287 VDD.t55 VSS 0.004472f
C1288 VDD.n225 VSS 0.007877f
C1289 VDD.n226 VSS 0.00348f
C1290 VDD.n227 VSS 0.002642f
C1291 VDD.n228 VSS 0.002498f
C1292 VDD.n229 VSS 0.004939f
C1293 VDD.n230 VSS 0.013871f
C1294 VDD.n231 VSS 0.019633f
C1295 VDD.t56 VSS 0.004472f
C1296 VDD.n232 VSS 0.007877f
C1297 VDD.n233 VSS 0.035693f
C1298 VDD.n234 VSS 0.00313f
C1299 VDD.n235 VSS 0.004796f
C1300 VDD.n236 VSS 0.002987f
C1301 VDD.n237 VSS 0.008233f
C1302 VDD.n238 VSS 0.00118f
C1303 VDD.n239 VSS 0.002786f
C1304 VDD.n240 VSS 0.002642f
C1305 VDD.n241 VSS 0.001085f
C1306 VDD.n242 VSS 0.001024f
C1307 VDD.t34 VSS 0.004921f
C1308 VDD.n243 VSS 0.003786f
C1309 VDD.n244 VSS 0.006238f
C1310 VDD.n245 VSS 0.005553f
C1311 VDD.n246 VSS 0.005274f
C1312 VDD.t105 VSS 9.3e-19
C1313 VDD.t128 VSS 0.003822f
C1314 VDD.n247 VSS 0.003518f
C1315 VDD.n248 VSS 0.002638f
C1316 VDD.n249 VSS 0.005017f
C1317 VDD.n250 VSS 0.005583f
C1318 VDD.n251 VSS 0.001838f
C1319 VDD.n252 VSS 0.002642f
C1320 VDD.n253 VSS 0.001771f
C1321 VDD.n254 VSS 0.002767f
C1322 VDD.n255 VSS 0.003054f
C1323 VDD.n256 VSS 0.114872f
C1324 VDD.n257 VSS 0.003054f
C1325 VDD.n258 VSS 0.002767f
C1326 VDD.n259 VSS 0.002646f
C1327 VDD.n260 VSS 0.004193f
C1328 VDD.n261 VSS 0.005284f
C1329 VDD.n262 VSS 0.00666f
C1330 VDD.n263 VSS 0.012423f
C1331 VDD.n264 VSS 0.005301f
C1332 VDD.n265 VSS 0.00313f
C1333 VDD.n266 VSS 0.002642f
C1334 VDD.n267 VSS 0.006595f
C1335 VDD.t14 VSS 0.004472f
C1336 VDD.n268 VSS 0.010271f
C1337 VDD.n269 VSS 0.018051f
C1338 VDD.n270 VSS 0.018051f
C1339 VDD.n271 VSS 0.005284f
C1340 VDD.n272 VSS 0.005284f
C1341 VDD.n273 VSS 0.006545f
C1342 VDD.n274 VSS 0.01473f
C1343 VDD.t186 VSS 0.033554f
C1344 VDD.n275 VSS 0.056186f
C1345 VDD.t15 VSS 0.004472f
C1346 VDD.n276 VSS 0.011514f
C1347 VDD.n277 VSS 0.019201f
C1348 VDD.t46 VSS 0.004509f
C1349 VDD.t196 VSS 0.009569f
C1350 VDD.n279 VSS 0.024536f
C1351 VDD.t47 VSS 0.004509f
C1352 VDD.n280 VSS 0.012134f
C1353 VDD.t191 VSS 0.018664f
C1354 VDD.n281 VSS 0.016882f
C1355 VDD.n282 VSS 0.002154f
C1356 VDD.n283 VSS 0.006059f
C1357 VDD.t64 VSS 0.004472f
C1358 VDD.n284 VSS 0.004409f
C1359 VDD.t57 VSS 0.004509f
C1360 VDD.t194 VSS 0.009569f
C1361 VDD.n286 VSS 0.024536f
C1362 VDD.t58 VSS 0.004509f
C1363 VDD.n287 VSS 0.013365f
C1364 VDD.t39 VSS 0.004509f
C1365 VDD.t176 VSS 0.009569f
C1366 VDD.n289 VSS 0.024536f
C1367 VDD.t40 VSS 0.004509f
C1368 VDD.n290 VSS 0.013365f
C1369 VDD.n291 VSS 0.011265f
C1370 VDD.n292 VSS 0.004909f
C1371 VDD.n293 VSS 0.006786f
C1372 VDD.n294 VSS 0.002474f
C1373 VDD.n295 VSS 0.001771f
C1374 VDD.n296 VSS 0.003159f
C1375 VDD.n297 VSS 0.001417f
C1376 VDD.n298 VSS 0.002767f
C1377 VDD.n299 VSS 0.001771f
C1378 VDD.n300 VSS 0.00201f
C1379 VDD.n301 VSS 0.001838f
C1380 VDD.n302 VSS 0.014674f
C1381 VDD.n303 VSS 0.011685f
C1382 VDD.n304 VSS 0.00135f
C1383 VDD.n305 VSS 0.002154f
C1384 VDD.n306 VSS 0.001771f
C1385 VDD.n307 VSS 0.002767f
C1386 VDD.n308 VSS 0.003054f
C1387 VDD.n309 VSS 0.114872f
C1388 VDD.n311 VSS 0.00308f
C1389 VDD.n312 VSS 0.003159f
C1390 VDD.n313 VSS 0.001771f
C1391 VDD.n314 VSS 0.00201f
C1392 VDD.n315 VSS 0.006059f
C1393 VDD.t36 VSS 0.045885f
C1394 VDD.t110 VSS 0.011175f
C1395 VDD.t161 VSS 0.016593f
C1396 VDD.t152 VSS 0.016085f
C1397 VDD.t141 VSS 0.0149f
C1398 VDD.t7 VSS 0.037927f
C1399 VDD.t173 VSS 0.030138f
C1400 VDD.t137 VSS 0.016085f
C1401 VDD.t75 VSS 0.026583f
C1402 VDD.t95 VSS 0.019641f
C1403 VDD.t131 VSS 0.0149f
C1404 VDD.t3 VSS 0.016085f
C1405 VDD.t156 VSS 0.026583f
C1406 VDD.t50 VSS 0.060277f
C1407 VDD.t22 VSS 0.022858f
C1408 VDD.t168 VSS 0.032001f
C1409 VDD.t93 VSS 0.047917f
C1410 VDD.t129 VSS 0.047917f
C1411 VDD.t116 VSS 0.040297f
C1412 VDD.t149 VSS 0.020487f
C1413 VDD.t25 VSS 0.016085f
C1414 VDD.t135 VSS 0.027091f
C1415 VDD.t41 VSS 0.072976f
C1416 VDD.t19 VSS 0.075007f
C1417 VDD.n316 VSS 0.036145f
C1418 VDD.n317 VSS 0.019586f
C1419 VDD.t48 VSS 0.004472f
C1420 VDD.t197 VSS 0.018829f
C1421 VDD.n319 VSS 0.032712f
C1422 VDD.t49 VSS 0.004472f
C1423 VDD.n320 VSS 0.01877f
C1424 VDD.n321 VSS 0.001838f
C1425 VDD.n322 VSS 0.001838f
C1426 VDD.n323 VSS 0.005284f
C1427 VDD.t184 VSS 0.018664f
C1428 VDD.t150 VSS 0.002858f
C1429 VDD.t136 VSS 8.29e-19
C1430 VDD.n324 VSS 0.00309f
C1431 VDD.t26 VSS 0.004472f
C1432 VDD.n325 VSS 0.007877f
C1433 VDD.n326 VSS 0.005284f
C1434 VDD.t130 VSS 0.002858f
C1435 VDD.t117 VSS 8.29e-19
C1436 VDD.n327 VSS 0.00309f
C1437 VDD.n328 VSS 0.00666f
C1438 VDD.n329 VSS 0.005284f
C1439 VDD.t185 VSS 0.065173f
C1440 VDD.t169 VSS 0.002858f
C1441 VDD.t94 VSS 8.29e-19
C1442 VDD.n330 VSS 0.00309f
C1443 VDD.n331 VSS 0.006347f
C1444 VDD.n332 VSS 0.001771f
C1445 VDD.n333 VSS 0.003159f
C1446 VDD.n334 VSS 0.001417f
C1447 VDD.n335 VSS 0.002642f
C1448 VDD.t187 VSS 0.018664f
C1449 VDD.n336 VSS 0.018051f
C1450 VDD.n337 VSS 0.002787f
C1451 VDD.n338 VSS 0.002817f
C1452 VDD.n339 VSS 0.005284f
C1453 VDD.t162 VSS 8.29e-19
C1454 VDD.t142 VSS 0.002858f
C1455 VDD.n340 VSS 0.00309f
C1456 VDD.n341 VSS 0.00481f
C1457 VDD.t111 VSS 6.78e-19
C1458 VDD.t153 VSS 0.00103f
C1459 VDD.n342 VSS 0.001759f
C1460 VDD.t65 VSS 0.004509f
C1461 VDD.t190 VSS 0.009569f
C1462 VDD.n344 VSS 0.024536f
C1463 VDD.t66 VSS 0.004509f
C1464 VDD.n345 VSS 0.013365f
C1465 VDD.t37 VSS 0.004509f
C1466 VDD.t195 VSS 0.009569f
C1467 VDD.n347 VSS 0.024536f
C1468 VDD.t38 VSS 0.004509f
C1469 VDD.n348 VSS 0.013365f
C1470 VDD.n349 VSS 0.011306f
C1471 VDD.n350 VSS 0.002642f
C1472 VDD.n351 VSS 0.001771f
C1473 VDD.n352 VSS 0.003159f
C1474 VDD.n353 VSS 0.001417f
C1475 VDD.n354 VSS 0.0021f
C1476 VDD.n355 VSS 0.003054f
C1477 VDD.n356 VSS 0.002767f
C1478 VDD.n357 VSS 0.001771f
C1479 VDD.n358 VSS 0.001895f
C1480 VDD.n359 VSS 0.001838f
C1481 VDD.n360 VSS 0.001838f
C1482 VDD.n361 VSS 0.002642f
C1483 VDD.n362 VSS 0.001771f
C1484 VDD.n363 VSS 0.001417f
C1485 VDD.n364 VSS 0.003159f
C1486 VDD.n365 VSS 0.003054f
C1487 VDD.n366 VSS 0.002767f
C1488 VDD.n367 VSS 3.49e-19
C1489 VDD.n368 VSS 0.001838f
C1490 VDD.n369 VSS 0.001556f
C1491 VDD.n370 VSS 0.00444f
C1492 VDD.n371 VSS 4.17e-19
C1493 VDD.n372 VSS 0.004796f
C1494 VDD.n373 VSS 0.005284f
C1495 VDD.n374 VSS 0.001368f
C1496 VDD.n375 VSS 0.002831f
C1497 VDD.n376 VSS 0.002987f
C1498 VDD.t8 VSS 9.3e-19
C1499 VDD.n377 VSS 0.002638f
C1500 VDD.t138 VSS 0.003822f
C1501 VDD.n378 VSS 0.003518f
C1502 VDD.n379 VSS 0.00314f
C1503 VDD.t174 VSS 8.29e-19
C1504 VDD.t76 VSS 0.002858f
C1505 VDD.n380 VSS 0.003049f
C1506 VDD.n381 VSS 0.003043f
C1507 VDD.n382 VSS 0.002625f
C1508 VDD.n383 VSS 0.005284f
C1509 VDD.n384 VSS 0.005284f
C1510 VDD.n385 VSS 0.00313f
C1511 VDD.n386 VSS 0.001434f
C1512 VDD.t96 VSS 0.001371f
C1513 VDD.t4 VSS 0.001371f
C1514 VDD.n387 VSS 0.003045f
C1515 VDD.t132 VSS 8.29e-19
C1516 VDD.t157 VSS 0.002858f
C1517 VDD.n388 VSS 0.003049f
C1518 VDD.n389 VSS 0.002437f
C1519 VDD.n390 VSS 0.008432f
C1520 VDD.n391 VSS 0.004796f
C1521 VDD.n392 VSS 0.005284f
C1522 VDD.n393 VSS 0.00313f
C1523 VDD.n394 VSS 0.002697f
C1524 VDD.t23 VSS 0.004921f
C1525 VDD.n395 VSS 0.003542f
C1526 VDD.t51 VSS 0.004472f
C1527 VDD.n396 VSS 0.010271f
C1528 VDD.n397 VSS 0.007784f
C1529 VDD.n398 VSS 0.002642f
C1530 VDD.n399 VSS 0.003819f
C1531 VDD.n400 VSS 0.001771f
C1532 VDD.n401 VSS 0.003054f
C1533 VDD.n402 VSS 0.002767f
C1534 VDD.n403 VSS 0.002646f
C1535 VDD.n404 VSS 0.001838f
C1536 VDD.n405 VSS 0.013995f
C1537 VDD.n406 VSS 0.01912f
C1538 VDD.t52 VSS 0.004472f
C1539 VDD.n407 VSS 0.005606f
C1540 VDD.n408 VSS 0.008033f
C1541 VDD.n409 VSS 0.001838f
C1542 VDD.n410 VSS 0.001091f
C1543 VDD.n411 VSS 0.002585f
C1544 VDD.n412 VSS 0.001895f
C1545 VDD.n413 VSS 0.001771f
C1546 VDD.n414 VSS 0.001417f
C1547 VDD.n415 VSS 0.003159f
C1548 VDD.n416 VSS 0.003054f
C1549 VDD.n417 VSS 0.001443f
C1550 VDD.n418 VSS 3.54e-19
C1551 VDD.n419 VSS 0.002297f
C1552 VDD.n420 VSS 0.004193f
C1553 VDD.n421 VSS 0.00666f
C1554 VDD.n422 VSS 0.003475f
C1555 VDD.n423 VSS 0.005431f
C1556 VDD.n424 VSS 0.030297f
C1557 VDD.n425 VSS 0.005103f
C1558 VDD.n426 VSS 0.005284f
C1559 VDD.n427 VSS 0.005284f
C1560 VDD.n428 VSS 0.005284f
C1561 VDD.n429 VSS 0.003728f
C1562 VDD.n430 VSS 0.006987f
C1563 VDD.t24 VSS 0.004921f
C1564 VDD.n431 VSS 0.003424f
C1565 VDD.n432 VSS 0.002582f
C1566 VDD.n433 VSS 0.005198f
C1567 VDD.n434 VSS 0.00313f
C1568 VDD.n435 VSS 0.004796f
C1569 VDD.n436 VSS 0.010554f
C1570 VDD.n437 VSS 0.01081f
C1571 VDD.n438 VSS 0.006332f
C1572 VDD.n439 VSS 0.016882f
C1573 VDD.t27 VSS 0.004472f
C1574 VDD.n440 VSS 0.004409f
C1575 VDD.n441 VSS 0.004909f
C1576 VDD.n442 VSS 0.003274f
C1577 VDD.n443 VSS 0.002843f
C1578 VDD.n444 VSS 0.001813f
C1579 VDD.n445 VSS 0.002741f
C1580 VDD.n446 VSS 0.001417f
C1581 VDD.n447 VSS 0.002642f
C1582 VDD.n448 VSS 0.001771f
C1583 VDD.n449 VSS 0.003159f
C1584 VDD.n450 VSS 0.001417f
C1585 VDD.n451 VSS 0.001771f
C1586 VDD.n452 VSS 0.002154f
C1587 VDD.n453 VSS 5.46e-19
C1588 VDD.t20 VSS 0.004472f
C1589 VDD.t179 VSS 0.018829f
C1590 VDD.n455 VSS 0.032712f
C1591 VDD.t21 VSS 0.004472f
C1592 VDD.n456 VSS 0.01877f
C1593 VDD.t42 VSS 0.004509f
C1594 VDD.t178 VSS 0.009569f
C1595 VDD.n458 VSS 0.024536f
C1596 VDD.t43 VSS 0.004509f
C1597 VDD.n459 VSS 0.013365f
C1598 VDD.t59 VSS 0.004509f
C1599 VDD.t183 VSS 0.009569f
C1600 VDD.n461 VSS 0.024536f
C1601 VDD.t60 VSS 0.004509f
C1602 VDD.n462 VSS 0.013365f
C1603 VDD.n463 VSS 0.011004f
C1604 VDD.n464 VSS 0.015879f
C1605 VDD.n465 VSS 0.006786f
C1606 VDD.n466 VSS 0.002474f
C1607 VDD.n467 VSS 0.002741f
C1608 VDD.n468 VSS 0.00308f
C1609 VDD.n469 VSS 0.115638f
C1610 VDD.n470 VSS 0.026229f
C1611 VDD.n471 VSS 0.075814f
C1612 VDD.n472 VSS 0.360185f
C1613 VDD.n473 VSS 0.075814f
C1614 VDD.n474 VSS 0.026229f
C1615 VDD.n475 VSS 0.384936f
C1616 VDD.n476 VSS 0.067851f
C1617 VDD.n477 VSS 0.075814f
C1618 VDD.n478 VSS 0.122169f
C1619 VDD.n479 VSS 0.100437f
C1620 VDD.n480 VSS 1.93e-19
C1621 VDD.n481 VSS 0.032316f
C1622 VDD.n482 VSS 0.060473f
C1623 VDD.n483 VSS 0.068782f
C1624 VDD.n484 VSS 0.050377f
C1625 VDD.t171 VSS 0.555684f
C1626 VDD.n485 VSS 0.102743f
C1627 VDD.n487 VSS 0.417917f
C1628 VDD.n488 VSS 0.050377f
C1629 VDD.n490 VSS 0.417917f
C1630 VDD.n491 VSS 0.049622f
C1631 VDD.n492 VSS 0.030592f
C1632 VDD.n493 VSS 0.005583f
C1633 VDD.n494 VSS 0.005464f
C1634 VDD.n495 VSS 0.082022f
C1635 VDD.n496 VSS 0.050682f
C1636 VDD.n497 VSS 0.030459f
C1637 VDD.n498 VSS 0.005613f
C1638 VDD.n499 VSS 0.417917f
C1639 VDD.n500 VSS 0.417917f
C1640 VDD.n501 VSS 0.049622f
C1641 VDD.n502 VSS 0.032078f
C1642 VDD.n503 VSS 0.060473f
C1643 VDD.n504 VSS 0.102743f
C1644 VDD.n505 VSS 0.068782f
C1645 VDD.n506 VSS 0.050377f
C1646 VDD.t85 VSS 0.555684f
C1647 VDD.n509 VSS 0.050377f
C1648 VDD.n510 VSS 0.00177f
C1649 VDD.n511 VSS 0.004f
C1650 VDD.n512 VSS 0.074678f
C1651 VDD.n513 VSS 0.051989f
C1652 VDD.n514 VSS 0.030561f
C1653 VDD.n515 VSS 0.005613f
C1654 VDD.n516 VSS 0.417917f
C1655 VDD.n517 VSS 0.417917f
C1656 VDD.n518 VSS 0.049622f
C1657 VDD.n519 VSS 0.032078f
C1658 VDD.n520 VSS 0.060473f
C1659 VDD.n521 VSS 0.102743f
C1660 VDD.n522 VSS 0.068782f
C1661 VDD.n523 VSS 0.050377f
C1662 VDD.t172 VSS 0.555684f
C1663 VDD.n526 VSS 0.050377f
C1664 VDD.n527 VSS 0.001668f
C1665 VDD.n528 VSS 0.003994f
C1666 VDD.n529 VSS 0.076174f
C1667 VDD.n530 VSS 0.06566f
C1668 VDD.n531 VSS 0.102743f
C1669 VDD.n532 VSS 0.023085f
C1670 VDD.n533 VSS 0.049622f
C1671 VDD.n534 VSS 0.417917f
C1672 VDD.n535 VSS 0.417917f
C1673 VDD.n536 VSS 0.068782f
C1674 VDD.n537 VSS 0.050377f
C1675 VDD.t163 VSS 0.555684f
C1676 VDD.n540 VSS 0.050377f
C1677 VDD.n541 VSS 2.14e-19
C1678 VDD.n542 VSS 0.030592f
C1679 VDD.n543 VSS 0.005562f
C1680 VDD.n544 VSS 0.060473f
C1681 VDD.n545 VSS 0.032334f
C1682 passgatesCtrl_0.net2.n0 VSS 0.241262f
C1683 passgatesCtrl_0.net2.t0 VSS 0.052358f
C1684 passgatesCtrl_0.net2.n1 VSS 0.013973f
C1685 passgatesCtrl_0.net2.t3 VSS 0.019097f
C1686 passgatesCtrl_0.net2.t7 VSS 0.012934f
C1687 passgatesCtrl_0.net2.n2 VSS 0.052064f
C1688 passgatesCtrl_0.net2.t1 VSS 0.032964f
C1689 passgatesCtrl_0.net2.n3 VSS 0.011845f
C1690 passgatesCtrl_0.net2.n4 VSS 0.031329f
C1691 passgatesCtrl_0.net2.t6 VSS 0.022133f
C1692 passgatesCtrl_0.net2.t15 VSS 0.05173f
C1693 passgatesCtrl_0.net2.n5 VSS 0.062148f
C1694 passgatesCtrl_0.net2.t10 VSS 0.014926f
C1695 passgatesCtrl_0.net2.t19 VSS 0.023903f
C1696 passgatesCtrl_0.net2.n6 VSS 0.04516f
C1697 passgatesCtrl_0.net2.n7 VSS 0.063372f
C1698 passgatesCtrl_0.net2.t16 VSS 0.010242f
C1699 passgatesCtrl_0.net2.t2 VSS 0.012844f
C1700 passgatesCtrl_0.net2.n8 VSS 0.047082f
C1701 passgatesCtrl_0.net2.n9 VSS 0.216971f
C1702 passgatesCtrl_0.net2.n10 VSS 0.157732f
C1703 passgatesCtrl_0.net2.t17 VSS 0.010314f
C1704 passgatesCtrl_0.net2.t9 VSS 0.012486f
C1705 passgatesCtrl_0.net2.n11 VSS 0.041569f
C1706 passgatesCtrl_0.net2.n12 VSS 0.009518f
C1707 passgatesCtrl_0.net2.t12 VSS 0.016063f
C1708 passgatesCtrl_0.net2.t8 VSS 0.011059f
C1709 passgatesCtrl_0.net2.n13 VSS 0.038188f
C1710 passgatesCtrl_0.net2.n14 VSS 0.010881f
C1711 passgatesCtrl_0.net2.t4 VSS 0.014893f
C1712 passgatesCtrl_0.net2.t11 VSS 0.023864f
C1713 passgatesCtrl_0.net2.n15 VSS 0.047068f
C1714 passgatesCtrl_0.net2.n16 VSS 0.061051f
C1715 passgatesCtrl_0.net2.n17 VSS 0.168444f
C1716 passgatesCtrl_0.net2.t18 VSS 0.01039f
C1717 passgatesCtrl_0.net2.t14 VSS 0.021912f
C1718 passgatesCtrl_0.net2.n18 VSS 0.078683f
C1719 passgatesCtrl_0.net2.n19 VSS 0.017108f
C1720 passgatesCtrl_0.net2.n20 VSS 0.16814f
C1721 passgatesCtrl_0.net2.t5 VSS 0.013096f
C1722 passgatesCtrl_0.net2.t13 VSS 0.019286f
C1723 passgatesCtrl_0.net2.n21 VSS 0.045566f
C1724 passgatesCtrl_0.net2.n22 VSS 0.010906f
C1725 passgatesCtrl_0.net2.n23 VSS 0.364405f
C1726 passgatesCtrl_0.net2.n24 VSS 0.041229f
.ends

